module miter ( 
    RI2b1c4342d4e0_65, RI2b1c4342c5e0_33, RI2b1c4342b6e0_1,
    RI2b1c4342d558_66, RI2b1c4342d5d0_67, RI2b1c4342d648_68,
    RI2b1c4342d6c0_69, RI2b1c4342d738_70, RI2b1c4342d7b0_71,
    RI2b1c4342d828_72, RI2b1c4342d8a0_73, RI2b1c4342d918_74,
    RI2b1c4342d990_75, RI2b1c4342da08_76, RI2b1c4342da80_77,
    RI2b1c4342daf8_78, RI2b1c4342db70_79, RI2b1c4342dbe8_80,
    RI2b1c4342dc60_81, RI2b1c4342dcd8_82, RI2b1c4342dd50_83,
    RI2b1c4342ddc8_84, RI2b1c4342de40_85, RI2b1c4342deb8_86,
    RI2b1c4342df30_87, RI2b1c4342dfa8_88, RI2b1c4342e020_89,
    RI2b1c4342e098_90, RI2b1c4342e110_91, RI2b1c4342e188_92,
    RI2b1c4342e200_93, RI2b1c4342e278_94, RI2b1c4342e2f0_95,
    RI2b1c4342e368_96, RI2b1c4342c658_34, RI2b1c4342b758_2,
    RI2b1c4342c6d0_35, RI2b1c4342b7d0_3, RI2b1c4342c748_36,
    RI2b1c4342b848_4, RI2b1c4342c7c0_37, RI2b1c4342b8c0_5,
    RI2b1c4342c838_38, RI2b1c4342b938_6, RI2b1c4342c8b0_39,
    RI2b1c4342b9b0_7, RI2b1c4342c928_40, RI2b1c4342ba28_8,
    RI2b1c4342c9a0_41, RI2b1c4342baa0_9, RI2b1c4342ca18_42,
    RI2b1c4342bb18_10, RI2b1c4342ca90_43, RI2b1c4342bb90_11,
    RI2b1c4342cb08_44, RI2b1c4342bc08_12, RI2b1c4342cb80_45,
    RI2b1c4342bc80_13, RI2b1c4342cbf8_46, RI2b1c4342bcf8_14,
    RI2b1c4342cc70_47, RI2b1c4342bd70_15, RI2b1c4342cce8_48,
    RI2b1c4342bde8_16, RI2b1c4342cd60_49, RI2b1c4342be60_17,
    RI2b1c4342cdd8_50, RI2b1c4342bed8_18, RI2b1c4342ce50_51,
    RI2b1c4342bf50_19, RI2b1c4342cec8_52, RI2b1c4342bfc8_20,
    RI2b1c4342cf40_53, RI2b1c4342c040_21, RI2b1c4342cfb8_54,
    RI2b1c4342c0b8_22, RI2b1c4342d030_55, RI2b1c4342c130_23,
    RI2b1c4342d0a8_56, RI2b1c4342c1a8_24, RI2b1c4342d120_57,
    RI2b1c4342c220_25, RI2b1c4342d198_58, RI2b1c4342c298_26,
    RI2b1c4342d210_59, RI2b1c4342c310_27, RI2b1c4342d288_60,
    RI2b1c4342c388_28, RI2b1c4342d300_61, RI2b1c4342c400_29,
    RI2b1c4342d378_62, RI2b1c4342c478_30, RI2b1c4342d3f0_63,
    RI2b1c4342c4f0_31, RI2b1c4342d468_64, RI2b1c4342c568_32,
    eq  );
  input  RI2b1c4342d4e0_65, RI2b1c4342c5e0_33, RI2b1c4342b6e0_1,
    RI2b1c4342d558_66, RI2b1c4342d5d0_67, RI2b1c4342d648_68,
    RI2b1c4342d6c0_69, RI2b1c4342d738_70, RI2b1c4342d7b0_71,
    RI2b1c4342d828_72, RI2b1c4342d8a0_73, RI2b1c4342d918_74,
    RI2b1c4342d990_75, RI2b1c4342da08_76, RI2b1c4342da80_77,
    RI2b1c4342daf8_78, RI2b1c4342db70_79, RI2b1c4342dbe8_80,
    RI2b1c4342dc60_81, RI2b1c4342dcd8_82, RI2b1c4342dd50_83,
    RI2b1c4342ddc8_84, RI2b1c4342de40_85, RI2b1c4342deb8_86,
    RI2b1c4342df30_87, RI2b1c4342dfa8_88, RI2b1c4342e020_89,
    RI2b1c4342e098_90, RI2b1c4342e110_91, RI2b1c4342e188_92,
    RI2b1c4342e200_93, RI2b1c4342e278_94, RI2b1c4342e2f0_95,
    RI2b1c4342e368_96, RI2b1c4342c658_34, RI2b1c4342b758_2,
    RI2b1c4342c6d0_35, RI2b1c4342b7d0_3, RI2b1c4342c748_36,
    RI2b1c4342b848_4, RI2b1c4342c7c0_37, RI2b1c4342b8c0_5,
    RI2b1c4342c838_38, RI2b1c4342b938_6, RI2b1c4342c8b0_39,
    RI2b1c4342b9b0_7, RI2b1c4342c928_40, RI2b1c4342ba28_8,
    RI2b1c4342c9a0_41, RI2b1c4342baa0_9, RI2b1c4342ca18_42,
    RI2b1c4342bb18_10, RI2b1c4342ca90_43, RI2b1c4342bb90_11,
    RI2b1c4342cb08_44, RI2b1c4342bc08_12, RI2b1c4342cb80_45,
    RI2b1c4342bc80_13, RI2b1c4342cbf8_46, RI2b1c4342bcf8_14,
    RI2b1c4342cc70_47, RI2b1c4342bd70_15, RI2b1c4342cce8_48,
    RI2b1c4342bde8_16, RI2b1c4342cd60_49, RI2b1c4342be60_17,
    RI2b1c4342cdd8_50, RI2b1c4342bed8_18, RI2b1c4342ce50_51,
    RI2b1c4342bf50_19, RI2b1c4342cec8_52, RI2b1c4342bfc8_20,
    RI2b1c4342cf40_53, RI2b1c4342c040_21, RI2b1c4342cfb8_54,
    RI2b1c4342c0b8_22, RI2b1c4342d030_55, RI2b1c4342c130_23,
    RI2b1c4342d0a8_56, RI2b1c4342c1a8_24, RI2b1c4342d120_57,
    RI2b1c4342c220_25, RI2b1c4342d198_58, RI2b1c4342c298_26,
    RI2b1c4342d210_59, RI2b1c4342c310_27, RI2b1c4342d288_60,
    RI2b1c4342c388_28, RI2b1c4342d300_61, RI2b1c4342c400_29,
    RI2b1c4342d378_62, RI2b1c4342c478_30, RI2b1c4342d3f0_63,
    RI2b1c4342c4f0_31, RI2b1c4342d468_64, RI2b1c4342c568_32;
  output eq;
  wire new_n98_, new_n99_, new_n100_, new_n101_, new_n102_, new_n103_,
    new_n104_, new_n105_, new_n106_, new_n107_, new_n108_, new_n109_,
    new_n110_, new_n111_, new_n112_, new_n113_, new_n114_, new_n115_,
    new_n116_, new_n117_, new_n118_, new_n119_, new_n120_, new_n121_,
    new_n122_, new_n123_, new_n124_, new_n125_, new_n126_, new_n127_,
    new_n128_, new_n129_, new_n130_, new_n131_, new_n132_, new_n133_,
    new_n134_, new_n135_, new_n136_, new_n137_, new_n138_, new_n139_,
    new_n140_, new_n141_, new_n142_, new_n143_, new_n144_, new_n145_,
    new_n146_, new_n147_, new_n148_, new_n149_, new_n150_, new_n151_,
    new_n152_, new_n153_, new_n154_, new_n155_, new_n156_, new_n157_,
    new_n158_, new_n159_, new_n160_, new_n161_, new_n162_, new_n163_,
    new_n164_, new_n165_, new_n166_, new_n167_, new_n168_, new_n169_,
    new_n170_, new_n171_, new_n172_, new_n173_, new_n174_, new_n175_,
    new_n176_, new_n177_, new_n178_, new_n179_, new_n180_, new_n181_,
    new_n182_, new_n183_, new_n184_, new_n185_, new_n186_, new_n187_,
    new_n188_, new_n189_, new_n190_, new_n191_, new_n192_, new_n193_,
    new_n194_, new_n195_, new_n196_, new_n197_, new_n198_, new_n199_,
    new_n200_, new_n201_, new_n202_, new_n203_, new_n204_, new_n205_,
    new_n206_, new_n207_, new_n208_, new_n209_, new_n210_, new_n211_,
    new_n212_, new_n213_, new_n214_, new_n215_, new_n216_, new_n217_,
    new_n218_, new_n219_, new_n220_, new_n221_, new_n222_, new_n223_,
    new_n224_, new_n225_, new_n226_, new_n227_, new_n228_, new_n229_,
    new_n230_, new_n231_, new_n232_, new_n233_, new_n234_, new_n235_,
    new_n236_, new_n237_, new_n238_, new_n239_, new_n240_, new_n241_,
    new_n242_, new_n243_, new_n244_, new_n245_, new_n246_, new_n247_,
    new_n248_, new_n249_, new_n250_, new_n251_, new_n252_, new_n253_,
    new_n254_, new_n255_, new_n256_, new_n257_, new_n258_, new_n259_,
    new_n260_, new_n261_, new_n262_, new_n263_, new_n264_, new_n265_,
    new_n266_, new_n267_, new_n268_, new_n269_, new_n270_, new_n271_,
    new_n272_, new_n273_, new_n274_, new_n275_, new_n276_, new_n277_,
    new_n278_, new_n279_, new_n280_, new_n281_, new_n282_, new_n283_,
    new_n284_, new_n285_, new_n286_, new_n287_, new_n288_, new_n289_,
    new_n290_, new_n291_, new_n292_, new_n293_, new_n294_, new_n295_,
    new_n296_, new_n297_, new_n298_, new_n299_, new_n300_, new_n301_,
    new_n302_, new_n303_, new_n304_, new_n305_, new_n306_, new_n307_,
    new_n308_, new_n309_, new_n310_, new_n311_, new_n312_, new_n313_,
    new_n314_, new_n315_, new_n316_, new_n317_, new_n318_, new_n319_,
    new_n320_, new_n321_, new_n322_, new_n323_, new_n324_, new_n325_,
    new_n326_, new_n327_, new_n328_, new_n329_, new_n330_, new_n331_,
    new_n332_, new_n333_, new_n334_, new_n335_, new_n336_, new_n337_,
    new_n338_, new_n339_, new_n340_, new_n341_, new_n342_, new_n343_,
    new_n344_, new_n345_, new_n346_, new_n347_, new_n348_, new_n349_,
    new_n350_, new_n351_, new_n352_, new_n353_, new_n354_, new_n355_,
    new_n356_, new_n357_, new_n358_, new_n359_, new_n360_, new_n361_,
    new_n362_, new_n363_, new_n364_, new_n365_, new_n366_, new_n367_,
    new_n368_, new_n369_, new_n370_, new_n371_, new_n372_, new_n373_,
    new_n374_, new_n375_, new_n376_, new_n377_, new_n378_, new_n379_,
    new_n380_, new_n381_, new_n382_, new_n383_, new_n384_, new_n385_,
    new_n386_, new_n387_, new_n388_, new_n389_, new_n390_, new_n391_,
    new_n392_, new_n393_, new_n394_, new_n395_, new_n396_, new_n397_,
    new_n398_, new_n399_, new_n400_, new_n401_, new_n402_, new_n403_,
    new_n404_, new_n405_, new_n406_, new_n407_, new_n408_, new_n409_,
    new_n410_, new_n411_, new_n412_, new_n413_, new_n414_, new_n415_,
    new_n416_, new_n417_, new_n418_, new_n419_, new_n420_, new_n421_,
    new_n422_, new_n423_, new_n424_, new_n425_, new_n426_, new_n427_,
    new_n428_, new_n429_, new_n430_, new_n431_, new_n432_, new_n433_,
    new_n434_, new_n435_, new_n436_, new_n437_, new_n438_, new_n439_,
    new_n440_, new_n441_, new_n442_, new_n443_, new_n444_, new_n445_,
    new_n446_, new_n447_, new_n448_, new_n449_, new_n450_, new_n451_,
    new_n452_, new_n453_, new_n454_, new_n455_, new_n456_, new_n457_,
    new_n458_, new_n459_, new_n460_, new_n461_, new_n462_, new_n463_,
    new_n464_, new_n465_, new_n466_, new_n467_, new_n468_, new_n469_,
    new_n470_, new_n471_, new_n472_, new_n473_, new_n474_, new_n475_,
    new_n476_, new_n477_, new_n478_, new_n479_, new_n480_, new_n481_,
    new_n482_, new_n483_, new_n484_, new_n485_, new_n486_, new_n487_,
    new_n488_, new_n489_, new_n490_, new_n491_, new_n492_, new_n493_,
    new_n494_, new_n495_, new_n496_, new_n497_, new_n498_, new_n499_,
    new_n500_, new_n501_, new_n502_, new_n503_, new_n504_, new_n505_,
    new_n506_, new_n507_, new_n508_, new_n509_, new_n510_, new_n511_,
    new_n512_, new_n513_, new_n514_, new_n515_, new_n516_, new_n517_,
    new_n518_, new_n519_, new_n520_, new_n521_, new_n522_, new_n523_,
    new_n524_, new_n525_, new_n526_, new_n527_, new_n528_, new_n529_,
    new_n530_, new_n531_, new_n532_, new_n533_, new_n534_, new_n535_,
    new_n536_, new_n537_, new_n538_, new_n539_, new_n540_, new_n541_,
    new_n542_, new_n543_, new_n544_, new_n545_, new_n546_, new_n547_,
    new_n548_, new_n549_, new_n550_, new_n551_, new_n552_, new_n553_,
    new_n554_, new_n555_, new_n556_, new_n557_, new_n558_, new_n559_,
    new_n560_, new_n561_, new_n562_, new_n563_, new_n564_, new_n565_,
    new_n566_, new_n567_, new_n568_, new_n569_, new_n570_, new_n571_,
    new_n572_, new_n573_, new_n574_, new_n575_, new_n576_, new_n577_,
    new_n578_, new_n579_, new_n580_, new_n581_, new_n582_, new_n583_,
    new_n584_, new_n585_, new_n586_, new_n587_, new_n588_, new_n589_,
    new_n590_, new_n591_, new_n592_, new_n593_, new_n594_, new_n595_,
    new_n596_, new_n597_, new_n598_, new_n599_, new_n600_, new_n601_,
    new_n602_, new_n603_, new_n604_, new_n605_, new_n606_, new_n607_,
    new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n917_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n922_, new_n923_, new_n924_, new_n925_,
    new_n926_, new_n927_, new_n928_, new_n929_, new_n930_, new_n931_,
    new_n932_, new_n933_, new_n934_, new_n935_, new_n936_, new_n937_,
    new_n938_, new_n939_, new_n940_, new_n941_, new_n942_, new_n943_,
    new_n944_, new_n945_, new_n946_, new_n947_, new_n948_, new_n949_,
    new_n950_, new_n951_, new_n952_, new_n953_, new_n954_, new_n955_,
    new_n956_, new_n957_, new_n958_, new_n959_, new_n960_, new_n961_,
    new_n962_, new_n963_, new_n964_, new_n965_, new_n966_, new_n967_,
    new_n968_, new_n969_, new_n970_, new_n971_, new_n972_, new_n973_,
    new_n974_, new_n975_, new_n976_, new_n977_, new_n978_, new_n979_,
    new_n980_, new_n981_, new_n982_, new_n983_, new_n984_, new_n985_,
    new_n986_, new_n987_, new_n988_, new_n989_, new_n990_, new_n991_,
    new_n992_, new_n993_, new_n994_, new_n995_, new_n996_, new_n997_,
    new_n998_, new_n999_, new_n1000_, new_n1001_, new_n1002_, new_n1003_,
    new_n1004_, new_n1005_, new_n1006_, new_n1007_, new_n1008_, new_n1009_,
    new_n1010_, new_n1011_, new_n1012_, new_n1013_, new_n1014_, new_n1015_,
    new_n1016_, new_n1017_, new_n1018_, new_n1019_, new_n1020_, new_n1021_,
    new_n1022_, new_n1023_, new_n1024_, new_n1025_, new_n1026_, new_n1027_,
    new_n1028_, new_n1029_, new_n1030_, new_n1031_, new_n1032_, new_n1033_,
    new_n1034_, new_n1035_, new_n1036_, new_n1037_, new_n1038_, new_n1039_,
    new_n1040_, new_n1041_, new_n1042_, new_n1043_, new_n1044_, new_n1045_,
    new_n1046_, new_n1047_, new_n1048_, new_n1049_, new_n1050_, new_n1051_,
    new_n1052_, new_n1053_, new_n1054_, new_n1055_, new_n1056_, new_n1057_,
    new_n1058_, new_n1059_, new_n1060_, new_n1061_, new_n1062_, new_n1063_,
    new_n1064_, new_n1065_, new_n1066_, new_n1067_, new_n1068_, new_n1069_,
    new_n1070_, new_n1071_, new_n1072_, new_n1073_, new_n1074_, new_n1075_,
    new_n1076_, new_n1077_, new_n1078_, new_n1079_, new_n1080_, new_n1081_,
    new_n1082_, new_n1083_, new_n1084_, new_n1085_, new_n1086_, new_n1087_,
    new_n1088_, new_n1089_, new_n1090_, new_n1091_, new_n1092_, new_n1093_,
    new_n1094_, new_n1095_, new_n1096_, new_n1097_, new_n1098_, new_n1099_,
    new_n1100_, new_n1101_, new_n1102_, new_n1103_, new_n1104_, new_n1105_,
    new_n1106_, new_n1107_, new_n1108_, new_n1109_, new_n1110_, new_n1111_,
    new_n1112_, new_n1113_, new_n1114_, new_n1115_, new_n1116_, new_n1117_,
    new_n1118_, new_n1119_, new_n1120_, new_n1121_, new_n1122_, new_n1123_,
    new_n1124_, new_n1125_, new_n1126_, new_n1127_, new_n1128_, new_n1129_,
    new_n1130_, new_n1131_, new_n1132_, new_n1133_, new_n1134_, new_n1135_,
    new_n1136_, new_n1137_, new_n1138_, new_n1139_, new_n1140_, new_n1141_,
    new_n1142_, new_n1143_, new_n1144_, new_n1145_, new_n1146_, new_n1147_,
    new_n1148_, new_n1149_, new_n1150_, new_n1151_, new_n1152_, new_n1153_,
    new_n1154_, new_n1155_, new_n1156_, new_n1157_, new_n1158_, new_n1159_,
    new_n1160_, new_n1161_, new_n1162_, new_n1163_, new_n1164_, new_n1165_,
    new_n1166_, new_n1167_, new_n1168_, new_n1169_, new_n1170_, new_n1171_,
    new_n1172_, new_n1173_, new_n1174_, new_n1175_, new_n1176_, new_n1177_,
    new_n1178_, new_n1179_, new_n1180_, new_n1181_, new_n1182_, new_n1183_,
    new_n1184_, new_n1185_, new_n1186_, new_n1187_, new_n1188_, new_n1189_,
    new_n1190_, new_n1191_, new_n1192_, new_n1193_, new_n1194_, new_n1195_,
    new_n1196_, new_n1197_, new_n1198_, new_n1199_, new_n1200_, new_n1201_,
    new_n1202_, new_n1203_, new_n1204_, new_n1205_, new_n1206_, new_n1207_,
    new_n1208_, new_n1209_, new_n1210_, new_n1211_, new_n1212_, new_n1213_,
    new_n1214_, new_n1215_, new_n1216_, new_n1217_, new_n1218_, new_n1219_,
    new_n1220_, new_n1221_, new_n1222_, new_n1223_, new_n1224_, new_n1225_,
    new_n1226_, new_n1227_, new_n1228_, new_n1229_, new_n1230_, new_n1231_,
    new_n1232_, new_n1233_, new_n1234_, new_n1235_, new_n1236_, new_n1237_,
    new_n1238_, new_n1239_, new_n1240_, new_n1241_, new_n1242_, new_n1243_,
    new_n1244_, new_n1245_, new_n1246_, new_n1247_, new_n1248_, new_n1249_,
    new_n1250_, new_n1251_, new_n1252_, new_n1253_, new_n1254_, new_n1255_,
    new_n1256_, new_n1257_, new_n1258_, new_n1259_, new_n1260_, new_n1261_,
    new_n1262_, new_n1263_, new_n1264_, new_n1265_, new_n1266_, new_n1267_,
    new_n1268_, new_n1269_, new_n1270_, new_n1271_, new_n1272_, new_n1273_,
    new_n1274_, new_n1275_, new_n1276_, new_n1277_, new_n1278_, new_n1279_,
    new_n1280_, new_n1281_, new_n1282_, new_n1283_, new_n1284_, new_n1285_,
    new_n1286_, new_n1287_, new_n1288_, new_n1289_, new_n1290_, new_n1291_,
    new_n1292_, new_n1293_, new_n1294_, new_n1295_, new_n1296_, new_n1297_,
    new_n1298_, new_n1299_, new_n1300_, new_n1301_, new_n1302_, new_n1303_,
    new_n1304_, new_n1305_, new_n1306_, new_n1307_, new_n1308_, new_n1309_,
    new_n1310_, new_n1311_, new_n1312_, new_n1313_, new_n1314_, new_n1315_,
    new_n1316_, new_n1317_, new_n1318_, new_n1319_, new_n1320_, new_n1321_,
    new_n1322_, new_n1323_, new_n1324_, new_n1325_, new_n1326_, new_n1327_,
    new_n1328_, new_n1329_, new_n1330_, new_n1331_, new_n1332_, new_n1333_,
    new_n1334_, new_n1335_, new_n1336_, new_n1337_, new_n1338_, new_n1339_,
    new_n1340_, new_n1341_, new_n1342_, new_n1343_, new_n1344_, new_n1345_,
    new_n1346_, new_n1347_, new_n1348_, new_n1349_, new_n1350_, new_n1351_,
    new_n1352_, new_n1353_, new_n1354_, new_n1355_, new_n1356_, new_n1357_,
    new_n1358_, new_n1359_, new_n1360_, new_n1361_, new_n1362_, new_n1363_,
    new_n1364_, new_n1365_, new_n1366_, new_n1367_, new_n1368_, new_n1369_,
    new_n1370_, new_n1371_, new_n1372_, new_n1373_, new_n1374_, new_n1375_,
    new_n1376_, new_n1377_, new_n1378_, new_n1379_, new_n1380_, new_n1381_,
    new_n1382_, new_n1383_, new_n1384_, new_n1385_, new_n1386_, new_n1387_,
    new_n1388_, new_n1389_, new_n1390_, new_n1391_, new_n1392_, new_n1393_,
    new_n1394_, new_n1395_, new_n1396_, new_n1397_, new_n1398_, new_n1399_,
    new_n1400_, new_n1401_, new_n1402_, new_n1403_, new_n1404_, new_n1405_,
    new_n1406_, new_n1407_, new_n1408_, new_n1409_, new_n1410_, new_n1411_,
    new_n1412_, new_n1413_, new_n1414_, new_n1415_, new_n1416_, new_n1417_,
    new_n1418_, new_n1419_, new_n1420_, new_n1421_, new_n1422_, new_n1423_,
    new_n1424_, new_n1425_, new_n1426_, new_n1427_, new_n1428_, new_n1429_,
    new_n1430_, new_n1431_, new_n1432_, new_n1433_, new_n1434_, new_n1435_,
    new_n1436_, new_n1437_, new_n1438_, new_n1439_, new_n1440_, new_n1441_,
    new_n1442_, new_n1443_, new_n1444_, new_n1445_, new_n1446_, new_n1447_,
    new_n1448_, new_n1449_, new_n1450_, new_n1451_, new_n1452_, new_n1453_,
    new_n1454_, new_n1455_, new_n1456_, new_n1457_, new_n1458_, new_n1459_,
    new_n1460_, new_n1461_, new_n1462_, new_n1463_, new_n1464_, new_n1465_,
    new_n1466_, new_n1467_, new_n1468_, new_n1469_, new_n1470_, new_n1471_,
    new_n1472_, new_n1473_, new_n1474_, new_n1475_, new_n1476_, new_n1477_,
    new_n1478_, new_n1479_, new_n1480_, new_n1481_, new_n1482_, new_n1483_,
    new_n1484_, new_n1485_, new_n1486_, new_n1487_, new_n1488_, new_n1489_,
    new_n1490_, new_n1491_, new_n1492_, new_n1493_, new_n1494_, new_n1495_,
    new_n1496_, new_n1497_, new_n1498_, new_n1499_, new_n1500_, new_n1501_,
    new_n1502_, new_n1503_, new_n1504_, new_n1505_, new_n1506_, new_n1507_,
    new_n1508_, new_n1509_, new_n1510_, new_n1511_, new_n1512_, new_n1513_,
    new_n1514_, new_n1515_, new_n1516_, new_n1517_, new_n1518_, new_n1519_,
    new_n1520_, new_n1521_, new_n1522_, new_n1523_, new_n1524_, new_n1525_,
    new_n1526_, new_n1527_, new_n1528_, new_n1529_, new_n1530_, new_n1531_,
    new_n1532_, new_n1533_, new_n1534_, new_n1535_, new_n1536_, new_n1537_,
    new_n1538_, new_n1539_, new_n1540_, new_n1541_, new_n1542_, new_n1543_,
    new_n1544_, new_n1545_, new_n1546_, new_n1547_, new_n1548_, new_n1549_,
    new_n1550_, new_n1551_, new_n1552_, new_n1553_, new_n1554_, new_n1555_,
    new_n1556_, new_n1557_, new_n1558_, new_n1559_, new_n1560_, new_n1561_,
    new_n1562_, new_n1563_, new_n1564_, new_n1565_, new_n1566_, new_n1567_,
    new_n1568_, new_n1569_, new_n1570_, new_n1571_, new_n1572_, new_n1573_,
    new_n1574_, new_n1575_, new_n1576_, new_n1577_, new_n1578_, new_n1579_,
    new_n1580_, new_n1581_, new_n1582_, new_n1583_, new_n1584_, new_n1585_,
    new_n1586_, new_n1587_, new_n1588_, new_n1589_, new_n1590_, new_n1591_,
    new_n1592_, new_n1593_, new_n1594_, new_n1595_, new_n1596_, new_n1597_,
    new_n1598_, new_n1599_, new_n1600_, new_n1601_, new_n1602_, new_n1603_,
    new_n1604_, new_n1605_, new_n1606_, new_n1607_, new_n1608_, new_n1609_,
    new_n1610_, new_n1611_, new_n1612_, new_n1613_, new_n1614_, new_n1615_,
    new_n1616_, new_n1617_, new_n1618_, new_n1619_, new_n1620_, new_n1621_,
    new_n1622_, new_n1623_, new_n1624_, new_n1625_, new_n1626_, new_n1627_,
    new_n1628_, new_n1629_, new_n1630_, new_n1631_, new_n1632_, new_n1633_,
    new_n1634_, new_n1635_, new_n1636_, new_n1637_, new_n1638_, new_n1639_,
    new_n1640_, new_n1641_, new_n1642_, new_n1643_, new_n1644_, new_n1645_,
    new_n1646_, new_n1647_, new_n1648_, new_n1649_, new_n1650_, new_n1651_,
    new_n1652_, new_n1653_, new_n1654_, new_n1655_, new_n1656_, new_n1657_,
    new_n1658_, new_n1659_, new_n1660_, new_n1661_, new_n1662_, new_n1663_,
    new_n1664_, new_n1665_, new_n1666_, new_n1667_, new_n1668_, new_n1669_,
    new_n1670_, new_n1671_, new_n1672_, new_n1673_, new_n1674_, new_n1675_,
    new_n1676_, new_n1677_, new_n1678_, new_n1679_, new_n1680_, new_n1681_,
    new_n1682_, new_n1683_, new_n1684_, new_n1685_, new_n1686_, new_n1687_,
    new_n1688_, new_n1689_, new_n1690_, new_n1691_, new_n1692_, new_n1693_,
    new_n1694_, new_n1695_, new_n1696_, new_n1697_, new_n1698_, new_n1699_,
    new_n1700_, new_n1701_, new_n1702_, new_n1703_, new_n1704_, new_n1705_,
    new_n1706_, new_n1707_, new_n1708_, new_n1709_, new_n1710_, new_n1711_,
    new_n1712_, new_n1713_, new_n1714_, new_n1715_, new_n1716_, new_n1717_,
    new_n1718_, new_n1719_, new_n1720_, new_n1721_, new_n1722_, new_n1723_,
    new_n1724_, new_n1725_, new_n1726_, new_n1727_, new_n1728_, new_n1729_,
    new_n1730_, new_n1731_, new_n1732_, new_n1733_, new_n1734_, new_n1735_,
    new_n1736_, new_n1737_, new_n1738_, new_n1739_, new_n1740_, new_n1741_,
    new_n1742_, new_n1743_, new_n1744_, new_n1745_, new_n1746_, new_n1747_,
    new_n1748_, new_n1749_, new_n1750_, new_n1751_, new_n1752_, new_n1753_,
    new_n1754_, new_n1755_, new_n1756_, new_n1757_, new_n1758_, new_n1759_,
    new_n1760_, new_n1761_, new_n1762_, new_n1763_, new_n1764_, new_n1765_,
    new_n1766_, new_n1767_, new_n1768_, new_n1769_, new_n1770_, new_n1771_,
    new_n1772_, new_n1773_, new_n1774_, new_n1775_, new_n1776_, new_n1777_,
    new_n1778_, new_n1779_, new_n1780_, new_n1781_, new_n1782_, new_n1783_,
    new_n1784_, new_n1785_, new_n1786_, new_n1787_, new_n1788_, new_n1789_,
    new_n1790_, new_n1791_, new_n1792_, new_n1793_, new_n1794_, new_n1795_,
    new_n1796_, new_n1797_, new_n1798_, new_n1799_, new_n1800_, new_n1801_,
    new_n1802_, new_n1803_, new_n1804_, new_n1805_, new_n1806_, new_n1807_,
    new_n1808_, new_n1809_, new_n1810_, new_n1811_, new_n1812_, new_n1813_,
    new_n1814_, new_n1815_, new_n1816_, new_n1817_, new_n1818_, new_n1819_,
    new_n1820_, new_n1821_, new_n1822_, new_n1823_, new_n1824_, new_n1825_,
    new_n1826_, new_n1827_, new_n1828_, new_n1829_, new_n1830_, new_n1831_,
    new_n1832_, new_n1833_, new_n1834_, new_n1835_, new_n1836_, new_n1837_,
    new_n1838_, new_n1839_, new_n1840_, new_n1841_, new_n1842_, new_n1843_,
    new_n1844_, new_n1845_, new_n1846_, new_n1847_, new_n1848_, new_n1849_,
    new_n1850_, new_n1851_, new_n1852_, new_n1853_, new_n1854_, new_n1855_,
    new_n1856_, new_n1857_, new_n1858_, new_n1859_, new_n1860_, new_n1861_,
    new_n1862_, new_n1863_, new_n1864_, new_n1865_, new_n1866_, new_n1867_,
    new_n1868_, new_n1869_, new_n1870_, new_n1871_, new_n1872_, new_n1873_,
    new_n1874_, new_n1875_, new_n1876_, new_n1877_, new_n1878_, new_n1879_,
    new_n1880_, new_n1881_, new_n1882_, new_n1883_, new_n1884_, new_n1885_,
    new_n1886_, new_n1887_, new_n1888_, new_n1889_, new_n1890_, new_n1891_,
    new_n1892_, new_n1893_, new_n1894_, new_n1895_, new_n1896_, new_n1897_,
    new_n1898_, new_n1899_, new_n1900_, new_n1901_, new_n1902_, new_n1903_,
    new_n1904_, new_n1905_, new_n1906_, new_n1907_, new_n1908_, new_n1909_,
    new_n1910_, new_n1911_, new_n1912_, new_n1913_, new_n1914_, new_n1915_,
    new_n1916_, new_n1917_, new_n1918_, new_n1919_, new_n1920_, new_n1921_,
    new_n1922_, new_n1923_, new_n1924_, new_n1925_, new_n1926_, new_n1927_,
    new_n1928_, new_n1929_, new_n1930_, new_n1931_, new_n1932_, new_n1933_,
    new_n1934_, new_n1935_, new_n1936_, new_n1937_, new_n1938_, new_n1939_,
    new_n1940_, new_n1941_, new_n1942_, new_n1943_, new_n1944_, new_n1945_,
    new_n1946_, new_n1947_, new_n1948_, new_n1949_, new_n1950_, new_n1951_,
    new_n1952_, new_n1953_, new_n1954_, new_n1955_, new_n1956_, new_n1957_,
    new_n1958_, new_n1959_, new_n1960_, new_n1961_, new_n1962_, new_n1963_,
    new_n1964_, new_n1965_, new_n1966_, new_n1967_, new_n1968_, new_n1969_,
    new_n1970_, new_n1971_, new_n1972_, new_n1973_, new_n1974_, new_n1975_,
    new_n1976_, new_n1977_, new_n1978_, new_n1979_, new_n1980_, new_n1981_,
    new_n1982_, new_n1983_, new_n1984_, new_n1985_, new_n1986_, new_n1987_,
    new_n1988_, new_n1989_, new_n1990_, new_n1991_, new_n1992_, new_n1993_,
    new_n1994_, new_n1995_, new_n1996_, new_n1997_, new_n1998_, new_n1999_,
    new_n2000_, new_n2001_, new_n2002_, new_n2003_, new_n2004_, new_n2005_,
    new_n2006_, new_n2007_, new_n2008_, new_n2009_, new_n2010_, new_n2011_,
    new_n2012_, new_n2013_, new_n2014_, new_n2015_, new_n2016_, new_n2017_,
    new_n2018_, new_n2019_, new_n2020_, new_n2021_, new_n2022_, new_n2023_,
    new_n2024_, new_n2025_, new_n2026_, new_n2027_, new_n2028_, new_n2029_,
    new_n2030_, new_n2031_, new_n2032_, new_n2033_, new_n2034_, new_n2035_,
    new_n2036_, new_n2037_, new_n2038_, new_n2039_, new_n2040_, new_n2041_,
    new_n2042_, new_n2043_, new_n2044_, new_n2045_, new_n2046_, new_n2047_,
    new_n2048_, new_n2049_, new_n2050_, new_n2051_, new_n2052_, new_n2053_,
    new_n2054_, new_n2055_, new_n2056_, new_n2057_, new_n2058_, new_n2059_,
    new_n2060_, new_n2061_, new_n2062_, new_n2063_, new_n2064_, new_n2065_,
    new_n2066_, new_n2067_, new_n2068_, new_n2069_, new_n2070_, new_n2071_,
    new_n2072_, new_n2073_, new_n2074_, new_n2075_, new_n2076_, new_n2077_,
    new_n2078_, new_n2079_, new_n2080_, new_n2081_, new_n2082_, new_n2083_,
    new_n2084_, new_n2085_, new_n2086_, new_n2087_, new_n2088_, new_n2089_,
    new_n2090_, new_n2091_, new_n2092_, new_n2093_, new_n2094_, new_n2095_,
    new_n2096_, new_n2097_, new_n2098_, new_n2099_, new_n2100_, new_n2101_,
    new_n2102_, new_n2103_, new_n2104_, new_n2105_, new_n2106_, new_n2107_,
    new_n2108_, new_n2109_, new_n2110_, new_n2111_, new_n2112_, new_n2113_,
    new_n2114_, new_n2115_, new_n2116_, new_n2117_, new_n2118_, new_n2119_,
    new_n2120_, new_n2121_, new_n2122_, new_n2123_, new_n2124_, new_n2125_,
    new_n2126_, new_n2127_, new_n2128_, new_n2129_, new_n2130_, new_n2131_,
    new_n2132_, new_n2133_, new_n2134_, new_n2135_, new_n2136_, new_n2137_,
    new_n2138_, new_n2139_, new_n2140_, new_n2141_, new_n2142_, new_n2143_,
    new_n2144_, new_n2145_, new_n2146_, new_n2147_, new_n2148_, new_n2149_,
    new_n2150_, new_n2151_, new_n2152_, new_n2153_, new_n2154_, new_n2155_,
    new_n2156_, new_n2157_, new_n2158_, new_n2159_, new_n2160_, new_n2161_,
    new_n2162_, new_n2163_, new_n2164_, new_n2165_, new_n2166_, new_n2167_,
    new_n2168_, new_n2169_, new_n2170_, new_n2171_, new_n2172_, new_n2173_,
    new_n2174_, new_n2175_, new_n2176_, new_n2177_, new_n2178_, new_n2179_,
    new_n2180_, new_n2181_, new_n2182_, new_n2183_, new_n2184_, new_n2185_,
    new_n2186_, new_n2187_, new_n2188_, new_n2189_, new_n2190_, new_n2191_,
    new_n2192_, new_n2193_, new_n2194_, new_n2195_, new_n2196_, new_n2197_,
    new_n2198_, new_n2199_, new_n2200_, new_n2201_, new_n2202_, new_n2203_,
    new_n2204_, new_n2205_, new_n2206_, new_n2207_, new_n2208_, new_n2209_,
    new_n2210_, new_n2211_, new_n2212_, new_n2213_, new_n2214_, new_n2215_,
    new_n2216_, new_n2217_, new_n2218_, new_n2219_, new_n2220_, new_n2221_,
    new_n2222_, new_n2223_, new_n2224_, new_n2225_, new_n2226_, new_n2227_,
    new_n2228_, new_n2229_, new_n2230_, new_n2231_, new_n2232_, new_n2233_,
    new_n2234_, new_n2235_, new_n2236_, new_n2237_, new_n2238_, new_n2239_,
    new_n2240_, new_n2241_, new_n2242_, new_n2243_, new_n2244_, new_n2245_,
    new_n2246_, new_n2247_, new_n2248_, new_n2249_, new_n2250_, new_n2251_,
    new_n2252_, new_n2253_, new_n2254_, new_n2255_, new_n2256_, new_n2257_,
    new_n2258_, new_n2259_, new_n2260_, new_n2261_, new_n2262_, new_n2263_,
    new_n2264_, new_n2265_, new_n2266_, new_n2267_, new_n2268_, new_n2269_,
    new_n2270_, new_n2271_, new_n2272_, new_n2273_, new_n2274_, new_n2275_,
    new_n2276_, new_n2277_, new_n2278_, new_n2279_, new_n2280_, new_n2281_,
    new_n2282_, new_n2283_, new_n2284_, new_n2285_, new_n2286_, new_n2287_,
    new_n2288_, new_n2289_, new_n2290_, new_n2291_, new_n2292_, new_n2293_,
    new_n2294_, new_n2295_, new_n2296_, new_n2297_, new_n2298_, new_n2299_,
    new_n2300_, new_n2301_, new_n2302_, new_n2303_, new_n2304_, new_n2305_,
    new_n2306_, new_n2307_, new_n2308_, new_n2309_, new_n2310_, new_n2311_,
    new_n2312_, new_n2313_, new_n2314_, new_n2315_, new_n2316_, new_n2317_,
    new_n2318_, new_n2319_, new_n2320_, new_n2321_, new_n2322_, new_n2323_,
    new_n2324_, new_n2325_, new_n2326_, new_n2327_, new_n2328_, new_n2329_,
    new_n2330_, new_n2331_, new_n2332_, new_n2333_, new_n2334_, new_n2335_,
    new_n2336_, new_n2337_, new_n2338_, new_n2339_, new_n2340_, new_n2341_,
    new_n2342_, new_n2343_, new_n2344_, new_n2345_, new_n2346_, new_n2347_,
    new_n2348_, new_n2349_, new_n2350_, new_n2351_, new_n2352_, new_n2353_,
    new_n2354_, new_n2355_, new_n2356_, new_n2357_, new_n2358_, new_n2359_,
    new_n2360_, new_n2361_, new_n2362_, new_n2363_, new_n2364_, new_n2365_,
    new_n2366_, new_n2367_, new_n2368_, new_n2369_, new_n2370_, new_n2371_,
    new_n2372_, new_n2373_, new_n2374_, new_n2375_, new_n2376_, new_n2377_,
    new_n2378_, new_n2379_, new_n2380_, new_n2381_, new_n2382_, new_n2383_,
    new_n2384_, new_n2385_, new_n2386_, new_n2387_, new_n2388_, new_n2389_,
    new_n2390_, new_n2391_, new_n2392_, new_n2393_, new_n2394_, new_n2395_,
    new_n2396_, new_n2397_, new_n2398_, new_n2399_, new_n2400_, new_n2401_,
    new_n2402_, new_n2403_, new_n2404_, new_n2405_, new_n2406_, new_n2407_,
    new_n2408_, new_n2409_, new_n2410_, new_n2411_, new_n2412_, new_n2413_,
    new_n2414_, new_n2415_, new_n2416_, new_n2417_, new_n2418_, new_n2419_,
    new_n2420_, new_n2421_, new_n2422_, new_n2423_, new_n2424_, new_n2425_,
    new_n2426_, new_n2427_, new_n2428_, new_n2429_, new_n2430_, new_n2431_,
    new_n2432_, new_n2433_, new_n2434_, new_n2435_, new_n2436_, new_n2437_,
    new_n2438_, new_n2439_, new_n2440_, new_n2441_, new_n2442_, new_n2443_,
    new_n2444_, new_n2445_, new_n2446_, new_n2447_, new_n2448_, new_n2449_,
    new_n2450_, new_n2451_, new_n2452_, new_n2453_, new_n2454_, new_n2455_,
    new_n2456_, new_n2457_, new_n2458_, new_n2459_, new_n2460_, new_n2461_,
    new_n2462_, new_n2463_, new_n2464_, new_n2465_, new_n2466_, new_n2467_,
    new_n2468_, new_n2469_, new_n2470_, new_n2471_, new_n2472_, new_n2473_,
    new_n2474_, new_n2475_, new_n2476_, new_n2477_, new_n2478_, new_n2479_,
    new_n2480_, new_n2481_, new_n2482_, new_n2483_, new_n2484_, new_n2485_,
    new_n2486_, new_n2487_, new_n2488_, new_n2489_, new_n2490_, new_n2491_,
    new_n2492_, new_n2493_, new_n2494_, new_n2495_, new_n2496_, new_n2497_,
    new_n2498_, new_n2499_, new_n2500_, new_n2501_, new_n2502_, new_n2503_,
    new_n2504_, new_n2505_, new_n2506_, new_n2507_, new_n2508_, new_n2509_,
    new_n2510_, new_n2511_, new_n2512_, new_n2513_, new_n2514_, new_n2515_,
    new_n2516_, new_n2517_, new_n2518_, new_n2519_, new_n2520_, new_n2521_,
    new_n2522_, new_n2523_, new_n2524_, new_n2525_, new_n2526_, new_n2527_,
    new_n2528_, new_n2529_, new_n2530_, new_n2531_, new_n2532_, new_n2533_,
    new_n2534_, new_n2535_, new_n2536_, new_n2537_, new_n2538_, new_n2539_,
    new_n2540_, new_n2541_, new_n2542_, new_n2543_, new_n2544_, new_n2545_,
    new_n2546_, new_n2547_, new_n2548_, new_n2549_, new_n2550_, new_n2551_,
    new_n2552_, new_n2553_, new_n2554_, new_n2555_, new_n2556_, new_n2557_,
    new_n2558_, new_n2559_, new_n2560_, new_n2561_, new_n2562_, new_n2563_,
    new_n2564_, new_n2565_, new_n2566_, new_n2567_, new_n2568_, new_n2569_,
    new_n2570_, new_n2571_, new_n2572_, new_n2573_, new_n2574_, new_n2575_,
    new_n2576_, new_n2577_, new_n2578_, new_n2579_, new_n2580_, new_n2581_,
    new_n2582_, new_n2583_, new_n2584_, new_n2585_, new_n2586_, new_n2587_,
    new_n2588_, new_n2589_, new_n2590_, new_n2591_, new_n2592_, new_n2593_,
    new_n2594_, new_n2595_, new_n2596_, new_n2597_, new_n2598_, new_n2599_,
    new_n2600_, new_n2601_, new_n2602_, new_n2603_, new_n2604_, new_n2605_,
    new_n2606_, new_n2607_, new_n2608_, new_n2609_, new_n2610_, new_n2611_,
    new_n2612_, new_n2613_, new_n2614_, new_n2615_, new_n2616_, new_n2617_,
    new_n2618_, new_n2619_, new_n2620_, new_n2621_, new_n2622_, new_n2623_,
    new_n2624_, new_n2625_, new_n2626_, new_n2627_, new_n2628_, new_n2629_,
    new_n2630_, new_n2631_, new_n2632_, new_n2633_, new_n2634_, new_n2635_,
    new_n2636_, new_n2637_, new_n2638_, new_n2639_, new_n2640_, new_n2641_,
    new_n2642_, new_n2643_, new_n2644_, new_n2645_, new_n2646_, new_n2647_,
    new_n2648_, new_n2649_, new_n2650_, new_n2651_, new_n2652_, new_n2653_,
    new_n2654_, new_n2655_, new_n2656_, new_n2657_, new_n2658_, new_n2659_,
    new_n2660_, new_n2661_, new_n2662_, new_n2663_, new_n2664_, new_n2665_,
    new_n2666_, new_n2667_, new_n2668_, new_n2669_, new_n2670_, new_n2671_,
    new_n2672_, new_n2673_, new_n2674_, new_n2675_, new_n2676_, new_n2677_,
    new_n2678_, new_n2679_, new_n2680_, new_n2681_, new_n2682_, new_n2683_,
    new_n2684_, new_n2685_, new_n2686_, new_n2687_, new_n2688_, new_n2689_,
    new_n2690_, new_n2691_, new_n2692_, new_n2693_, new_n2694_, new_n2695_,
    new_n2696_, new_n2697_, new_n2698_, new_n2699_, new_n2700_, new_n2701_,
    new_n2702_, new_n2703_, new_n2704_, new_n2705_, new_n2706_, new_n2707_,
    new_n2708_, new_n2709_, new_n2710_, new_n2711_, new_n2712_, new_n2713_,
    new_n2714_, new_n2715_, new_n2716_, new_n2717_, new_n2718_, new_n2719_,
    new_n2720_, new_n2721_, new_n2722_, new_n2723_, new_n2724_, new_n2725_,
    new_n2726_, new_n2727_, new_n2728_, new_n2729_, new_n2730_, new_n2731_,
    new_n2732_, new_n2733_, new_n2734_, new_n2735_, new_n2736_, new_n2737_,
    new_n2738_, new_n2739_, new_n2740_, new_n2741_, new_n2742_, new_n2743_,
    new_n2744_, new_n2745_, new_n2746_, new_n2747_, new_n2748_, new_n2749_,
    new_n2750_, new_n2751_, new_n2752_, new_n2753_, new_n2754_, new_n2755_,
    new_n2756_, new_n2757_, new_n2758_, new_n2759_, new_n2760_, new_n2761_,
    new_n2762_, new_n2763_, new_n2764_, new_n2765_, new_n2766_, new_n2767_,
    new_n2768_, new_n2769_, new_n2770_, new_n2771_, new_n2772_, new_n2773_,
    new_n2774_, new_n2775_, new_n2776_, new_n2777_, new_n2778_, new_n2779_,
    new_n2780_, new_n2781_, new_n2782_, new_n2783_, new_n2784_, new_n2785_,
    new_n2786_, new_n2787_, new_n2788_, new_n2789_, new_n2790_, new_n2791_,
    new_n2792_, new_n2793_, new_n2794_, new_n2795_, new_n2796_, new_n2797_,
    new_n2798_, new_n2799_, new_n2800_, new_n2801_, new_n2802_, new_n2803_,
    new_n2804_, new_n2805_, new_n2806_, new_n2807_, new_n2808_, new_n2809_,
    new_n2810_, new_n2811_, new_n2812_, new_n2813_, new_n2814_, new_n2815_,
    new_n2816_, new_n2817_, new_n2818_, new_n2819_, new_n2820_, new_n2821_,
    new_n2822_, new_n2823_, new_n2824_, new_n2825_, new_n2826_, new_n2827_,
    new_n2828_, new_n2829_, new_n2830_, new_n2831_, new_n2832_, new_n2833_,
    new_n2834_, new_n2835_, new_n2836_, new_n2837_, new_n2838_, new_n2839_,
    new_n2840_, new_n2841_, new_n2842_, new_n2843_, new_n2844_, new_n2845_,
    new_n2846_, new_n2847_, new_n2848_, new_n2849_, new_n2850_, new_n2851_,
    new_n2852_, new_n2853_, new_n2854_, new_n2855_, new_n2856_, new_n2857_,
    new_n2858_, new_n2859_, new_n2860_, new_n2861_, new_n2862_, new_n2863_,
    new_n2864_, new_n2865_, new_n2866_, new_n2867_, new_n2868_, new_n2869_,
    new_n2870_, new_n2871_, new_n2872_, new_n2873_, new_n2874_, new_n2875_,
    new_n2876_, new_n2877_, new_n2878_, new_n2879_, new_n2880_, new_n2881_,
    new_n2882_, new_n2883_, new_n2884_, new_n2885_, new_n2886_, new_n2887_,
    new_n2888_, new_n2889_, new_n2890_, new_n2891_, new_n2892_, new_n2893_,
    new_n2894_, new_n2895_, new_n2896_, new_n2897_, new_n2898_, new_n2899_,
    new_n2900_, new_n2901_, new_n2902_, new_n2903_, new_n2904_, new_n2905_,
    new_n2906_, new_n2907_, new_n2908_, new_n2909_, new_n2910_, new_n2911_,
    new_n2912_, new_n2913_, new_n2914_, new_n2915_, new_n2916_, new_n2917_,
    new_n2918_, new_n2919_, new_n2920_, new_n2921_, new_n2922_, new_n2923_,
    new_n2924_, new_n2925_, new_n2926_, new_n2927_, new_n2928_, new_n2929_,
    new_n2930_, new_n2931_, new_n2932_, new_n2933_, new_n2934_, new_n2935_,
    new_n2936_, new_n2937_, new_n2938_, new_n2939_, new_n2940_, new_n2941_,
    new_n2942_, new_n2943_, new_n2944_, new_n2945_, new_n2946_, new_n2947_,
    new_n2948_, new_n2949_, new_n2950_, new_n2951_, new_n2952_, new_n2953_,
    new_n2954_, new_n2955_, new_n2956_, new_n2957_, new_n2958_, new_n2959_,
    new_n2960_, new_n2961_, new_n2962_, new_n2963_, new_n2964_, new_n2965_,
    new_n2966_, new_n2967_, new_n2968_, new_n2969_, new_n2970_, new_n2971_,
    new_n2972_, new_n2973_, new_n2974_, new_n2975_, new_n2976_, new_n2977_,
    new_n2978_, new_n2979_, new_n2980_, new_n2981_, new_n2982_, new_n2983_,
    new_n2984_, new_n2985_, new_n2986_, new_n2987_, new_n2988_, new_n2989_,
    new_n2990_, new_n2991_, new_n2992_, new_n2993_, new_n2994_, new_n2995_,
    new_n2996_, new_n2997_, new_n2998_, new_n2999_, new_n3000_, new_n3001_,
    new_n3002_, new_n3003_, new_n3004_, new_n3005_, new_n3006_, new_n3007_,
    new_n3008_, new_n3009_, new_n3010_, new_n3011_, new_n3012_, new_n3013_,
    new_n3014_, new_n3015_, new_n3016_, new_n3017_, new_n3018_, new_n3019_,
    new_n3020_, new_n3021_, new_n3022_, new_n3023_, new_n3024_, new_n3025_,
    new_n3026_, new_n3027_, new_n3028_, new_n3029_, new_n3030_, new_n3031_,
    new_n3032_, new_n3033_, new_n3034_, new_n3035_, new_n3036_, new_n3037_,
    new_n3038_, new_n3039_, new_n3040_, new_n3041_, new_n3042_, new_n3043_,
    new_n3044_, new_n3045_, new_n3046_, new_n3047_, new_n3048_, new_n3049_,
    new_n3050_, new_n3051_, new_n3052_, new_n3053_, new_n3054_, new_n3055_,
    new_n3056_, new_n3057_, new_n3058_, new_n3059_, new_n3060_, new_n3061_,
    new_n3062_, new_n3063_, new_n3064_, new_n3065_, new_n3066_, new_n3067_,
    new_n3068_, new_n3069_, new_n3070_, new_n3071_, new_n3072_, new_n3073_,
    new_n3074_, new_n3075_, new_n3076_, new_n3077_, new_n3078_, new_n3079_,
    new_n3080_, new_n3081_, new_n3082_, new_n3083_, new_n3084_, new_n3085_,
    new_n3086_, new_n3087_, new_n3088_, new_n3089_, new_n3090_, new_n3091_,
    new_n3092_, new_n3093_, new_n3094_, new_n3095_, new_n3096_, new_n3097_,
    new_n3098_, new_n3099_, new_n3100_, new_n3101_, new_n3102_, new_n3103_,
    new_n3104_, new_n3105_, new_n3106_, new_n3107_, new_n3108_, new_n3109_,
    new_n3110_, new_n3111_, new_n3112_, new_n3113_, new_n3114_, new_n3115_,
    new_n3116_, new_n3117_, new_n3118_, new_n3119_, new_n3120_, new_n3121_,
    new_n3122_, new_n3123_, new_n3124_, new_n3125_, new_n3126_, new_n3127_,
    new_n3128_, new_n3129_, new_n3130_, new_n3131_, new_n3132_, new_n3133_,
    new_n3134_, new_n3135_, new_n3136_, new_n3137_, new_n3138_, new_n3139_,
    new_n3140_, new_n3141_, new_n3142_, new_n3143_, new_n3144_, new_n3145_,
    new_n3146_, new_n3147_, new_n3148_, new_n3149_, new_n3150_, new_n3151_,
    new_n3152_, new_n3153_, new_n3154_, new_n3155_, new_n3156_, new_n3157_,
    new_n3158_, new_n3159_, new_n3160_, new_n3161_, new_n3162_, new_n3163_,
    new_n3164_, new_n3165_, new_n3166_, new_n3167_, new_n3168_, new_n3169_,
    new_n3170_, new_n3171_, new_n3172_, new_n3173_, new_n3174_, new_n3175_,
    new_n3176_, new_n3177_, new_n3178_, new_n3179_, new_n3180_, new_n3181_,
    new_n3182_, new_n3183_, new_n3184_, new_n3185_, new_n3186_, new_n3187_,
    new_n3188_, new_n3189_, new_n3190_, new_n3191_, new_n3192_, new_n3193_,
    new_n3194_, new_n3195_, new_n3196_, new_n3197_, new_n3198_, new_n3199_,
    new_n3200_, new_n3201_, new_n3202_, new_n3203_, new_n3204_, new_n3205_,
    new_n3206_, new_n3207_, new_n3208_, new_n3209_, new_n3210_, new_n3211_,
    new_n3212_, new_n3213_, new_n3214_, new_n3215_, new_n3216_, new_n3217_,
    new_n3218_, new_n3219_, new_n3220_, new_n3221_, new_n3222_, new_n3223_,
    new_n3224_, new_n3225_, new_n3226_, new_n3227_, new_n3228_, new_n3229_,
    new_n3230_, new_n3231_, new_n3232_, new_n3233_, new_n3234_, new_n3235_,
    new_n3236_, new_n3237_, new_n3238_, new_n3239_, new_n3240_, new_n3241_,
    new_n3242_, new_n3243_, new_n3244_, new_n3245_, new_n3246_, new_n3247_,
    new_n3248_, new_n3249_, new_n3250_, new_n3251_, new_n3252_, new_n3253_,
    new_n3254_, new_n3255_, new_n3256_, new_n3257_, new_n3258_, new_n3259_,
    new_n3260_, new_n3261_, new_n3262_, new_n3263_, new_n3264_, new_n3265_,
    new_n3266_, new_n3267_, new_n3268_, new_n3269_, new_n3270_, new_n3271_,
    new_n3272_, new_n3273_, new_n3274_, new_n3275_, new_n3276_, new_n3277_,
    new_n3278_, new_n3279_, new_n3280_, new_n3281_, new_n3282_, new_n3283_,
    new_n3284_, new_n3285_, new_n3286_, new_n3287_, new_n3288_, new_n3289_,
    new_n3290_, new_n3291_, new_n3292_, new_n3293_, new_n3294_, new_n3295_,
    new_n3296_, new_n3297_, new_n3298_, new_n3299_, new_n3300_, new_n3301_,
    new_n3302_, new_n3303_, new_n3304_, new_n3305_, new_n3306_, new_n3307_,
    new_n3308_, new_n3309_, new_n3310_, new_n3311_, new_n3312_, new_n3313_,
    new_n3314_, new_n3315_, new_n3316_, new_n3317_, new_n3318_, new_n3319_,
    new_n3320_, new_n3321_, new_n3322_, new_n3323_, new_n3324_, new_n3325_,
    new_n3326_, new_n3327_, new_n3328_, new_n3329_, new_n3330_, new_n3331_,
    new_n3332_, new_n3333_, new_n3334_, new_n3335_, new_n3336_, new_n3337_,
    new_n3338_, new_n3339_, new_n3340_, new_n3341_, new_n3342_, new_n3343_,
    new_n3344_, new_n3345_, new_n3346_, new_n3347_, new_n3348_, new_n3349_,
    new_n3350_, new_n3351_, new_n3352_, new_n3353_, new_n3354_, new_n3355_,
    new_n3356_, new_n3357_, new_n3358_, new_n3359_, new_n3360_, new_n3361_,
    new_n3362_, new_n3363_, new_n3364_, new_n3365_, new_n3366_, new_n3367_,
    new_n3368_, new_n3369_, new_n3370_, new_n3371_, new_n3372_, new_n3373_,
    new_n3374_, new_n3375_, new_n3376_, new_n3377_, new_n3378_, new_n3379_,
    new_n3380_, new_n3381_, new_n3382_, new_n3383_, new_n3384_, new_n3385_,
    new_n3386_, new_n3387_, new_n3388_, new_n3389_, new_n3390_, new_n3391_,
    new_n3392_, new_n3393_, new_n3394_, new_n3395_, new_n3396_, new_n3397_,
    new_n3398_, new_n3399_, new_n3400_, new_n3401_, new_n3402_, new_n3403_,
    new_n3404_, new_n3405_, new_n3406_, new_n3407_, new_n3408_, new_n3409_,
    new_n3410_, new_n3411_, new_n3412_, new_n3413_, new_n3414_, new_n3415_,
    new_n3416_, new_n3417_, new_n3418_, new_n3419_, new_n3420_, new_n3421_,
    new_n3422_, new_n3423_, new_n3424_, new_n3425_, new_n3426_, new_n3427_,
    new_n3428_, new_n3429_, new_n3430_, new_n3431_, new_n3432_, new_n3433_,
    new_n3434_, new_n3435_, new_n3436_, new_n3437_, new_n3438_, new_n3439_,
    new_n3440_, new_n3441_, new_n3442_, new_n3443_, new_n3444_, new_n3445_,
    new_n3446_, new_n3447_, new_n3448_, new_n3449_, new_n3450_, new_n3451_,
    new_n3452_, new_n3453_, new_n3454_, new_n3455_, new_n3456_, new_n3457_,
    new_n3458_, new_n3459_, new_n3460_, new_n3461_, new_n3462_, new_n3463_,
    new_n3464_, new_n3465_, new_n3466_, new_n3467_, new_n3468_, new_n3469_,
    new_n3470_, new_n3471_, new_n3472_, new_n3473_, new_n3474_, new_n3475_,
    new_n3476_, new_n3477_, new_n3478_, new_n3479_, new_n3480_, new_n3481_,
    new_n3482_, new_n3483_, new_n3484_, new_n3485_, new_n3486_, new_n3487_,
    new_n3488_, new_n3489_, new_n3490_, new_n3491_, new_n3492_, new_n3493_,
    new_n3494_, new_n3495_, new_n3496_, new_n3497_, new_n3498_, new_n3499_,
    new_n3500_, new_n3501_, new_n3502_, new_n3503_, new_n3504_, new_n3505_,
    new_n3506_, new_n3507_, new_n3508_, new_n3509_, new_n3510_, new_n3511_,
    new_n3512_, new_n3513_, new_n3514_, new_n3515_, new_n3516_, new_n3517_,
    new_n3518_, new_n3519_, new_n3520_, new_n3521_, new_n3522_, new_n3523_,
    new_n3524_, new_n3525_, new_n3526_, new_n3527_, new_n3528_, new_n3529_,
    new_n3530_, new_n3531_, new_n3532_, new_n3533_, new_n3534_, new_n3535_,
    new_n3536_, new_n3537_, new_n3538_, new_n3539_, new_n3540_, new_n3541_,
    new_n3542_, new_n3543_, new_n3544_, new_n3545_, new_n3546_, new_n3547_,
    new_n3548_, new_n3549_, new_n3550_, new_n3551_, new_n3552_, new_n3553_,
    new_n3554_, new_n3555_, new_n3556_, new_n3557_, new_n3558_, new_n3559_,
    new_n3560_, new_n3561_, new_n3562_, new_n3563_, new_n3564_, new_n3565_,
    new_n3566_, new_n3567_, new_n3568_, new_n3569_, new_n3570_, new_n3571_,
    new_n3572_, new_n3573_, new_n3574_, new_n3575_, new_n3576_, new_n3577_,
    new_n3578_, new_n3579_, new_n3580_, new_n3581_, new_n3582_, new_n3583_,
    new_n3584_, new_n3585_, new_n3586_, new_n3587_, new_n3588_, new_n3589_,
    new_n3590_, new_n3591_, new_n3592_, new_n3593_, new_n3594_, new_n3595_,
    new_n3596_, new_n3597_, new_n3598_, new_n3599_, new_n3600_, new_n3601_,
    new_n3602_, new_n3603_, new_n3604_, new_n3605_, new_n3606_, new_n3607_,
    new_n3608_, new_n3609_, new_n3610_, new_n3611_, new_n3612_, new_n3613_,
    new_n3614_, new_n3615_, new_n3616_, new_n3617_, new_n3618_, new_n3619_,
    new_n3620_, new_n3621_, new_n3622_, new_n3623_, new_n3624_, new_n3625_,
    new_n3626_, new_n3627_, new_n3628_, new_n3629_, new_n3630_, new_n3631_,
    new_n3632_, new_n3633_, new_n3634_, new_n3635_, new_n3636_, new_n3637_,
    new_n3638_, new_n3639_, new_n3640_, new_n3641_, new_n3642_, new_n3643_,
    new_n3644_, new_n3645_, new_n3646_, new_n3647_, new_n3648_, new_n3649_,
    new_n3650_, new_n3651_, new_n3652_, new_n3653_, new_n3654_, new_n3655_,
    new_n3656_, new_n3657_, new_n3658_, new_n3659_, new_n3660_, new_n3661_,
    new_n3662_, new_n3663_, new_n3664_, new_n3665_, new_n3666_, new_n3667_,
    new_n3668_, new_n3669_, new_n3670_, new_n3671_, new_n3672_, new_n3673_,
    new_n3674_, new_n3675_, new_n3676_, new_n3677_, new_n3678_, new_n3679_,
    new_n3680_, new_n3681_, new_n3682_, new_n3683_, new_n3684_, new_n3685_,
    new_n3686_, new_n3687_, new_n3688_, new_n3689_, new_n3690_, new_n3691_,
    new_n3692_, new_n3693_, new_n3694_, new_n3695_, new_n3696_, new_n3697_,
    new_n3698_, new_n3699_, new_n3700_, new_n3701_, new_n3702_, new_n3703_,
    new_n3704_, new_n3705_, new_n3706_, new_n3707_, new_n3708_, new_n3709_,
    new_n3710_, new_n3711_, new_n3712_, new_n3713_, new_n3714_, new_n3715_,
    new_n3716_, new_n3717_, new_n3718_, new_n3719_, new_n3720_, new_n3721_,
    new_n3722_, new_n3723_, new_n3724_, new_n3725_, new_n3726_, new_n3727_,
    new_n3728_, new_n3729_, new_n3730_, new_n3731_, new_n3732_, new_n3733_,
    new_n3734_, new_n3735_, new_n3736_, new_n3737_, new_n3738_, new_n3739_,
    new_n3740_, new_n3741_, new_n3742_, new_n3743_, new_n3744_, new_n3745_,
    new_n3746_, new_n3747_, new_n3748_, new_n3749_, new_n3750_, new_n3751_,
    new_n3752_, new_n3753_, new_n3754_, new_n3755_, new_n3756_, new_n3757_,
    new_n3758_, new_n3759_, new_n3760_, new_n3761_, new_n3762_, new_n3763_,
    new_n3764_, new_n3765_, new_n3766_, new_n3767_, new_n3768_, new_n3769_,
    new_n3770_, new_n3771_, new_n3772_, new_n3773_, new_n3774_, new_n3775_,
    new_n3776_, new_n3777_, new_n3778_, new_n3779_, new_n3780_, new_n3781_,
    new_n3782_, new_n3783_, new_n3784_, new_n3785_, new_n3786_, new_n3787_,
    new_n3788_, new_n3789_, new_n3790_, new_n3791_, new_n3792_, new_n3793_,
    new_n3794_, new_n3795_, new_n3796_, new_n3797_, new_n3798_, new_n3799_,
    new_n3800_, new_n3801_, new_n3802_, new_n3803_, new_n3804_, new_n3805_,
    new_n3806_, new_n3807_, new_n3808_, new_n3809_, new_n3810_, new_n3811_,
    new_n3812_, new_n3813_, new_n3814_, new_n3815_, new_n3816_, new_n3817_,
    new_n3818_, new_n3819_, new_n3820_, new_n3821_, new_n3822_, new_n3823_,
    new_n3824_, new_n3825_, new_n3826_, new_n3827_, new_n3828_, new_n3829_,
    new_n3830_, new_n3831_, new_n3832_, new_n3833_, new_n3834_, new_n3835_,
    new_n3836_, new_n3837_, new_n3838_, new_n3839_, new_n3840_, new_n3841_,
    new_n3842_, new_n3843_, new_n3844_, new_n3845_, new_n3846_, new_n3847_,
    new_n3848_, new_n3849_, new_n3850_, new_n3851_, new_n3852_, new_n3853_,
    new_n3854_, new_n3855_, new_n3856_, new_n3857_, new_n3858_, new_n3859_,
    new_n3860_, new_n3861_, new_n3862_, new_n3863_, new_n3864_, new_n3865_,
    new_n3866_, new_n3867_, new_n3868_, new_n3869_, new_n3870_, new_n3871_,
    new_n3872_, new_n3873_, new_n3874_, new_n3875_, new_n3876_, new_n3877_,
    new_n3878_, new_n3879_, new_n3880_, new_n3881_, new_n3882_, new_n3883_,
    new_n3884_, new_n3885_, new_n3886_, new_n3887_, new_n3888_, new_n3889_,
    new_n3890_, new_n3891_, new_n3892_, new_n3893_, new_n3894_, new_n3895_,
    new_n3896_, new_n3897_, new_n3898_, new_n3899_, new_n3900_, new_n3901_,
    new_n3902_, new_n3903_, new_n3904_, new_n3905_, new_n3906_, new_n3907_,
    new_n3908_, new_n3909_, new_n3910_, new_n3911_, new_n3912_, new_n3913_,
    new_n3914_, new_n3915_, new_n3916_, new_n3917_, new_n3918_, new_n3919_,
    new_n3920_, new_n3921_, new_n3922_, new_n3923_, new_n3924_, new_n3925_,
    new_n3926_, new_n3927_, new_n3928_, new_n3929_, new_n3930_, new_n3931_,
    new_n3932_, new_n3933_, new_n3934_, new_n3935_, new_n3936_, new_n3937_,
    new_n3938_, new_n3939_, new_n3940_, new_n3941_, new_n3942_, new_n3943_,
    new_n3944_, new_n3945_, new_n3946_, new_n3947_, new_n3948_, new_n3949_,
    new_n3950_, new_n3951_, new_n3952_, new_n3953_, new_n3954_, new_n3955_,
    new_n3956_, new_n3957_, new_n3958_, new_n3959_, new_n3960_, new_n3961_,
    new_n3962_, new_n3963_, new_n3964_, new_n3965_, new_n3966_, new_n3967_,
    new_n3968_, new_n3969_, new_n3970_, new_n3971_, new_n3972_, new_n3973_,
    new_n3974_, new_n3975_, new_n3976_, new_n3977_, new_n3978_, new_n3979_,
    new_n3980_, new_n3981_, new_n3982_, new_n3983_, new_n3984_, new_n3985_,
    new_n3986_, new_n3987_, new_n3988_, new_n3989_, new_n3990_, new_n3991_,
    new_n3992_, new_n3993_, new_n3994_, new_n3995_, new_n3996_, new_n3997_,
    new_n3998_, new_n3999_, new_n4000_, new_n4001_, new_n4002_, new_n4003_,
    new_n4004_, new_n4005_, new_n4006_, new_n4007_, new_n4008_, new_n4009_,
    new_n4010_, new_n4011_, new_n4012_, new_n4013_, new_n4014_, new_n4015_,
    new_n4016_, new_n4017_, new_n4018_, new_n4019_, new_n4020_, new_n4021_,
    new_n4022_, new_n4023_, new_n4024_, new_n4025_, new_n4026_, new_n4027_,
    new_n4028_, new_n4029_, new_n4030_, new_n4031_, new_n4032_, new_n4033_,
    new_n4034_, new_n4035_, new_n4036_, new_n4037_, new_n4038_, new_n4039_,
    new_n4040_, new_n4041_, new_n4042_, new_n4043_, new_n4044_, new_n4045_,
    new_n4046_, new_n4047_, new_n4048_, new_n4049_, new_n4050_, new_n4051_,
    new_n4052_, new_n4053_, new_n4054_, new_n4055_, new_n4056_, new_n4057_,
    new_n4058_, new_n4059_, new_n4060_, new_n4061_, new_n4062_, new_n4063_,
    new_n4064_, new_n4065_, new_n4066_, new_n4067_, new_n4068_, new_n4069_,
    new_n4070_, new_n4071_, new_n4072_, new_n4073_, new_n4074_, new_n4075_,
    new_n4076_, new_n4077_, new_n4078_, new_n4079_, new_n4080_, new_n4081_,
    new_n4082_, new_n4083_, new_n4084_, new_n4085_, new_n4086_, new_n4087_,
    new_n4088_, new_n4089_, new_n4090_, new_n4091_, new_n4092_, new_n4093_,
    new_n4094_, new_n4095_, new_n4096_, new_n4097_, new_n4098_, new_n4099_,
    new_n4100_, new_n4101_, new_n4102_, new_n4103_, new_n4104_, new_n4105_,
    new_n4106_, new_n4107_, new_n4108_, new_n4109_, new_n4110_, new_n4111_,
    new_n4112_, new_n4113_, new_n4114_, new_n4115_, new_n4116_, new_n4117_,
    new_n4118_, new_n4119_, new_n4120_, new_n4121_, new_n4122_, new_n4123_,
    new_n4124_, new_n4125_, new_n4126_, new_n4127_, new_n4128_, new_n4129_,
    new_n4130_, new_n4131_, new_n4132_, new_n4133_, new_n4134_, new_n4135_,
    new_n4136_, new_n4137_, new_n4138_, new_n4139_, new_n4140_, new_n4141_,
    new_n4142_, new_n4143_, new_n4144_, new_n4145_, new_n4146_, new_n4147_,
    new_n4148_, new_n4149_, new_n4150_, new_n4151_, new_n4152_, new_n4153_,
    new_n4154_, new_n4155_, new_n4156_, new_n4157_, new_n4158_, new_n4159_,
    new_n4160_, new_n4161_, new_n4162_, new_n4163_, new_n4164_, new_n4165_,
    new_n4166_, new_n4167_, new_n4168_, new_n4169_, new_n4170_, new_n4171_,
    new_n4172_, new_n4173_, new_n4174_, new_n4175_, new_n4176_, new_n4177_,
    new_n4178_, new_n4179_, new_n4180_, new_n4181_, new_n4182_, new_n4183_,
    new_n4184_, new_n4185_, new_n4186_, new_n4187_, new_n4188_, new_n4189_,
    new_n4190_, new_n4191_, new_n4192_, new_n4193_, new_n4194_, new_n4195_,
    new_n4196_, new_n4197_, new_n4198_, new_n4199_, new_n4200_, new_n4201_,
    new_n4202_, new_n4203_, new_n4204_, new_n4205_, new_n4206_, new_n4207_,
    new_n4208_, new_n4209_, new_n4210_, new_n4211_, new_n4212_, new_n4213_,
    new_n4214_, new_n4215_, new_n4216_, new_n4217_, new_n4218_, new_n4219_,
    new_n4220_, new_n4221_, new_n4222_, new_n4223_, new_n4224_, new_n4225_,
    new_n4226_, new_n4227_, new_n4228_, new_n4229_, new_n4230_, new_n4231_,
    new_n4232_, new_n4233_, new_n4234_, new_n4235_, new_n4236_, new_n4237_,
    new_n4238_, new_n4239_, new_n4240_, new_n4241_, new_n4242_, new_n4243_,
    new_n4244_, new_n4245_, new_n4246_, new_n4247_, new_n4248_, new_n4249_,
    new_n4250_, new_n4251_, new_n4252_, new_n4253_, new_n4254_, new_n4255_,
    new_n4256_, new_n4257_, new_n4258_, new_n4259_, new_n4260_, new_n4261_,
    new_n4262_, new_n4263_, new_n4264_, new_n4265_, new_n4266_, new_n4267_,
    new_n4268_, new_n4269_, new_n4270_, new_n4271_, new_n4272_, new_n4273_,
    new_n4274_, new_n4275_, new_n4276_, new_n4277_, new_n4278_, new_n4279_,
    new_n4280_, new_n4281_, new_n4282_, new_n4283_, new_n4284_, new_n4285_,
    new_n4286_, new_n4287_, new_n4288_, new_n4289_, new_n4290_, new_n4291_,
    new_n4292_, new_n4293_, new_n4294_, new_n4295_, new_n4296_, new_n4297_,
    new_n4298_, new_n4299_, new_n4300_, new_n4301_, new_n4302_, new_n4303_,
    new_n4304_, new_n4305_, new_n4306_, new_n4307_, new_n4308_, new_n4309_,
    new_n4310_, new_n4311_, new_n4312_, new_n4313_, new_n4314_, new_n4315_,
    new_n4316_, new_n4317_, new_n4318_, new_n4319_, new_n4320_, new_n4321_,
    new_n4322_, new_n4323_, new_n4324_, new_n4325_, new_n4326_, new_n4327_,
    new_n4328_, new_n4329_, new_n4330_, new_n4331_, new_n4332_, new_n4333_,
    new_n4334_, new_n4335_, new_n4336_, new_n4337_, new_n4338_, new_n4339_,
    new_n4340_, new_n4341_, new_n4342_, new_n4343_, new_n4344_, new_n4345_,
    new_n4346_, new_n4347_, new_n4348_, new_n4349_, new_n4350_, new_n4351_,
    new_n4352_, new_n4353_, new_n4354_, new_n4355_, new_n4356_, new_n4357_,
    new_n4358_, new_n4359_, new_n4360_, new_n4361_, new_n4362_, new_n4363_,
    new_n4364_, new_n4365_, new_n4366_, new_n4367_, new_n4368_, new_n4369_,
    new_n4370_, new_n4371_, new_n4372_, new_n4373_, new_n4374_, new_n4375_,
    new_n4376_, new_n4377_, new_n4378_, new_n4379_, new_n4380_, new_n4381_,
    new_n4382_, new_n4383_, new_n4384_, new_n4385_, new_n4386_, new_n4387_,
    new_n4388_, new_n4389_, new_n4390_, new_n4391_, new_n4392_, new_n4393_,
    new_n4394_, new_n4395_, new_n4396_, new_n4397_, new_n4398_, new_n4399_,
    new_n4400_, new_n4401_, new_n4402_, new_n4403_, new_n4404_, new_n4405_,
    new_n4406_, new_n4407_, new_n4408_, new_n4409_, new_n4410_, new_n4411_,
    new_n4412_, new_n4413_, new_n4414_, new_n4415_, new_n4416_, new_n4417_,
    new_n4418_, new_n4419_, new_n4420_, new_n4421_, new_n4422_, new_n4423_,
    new_n4424_, new_n4425_, new_n4426_, new_n4427_, new_n4428_, new_n4429_,
    new_n4430_, new_n4431_, new_n4432_, new_n4433_, new_n4434_, new_n4435_,
    new_n4436_, new_n4437_, new_n4438_, new_n4439_, new_n4440_, new_n4441_,
    new_n4442_, new_n4443_, new_n4444_, new_n4445_, new_n4446_, new_n4447_,
    new_n4448_, new_n4449_, new_n4450_, new_n4451_, new_n4452_, new_n4453_,
    new_n4454_, new_n4455_, new_n4456_, new_n4457_, new_n4458_, new_n4459_,
    new_n4460_, new_n4461_, new_n4462_, new_n4463_, new_n4464_, new_n4465_,
    new_n4466_, new_n4467_, new_n4468_, new_n4469_, new_n4470_, new_n4471_,
    new_n4472_, new_n4473_, new_n4474_, new_n4475_, new_n4476_, new_n4477_,
    new_n4478_, new_n4479_, new_n4480_, new_n4481_, new_n4482_, new_n4483_,
    new_n4484_, new_n4485_, new_n4486_, new_n4487_, new_n4488_, new_n4489_,
    new_n4490_, new_n4491_, new_n4492_, new_n4493_, new_n4494_, new_n4495_,
    new_n4496_, new_n4497_, new_n4498_, new_n4499_, new_n4500_, new_n4501_,
    new_n4502_, new_n4503_, new_n4504_, new_n4505_, new_n4506_, new_n4507_,
    new_n4508_, new_n4509_, new_n4510_, new_n4511_, new_n4512_, new_n4513_,
    new_n4514_, new_n4515_, new_n4516_, new_n4517_, new_n4518_, new_n4519_,
    new_n4520_, new_n4521_, new_n4522_, new_n4523_, new_n4524_, new_n4525_,
    new_n4526_, new_n4527_, new_n4528_, new_n4529_, new_n4530_, new_n4531_,
    new_n4532_, new_n4533_, new_n4534_, new_n4535_, new_n4536_, new_n4537_,
    new_n4538_, new_n4539_, new_n4540_, new_n4541_, new_n4542_, new_n4543_,
    new_n4544_, new_n4545_, new_n4546_, new_n4547_, new_n4548_, new_n4549_,
    new_n4550_, new_n4551_, new_n4552_, new_n4553_, new_n4554_, new_n4555_,
    new_n4556_, new_n4557_, new_n4558_, new_n4559_, new_n4560_, new_n4561_,
    new_n4562_, new_n4563_, new_n4564_, new_n4565_, new_n4566_, new_n4567_,
    new_n4568_, new_n4569_, new_n4570_, new_n4571_, new_n4572_, new_n4573_,
    new_n4574_, new_n4575_, new_n4576_, new_n4577_, new_n4578_, new_n4579_,
    new_n4580_, new_n4581_, new_n4582_, new_n4583_, new_n4584_, new_n4585_,
    new_n4586_, new_n4587_, new_n4588_, new_n4589_, new_n4590_, new_n4591_,
    new_n4592_, new_n4593_, new_n4594_, new_n4595_, new_n4596_, new_n4597_,
    new_n4598_, new_n4599_, new_n4600_, new_n4601_, new_n4602_, new_n4603_,
    new_n4604_, new_n4605_, new_n4606_, new_n4607_, new_n4608_, new_n4609_,
    new_n4610_, new_n4611_, new_n4612_, new_n4613_, new_n4614_, new_n4615_,
    new_n4616_, new_n4617_, new_n4618_, new_n4619_, new_n4620_, new_n4621_,
    new_n4622_, new_n4623_, new_n4624_, new_n4625_, new_n4626_, new_n4627_,
    new_n4628_, new_n4629_, new_n4630_, new_n4631_, new_n4632_, new_n4633_,
    new_n4634_, new_n4635_, new_n4636_, new_n4637_, new_n4638_, new_n4639_,
    new_n4640_, new_n4641_, new_n4642_, new_n4643_, new_n4644_, new_n4645_,
    new_n4646_, new_n4647_, new_n4648_, new_n4649_, new_n4650_, new_n4651_,
    new_n4652_, new_n4653_, new_n4654_, new_n4655_, new_n4656_, new_n4657_,
    new_n4658_, new_n4659_, new_n4660_, new_n4661_, new_n4662_, new_n4663_,
    new_n4664_, new_n4665_, new_n4666_, new_n4667_, new_n4668_, new_n4669_,
    new_n4670_, new_n4671_, new_n4672_, new_n4673_, new_n4674_, new_n4675_,
    new_n4676_, new_n4677_, new_n4678_, new_n4679_, new_n4680_, new_n4681_,
    new_n4682_, new_n4683_, new_n4684_, new_n4685_, new_n4686_, new_n4687_,
    new_n4688_, new_n4689_, new_n4690_, new_n4691_, new_n4692_, new_n4693_,
    new_n4694_, new_n4695_, new_n4696_, new_n4697_, new_n4698_, new_n4699_,
    new_n4700_, new_n4701_, new_n4702_, new_n4703_, new_n4704_, new_n4705_,
    new_n4706_, new_n4707_, new_n4708_, new_n4709_, new_n4710_, new_n4711_,
    new_n4712_, new_n4713_, new_n4714_, new_n4715_, new_n4716_, new_n4717_,
    new_n4718_, new_n4719_, new_n4720_, new_n4721_, new_n4722_, new_n4723_,
    new_n4724_, new_n4725_, new_n4726_, new_n4727_, new_n4728_, new_n4729_,
    new_n4730_, new_n4731_, new_n4732_, new_n4733_, new_n4734_, new_n4735_,
    new_n4736_, new_n4737_, new_n4738_, new_n4739_, new_n4740_, new_n4741_,
    new_n4742_, new_n4743_, new_n4744_, new_n4745_, new_n4746_, new_n4747_,
    new_n4748_, new_n4749_, new_n4750_, new_n4751_, new_n4752_, new_n4753_,
    new_n4754_, new_n4755_, new_n4756_, new_n4757_, new_n4758_, new_n4759_,
    new_n4760_, new_n4761_, new_n4762_, new_n4763_, new_n4764_, new_n4765_,
    new_n4766_, new_n4767_, new_n4768_, new_n4769_, new_n4770_, new_n4771_,
    new_n4772_, new_n4773_, new_n4774_, new_n4775_, new_n4776_, new_n4777_,
    new_n4778_, new_n4779_, new_n4780_, new_n4781_, new_n4782_, new_n4783_,
    new_n4784_, new_n4785_, new_n4786_, new_n4787_, new_n4788_, new_n4789_,
    new_n4790_, new_n4791_, new_n4792_, new_n4793_, new_n4794_, new_n4795_,
    new_n4796_, new_n4797_, new_n4798_, new_n4799_, new_n4800_, new_n4801_,
    new_n4802_, new_n4803_, new_n4804_, new_n4805_, new_n4806_, new_n4807_,
    new_n4808_, new_n4809_, new_n4810_, new_n4811_, new_n4812_, new_n4813_,
    new_n4814_, new_n4815_, new_n4816_, new_n4817_, new_n4818_, new_n4819_,
    new_n4820_, new_n4821_, new_n4822_, new_n4823_, new_n4824_, new_n4825_,
    new_n4826_, new_n4827_, new_n4828_, new_n4829_, new_n4830_, new_n4831_,
    new_n4832_, new_n4833_, new_n4834_, new_n4835_, new_n4836_, new_n4837_,
    new_n4838_, new_n4839_, new_n4840_, new_n4841_, new_n4842_, new_n4843_,
    new_n4844_, new_n4845_, new_n4846_, new_n4847_, new_n4848_, new_n4849_,
    new_n4850_, new_n4851_, new_n4852_, new_n4853_, new_n4854_, new_n4855_,
    new_n4856_, new_n4857_, new_n4858_, new_n4859_, new_n4860_, new_n4861_,
    new_n4862_, new_n4863_, new_n4864_, new_n4865_, new_n4866_, new_n4867_,
    new_n4868_, new_n4869_, new_n4870_, new_n4871_, new_n4872_, new_n4873_,
    new_n4874_, new_n4875_, new_n4876_, new_n4877_, new_n4878_, new_n4879_,
    new_n4880_, new_n4881_, new_n4882_, new_n4883_, new_n4884_, new_n4885_,
    new_n4886_, new_n4887_, new_n4888_, new_n4889_, new_n4890_, new_n4891_,
    new_n4892_, new_n4893_, new_n4894_, new_n4895_, new_n4896_, new_n4897_,
    new_n4898_, new_n4899_, new_n4900_, new_n4901_, new_n4902_, new_n4903_,
    new_n4904_, new_n4905_, new_n4906_, new_n4907_, new_n4908_, new_n4909_,
    new_n4910_, new_n4911_, new_n4912_, new_n4913_, new_n4914_, new_n4915_,
    new_n4916_, new_n4917_, new_n4918_, new_n4919_, new_n4920_, new_n4921_,
    new_n4922_, new_n4923_, new_n4924_, new_n4925_, new_n4926_, new_n4927_,
    new_n4928_, new_n4929_, new_n4930_, new_n4931_, new_n4932_, new_n4933_,
    new_n4934_, new_n4935_, new_n4936_, new_n4937_, new_n4938_, new_n4939_,
    new_n4940_, new_n4941_, new_n4942_, new_n4943_, new_n4944_, new_n4945_,
    new_n4946_, new_n4947_, new_n4948_, new_n4949_, new_n4950_, new_n4951_,
    new_n4952_, new_n4953_, new_n4954_, new_n4955_, new_n4956_, new_n4957_,
    new_n4958_, new_n4959_, new_n4960_, new_n4961_, new_n4962_, new_n4963_,
    new_n4964_, new_n4965_, new_n4966_, new_n4967_, new_n4968_, new_n4969_,
    new_n4970_, new_n4971_, new_n4972_, new_n4973_, new_n4974_, new_n4975_,
    new_n4976_, new_n4977_, new_n4978_, new_n4979_, new_n4980_, new_n4981_,
    new_n4982_, new_n4983_, new_n4984_, new_n4985_, new_n4986_, new_n4987_,
    new_n4988_, new_n4989_, new_n4990_, new_n4991_, new_n4992_, new_n4993_,
    new_n4994_, new_n4995_, new_n4996_, new_n4997_, new_n4998_, new_n4999_,
    new_n5000_, new_n5001_, new_n5002_, new_n5003_, new_n5004_, new_n5005_,
    new_n5006_, new_n5007_, new_n5008_, new_n5009_, new_n5010_, new_n5011_,
    new_n5012_, new_n5013_, new_n5014_, new_n5015_, new_n5016_, new_n5017_,
    new_n5018_, new_n5019_, new_n5020_, new_n5021_, new_n5022_, new_n5023_,
    new_n5024_, new_n5025_, new_n5026_, new_n5027_, new_n5028_, new_n5029_,
    new_n5030_, new_n5031_, new_n5032_, new_n5033_, new_n5034_, new_n5035_,
    new_n5036_, new_n5037_, new_n5038_, new_n5039_, new_n5040_, new_n5041_,
    new_n5042_, new_n5043_, new_n5044_, new_n5045_, new_n5046_, new_n5047_,
    new_n5048_, new_n5049_, new_n5050_, new_n5051_, new_n5052_, new_n5053_,
    new_n5054_, new_n5055_, new_n5056_, new_n5057_, new_n5058_, new_n5059_,
    new_n5060_, new_n5061_, new_n5062_, new_n5063_, new_n5064_, new_n5065_,
    new_n5066_, new_n5067_, new_n5068_, new_n5069_, new_n5070_, new_n5071_,
    new_n5072_, new_n5073_, new_n5074_, new_n5075_, new_n5076_, new_n5077_,
    new_n5078_, new_n5079_, new_n5080_, new_n5081_, new_n5082_, new_n5083_,
    new_n5084_, new_n5085_, new_n5086_, new_n5087_, new_n5088_, new_n5089_,
    new_n5090_, new_n5091_, new_n5092_, new_n5093_, new_n5094_, new_n5095_,
    new_n5096_, new_n5097_, new_n5098_, new_n5099_, new_n5100_, new_n5101_,
    new_n5102_, new_n5103_, new_n5104_, new_n5105_, new_n5106_, new_n5107_,
    new_n5108_, new_n5109_, new_n5110_, new_n5111_, new_n5112_, new_n5113_,
    new_n5114_, new_n5115_, new_n5116_, new_n5117_, new_n5118_, new_n5119_,
    new_n5120_, new_n5121_, new_n5122_, new_n5123_, new_n5124_, new_n5125_,
    new_n5126_, new_n5127_, new_n5128_, new_n5129_, new_n5130_, new_n5131_,
    new_n5132_, new_n5133_, new_n5134_, new_n5135_, new_n5136_, new_n5137_,
    new_n5138_, new_n5139_, new_n5140_, new_n5141_, new_n5142_, new_n5143_,
    new_n5144_, new_n5145_, new_n5146_, new_n5147_, new_n5148_, new_n5149_,
    new_n5150_, new_n5151_, new_n5152_, new_n5153_, new_n5154_, new_n5155_,
    new_n5156_, new_n5157_, new_n5158_, new_n5159_, new_n5160_, new_n5161_,
    new_n5162_, new_n5163_, new_n5164_, new_n5165_, new_n5166_, new_n5167_,
    new_n5168_, new_n5169_, new_n5170_, new_n5171_, new_n5172_, new_n5173_,
    new_n5174_, new_n5175_, new_n5176_, new_n5177_, new_n5178_, new_n5179_,
    new_n5180_, new_n5181_, new_n5182_, new_n5183_, new_n5184_, new_n5185_,
    new_n5186_, new_n5187_, new_n5188_, new_n5189_, new_n5190_, new_n5191_,
    new_n5192_, new_n5193_, new_n5194_, new_n5195_, new_n5196_, new_n5197_,
    new_n5198_, new_n5199_, new_n5200_, new_n5201_, new_n5202_, new_n5203_,
    new_n5204_, new_n5205_, new_n5206_, new_n5207_, new_n5208_, new_n5209_,
    new_n5210_, new_n5211_, new_n5212_, new_n5213_, new_n5214_, new_n5215_,
    new_n5216_, new_n5217_, new_n5218_, new_n5219_, new_n5220_, new_n5221_,
    new_n5222_, new_n5223_, new_n5224_, new_n5225_, new_n5226_, new_n5227_,
    new_n5228_, new_n5229_, new_n5230_, new_n5231_, new_n5232_, new_n5233_,
    new_n5234_, new_n5235_, new_n5236_, new_n5237_, new_n5238_, new_n5239_,
    new_n5240_, new_n5241_, new_n5242_, new_n5243_, new_n5244_, new_n5245_,
    new_n5246_, new_n5247_, new_n5248_, new_n5249_, new_n5250_, new_n5251_,
    new_n5252_, new_n5253_, new_n5254_, new_n5255_, new_n5256_, new_n5257_,
    new_n5258_, new_n5259_, new_n5260_, new_n5261_, new_n5262_, new_n5263_,
    new_n5264_, new_n5265_, new_n5266_, new_n5267_, new_n5268_, new_n5269_,
    new_n5270_, new_n5271_, new_n5272_, new_n5273_, new_n5274_, new_n5275_,
    new_n5276_, new_n5277_, new_n5278_, new_n5279_, new_n5280_, new_n5281_,
    new_n5282_, new_n5283_, new_n5284_, new_n5285_, new_n5286_, new_n5287_,
    new_n5288_, new_n5289_, new_n5290_, new_n5291_, new_n5292_, new_n5293_,
    new_n5294_, new_n5295_, new_n5296_, new_n5297_, new_n5298_, new_n5299_,
    new_n5300_, new_n5301_, new_n5302_, new_n5303_, new_n5304_, new_n5305_,
    new_n5306_, new_n5307_, new_n5308_, new_n5309_, new_n5310_, new_n5311_,
    new_n5312_, new_n5313_, new_n5314_, new_n5315_, new_n5316_, new_n5317_,
    new_n5318_, new_n5319_, new_n5320_, new_n5321_, new_n5322_, new_n5323_,
    new_n5324_, new_n5325_, new_n5326_, new_n5327_, new_n5328_, new_n5329_,
    new_n5330_, new_n5331_, new_n5332_, new_n5333_, new_n5334_, new_n5335_,
    new_n5336_, new_n5337_, new_n5338_, new_n5339_, new_n5340_, new_n5341_,
    new_n5342_, new_n5343_, new_n5344_, new_n5345_, new_n5346_, new_n5347_,
    new_n5348_, new_n5349_, new_n5350_, new_n5351_, new_n5352_, new_n5353_,
    new_n5354_, new_n5355_, new_n5356_, new_n5357_, new_n5358_, new_n5359_,
    new_n5360_, new_n5361_, new_n5362_, new_n5363_, new_n5364_, new_n5365_,
    new_n5366_, new_n5367_, new_n5368_, new_n5369_, new_n5370_, new_n5371_,
    new_n5372_, new_n5373_, new_n5374_, new_n5375_, new_n5376_, new_n5377_,
    new_n5378_, new_n5379_, new_n5380_, new_n5381_, new_n5382_, new_n5383_,
    new_n5384_, new_n5385_, new_n5386_, new_n5387_, new_n5388_, new_n5389_,
    new_n5390_, new_n5391_, new_n5392_, new_n5393_, new_n5394_, new_n5395_,
    new_n5396_, new_n5397_, new_n5398_, new_n5399_, new_n5400_, new_n5401_,
    new_n5402_, new_n5403_, new_n5404_, new_n5405_, new_n5406_, new_n5407_,
    new_n5408_, new_n5409_, new_n5410_, new_n5411_, new_n5412_, new_n5413_,
    new_n5414_, new_n5415_, new_n5416_, new_n5417_, new_n5418_, new_n5419_,
    new_n5420_, new_n5421_, new_n5422_, new_n5423_, new_n5424_, new_n5425_,
    new_n5426_, new_n5427_, new_n5428_, new_n5429_, new_n5430_, new_n5431_,
    new_n5432_, new_n5433_, new_n5434_, new_n5435_, new_n5436_, new_n5437_,
    new_n5438_, new_n5439_, new_n5440_, new_n5441_, new_n5442_, new_n5443_,
    new_n5444_, new_n5445_, new_n5446_, new_n5447_, new_n5448_, new_n5449_,
    new_n5450_, new_n5451_, new_n5452_, new_n5453_, new_n5454_, new_n5455_,
    new_n5456_, new_n5457_, new_n5458_, new_n5459_, new_n5460_, new_n5461_,
    new_n5462_, new_n5463_, new_n5464_, new_n5465_, new_n5466_, new_n5467_,
    new_n5468_, new_n5469_, new_n5470_, new_n5471_, new_n5472_, new_n5473_,
    new_n5474_, new_n5475_, new_n5476_, new_n5477_, new_n5478_, new_n5479_,
    new_n5480_, new_n5481_, new_n5482_, new_n5483_, new_n5484_, new_n5485_,
    new_n5486_, new_n5487_, new_n5488_, new_n5489_, new_n5490_, new_n5491_,
    new_n5492_, new_n5493_, new_n5494_, new_n5495_, new_n5496_, new_n5497_,
    new_n5498_, new_n5499_, new_n5500_, new_n5501_, new_n5502_, new_n5503_,
    new_n5504_, new_n5505_, new_n5506_, new_n5507_, new_n5508_, new_n5509_,
    new_n5510_, new_n5511_, new_n5512_, new_n5513_, new_n5514_, new_n5515_,
    new_n5516_, new_n5517_, new_n5518_, new_n5519_, new_n5520_, new_n5521_,
    new_n5522_, new_n5523_, new_n5524_, new_n5525_, new_n5526_, new_n5527_,
    new_n5528_, new_n5529_, new_n5530_, new_n5531_, new_n5532_, new_n5533_,
    new_n5534_, new_n5535_, new_n5536_, new_n5537_, new_n5538_, new_n5539_,
    new_n5540_, new_n5541_, new_n5542_, new_n5543_, new_n5544_, new_n5545_,
    new_n5546_, new_n5547_, new_n5548_, new_n5549_, new_n5550_, new_n5551_,
    new_n5552_, new_n5553_, new_n5554_, new_n5555_, new_n5556_, new_n5557_,
    new_n5558_, new_n5559_, new_n5560_, new_n5561_, new_n5562_, new_n5563_,
    new_n5564_, new_n5565_, new_n5566_, new_n5567_, new_n5568_, new_n5569_,
    new_n5570_, new_n5571_, new_n5572_, new_n5573_, new_n5574_, new_n5575_,
    new_n5576_, new_n5577_, new_n5578_, new_n5579_, new_n5580_, new_n5581_,
    new_n5582_, new_n5583_, new_n5584_, new_n5585_, new_n5586_, new_n5587_,
    new_n5588_, new_n5589_, new_n5590_, new_n5591_, new_n5592_, new_n5593_,
    new_n5594_, new_n5595_, new_n5596_, new_n5597_, new_n5598_, new_n5599_,
    new_n5600_, new_n5601_, new_n5602_, new_n5603_, new_n5604_, new_n5605_,
    new_n5606_, new_n5607_, new_n5608_, new_n5609_, new_n5610_, new_n5611_,
    new_n5612_, new_n5613_, new_n5614_, new_n5615_, new_n5616_, new_n5617_,
    new_n5618_, new_n5619_, new_n5620_, new_n5621_, new_n5622_, new_n5623_,
    new_n5624_, new_n5625_, new_n5626_, new_n5627_, new_n5628_, new_n5629_,
    new_n5630_, new_n5631_, new_n5632_, new_n5633_, new_n5634_, new_n5635_,
    new_n5636_, new_n5637_, new_n5638_, new_n5639_, new_n5640_, new_n5641_,
    new_n5642_, new_n5643_, new_n5644_, new_n5645_, new_n5646_, new_n5647_,
    new_n5648_, new_n5649_, new_n5650_, new_n5651_, new_n5652_, new_n5653_,
    new_n5654_, new_n5655_, new_n5656_, new_n5657_, new_n5658_, new_n5659_,
    new_n5660_, new_n5661_, new_n5662_, new_n5663_, new_n5664_, new_n5665_,
    new_n5666_, new_n5667_, new_n5668_, new_n5669_, new_n5670_, new_n5671_,
    new_n5672_, new_n5673_, new_n5674_, new_n5675_, new_n5676_, new_n5677_,
    new_n5678_, new_n5679_, new_n5680_, new_n5681_, new_n5682_, new_n5683_,
    new_n5684_, new_n5685_, new_n5686_, new_n5687_, new_n5688_, new_n5689_,
    new_n5690_, new_n5691_, new_n5692_, new_n5693_, new_n5694_, new_n5695_,
    new_n5696_, new_n5697_, new_n5698_, new_n5699_, new_n5700_, new_n5701_,
    new_n5702_, new_n5703_, new_n5704_, new_n5705_, new_n5706_, new_n5707_,
    new_n5708_, new_n5709_, new_n5710_, new_n5711_, new_n5712_, new_n5713_,
    new_n5714_, new_n5715_, new_n5716_, new_n5717_, new_n5718_, new_n5719_,
    new_n5720_, new_n5721_, new_n5722_, new_n5723_, new_n5724_, new_n5725_,
    new_n5726_, new_n5727_, new_n5728_, new_n5729_, new_n5730_, new_n5731_,
    new_n5732_, new_n5733_, new_n5734_, new_n5735_, new_n5736_, new_n5737_,
    new_n5738_, new_n5739_, new_n5740_, new_n5741_, new_n5742_, new_n5743_,
    new_n5744_, new_n5745_, new_n5746_, new_n5747_, new_n5748_, new_n5749_,
    new_n5750_, new_n5751_, new_n5752_, new_n5753_, new_n5754_, new_n5755_,
    new_n5756_, new_n5757_, new_n5758_, new_n5759_, new_n5760_, new_n5761_,
    new_n5762_, new_n5763_, new_n5764_, new_n5765_, new_n5766_, new_n5767_,
    new_n5768_, new_n5769_, new_n5770_, new_n5771_, new_n5772_, new_n5773_,
    new_n5774_, new_n5775_, new_n5776_, new_n5777_, new_n5778_, new_n5779_,
    new_n5780_, new_n5781_, new_n5782_, new_n5783_, new_n5784_, new_n5785_,
    new_n5786_, new_n5787_, new_n5788_, new_n5789_, new_n5790_, new_n5791_,
    new_n5792_, new_n5793_, new_n5794_, new_n5795_, new_n5796_, new_n5797_,
    new_n5798_, new_n5799_, new_n5800_, new_n5801_, new_n5802_, new_n5803_,
    new_n5804_, new_n5805_, new_n5806_, new_n5807_, new_n5808_, new_n5809_,
    new_n5810_, new_n5811_, new_n5812_, new_n5813_, new_n5814_, new_n5815_,
    new_n5816_, new_n5817_, new_n5818_, new_n5819_, new_n5820_, new_n5821_,
    new_n5822_, new_n5823_, new_n5824_, new_n5825_, new_n5826_, new_n5827_,
    new_n5828_, new_n5829_, new_n5830_, new_n5831_, new_n5832_, new_n5833_,
    new_n5834_, new_n5835_, new_n5836_, new_n5837_, new_n5838_, new_n5839_,
    new_n5840_, new_n5841_, new_n5842_, new_n5843_, new_n5844_, new_n5845_,
    new_n5846_, new_n5847_, new_n5848_, new_n5849_, new_n5850_, new_n5851_,
    new_n5852_, new_n5853_, new_n5854_, new_n5855_, new_n5856_, new_n5857_,
    new_n5858_, new_n5859_, new_n5860_, new_n5861_, new_n5862_, new_n5863_,
    new_n5864_, new_n5865_, new_n5866_, new_n5867_, new_n5868_, new_n5869_,
    new_n5870_, new_n5871_, new_n5872_, new_n5873_, new_n5874_, new_n5875_,
    new_n5876_, new_n5877_, new_n5878_, new_n5879_, new_n5880_, new_n5881_,
    new_n5882_, new_n5883_, new_n5884_, new_n5885_, new_n5886_, new_n5887_,
    new_n5888_, new_n5889_, new_n5890_, new_n5891_, new_n5892_, new_n5893_,
    new_n5894_, new_n5895_, new_n5896_, new_n5897_, new_n5898_, new_n5899_,
    new_n5900_, new_n5901_, new_n5902_, new_n5903_, new_n5904_, new_n5905_,
    new_n5906_, new_n5907_, new_n5908_, new_n5909_, new_n5910_, new_n5911_,
    new_n5912_, new_n5913_, new_n5914_, new_n5915_, new_n5916_, new_n5917_,
    new_n5918_, new_n5919_, new_n5920_, new_n5921_, new_n5922_, new_n5923_,
    new_n5924_, new_n5925_, new_n5926_, new_n5927_, new_n5928_, new_n5929_,
    new_n5930_, new_n5931_, new_n5932_, new_n5933_, new_n5934_, new_n5935_,
    new_n5936_, new_n5937_, new_n5938_, new_n5939_, new_n5940_, new_n5941_,
    new_n5942_, new_n5943_, new_n5944_, new_n5945_, new_n5946_, new_n5947_,
    new_n5948_, new_n5949_, new_n5950_, new_n5951_, new_n5952_, new_n5953_,
    new_n5954_, new_n5955_, new_n5956_, new_n5957_, new_n5958_, new_n5959_,
    new_n5960_, new_n5961_, new_n5962_, new_n5963_, new_n5964_, new_n5965_,
    new_n5966_, new_n5967_, new_n5968_, new_n5969_, new_n5970_, new_n5971_,
    new_n5972_, new_n5973_, new_n5974_, new_n5975_, new_n5976_, new_n5977_,
    new_n5978_, new_n5979_, new_n5980_, new_n5981_, new_n5982_, new_n5983_,
    new_n5984_, new_n5985_, new_n5986_, new_n5987_, new_n5988_, new_n5989_,
    new_n5990_, new_n5991_, new_n5992_, new_n5993_, new_n5994_, new_n5995_,
    new_n5996_, new_n5997_, new_n5998_, new_n5999_, new_n6000_, new_n6001_,
    new_n6002_, new_n6003_, new_n6004_, new_n6005_, new_n6006_, new_n6007_,
    new_n6008_, new_n6009_, new_n6010_, new_n6011_, new_n6012_, new_n6013_,
    new_n6014_, new_n6015_, new_n6016_, new_n6017_, new_n6018_, new_n6019_,
    new_n6020_, new_n6021_, new_n6022_, new_n6023_, new_n6024_, new_n6025_,
    new_n6026_, new_n6027_, new_n6028_, new_n6029_, new_n6030_, new_n6031_,
    new_n6032_, new_n6033_, new_n6034_, new_n6035_, new_n6036_, new_n6037_,
    new_n6038_, new_n6039_, new_n6040_, new_n6041_, new_n6042_, new_n6043_,
    new_n6044_, new_n6045_, new_n6046_, new_n6047_, new_n6048_, new_n6049_,
    new_n6050_, new_n6051_, new_n6052_, new_n6053_, new_n6054_, new_n6055_,
    new_n6056_, new_n6057_, new_n6058_, new_n6059_, new_n6060_, new_n6061_,
    new_n6062_, new_n6063_, new_n6064_, new_n6065_, new_n6066_, new_n6067_,
    new_n6068_, new_n6069_, new_n6070_, new_n6071_, new_n6072_, new_n6073_,
    new_n6074_, new_n6075_, new_n6076_, new_n6077_, new_n6078_, new_n6079_,
    new_n6080_, new_n6081_, new_n6082_, new_n6083_, new_n6084_, new_n6085_,
    new_n6086_, new_n6087_, new_n6088_, new_n6089_, new_n6090_, new_n6091_,
    new_n6092_, new_n6093_, new_n6094_, new_n6095_, new_n6096_, new_n6097_,
    new_n6098_, new_n6099_, new_n6100_, new_n6101_, new_n6102_, new_n6103_,
    new_n6104_, new_n6105_, new_n6106_, new_n6107_, new_n6108_, new_n6109_,
    new_n6110_, new_n6111_, new_n6112_, new_n6113_, new_n6114_, new_n6115_,
    new_n6116_, new_n6117_, new_n6118_, new_n6119_, new_n6120_, new_n6121_,
    new_n6122_, new_n6123_, new_n6124_, new_n6125_, new_n6126_, new_n6127_,
    new_n6128_, new_n6129_, new_n6130_, new_n6131_, new_n6132_, new_n6133_,
    new_n6134_, new_n6135_, new_n6136_, new_n6137_, new_n6138_, new_n6139_,
    new_n6140_, new_n6141_, new_n6142_, new_n6143_, new_n6144_, new_n6145_,
    new_n6146_, new_n6147_, new_n6148_, new_n6149_, new_n6150_, new_n6151_,
    new_n6152_, new_n6153_, new_n6154_, new_n6155_, new_n6156_, new_n6157_,
    new_n6158_, new_n6159_, new_n6160_, new_n6161_, new_n6162_, new_n6163_,
    new_n6164_, new_n6165_, new_n6166_, new_n6167_, new_n6168_, new_n6169_,
    new_n6170_, new_n6171_, new_n6172_, new_n6173_, new_n6174_, new_n6175_,
    new_n6176_, new_n6177_, new_n6178_, new_n6179_, new_n6180_, new_n6181_,
    new_n6182_, new_n6183_, new_n6184_, new_n6185_, new_n6186_, new_n6187_,
    new_n6188_, new_n6189_, new_n6190_, new_n6191_, new_n6192_, new_n6193_,
    new_n6194_, new_n6195_, new_n6196_, new_n6197_, new_n6198_, new_n6199_,
    new_n6200_, new_n6201_, new_n6202_, new_n6203_, new_n6204_, new_n6205_,
    new_n6206_, new_n6207_, new_n6208_, new_n6209_, new_n6210_, new_n6211_,
    new_n6212_, new_n6213_, new_n6214_, new_n6215_, new_n6216_, new_n6217_,
    new_n6218_, new_n6219_, new_n6220_, new_n6221_, new_n6222_, new_n6223_,
    new_n6224_, new_n6225_, new_n6226_, new_n6227_, new_n6228_, new_n6229_,
    new_n6230_, new_n6231_, new_n6232_, new_n6233_, new_n6234_, new_n6235_,
    new_n6236_, new_n6237_, new_n6238_, new_n6239_, new_n6240_, new_n6241_,
    new_n6242_, new_n6243_, new_n6244_, new_n6245_, new_n6246_, new_n6247_,
    new_n6248_, new_n6249_, new_n6250_, new_n6251_, new_n6252_, new_n6253_,
    new_n6254_, new_n6255_, new_n6256_, new_n6257_, new_n6258_, new_n6259_,
    new_n6260_, new_n6261_, new_n6262_, new_n6263_, new_n6264_, new_n6265_,
    new_n6266_, new_n6267_, new_n6268_, new_n6269_, new_n6270_, new_n6271_,
    new_n6272_, new_n6273_, new_n6274_, new_n6275_, new_n6276_, new_n6277_,
    new_n6278_, new_n6279_, new_n6280_, new_n6281_, new_n6282_, new_n6283_,
    new_n6284_, new_n6285_, new_n6286_, new_n6287_, new_n6288_, new_n6289_,
    new_n6290_, new_n6291_, new_n6292_, new_n6293_, new_n6294_, new_n6295_,
    new_n6296_, new_n6297_, new_n6298_, new_n6299_, new_n6300_, new_n6301_,
    new_n6302_, new_n6303_, new_n6304_, new_n6305_, new_n6306_, new_n6307_,
    new_n6308_, new_n6309_, new_n6310_, new_n6311_, new_n6312_, new_n6313_,
    new_n6314_, new_n6315_, new_n6316_, new_n6317_, new_n6318_, new_n6319_,
    new_n6320_, new_n6321_, new_n6322_, new_n6323_, new_n6324_, new_n6325_,
    new_n6326_, new_n6327_, new_n6328_, new_n6329_, new_n6330_, new_n6331_,
    new_n6332_, new_n6333_, new_n6334_, new_n6335_, new_n6336_, new_n6337_,
    new_n6338_, new_n6339_, new_n6340_, new_n6341_, new_n6342_, new_n6343_,
    new_n6344_, new_n6345_, new_n6346_, new_n6347_, new_n6348_, new_n6349_,
    new_n6350_, new_n6351_, new_n6352_, new_n6353_, new_n6354_, new_n6355_,
    new_n6356_, new_n6357_, new_n6358_, new_n6359_, new_n6360_, new_n6361_,
    new_n6362_, new_n6363_, new_n6364_, new_n6365_, new_n6366_, new_n6367_,
    new_n6368_, new_n6369_, new_n6370_, new_n6371_, new_n6372_, new_n6373_,
    new_n6374_, new_n6375_, new_n6376_, new_n6377_, new_n6378_, new_n6379_,
    new_n6380_, new_n6381_, new_n6382_, new_n6383_, new_n6384_, new_n6385_,
    new_n6386_, new_n6387_, new_n6388_, new_n6389_, new_n6390_, new_n6391_,
    new_n6392_, new_n6393_, new_n6394_, new_n6395_, new_n6396_, new_n6397_,
    new_n6398_, new_n6399_, new_n6400_, new_n6401_, new_n6402_, new_n6403_,
    new_n6404_, new_n6405_, new_n6406_, new_n6407_, new_n6408_, new_n6409_,
    new_n6410_, new_n6411_, new_n6412_, new_n6413_, new_n6414_, new_n6415_,
    new_n6416_, new_n6417_, new_n6418_, new_n6419_, new_n6420_, new_n6421_,
    new_n6422_, new_n6423_, new_n6424_, new_n6425_, new_n6426_, new_n6427_,
    new_n6428_, new_n6429_, new_n6430_, new_n6431_, new_n6432_, new_n6433_,
    new_n6434_, new_n6435_, new_n6436_, new_n6437_, new_n6438_, new_n6439_,
    new_n6440_, new_n6441_, new_n6442_, new_n6443_, new_n6444_, new_n6445_,
    new_n6446_, new_n6447_, new_n6448_, new_n6449_, new_n6450_, new_n6451_,
    new_n6452_, new_n6453_, new_n6454_, new_n6455_, new_n6456_, new_n6457_,
    new_n6458_, new_n6459_, new_n6460_, new_n6461_, new_n6462_, new_n6463_,
    new_n6464_, new_n6465_, new_n6466_, new_n6467_, new_n6468_, new_n6469_,
    new_n6470_, new_n6471_, new_n6472_, new_n6473_, new_n6474_, new_n6475_,
    new_n6476_, new_n6477_, new_n6478_, new_n6479_, new_n6480_, new_n6481_,
    new_n6482_, new_n6483_, new_n6484_, new_n6485_, new_n6486_, new_n6487_,
    new_n6488_, new_n6489_, new_n6490_, new_n6491_, new_n6492_, new_n6493_,
    new_n6494_, new_n6495_, new_n6496_, new_n6497_, new_n6498_, new_n6499_,
    new_n6500_, new_n6501_, new_n6502_, new_n6503_, new_n6504_, new_n6505_,
    new_n6506_, new_n6507_, new_n6508_, new_n6509_, new_n6510_, new_n6511_,
    new_n6512_, new_n6513_, new_n6514_, new_n6515_, new_n6516_, new_n6517_,
    new_n6518_, new_n6519_, new_n6520_, new_n6521_, new_n6522_, new_n6523_,
    new_n6524_, new_n6525_, new_n6526_, new_n6527_, new_n6528_, new_n6529_,
    new_n6530_, new_n6531_, new_n6532_, new_n6533_, new_n6534_, new_n6535_,
    new_n6536_, new_n6537_, new_n6538_, new_n6539_, new_n6540_, new_n6541_,
    new_n6542_, new_n6543_, new_n6544_, new_n6545_, new_n6546_, new_n6547_,
    new_n6548_, new_n6549_, new_n6550_, new_n6551_, new_n6552_, new_n6553_,
    new_n6554_, new_n6555_, new_n6556_, new_n6557_, new_n6558_, new_n6559_,
    new_n6560_, new_n6561_, new_n6562_, new_n6563_, new_n6564_, new_n6565_,
    new_n6566_, new_n6567_, new_n6568_, new_n6569_, new_n6570_, new_n6571_,
    new_n6572_, new_n6573_, new_n6574_, new_n6575_, new_n6576_, new_n6577_,
    new_n6578_, new_n6579_, new_n6580_, new_n6581_, new_n6582_, new_n6583_,
    new_n6584_, new_n6585_, new_n6586_, new_n6587_, new_n6588_, new_n6589_,
    new_n6590_, new_n6591_, new_n6592_, new_n6593_, new_n6594_, new_n6595_,
    new_n6596_, new_n6597_, new_n6598_, new_n6599_, new_n6600_, new_n6601_,
    new_n6602_, new_n6603_, new_n6604_, new_n6605_, new_n6606_, new_n6607_,
    new_n6608_, new_n6609_, new_n6610_, new_n6611_, new_n6612_, new_n6613_,
    new_n6614_, new_n6615_, new_n6616_, new_n6617_, new_n6618_, new_n6619_,
    new_n6620_, new_n6621_, new_n6622_, new_n6623_, new_n6624_, new_n6625_,
    new_n6626_, new_n6627_, new_n6628_, new_n6629_, new_n6630_, new_n6631_,
    new_n6632_, new_n6633_, new_n6634_, new_n6635_, new_n6636_, new_n6637_,
    new_n6638_, new_n6639_, new_n6640_, new_n6641_, new_n6642_, new_n6643_,
    new_n6644_, new_n6645_, new_n6646_, new_n6647_, new_n6648_, new_n6649_,
    new_n6650_, new_n6651_, new_n6652_, new_n6653_, new_n6654_, new_n6655_,
    new_n6656_, new_n6657_, new_n6658_, new_n6659_, new_n6660_, new_n6661_,
    new_n6662_, new_n6663_, new_n6664_, new_n6665_, new_n6666_, new_n6667_,
    new_n6668_, new_n6669_, new_n6670_, new_n6671_, new_n6672_, new_n6673_,
    new_n6674_, new_n6675_, new_n6676_, new_n6677_, new_n6678_, new_n6679_,
    new_n6680_, new_n6681_, new_n6682_, new_n6683_, new_n6684_, new_n6685_,
    new_n6686_, new_n6687_, new_n6688_, new_n6689_, new_n6690_, new_n6691_,
    new_n6692_, new_n6693_, new_n6694_, new_n6695_, new_n6696_, new_n6697_,
    new_n6698_, new_n6699_, new_n6700_, new_n6701_, new_n6702_, new_n6703_,
    new_n6704_, new_n6705_, new_n6706_, new_n6707_, new_n6708_, new_n6709_,
    new_n6710_, new_n6711_, new_n6712_, new_n6713_, new_n6714_, new_n6715_,
    new_n6716_, new_n6717_, new_n6718_, new_n6719_, new_n6720_, new_n6721_,
    new_n6722_, new_n6723_, new_n6724_, new_n6725_, new_n6726_, new_n6727_,
    new_n6728_, new_n6729_, new_n6730_, new_n6731_, new_n6732_, new_n6733_,
    new_n6734_, new_n6735_, new_n6736_, new_n6737_, new_n6738_, new_n6739_,
    new_n6740_, new_n6741_, new_n6742_, new_n6743_, new_n6744_, new_n6745_,
    new_n6746_, new_n6747_, new_n6748_, new_n6749_, new_n6750_, new_n6751_,
    new_n6752_, new_n6753_, new_n6754_, new_n6755_, new_n6756_, new_n6757_,
    new_n6758_, new_n6759_, new_n6760_, new_n6761_, new_n6762_, new_n6763_,
    new_n6764_, new_n6765_, new_n6766_, new_n6767_, new_n6768_, new_n6769_,
    new_n6770_, new_n6771_, new_n6772_, new_n6773_, new_n6774_, new_n6775_,
    new_n6776_, new_n6777_, new_n6778_, new_n6779_, new_n6780_, new_n6781_,
    new_n6782_, new_n6783_, new_n6784_, new_n6785_, new_n6786_, new_n6787_,
    new_n6788_, new_n6789_, new_n6790_, new_n6791_, new_n6792_, new_n6793_,
    new_n6794_, new_n6795_, new_n6796_, new_n6797_, new_n6798_, new_n6799_,
    new_n6800_, new_n6801_, new_n6802_, new_n6803_, new_n6804_, new_n6805_,
    new_n6806_, new_n6807_, new_n6808_, new_n6809_, new_n6810_, new_n6811_,
    new_n6812_, new_n6813_, new_n6814_, new_n6815_, new_n6816_, new_n6817_,
    new_n6818_, new_n6819_, new_n6820_, new_n6821_, new_n6822_, new_n6823_,
    new_n6824_, new_n6825_, new_n6826_, new_n6827_, new_n6828_, new_n6829_,
    new_n6830_, new_n6831_, new_n6832_, new_n6833_, new_n6834_, new_n6835_,
    new_n6836_, new_n6837_, new_n6838_, new_n6839_, new_n6840_, new_n6841_,
    new_n6842_, new_n6843_, new_n6844_, new_n6845_, new_n6846_, new_n6847_,
    new_n6848_, new_n6849_, new_n6850_, new_n6851_, new_n6852_, new_n6853_,
    new_n6854_, new_n6855_, new_n6856_, new_n6857_, new_n6858_, new_n6859_,
    new_n6860_, new_n6861_, new_n6862_, new_n6863_, new_n6864_, new_n6865_,
    new_n6866_, new_n6867_, new_n6868_, new_n6869_, new_n6870_, new_n6871_,
    new_n6872_, new_n6873_, new_n6874_, new_n6875_, new_n6876_, new_n6877_,
    new_n6878_, new_n6879_, new_n6880_, new_n6881_, new_n6882_, new_n6883_,
    new_n6884_, new_n6885_, new_n6886_, new_n6887_, new_n6888_, new_n6889_,
    new_n6890_, new_n6891_, new_n6892_, new_n6893_, new_n6894_, new_n6895_,
    new_n6896_, new_n6897_, new_n6898_, new_n6899_, new_n6900_, new_n6901_,
    new_n6902_, new_n6903_, new_n6904_, new_n6905_, new_n6906_, new_n6907_,
    new_n6908_, new_n6909_, new_n6910_, new_n6911_, new_n6912_, new_n6913_,
    new_n6914_, new_n6915_, new_n6916_, new_n6917_, new_n6918_, new_n6919_,
    new_n6920_, new_n6921_, new_n6922_, new_n6923_, new_n6924_, new_n6925_,
    new_n6926_, new_n6927_, new_n6928_, new_n6929_, new_n6930_, new_n6931_,
    new_n6932_, new_n6933_, new_n6934_, new_n6935_, new_n6936_, new_n6937_,
    new_n6938_, new_n6939_, new_n6940_, new_n6941_, new_n6942_, new_n6943_,
    new_n6944_, new_n6945_, new_n6946_, new_n6947_, new_n6948_, new_n6949_,
    new_n6950_, new_n6951_, new_n6952_, new_n6953_, new_n6954_, new_n6955_,
    new_n6956_, new_n6957_, new_n6958_, new_n6959_, new_n6960_, new_n6961_,
    new_n6962_, new_n6963_, new_n6964_, new_n6965_, new_n6966_, new_n6967_,
    new_n6968_, new_n6969_, new_n6970_, new_n6971_, new_n6972_, new_n6973_,
    new_n6974_, new_n6975_, new_n6976_, new_n6977_, new_n6978_, new_n6979_,
    new_n6980_, new_n6981_, new_n6982_, new_n6983_, new_n6984_, new_n6985_,
    new_n6986_, new_n6987_, new_n6988_, new_n6989_, new_n6990_, new_n6991_,
    new_n6992_, new_n6993_, new_n6994_, new_n6995_, new_n6996_, new_n6997_,
    new_n6998_, new_n6999_, new_n7000_, new_n7001_, new_n7002_, new_n7003_,
    new_n7004_, new_n7005_, new_n7006_, new_n7007_, new_n7008_, new_n7009_,
    new_n7010_, new_n7011_, new_n7012_, new_n7013_, new_n7014_, new_n7015_,
    new_n7016_, new_n7017_, new_n7018_, new_n7019_, new_n7020_, new_n7021_,
    new_n7022_, new_n7023_, new_n7024_, new_n7025_, new_n7026_, new_n7027_,
    new_n7028_, new_n7029_, new_n7030_, new_n7031_, new_n7032_, new_n7033_,
    new_n7034_, new_n7035_, new_n7036_, new_n7037_, new_n7038_, new_n7039_,
    new_n7040_, new_n7041_, new_n7042_, new_n7043_, new_n7044_, new_n7045_,
    new_n7046_, new_n7047_, new_n7048_, new_n7049_, new_n7050_, new_n7051_,
    new_n7052_, new_n7053_, new_n7054_, new_n7055_, new_n7056_, new_n7057_,
    new_n7058_, new_n7059_, new_n7060_, new_n7061_, new_n7062_, new_n7063_,
    new_n7064_, new_n7065_, new_n7066_, new_n7067_, new_n7068_, new_n7069_,
    new_n7070_, new_n7071_, new_n7072_, new_n7073_, new_n7074_, new_n7075_,
    new_n7076_, new_n7077_, new_n7078_, new_n7079_, new_n7080_, new_n7081_,
    new_n7082_, new_n7083_, new_n7084_, new_n7085_, new_n7086_, new_n7087_,
    new_n7088_, new_n7089_, new_n7090_, new_n7091_, new_n7092_, new_n7093_,
    new_n7094_, new_n7095_, new_n7096_, new_n7097_, new_n7098_, new_n7099_,
    new_n7100_, new_n7101_, new_n7102_, new_n7103_, new_n7104_, new_n7105_,
    new_n7106_, new_n7107_, new_n7108_, new_n7109_, new_n7110_, new_n7111_,
    new_n7112_, new_n7113_, new_n7114_, new_n7115_, new_n7116_, new_n7117_,
    new_n7118_, new_n7119_, new_n7120_, new_n7121_, new_n7122_, new_n7123_,
    new_n7124_, new_n7125_, new_n7126_, new_n7127_, new_n7128_, new_n7129_,
    new_n7130_, new_n7131_, new_n7132_, new_n7133_, new_n7134_, new_n7135_,
    new_n7136_, new_n7137_, new_n7138_, new_n7139_, new_n7140_, new_n7141_,
    new_n7142_, new_n7143_, new_n7144_, new_n7145_, new_n7146_, new_n7147_,
    new_n7148_, new_n7149_, new_n7150_, new_n7151_, new_n7152_, new_n7153_,
    new_n7154_, new_n7155_, new_n7156_, new_n7157_, new_n7158_, new_n7159_,
    new_n7160_, new_n7161_, new_n7162_, new_n7163_, new_n7164_, new_n7165_,
    new_n7166_, new_n7167_, new_n7168_, new_n7169_, new_n7170_, new_n7171_,
    new_n7172_, new_n7173_, new_n7174_, new_n7175_, new_n7176_, new_n7177_,
    new_n7178_, new_n7179_, new_n7180_, new_n7181_, new_n7182_, new_n7183_,
    new_n7184_, new_n7185_, new_n7186_, new_n7187_, new_n7188_, new_n7189_,
    new_n7190_, new_n7191_, new_n7192_, new_n7193_, new_n7194_, new_n7195_,
    new_n7196_, new_n7197_, new_n7198_, new_n7199_, new_n7200_, new_n7201_,
    new_n7202_, new_n7203_, new_n7204_, new_n7205_, new_n7206_, new_n7207_,
    new_n7208_, new_n7209_, new_n7210_, new_n7211_, new_n7212_, new_n7213_,
    new_n7214_, new_n7215_, new_n7216_, new_n7217_, new_n7218_, new_n7219_,
    new_n7220_, new_n7221_, new_n7222_, new_n7223_, new_n7224_, new_n7225_,
    new_n7226_, new_n7227_, new_n7228_, new_n7229_, new_n7230_, new_n7231_,
    new_n7232_, new_n7233_, new_n7234_, new_n7235_, new_n7236_, new_n7237_,
    new_n7238_, new_n7239_, new_n7240_, new_n7241_, new_n7242_, new_n7243_,
    new_n7244_, new_n7245_, new_n7246_, new_n7247_, new_n7248_, new_n7249_,
    new_n7250_, new_n7251_, new_n7252_, new_n7253_, new_n7254_, new_n7255_,
    new_n7256_, new_n7257_, new_n7258_, new_n7259_, new_n7260_, new_n7261_,
    new_n7262_, new_n7263_, new_n7264_, new_n7265_, new_n7266_, new_n7267_,
    new_n7268_, new_n7269_, new_n7270_, new_n7271_, new_n7272_, new_n7273_,
    new_n7274_, new_n7275_, new_n7276_, new_n7277_, new_n7278_, new_n7279_,
    new_n7280_, new_n7281_, new_n7282_, new_n7283_, new_n7284_, new_n7285_,
    new_n7286_, new_n7287_, new_n7288_, new_n7289_, new_n7290_, new_n7291_,
    new_n7292_, new_n7293_, new_n7294_, new_n7295_, new_n7296_, new_n7297_,
    new_n7298_, new_n7299_, new_n7300_, new_n7301_, new_n7302_, new_n7303_,
    new_n7304_, new_n7305_, new_n7306_, new_n7307_, new_n7308_, new_n7309_,
    new_n7310_, new_n7311_, new_n7312_, new_n7313_, new_n7314_, new_n7315_,
    new_n7316_, new_n7317_, new_n7318_, new_n7319_, new_n7320_, new_n7321_,
    new_n7322_, new_n7323_, new_n7324_, new_n7325_, new_n7326_, new_n7327_,
    new_n7328_, new_n7329_, new_n7330_, new_n7331_, new_n7332_, new_n7333_,
    new_n7334_, new_n7335_, new_n7336_, new_n7337_, new_n7338_, new_n7339_,
    new_n7340_, new_n7341_, new_n7342_, new_n7343_, new_n7344_, new_n7345_,
    new_n7346_, new_n7347_, new_n7348_, new_n7349_, new_n7350_, new_n7351_,
    new_n7352_, new_n7353_, new_n7354_, new_n7355_, new_n7356_, new_n7357_,
    new_n7358_, new_n7359_, new_n7360_, new_n7361_, new_n7362_, new_n7363_,
    new_n7364_, new_n7365_, new_n7366_, new_n7367_, new_n7368_, new_n7369_,
    new_n7370_, new_n7371_, new_n7372_, new_n7373_, new_n7374_, new_n7375_,
    new_n7376_, new_n7377_, new_n7378_, new_n7379_, new_n7380_, new_n7381_,
    new_n7382_, new_n7383_, new_n7384_, new_n7385_, new_n7386_, new_n7387_,
    new_n7388_, new_n7389_, new_n7390_, new_n7391_, new_n7392_, new_n7393_,
    new_n7394_, new_n7395_, new_n7396_, new_n7397_, new_n7398_, new_n7399_,
    new_n7400_, new_n7401_, new_n7402_, new_n7403_, new_n7404_, new_n7405_,
    new_n7406_, new_n7407_, new_n7408_, new_n7409_, new_n7410_, new_n7411_,
    new_n7412_, new_n7413_, new_n7414_, new_n7415_, new_n7416_, new_n7417_,
    new_n7418_, new_n7419_, new_n7420_, new_n7421_, new_n7422_, new_n7423_,
    new_n7424_, new_n7425_, new_n7426_, new_n7427_, new_n7428_, new_n7429_,
    new_n7430_, new_n7431_, new_n7432_, new_n7433_, new_n7434_, new_n7435_,
    new_n7436_, new_n7437_, new_n7438_, new_n7439_, new_n7440_, new_n7441_,
    new_n7442_, new_n7443_, new_n7444_, new_n7445_, new_n7446_, new_n7447_,
    new_n7448_, new_n7449_, new_n7450_, new_n7451_, new_n7452_, new_n7453_,
    new_n7454_, new_n7455_, new_n7456_, new_n7457_, new_n7458_, new_n7459_,
    new_n7460_, new_n7461_, new_n7462_, new_n7463_, new_n7464_, new_n7465_,
    new_n7466_, new_n7467_, new_n7468_, new_n7469_, new_n7470_, new_n7471_,
    new_n7472_, new_n7473_, new_n7474_, new_n7475_, new_n7476_, new_n7477_,
    new_n7478_, new_n7479_, new_n7480_, new_n7481_, new_n7482_, new_n7483_,
    new_n7484_, new_n7485_, new_n7486_, new_n7487_, new_n7488_, new_n7489_,
    new_n7490_, new_n7491_, new_n7492_, new_n7493_, new_n7494_, new_n7495_,
    new_n7496_, new_n7497_, new_n7498_, new_n7499_, new_n7500_, new_n7501_,
    new_n7502_, new_n7503_, new_n7504_, new_n7505_, new_n7506_, new_n7507_,
    new_n7508_, new_n7509_, new_n7510_, new_n7511_, new_n7512_, new_n7513_,
    new_n7514_, new_n7515_, new_n7516_, new_n7517_, new_n7518_, new_n7519_,
    new_n7520_, new_n7521_, new_n7522_, new_n7523_, new_n7524_, new_n7525_,
    new_n7526_, new_n7527_, new_n7528_, new_n7529_, new_n7530_, new_n7531_,
    new_n7532_, new_n7533_, new_n7534_, new_n7535_, new_n7536_, new_n7537_,
    new_n7538_, new_n7539_, new_n7540_, new_n7541_, new_n7542_, new_n7543_,
    new_n7544_, new_n7545_, new_n7546_, new_n7547_, new_n7548_, new_n7549_,
    new_n7550_, new_n7551_, new_n7552_, new_n7553_, new_n7554_, new_n7555_,
    new_n7556_, new_n7557_, new_n7558_, new_n7559_, new_n7560_, new_n7561_,
    new_n7562_, new_n7563_, new_n7564_, new_n7565_, new_n7566_, new_n7567_,
    new_n7568_, new_n7569_, new_n7570_, new_n7571_, new_n7572_, new_n7573_,
    new_n7574_, new_n7575_, new_n7576_, new_n7577_, new_n7578_, new_n7579_,
    new_n7580_, new_n7581_, new_n7582_, new_n7583_, new_n7584_, new_n7585_,
    new_n7586_, new_n7587_, new_n7588_, new_n7589_, new_n7590_, new_n7591_,
    new_n7592_, new_n7593_, new_n7594_, new_n7595_, new_n7596_, new_n7597_,
    new_n7598_, new_n7599_, new_n7600_, new_n7601_, new_n7602_, new_n7603_,
    new_n7604_, new_n7605_, new_n7606_, new_n7607_, new_n7608_, new_n7609_,
    new_n7610_, new_n7611_, new_n7612_, new_n7613_, new_n7614_, new_n7615_,
    new_n7616_, new_n7617_, new_n7618_, new_n7619_, new_n7620_, new_n7621_,
    new_n7622_, new_n7623_, new_n7624_, new_n7625_, new_n7626_, new_n7627_,
    new_n7628_, new_n7629_, new_n7630_, new_n7631_, new_n7632_, new_n7633_,
    new_n7634_, new_n7635_, new_n7636_, new_n7637_, new_n7638_, new_n7639_,
    new_n7640_, new_n7641_, new_n7642_, new_n7643_, new_n7644_, new_n7645_,
    new_n7646_, new_n7647_, new_n7648_, new_n7649_, new_n7650_, new_n7651_,
    new_n7652_, new_n7653_, new_n7654_, new_n7655_, new_n7656_, new_n7657_,
    new_n7658_, new_n7659_, new_n7660_, new_n7661_, new_n7662_, new_n7663_,
    new_n7664_, new_n7665_, new_n7666_, new_n7667_, new_n7668_, new_n7669_,
    new_n7670_, new_n7671_, new_n7672_, new_n7673_, new_n7674_, new_n7675_,
    new_n7676_, new_n7677_, new_n7678_, new_n7679_, new_n7680_, new_n7681_,
    new_n7682_, new_n7683_, new_n7684_, new_n7685_, new_n7686_, new_n7687_,
    new_n7688_, new_n7689_, new_n7690_, new_n7691_, new_n7692_, new_n7693_,
    new_n7694_, new_n7695_, new_n7696_, new_n7697_, new_n7698_, new_n7699_,
    new_n7700_, new_n7701_, new_n7702_, new_n7703_, new_n7704_, new_n7705_,
    new_n7706_, new_n7707_, new_n7708_, new_n7709_, new_n7710_, new_n7711_,
    new_n7712_, new_n7713_, new_n7714_, new_n7715_, new_n7716_, new_n7717_,
    new_n7718_, new_n7719_, new_n7720_, new_n7721_, new_n7722_, new_n7723_,
    new_n7724_, new_n7725_, new_n7726_, new_n7727_, new_n7728_, new_n7729_,
    new_n7730_, new_n7731_, new_n7732_, new_n7733_, new_n7734_, new_n7735_,
    new_n7736_, new_n7737_, new_n7738_, new_n7739_, new_n7740_, new_n7741_,
    new_n7742_, new_n7743_, new_n7744_, new_n7745_, new_n7746_, new_n7747_,
    new_n7748_, new_n7749_, new_n7750_, new_n7751_, new_n7752_, new_n7753_,
    new_n7754_, new_n7755_, new_n7756_, new_n7757_, new_n7758_, new_n7759_,
    new_n7760_, new_n7761_, new_n7762_, new_n7763_, new_n7764_, new_n7765_,
    new_n7766_, new_n7767_, new_n7768_, new_n7769_, new_n7770_, new_n7771_,
    new_n7772_, new_n7773_, new_n7774_, new_n7775_, new_n7776_, new_n7777_,
    new_n7778_, new_n7779_, new_n7780_, new_n7781_, new_n7782_, new_n7783_,
    new_n7784_, new_n7785_, new_n7786_, new_n7787_, new_n7788_, new_n7789_,
    new_n7790_, new_n7791_, new_n7792_, new_n7793_, new_n7794_, new_n7795_,
    new_n7796_, new_n7797_, new_n7798_, new_n7799_, new_n7800_, new_n7801_,
    new_n7802_, new_n7803_, new_n7804_, new_n7805_, new_n7806_, new_n7807_,
    new_n7808_, new_n7809_, new_n7810_, new_n7811_, new_n7812_, new_n7813_,
    new_n7814_, new_n7815_, new_n7816_, new_n7817_, new_n7818_, new_n7819_,
    new_n7820_, new_n7821_, new_n7822_, new_n7823_, new_n7824_, new_n7825_,
    new_n7826_, new_n7827_, new_n7828_, new_n7829_, new_n7830_, new_n7831_,
    new_n7832_, new_n7833_, new_n7834_, new_n7835_, new_n7836_, new_n7837_,
    new_n7838_, new_n7839_, new_n7840_, new_n7841_, new_n7842_, new_n7843_,
    new_n7844_, new_n7845_, new_n7846_, new_n7847_, new_n7848_, new_n7849_,
    new_n7850_, new_n7851_, new_n7852_, new_n7853_, new_n7854_, new_n7855_,
    new_n7856_, new_n7857_, new_n7858_, new_n7859_, new_n7860_, new_n7861_,
    new_n7862_, new_n7863_, new_n7864_, new_n7865_, new_n7866_, new_n7867_,
    new_n7868_, new_n7869_, new_n7870_, new_n7871_, new_n7872_, new_n7873_,
    new_n7874_, new_n7875_, new_n7876_, new_n7877_, new_n7878_, new_n7879_,
    new_n7880_, new_n7881_, new_n7882_, new_n7883_, new_n7884_, new_n7885_,
    new_n7886_, new_n7887_, new_n7888_, new_n7889_, new_n7890_, new_n7891_,
    new_n7892_, new_n7893_, new_n7894_, new_n7895_, new_n7896_, new_n7897_,
    new_n7898_, new_n7899_, new_n7900_, new_n7901_, new_n7902_, new_n7903_,
    new_n7904_, new_n7905_, new_n7906_, new_n7907_, new_n7908_, new_n7909_,
    new_n7910_, new_n7911_, new_n7912_, new_n7913_, new_n7914_, new_n7915_,
    new_n7916_, new_n7917_, new_n7918_, new_n7919_, new_n7920_, new_n7921_,
    new_n7922_, new_n7923_, new_n7924_, new_n7925_, new_n7926_, new_n7927_,
    new_n7928_, new_n7929_, new_n7930_, new_n7931_, new_n7932_, new_n7933_,
    new_n7934_, new_n7935_, new_n7936_, new_n7937_, new_n7938_, new_n7939_,
    new_n7940_, new_n7941_, new_n7942_, new_n7943_, new_n7944_, new_n7945_,
    new_n7946_, new_n7947_, new_n7948_, new_n7949_, new_n7950_, new_n7951_,
    new_n7952_, new_n7953_, new_n7954_, new_n7955_, new_n7956_, new_n7957_,
    new_n7958_, new_n7959_, new_n7960_, new_n7961_, new_n7962_, new_n7963_,
    new_n7964_, new_n7965_, new_n7966_, new_n7967_, new_n7968_, new_n7969_,
    new_n7970_, new_n7971_, new_n7972_, new_n7973_, new_n7974_, new_n7975_,
    new_n7976_, new_n7977_, new_n7978_, new_n7979_, new_n7980_, new_n7981_,
    new_n7982_, new_n7983_, new_n7984_, new_n7985_, new_n7986_, new_n7987_,
    new_n7988_, new_n7989_, new_n7990_, new_n7991_, new_n7992_, new_n7993_,
    new_n7994_, new_n7995_, new_n7996_, new_n7997_, new_n7998_, new_n7999_,
    new_n8000_, new_n8001_, new_n8002_, new_n8003_, new_n8004_, new_n8005_,
    new_n8006_, new_n8007_, new_n8008_, new_n8009_, new_n8010_, new_n8011_,
    new_n8012_, new_n8013_, new_n8014_, new_n8015_, new_n8016_, new_n8017_,
    new_n8018_, new_n8019_, new_n8020_, new_n8021_, new_n8022_, new_n8023_,
    new_n8024_, new_n8025_, new_n8026_, new_n8027_, new_n8028_, new_n8029_,
    new_n8030_, new_n8031_, new_n8032_, new_n8033_, new_n8034_, new_n8035_,
    new_n8036_, new_n8037_, new_n8038_, new_n8039_, new_n8040_, new_n8041_,
    new_n8042_, new_n8043_, new_n8044_, new_n8045_, new_n8046_, new_n8047_,
    new_n8048_, new_n8049_, new_n8050_, new_n8051_, new_n8052_, new_n8053_,
    new_n8054_, new_n8055_, new_n8056_, new_n8057_, new_n8058_, new_n8059_,
    new_n8060_, new_n8061_, new_n8062_, new_n8063_, new_n8064_, new_n8065_,
    new_n8066_, new_n8067_, new_n8068_, new_n8069_, new_n8070_, new_n8071_,
    new_n8072_, new_n8073_, new_n8074_, new_n8075_, new_n8076_, new_n8077_,
    new_n8078_, new_n8079_, new_n8080_, new_n8081_, new_n8082_, new_n8083_,
    new_n8084_, new_n8085_, new_n8086_, new_n8087_, new_n8088_, new_n8089_,
    new_n8090_, new_n8091_, new_n8092_, new_n8093_, new_n8094_, new_n8095_,
    new_n8096_, new_n8097_, new_n8098_, new_n8099_, new_n8100_, new_n8101_,
    new_n8102_, new_n8103_, new_n8104_, new_n8105_, new_n8106_, new_n8107_,
    new_n8108_, new_n8109_, new_n8110_, new_n8111_, new_n8112_, new_n8113_,
    new_n8114_, new_n8115_, new_n8116_, new_n8117_, new_n8118_, new_n8119_,
    new_n8120_, new_n8121_, new_n8122_, new_n8123_, new_n8124_, new_n8125_,
    new_n8126_, new_n8127_, new_n8128_, new_n8129_, new_n8130_, new_n8131_,
    new_n8132_, new_n8133_, new_n8134_, new_n8135_, new_n8136_, new_n8137_,
    new_n8138_, new_n8139_, new_n8140_, new_n8141_, new_n8142_, new_n8143_,
    new_n8144_, new_n8145_, new_n8146_, new_n8147_, new_n8148_, new_n8149_,
    new_n8150_, new_n8151_, new_n8152_, new_n8153_, new_n8154_, new_n8155_,
    new_n8156_, new_n8157_, new_n8158_, new_n8159_, new_n8160_, new_n8161_,
    new_n8162_, new_n8163_, new_n8164_, new_n8165_, new_n8166_, new_n8167_,
    new_n8168_, new_n8169_, new_n8170_, new_n8171_, new_n8172_, new_n8173_,
    new_n8174_, new_n8175_, new_n8176_, new_n8177_, new_n8178_, new_n8179_,
    new_n8180_, new_n8181_, new_n8182_, new_n8183_, new_n8184_, new_n8185_,
    new_n8186_, new_n8187_, new_n8188_, new_n8189_, new_n8190_, new_n8191_,
    new_n8192_, new_n8193_, new_n8194_, new_n8195_, new_n8196_, new_n8197_,
    new_n8198_, new_n8199_, new_n8200_, new_n8201_, new_n8202_, new_n8203_,
    new_n8204_, new_n8205_, new_n8206_, new_n8207_, new_n8208_, new_n8209_,
    new_n8210_, new_n8211_, new_n8212_, new_n8213_, new_n8214_, new_n8215_,
    new_n8216_, new_n8217_, new_n8218_, new_n8219_, new_n8220_, new_n8221_,
    new_n8222_, new_n8223_, new_n8224_, new_n8225_, new_n8226_, new_n8227_,
    new_n8228_, new_n8229_, new_n8230_, new_n8231_, new_n8232_, new_n8233_,
    new_n8234_, new_n8235_, new_n8236_, new_n8237_, new_n8238_, new_n8239_,
    new_n8240_, new_n8241_, new_n8242_, new_n8243_, new_n8244_, new_n8245_,
    new_n8246_, new_n8247_, new_n8248_, new_n8249_, new_n8250_, new_n8251_,
    new_n8252_, new_n8253_, new_n8254_, new_n8255_, new_n8256_, new_n8257_,
    new_n8258_, new_n8259_, new_n8260_, new_n8261_, new_n8262_, new_n8263_,
    new_n8264_, new_n8265_, new_n8266_, new_n8267_, new_n8268_, new_n8269_,
    new_n8270_, new_n8271_, new_n8272_, new_n8273_, new_n8274_, new_n8275_,
    new_n8276_, new_n8277_, new_n8278_, new_n8279_, new_n8280_, new_n8281_,
    new_n8282_, new_n8283_, new_n8284_, new_n8285_, new_n8286_, new_n8287_,
    new_n8288_, new_n8289_, new_n8290_, new_n8291_, new_n8292_, new_n8293_,
    new_n8294_, new_n8295_, new_n8296_, new_n8297_, new_n8298_, new_n8299_,
    new_n8300_, new_n8301_, new_n8302_, new_n8303_, new_n8304_, new_n8305_,
    new_n8306_, new_n8307_, new_n8308_, new_n8309_, new_n8310_, new_n8311_,
    new_n8312_, new_n8313_, new_n8314_, new_n8315_, new_n8316_, new_n8317_,
    new_n8318_, new_n8319_, new_n8320_, new_n8321_, new_n8322_, new_n8323_,
    new_n8324_, new_n8325_, new_n8326_, new_n8327_, new_n8328_, new_n8329_,
    new_n8330_, new_n8331_, new_n8332_, new_n8333_, new_n8334_, new_n8335_,
    new_n8336_, new_n8337_, new_n8338_, new_n8339_, new_n8340_, new_n8341_,
    new_n8342_, new_n8343_, new_n8344_, new_n8345_, new_n8346_, new_n8347_,
    new_n8348_, new_n8349_, new_n8350_, new_n8351_, new_n8352_, new_n8353_,
    new_n8354_, new_n8355_, new_n8356_, new_n8357_, new_n8358_, new_n8359_,
    new_n8360_, new_n8361_, new_n8362_, new_n8363_, new_n8364_, new_n8365_,
    new_n8366_, new_n8367_, new_n8368_, new_n8369_, new_n8370_, new_n8371_,
    new_n8372_, new_n8373_, new_n8374_, new_n8375_, new_n8376_, new_n8377_,
    new_n8378_, new_n8379_, new_n8380_, new_n8381_, new_n8382_, new_n8383_,
    new_n8384_, new_n8385_, new_n8386_, new_n8387_, new_n8388_, new_n8389_,
    new_n8390_, new_n8391_, new_n8392_, new_n8393_, new_n8394_, new_n8395_,
    new_n8396_, new_n8397_, new_n8398_, new_n8399_, new_n8400_, new_n8401_,
    new_n8402_, new_n8403_, new_n8404_, new_n8405_, new_n8406_, new_n8407_,
    new_n8408_, new_n8409_, new_n8410_, new_n8411_, new_n8412_, new_n8413_,
    new_n8414_, new_n8415_, new_n8416_, new_n8417_, new_n8418_, new_n8419_,
    new_n8420_, new_n8421_, new_n8422_, new_n8423_, new_n8424_, new_n8425_,
    new_n8426_, new_n8427_, new_n8428_, new_n8429_, new_n8430_, new_n8431_,
    new_n8432_, new_n8433_, new_n8434_, new_n8435_, new_n8436_, new_n8437_,
    new_n8438_, new_n8439_, new_n8440_, new_n8441_, new_n8442_, new_n8443_,
    new_n8444_, new_n8445_, new_n8446_, new_n8447_, new_n8448_, new_n8449_,
    new_n8450_, new_n8451_, new_n8452_, new_n8453_, new_n8454_, new_n8455_,
    new_n8456_, new_n8457_, new_n8458_, new_n8459_, new_n8460_, new_n8461_,
    new_n8462_, new_n8463_, new_n8464_, new_n8465_, new_n8466_, new_n8467_,
    new_n8468_, new_n8469_, new_n8470_, new_n8471_, new_n8472_, new_n8473_,
    new_n8474_, new_n8475_, new_n8476_, new_n8477_, new_n8478_, new_n8479_,
    new_n8480_, new_n8481_, new_n8482_, new_n8483_, new_n8484_, new_n8485_,
    new_n8486_, new_n8487_, new_n8488_, new_n8489_, new_n8490_, new_n8491_,
    new_n8492_, new_n8493_, new_n8494_, new_n8495_, new_n8496_, new_n8497_,
    new_n8498_, new_n8499_, new_n8500_, new_n8501_, new_n8502_, new_n8503_,
    new_n8504_, new_n8505_, new_n8506_, new_n8507_, new_n8508_, new_n8509_,
    new_n8510_, new_n8511_, new_n8512_, new_n8513_, new_n8514_, new_n8515_,
    new_n8516_, new_n8517_, new_n8518_, new_n8519_, new_n8520_, new_n8521_,
    new_n8522_, new_n8523_, new_n8524_, new_n8525_, new_n8526_, new_n8527_,
    new_n8528_, new_n8529_, new_n8530_, new_n8531_, new_n8532_, new_n8533_,
    new_n8534_, new_n8535_, new_n8536_, new_n8537_, new_n8538_, new_n8539_,
    new_n8540_, new_n8541_, new_n8542_, new_n8543_, new_n8544_, new_n8545_,
    new_n8546_, new_n8547_, new_n8548_, new_n8549_, new_n8550_, new_n8551_,
    new_n8552_, new_n8553_, new_n8554_, new_n8555_, new_n8556_, new_n8557_,
    new_n8558_, new_n8559_, new_n8560_, new_n8561_, new_n8562_, new_n8563_,
    new_n8564_, new_n8565_, new_n8566_, new_n8567_, new_n8568_, new_n8569_,
    new_n8570_, new_n8571_, new_n8572_, new_n8573_, new_n8574_, new_n8575_,
    new_n8576_, new_n8577_, new_n8578_, new_n8579_, new_n8580_, new_n8581_,
    new_n8582_, new_n8583_, new_n8584_, new_n8585_, new_n8586_, new_n8587_,
    new_n8588_, new_n8589_, new_n8590_, new_n8591_, new_n8592_, new_n8593_,
    new_n8594_, new_n8595_, new_n8596_, new_n8597_, new_n8598_, new_n8599_,
    new_n8600_, new_n8601_, new_n8602_, new_n8603_, new_n8604_, new_n8605_,
    new_n8606_, new_n8607_, new_n8608_, new_n8609_, new_n8610_, new_n8611_,
    new_n8612_, new_n8613_, new_n8614_, new_n8615_, new_n8616_, new_n8617_,
    new_n8618_, new_n8619_, new_n8620_, new_n8621_, new_n8622_, new_n8623_,
    new_n8624_, new_n8625_, new_n8626_, new_n8627_, new_n8628_, new_n8629_,
    new_n8630_, new_n8631_, new_n8632_, new_n8633_, new_n8634_, new_n8635_,
    new_n8636_, new_n8637_, new_n8638_, new_n8639_, new_n8640_, new_n8641_,
    new_n8642_, new_n8643_, new_n8644_, new_n8645_, new_n8646_, new_n8647_,
    new_n8648_, new_n8649_, new_n8650_, new_n8651_, new_n8652_, new_n8653_,
    new_n8654_, new_n8655_, new_n8656_, new_n8657_, new_n8658_, new_n8659_,
    new_n8660_, new_n8661_, new_n8662_, new_n8663_, new_n8664_, new_n8665_,
    new_n8666_, new_n8667_, new_n8668_, new_n8669_, new_n8670_, new_n8671_,
    new_n8672_, new_n8673_, new_n8674_, new_n8675_, new_n8676_, new_n8677_,
    new_n8678_, new_n8679_, new_n8680_, new_n8681_, new_n8682_, new_n8683_,
    new_n8684_, new_n8685_, new_n8686_, new_n8687_, new_n8688_, new_n8689_,
    new_n8690_, new_n8691_, new_n8692_, new_n8693_, new_n8694_, new_n8695_,
    new_n8696_, new_n8697_, new_n8698_, new_n8699_, new_n8700_, new_n8701_,
    new_n8702_, new_n8703_, new_n8704_, new_n8705_, new_n8706_, new_n8707_,
    new_n8708_, new_n8709_, new_n8710_, new_n8711_, new_n8712_, new_n8713_,
    new_n8714_, new_n8715_, new_n8716_, new_n8717_, new_n8718_, new_n8719_,
    new_n8720_, new_n8721_, new_n8722_, new_n8723_, new_n8724_, new_n8725_,
    new_n8726_, new_n8727_, new_n8728_, new_n8729_, new_n8730_, new_n8731_,
    new_n8732_, new_n8733_, new_n8734_, new_n8735_, new_n8736_, new_n8737_,
    new_n8738_, new_n8739_, new_n8740_, new_n8741_, new_n8742_, new_n8743_,
    new_n8744_, new_n8745_, new_n8746_, new_n8747_, new_n8748_, new_n8749_,
    new_n8750_, new_n8751_, new_n8752_, new_n8753_, new_n8754_, new_n8755_,
    new_n8756_, new_n8757_, new_n8758_, new_n8759_, new_n8760_, new_n8761_,
    new_n8762_, new_n8763_, new_n8764_, new_n8765_, new_n8766_, new_n8767_,
    new_n8768_, new_n8769_, new_n8770_, new_n8771_, new_n8772_, new_n8773_,
    new_n8774_, new_n8775_, new_n8776_, new_n8777_, new_n8778_, new_n8779_,
    new_n8780_, new_n8781_, new_n8782_, new_n8783_, new_n8784_, new_n8785_,
    new_n8786_, new_n8787_, new_n8788_, new_n8789_, new_n8790_, new_n8791_,
    new_n8792_, new_n8793_, new_n8794_, new_n8795_, new_n8796_, new_n8797_,
    new_n8798_, new_n8799_, new_n8800_, new_n8801_, new_n8802_, new_n8803_,
    new_n8804_, new_n8805_, new_n8806_, new_n8807_, new_n8808_, new_n8809_,
    new_n8810_, new_n8811_, new_n8812_, new_n8813_, new_n8814_, new_n8815_,
    new_n8816_, new_n8817_, new_n8818_, new_n8819_, new_n8820_, new_n8821_,
    new_n8822_, new_n8823_, new_n8824_, new_n8825_, new_n8826_, new_n8827_,
    new_n8828_, new_n8829_, new_n8830_, new_n8831_, new_n8832_, new_n8833_,
    new_n8834_, new_n8835_, new_n8836_, new_n8837_, new_n8838_, new_n8839_,
    new_n8840_, new_n8841_, new_n8842_, new_n8843_, new_n8844_, new_n8845_,
    new_n8846_, new_n8847_, new_n8848_, new_n8849_, new_n8850_, new_n8851_,
    new_n8852_, new_n8853_, new_n8854_, new_n8855_, new_n8856_, new_n8857_,
    new_n8858_, new_n8859_, new_n8860_, new_n8861_, new_n8862_, new_n8863_,
    new_n8864_, new_n8865_, new_n8866_, new_n8867_, new_n8868_, new_n8869_,
    new_n8870_, new_n8871_, new_n8872_, new_n8873_, new_n8874_, new_n8875_,
    new_n8876_, new_n8877_, new_n8878_, new_n8879_, new_n8880_, new_n8881_,
    new_n8882_, new_n8883_, new_n8884_, new_n8885_, new_n8886_, new_n8887_,
    new_n8888_, new_n8889_, new_n8890_, new_n8891_, new_n8892_, new_n8893_,
    new_n8894_, new_n8895_, new_n8896_, new_n8897_, new_n8898_, new_n8899_,
    new_n8900_, new_n8901_, new_n8902_, new_n8903_, new_n8904_, new_n8905_,
    new_n8906_, new_n8907_, new_n8908_, new_n8909_, new_n8910_, new_n8911_,
    new_n8912_, new_n8913_, new_n8914_, new_n8915_, new_n8916_, new_n8917_,
    new_n8918_, new_n8919_, new_n8920_, new_n8921_, new_n8922_, new_n8923_,
    new_n8924_, new_n8925_, new_n8926_, new_n8927_, new_n8928_, new_n8929_,
    new_n8930_, new_n8931_, new_n8932_, new_n8933_, new_n8934_, new_n8935_,
    new_n8936_, new_n8937_, new_n8938_, new_n8939_, new_n8940_, new_n8941_,
    new_n8942_, new_n8943_, new_n8944_, new_n8945_, new_n8946_, new_n8947_,
    new_n8948_, new_n8949_, new_n8950_, new_n8951_, new_n8952_, new_n8953_,
    new_n8954_, new_n8955_, new_n8956_, new_n8957_, new_n8958_, new_n8959_,
    new_n8960_, new_n8961_, new_n8962_, new_n8963_, new_n8964_, new_n8965_,
    new_n8966_, new_n8967_, new_n8968_, new_n8969_, new_n8970_, new_n8971_,
    new_n8972_, new_n8973_, new_n8974_, new_n8975_, new_n8976_, new_n8977_,
    new_n8978_, new_n8979_, new_n8980_, new_n8981_, new_n8982_, new_n8983_,
    new_n8984_, new_n8985_, new_n8986_, new_n8987_, new_n8988_, new_n8989_,
    new_n8990_, new_n8991_, new_n8992_, new_n8993_, new_n8994_, new_n8995_,
    new_n8996_, new_n8997_, new_n8998_, new_n8999_, new_n9000_, new_n9001_,
    new_n9002_, new_n9003_, new_n9004_, new_n9005_, new_n9006_, new_n9007_,
    new_n9008_, new_n9009_, new_n9010_, new_n9011_, new_n9012_, new_n9013_,
    new_n9014_, new_n9015_, new_n9016_, new_n9017_, new_n9018_, new_n9019_,
    new_n9020_, new_n9021_, new_n9022_, new_n9023_, new_n9024_, new_n9025_,
    new_n9026_, new_n9027_, new_n9028_, new_n9029_, new_n9030_, new_n9031_,
    new_n9032_, new_n9033_, new_n9034_, new_n9035_, new_n9036_, new_n9037_,
    new_n9038_, new_n9039_, new_n9040_, new_n9041_, new_n9042_, new_n9043_,
    new_n9044_, new_n9045_, new_n9046_, new_n9047_, new_n9048_, new_n9049_,
    new_n9050_, new_n9051_, new_n9052_, new_n9053_, new_n9054_, new_n9055_,
    new_n9056_, new_n9057_, new_n9058_, new_n9059_, new_n9060_, new_n9061_,
    new_n9062_, new_n9063_, new_n9064_, new_n9065_, new_n9066_, new_n9067_,
    new_n9068_, new_n9069_, new_n9070_, new_n9071_, new_n9072_, new_n9073_,
    new_n9074_, new_n9075_, new_n9076_, new_n9077_, new_n9078_, new_n9079_,
    new_n9080_, new_n9081_, new_n9082_, new_n9083_, new_n9084_, new_n9085_,
    new_n9086_, new_n9087_, new_n9088_, new_n9089_, new_n9090_, new_n9091_,
    new_n9092_, new_n9093_, new_n9094_, new_n9095_, new_n9096_, new_n9097_,
    new_n9098_, new_n9099_, new_n9100_, new_n9101_, new_n9102_, new_n9103_,
    new_n9104_, new_n9105_, new_n9106_, new_n9107_, new_n9108_, new_n9109_,
    new_n9110_, new_n9111_, new_n9112_, new_n9113_, new_n9114_, new_n9115_,
    new_n9116_, new_n9117_, new_n9118_, new_n9119_, new_n9120_, new_n9121_,
    new_n9122_, new_n9123_, new_n9124_, new_n9125_, new_n9126_, new_n9127_,
    new_n9128_, new_n9129_, new_n9130_, new_n9131_, new_n9132_, new_n9133_,
    new_n9134_, new_n9135_, new_n9136_, new_n9137_, new_n9138_, new_n9139_,
    new_n9140_, new_n9141_, new_n9142_, new_n9143_, new_n9144_, new_n9145_,
    new_n9146_, new_n9147_, new_n9148_, new_n9149_, new_n9150_, new_n9151_,
    new_n9152_, new_n9153_, new_n9154_, new_n9155_, new_n9156_, new_n9157_,
    new_n9158_, new_n9159_, new_n9160_, new_n9161_, new_n9162_, new_n9163_,
    new_n9164_, new_n9165_, new_n9166_, new_n9167_, new_n9168_, new_n9169_,
    new_n9170_, new_n9171_, new_n9172_, new_n9173_, new_n9174_, new_n9175_,
    new_n9176_, new_n9177_, new_n9178_, new_n9179_, new_n9180_, new_n9181_,
    new_n9182_, new_n9183_, new_n9184_, new_n9185_, new_n9186_, new_n9187_,
    new_n9188_, new_n9189_, new_n9190_, new_n9191_, new_n9192_, new_n9193_,
    new_n9194_, new_n9195_, new_n9196_, new_n9197_, new_n9198_, new_n9199_,
    new_n9200_, new_n9201_, new_n9202_, new_n9203_, new_n9204_, new_n9205_,
    new_n9206_, new_n9207_, new_n9208_, new_n9209_, new_n9210_, new_n9211_,
    new_n9212_, new_n9213_, new_n9214_, new_n9215_, new_n9216_, new_n9217_,
    new_n9218_, new_n9219_, new_n9220_, new_n9221_, new_n9222_, new_n9223_,
    new_n9224_, new_n9225_, new_n9226_, new_n9227_, new_n9228_, new_n9229_,
    new_n9230_, new_n9231_, new_n9232_, new_n9233_, new_n9234_, new_n9235_,
    new_n9236_, new_n9237_, new_n9238_, new_n9239_, new_n9240_, new_n9241_,
    new_n9242_, new_n9243_, new_n9244_, new_n9245_, new_n9246_, new_n9247_,
    new_n9248_, new_n9249_, new_n9250_, new_n9251_, new_n9252_, new_n9253_,
    new_n9254_, new_n9255_, new_n9256_, new_n9257_, new_n9258_, new_n9259_,
    new_n9260_, new_n9261_, new_n9262_, new_n9263_, new_n9264_, new_n9265_,
    new_n9266_, new_n9267_, new_n9268_, new_n9269_, new_n9270_, new_n9271_,
    new_n9272_, new_n9273_, new_n9274_, new_n9275_, new_n9276_, new_n9277_,
    new_n9278_, new_n9279_, new_n9280_, new_n9281_, new_n9282_, new_n9283_,
    new_n9284_, new_n9285_, new_n9286_, new_n9287_, new_n9288_, new_n9289_,
    new_n9290_, new_n9291_, new_n9292_, new_n9293_, new_n9294_, new_n9295_,
    new_n9296_, new_n9297_, new_n9298_, new_n9299_, new_n9300_, new_n9301_,
    new_n9302_, new_n9303_, new_n9304_, new_n9305_, new_n9306_, new_n9307_,
    new_n9308_, new_n9309_, new_n9310_, new_n9311_, new_n9312_, new_n9313_,
    new_n9314_, new_n9315_, new_n9316_, new_n9317_, new_n9318_, new_n9319_,
    new_n9320_, new_n9321_, new_n9322_, new_n9323_, new_n9324_, new_n9325_,
    new_n9326_, new_n9327_, new_n9328_, new_n9329_, new_n9330_, new_n9331_,
    new_n9332_, new_n9333_, new_n9334_, new_n9335_, new_n9336_, new_n9337_,
    new_n9338_, new_n9339_, new_n9340_, new_n9341_, new_n9342_, new_n9343_,
    new_n9344_, new_n9345_, new_n9346_, new_n9347_, new_n9348_, new_n9349_,
    new_n9350_, new_n9351_, new_n9352_, new_n9353_, new_n9354_, new_n9355_,
    new_n9356_, new_n9357_, new_n9358_, new_n9359_, new_n9360_, new_n9361_,
    new_n9362_, new_n9363_, new_n9364_, new_n9365_, new_n9366_, new_n9367_,
    new_n9368_, new_n9369_, new_n9370_, new_n9371_, new_n9372_, new_n9373_,
    new_n9374_, new_n9375_, new_n9376_, new_n9377_, new_n9378_, new_n9379_,
    new_n9380_, new_n9381_, new_n9382_, new_n9383_, new_n9384_, new_n9385_,
    new_n9386_, new_n9387_, new_n9388_, new_n9389_, new_n9390_, new_n9391_,
    new_n9392_, new_n9393_, new_n9394_, new_n9395_, new_n9396_, new_n9397_,
    new_n9398_, new_n9399_, new_n9400_, new_n9401_, new_n9402_, new_n9403_,
    new_n9404_, new_n9405_, new_n9406_, new_n9407_, new_n9408_, new_n9409_,
    new_n9410_, new_n9411_, new_n9412_, new_n9413_, new_n9414_, new_n9415_,
    new_n9416_, new_n9417_, new_n9418_, new_n9419_, new_n9420_, new_n9421_,
    new_n9422_, new_n9423_, new_n9424_, new_n9425_, new_n9426_, new_n9427_,
    new_n9428_, new_n9429_, new_n9430_, new_n9431_, new_n9432_, new_n9433_,
    new_n9434_, new_n9435_, new_n9436_, new_n9437_, new_n9438_, new_n9439_,
    new_n9440_, new_n9441_, new_n9442_, new_n9443_, new_n9444_, new_n9445_,
    new_n9446_, new_n9447_, new_n9448_, new_n9449_, new_n9450_, new_n9451_,
    new_n9452_, new_n9453_, new_n9454_, new_n9455_, new_n9456_, new_n9457_,
    new_n9458_, new_n9459_, new_n9460_, new_n9461_, new_n9462_, new_n9463_,
    new_n9464_, new_n9465_, new_n9466_, new_n9467_, new_n9468_, new_n9469_,
    new_n9470_, new_n9471_, new_n9472_, new_n9473_, new_n9474_, new_n9475_,
    new_n9476_, new_n9477_, new_n9478_, new_n9479_, new_n9480_, new_n9481_,
    new_n9482_, new_n9483_, new_n9484_, new_n9485_, new_n9486_, new_n9487_,
    new_n9488_, new_n9489_, new_n9490_, new_n9491_, new_n9492_, new_n9493_,
    new_n9494_, new_n9495_, new_n9496_, new_n9497_, new_n9498_, new_n9499_,
    new_n9500_, new_n9501_, new_n9502_, new_n9503_, new_n9504_, new_n9505_,
    new_n9506_, new_n9507_, new_n9508_, new_n9509_, new_n9510_, new_n9511_,
    new_n9512_, new_n9513_, new_n9514_, new_n9515_, new_n9516_, new_n9517_,
    new_n9518_, new_n9519_, new_n9520_, new_n9521_, new_n9522_, new_n9523_,
    new_n9524_, new_n9525_, new_n9526_, new_n9527_, new_n9528_, new_n9529_,
    new_n9530_, new_n9531_, new_n9532_, new_n9533_, new_n9534_, new_n9535_,
    new_n9536_, new_n9537_, new_n9538_, new_n9539_, new_n9540_, new_n9541_,
    new_n9542_, new_n9543_, new_n9544_, new_n9545_, new_n9546_, new_n9547_,
    new_n9548_, new_n9549_, new_n9550_, new_n9551_, new_n9552_, new_n9553_,
    new_n9554_, new_n9555_, new_n9556_, new_n9557_, new_n9558_, new_n9559_,
    new_n9560_, new_n9561_, new_n9562_, new_n9563_, new_n9564_, new_n9565_,
    new_n9566_, new_n9567_, new_n9568_, new_n9569_, new_n9570_, new_n9571_,
    new_n9572_, new_n9573_, new_n9574_, new_n9575_, new_n9576_, new_n9577_,
    new_n9578_, new_n9579_, new_n9580_, new_n9581_, new_n9582_, new_n9583_,
    new_n9584_, new_n9585_, new_n9586_, new_n9587_, new_n9588_, new_n9589_,
    new_n9590_, new_n9591_, new_n9592_, new_n9593_, new_n9594_, new_n9595_,
    new_n9596_, new_n9597_, new_n9598_, new_n9599_, new_n9600_, new_n9601_,
    new_n9602_, new_n9603_, new_n9604_, new_n9605_, new_n9606_, new_n9607_,
    new_n9608_, new_n9609_, new_n9610_, new_n9611_, new_n9612_, new_n9613_,
    new_n9614_, new_n9615_, new_n9616_, new_n9617_, new_n9618_, new_n9619_,
    new_n9620_, new_n9621_, new_n9622_, new_n9623_, new_n9624_, new_n9625_,
    new_n9626_, new_n9627_, new_n9628_, new_n9629_, new_n9630_, new_n9631_,
    new_n9632_, new_n9633_, new_n9634_, new_n9635_, new_n9636_, new_n9637_,
    new_n9638_, new_n9639_, new_n9640_, new_n9641_, new_n9642_, new_n9643_,
    new_n9644_, new_n9645_, new_n9646_, new_n9647_, new_n9648_, new_n9649_,
    new_n9650_, new_n9651_, new_n9652_, new_n9653_, new_n9654_, new_n9655_,
    new_n9656_, new_n9657_, new_n9658_, new_n9659_, new_n9660_, new_n9661_,
    new_n9662_, new_n9663_, new_n9664_, new_n9665_, new_n9666_, new_n9667_,
    new_n9668_, new_n9669_, new_n9670_, new_n9671_, new_n9672_, new_n9673_,
    new_n9674_, new_n9675_, new_n9676_, new_n9677_, new_n9678_, new_n9679_,
    new_n9680_, new_n9681_, new_n9682_, new_n9683_, new_n9684_, new_n9685_,
    new_n9686_, new_n9687_, new_n9688_, new_n9689_, new_n9690_, new_n9691_,
    new_n9692_, new_n9693_, new_n9694_, new_n9695_, new_n9696_, new_n9697_,
    new_n9698_, new_n9699_, new_n9700_, new_n9701_, new_n9702_, new_n9703_,
    new_n9704_, new_n9705_, new_n9706_, new_n9707_, new_n9708_, new_n9709_,
    new_n9710_, new_n9711_, new_n9712_, new_n9713_, new_n9714_, new_n9715_,
    new_n9716_, new_n9717_, new_n9718_, new_n9719_, new_n9720_, new_n9721_,
    new_n9722_, new_n9723_, new_n9724_, new_n9725_, new_n9726_, new_n9727_,
    new_n9728_, new_n9729_, new_n9730_, new_n9731_, new_n9732_, new_n9733_,
    new_n9734_, new_n9735_, new_n9736_, new_n9737_, new_n9738_, new_n9739_,
    new_n9740_, new_n9741_, new_n9742_, new_n9743_, new_n9744_, new_n9745_,
    new_n9746_, new_n9747_, new_n9748_, new_n9749_, new_n9750_, new_n9751_,
    new_n9752_, new_n9753_, new_n9754_, new_n9755_, new_n9756_, new_n9757_,
    new_n9758_, new_n9759_, new_n9760_, new_n9761_, new_n9762_, new_n9763_,
    new_n9764_, new_n9765_, new_n9766_, new_n9767_, new_n9768_, new_n9769_,
    new_n9770_, new_n9771_, new_n9772_, new_n9773_, new_n9774_, new_n9775_,
    new_n9776_, new_n9777_, new_n9778_, new_n9779_, new_n9780_, new_n9781_,
    new_n9782_, new_n9783_, new_n9784_, new_n9785_, new_n9786_, new_n9787_,
    new_n9788_, new_n9789_, new_n9790_, new_n9791_, new_n9792_, new_n9793_,
    new_n9794_, new_n9795_, new_n9796_, new_n9797_, new_n9798_, new_n9799_,
    new_n9800_, new_n9801_, new_n9802_, new_n9803_, new_n9804_, new_n9805_,
    new_n9806_, new_n9807_, new_n9808_, new_n9809_, new_n9810_, new_n9811_,
    new_n9812_, new_n9813_, new_n9814_, new_n9815_, new_n9816_, new_n9817_,
    new_n9818_, new_n9819_, new_n9820_, new_n9821_, new_n9822_, new_n9823_,
    new_n9824_, new_n9825_, new_n9826_, new_n9827_, new_n9828_, new_n9829_,
    new_n9830_, new_n9831_, new_n9832_, new_n9833_, new_n9834_, new_n9835_,
    new_n9836_, new_n9837_, new_n9838_, new_n9839_, new_n9840_, new_n9841_,
    new_n9842_, new_n9843_, new_n9844_, new_n9845_, new_n9846_, new_n9847_,
    new_n9848_, new_n9849_, new_n9850_, new_n9851_, new_n9852_, new_n9853_,
    new_n9854_, new_n9855_, new_n9856_, new_n9857_, new_n9858_, new_n9859_,
    new_n9860_, new_n9861_, new_n9862_, new_n9863_, new_n9864_, new_n9865_,
    new_n9866_, new_n9867_, new_n9868_, new_n9869_, new_n9870_, new_n9871_,
    new_n9872_, new_n9873_, new_n9874_, new_n9875_, new_n9876_, new_n9877_,
    new_n9878_, new_n9879_, new_n9880_, new_n9881_, new_n9882_, new_n9883_,
    new_n9884_, new_n9885_, new_n9886_, new_n9887_, new_n9888_, new_n9889_,
    new_n9890_, new_n9891_, new_n9892_, new_n9893_, new_n9894_, new_n9895_,
    new_n9896_, new_n9897_, new_n9898_, new_n9899_, new_n9900_, new_n9901_,
    new_n9902_, new_n9903_, new_n9904_, new_n9905_, new_n9906_, new_n9907_,
    new_n9908_, new_n9909_, new_n9910_, new_n9911_, new_n9912_, new_n9913_,
    new_n9914_, new_n9915_, new_n9916_, new_n9917_, new_n9918_, new_n9919_,
    new_n9920_, new_n9921_, new_n9922_, new_n9923_, new_n9924_, new_n9925_,
    new_n9926_, new_n9927_, new_n9928_, new_n9929_, new_n9930_, new_n9931_,
    new_n9932_, new_n9933_, new_n9934_, new_n9935_, new_n9936_, new_n9937_,
    new_n9938_, new_n9939_, new_n9940_, new_n9941_, new_n9942_, new_n9943_,
    new_n9944_, new_n9945_, new_n9946_, new_n9947_, new_n9948_, new_n9949_,
    new_n9950_, new_n9951_, new_n9952_, new_n9953_, new_n9954_, new_n9955_,
    new_n9956_, new_n9957_, new_n9958_, new_n9959_, new_n9960_, new_n9961_,
    new_n9962_, new_n9963_, new_n9964_, new_n9965_, new_n9966_, new_n9967_,
    new_n9968_, new_n9969_, new_n9970_, new_n9971_, new_n9972_, new_n9973_,
    new_n9974_, new_n9975_, new_n9976_, new_n9977_, new_n9978_, new_n9979_,
    new_n9980_, new_n9981_, new_n9982_, new_n9983_, new_n9984_, new_n9985_,
    new_n9986_, new_n9987_, new_n9988_, new_n9989_, new_n9990_, new_n9991_,
    new_n9992_, new_n9993_, new_n9994_, new_n9995_, new_n9996_, new_n9997_,
    new_n9998_, new_n9999_, new_n10000_, new_n10001_, new_n10002_,
    new_n10003_, new_n10004_, new_n10005_, new_n10006_, new_n10007_,
    new_n10008_, new_n10009_, new_n10010_, new_n10011_, new_n10012_,
    new_n10013_, new_n10014_, new_n10015_, new_n10016_, new_n10017_,
    new_n10018_, new_n10019_, new_n10020_, new_n10021_, new_n10022_,
    new_n10023_, new_n10024_, new_n10025_, new_n10026_, new_n10027_,
    new_n10028_, new_n10029_, new_n10030_, new_n10031_, new_n10032_,
    new_n10033_, new_n10034_, new_n10035_, new_n10036_, new_n10037_,
    new_n10038_, new_n10039_, new_n10040_, new_n10041_, new_n10042_,
    new_n10043_, new_n10044_, new_n10045_, new_n10046_, new_n10047_,
    new_n10048_, new_n10049_, new_n10050_, new_n10051_, new_n10052_,
    new_n10053_, new_n10054_, new_n10055_, new_n10056_, new_n10057_,
    new_n10058_, new_n10059_, new_n10060_, new_n10061_, new_n10062_,
    new_n10063_, new_n10064_, new_n10065_, new_n10066_, new_n10067_,
    new_n10068_, new_n10069_, new_n10070_, new_n10071_, new_n10072_,
    new_n10073_, new_n10074_, new_n10075_, new_n10076_, new_n10077_,
    new_n10078_, new_n10079_, new_n10080_, new_n10081_, new_n10082_,
    new_n10083_, new_n10084_, new_n10085_, new_n10086_, new_n10087_,
    new_n10088_, new_n10089_, new_n10090_, new_n10091_, new_n10092_,
    new_n10093_, new_n10094_, new_n10095_, new_n10096_, new_n10097_,
    new_n10098_, new_n10099_, new_n10100_, new_n10101_, new_n10102_,
    new_n10103_, new_n10104_, new_n10105_, new_n10106_, new_n10107_,
    new_n10108_, new_n10109_, new_n10110_, new_n10111_, new_n10112_,
    new_n10113_, new_n10114_, new_n10115_, new_n10116_, new_n10117_,
    new_n10118_, new_n10119_, new_n10120_, new_n10121_, new_n10122_,
    new_n10123_, new_n10124_, new_n10125_, new_n10126_, new_n10127_,
    new_n10128_, new_n10129_, new_n10130_, new_n10131_, new_n10132_,
    new_n10133_, new_n10134_, new_n10135_, new_n10136_, new_n10137_,
    new_n10138_, new_n10139_, new_n10140_, new_n10141_, new_n10142_,
    new_n10143_, new_n10144_, new_n10145_, new_n10146_, new_n10147_,
    new_n10148_, new_n10149_, new_n10150_, new_n10151_, new_n10152_,
    new_n10153_, new_n10154_, new_n10155_, new_n10156_, new_n10157_,
    new_n10158_, new_n10159_, new_n10160_, new_n10161_, new_n10162_,
    new_n10163_, new_n10164_, new_n10165_, new_n10166_, new_n10167_,
    new_n10168_, new_n10169_, new_n10170_, new_n10171_, new_n10172_,
    new_n10173_, new_n10174_, new_n10175_, new_n10176_, new_n10177_,
    new_n10178_, new_n10179_, new_n10180_, new_n10181_, new_n10182_,
    new_n10183_, new_n10184_, new_n10185_, new_n10186_, new_n10187_,
    new_n10188_, new_n10189_, new_n10190_, new_n10191_, new_n10192_,
    new_n10193_, new_n10194_, new_n10195_, new_n10196_, new_n10197_,
    new_n10198_, new_n10199_, new_n10200_, new_n10201_, new_n10202_,
    new_n10203_, new_n10204_, new_n10205_, new_n10206_, new_n10207_,
    new_n10208_, new_n10209_, new_n10210_, new_n10211_, new_n10212_,
    new_n10213_, new_n10214_, new_n10215_, new_n10216_, new_n10217_,
    new_n10218_, new_n10219_, new_n10220_, new_n10221_, new_n10222_,
    new_n10223_, new_n10224_, new_n10225_, new_n10226_, new_n10227_,
    new_n10228_, new_n10229_, new_n10230_, new_n10231_, new_n10232_,
    new_n10233_, new_n10234_, new_n10235_, new_n10236_, new_n10237_,
    new_n10238_, new_n10239_, new_n10240_, new_n10241_, new_n10242_,
    new_n10243_, new_n10244_, new_n10245_, new_n10246_, new_n10247_,
    new_n10248_, new_n10249_, new_n10250_, new_n10251_, new_n10252_,
    new_n10253_, new_n10254_, new_n10255_, new_n10256_, new_n10257_,
    new_n10258_, new_n10259_, new_n10260_, new_n10261_, new_n10262_,
    new_n10263_, new_n10264_, new_n10265_, new_n10266_, new_n10267_,
    new_n10268_, new_n10269_, new_n10270_, new_n10271_, new_n10272_,
    new_n10273_, new_n10274_, new_n10275_, new_n10276_, new_n10277_,
    new_n10278_, new_n10279_, new_n10280_, new_n10281_, new_n10282_,
    new_n10283_, new_n10284_, new_n10285_, new_n10286_, new_n10287_,
    new_n10288_, new_n10289_, new_n10290_, new_n10291_, new_n10292_,
    new_n10293_, new_n10294_, new_n10295_, new_n10296_, new_n10297_,
    new_n10298_, new_n10299_, new_n10300_, new_n10301_, new_n10302_,
    new_n10303_, new_n10304_, new_n10305_, new_n10306_, new_n10307_,
    new_n10308_, new_n10309_, new_n10310_, new_n10311_, new_n10312_,
    new_n10313_, new_n10314_, new_n10315_, new_n10316_, new_n10317_,
    new_n10318_, new_n10319_, new_n10320_, new_n10321_, new_n10322_,
    new_n10323_, new_n10324_, new_n10325_, new_n10326_, new_n10327_,
    new_n10328_, new_n10329_, new_n10330_, new_n10331_, new_n10332_,
    new_n10333_, new_n10334_, new_n10335_, new_n10336_, new_n10337_,
    new_n10338_, new_n10339_, new_n10340_, new_n10341_, new_n10342_,
    new_n10343_, new_n10344_, new_n10345_, new_n10346_, new_n10347_,
    new_n10348_, new_n10349_, new_n10350_, new_n10351_, new_n10352_,
    new_n10353_, new_n10354_, new_n10355_, new_n10356_, new_n10357_,
    new_n10358_, new_n10359_, new_n10360_, new_n10361_, new_n10362_,
    new_n10363_, new_n10364_, new_n10365_, new_n10366_, new_n10367_,
    new_n10368_, new_n10369_, new_n10370_, new_n10371_, new_n10372_,
    new_n10373_, new_n10374_, new_n10375_, new_n10376_, new_n10377_,
    new_n10378_, new_n10379_, new_n10380_, new_n10381_, new_n10382_,
    new_n10383_, new_n10384_, new_n10385_, new_n10386_, new_n10387_,
    new_n10388_, new_n10389_, new_n10390_, new_n10391_, new_n10392_,
    new_n10393_, new_n10394_, new_n10395_, new_n10396_, new_n10397_,
    new_n10398_, new_n10399_, new_n10400_, new_n10401_, new_n10402_,
    new_n10403_, new_n10404_, new_n10405_, new_n10406_, new_n10407_,
    new_n10408_, new_n10409_, new_n10410_, new_n10411_, new_n10412_,
    new_n10413_, new_n10414_, new_n10415_, new_n10416_, new_n10417_,
    new_n10418_, new_n10419_, new_n10420_, new_n10421_, new_n10422_,
    new_n10423_, new_n10424_, new_n10425_, new_n10426_, new_n10427_,
    new_n10428_, new_n10429_, new_n10430_, new_n10431_, new_n10432_,
    new_n10433_, new_n10434_, new_n10435_, new_n10436_, new_n10437_,
    new_n10438_, new_n10439_, new_n10440_, new_n10441_, new_n10442_,
    new_n10443_, new_n10444_, new_n10445_, new_n10446_, new_n10447_,
    new_n10448_, new_n10449_, new_n10450_, new_n10451_, new_n10452_,
    new_n10453_, new_n10454_, new_n10455_, new_n10456_, new_n10457_,
    new_n10458_, new_n10459_, new_n10460_, new_n10461_, new_n10462_,
    new_n10463_, new_n10464_, new_n10465_, new_n10466_, new_n10467_,
    new_n10468_, new_n10469_, new_n10470_, new_n10471_, new_n10472_,
    new_n10473_, new_n10474_, new_n10475_, new_n10476_, new_n10477_,
    new_n10478_, new_n10479_, new_n10480_, new_n10481_, new_n10482_,
    new_n10483_, new_n10484_, new_n10485_, new_n10486_, new_n10487_,
    new_n10488_, new_n10489_, new_n10490_, new_n10491_, new_n10492_,
    new_n10493_, new_n10494_, new_n10495_, new_n10496_, new_n10497_,
    new_n10498_, new_n10499_, new_n10500_, new_n10501_, new_n10502_,
    new_n10503_, new_n10504_, new_n10505_, new_n10506_, new_n10507_,
    new_n10508_, new_n10509_, new_n10510_, new_n10511_, new_n10512_,
    new_n10513_, new_n10514_, new_n10515_, new_n10516_, new_n10517_,
    new_n10518_, new_n10519_, new_n10520_, new_n10521_, new_n10522_,
    new_n10523_, new_n10524_, new_n10525_, new_n10526_, new_n10527_,
    new_n10528_, new_n10529_, new_n10530_, new_n10531_, new_n10532_,
    new_n10533_, new_n10534_, new_n10535_, new_n10536_, new_n10537_,
    new_n10538_, new_n10539_, new_n10540_, new_n10541_, new_n10542_,
    new_n10543_, new_n10544_, new_n10545_, new_n10546_, new_n10547_,
    new_n10548_, new_n10549_, new_n10550_, new_n10551_, new_n10552_,
    new_n10553_, new_n10554_, new_n10555_, new_n10556_, new_n10557_,
    new_n10558_, new_n10559_, new_n10560_, new_n10561_, new_n10562_,
    new_n10563_, new_n10564_, new_n10565_, new_n10566_, new_n10567_,
    new_n10568_, new_n10569_, new_n10570_, new_n10571_, new_n10572_,
    new_n10573_, new_n10574_, new_n10575_, new_n10576_, new_n10577_,
    new_n10578_, new_n10579_, new_n10580_, new_n10581_, new_n10582_,
    new_n10583_, new_n10584_, new_n10585_, new_n10586_, new_n10587_,
    new_n10588_, new_n10589_, new_n10590_, new_n10591_, new_n10592_,
    new_n10593_, new_n10594_, new_n10595_, new_n10596_, new_n10597_,
    new_n10598_, new_n10599_, new_n10600_, new_n10601_, new_n10602_,
    new_n10603_, new_n10604_, new_n10605_, new_n10606_, new_n10607_,
    new_n10608_, new_n10609_, new_n10610_, new_n10611_, new_n10612_,
    new_n10613_, new_n10614_, new_n10615_, new_n10616_, new_n10617_,
    new_n10618_, new_n10619_, new_n10620_, new_n10621_, new_n10622_,
    new_n10623_, new_n10624_, new_n10625_, new_n10626_, new_n10627_,
    new_n10628_, new_n10629_, new_n10630_, new_n10631_, new_n10632_,
    new_n10633_, new_n10634_, new_n10635_, new_n10636_, new_n10637_,
    new_n10638_, new_n10639_, new_n10640_, new_n10641_, new_n10642_,
    new_n10643_, new_n10644_, new_n10645_, new_n10646_, new_n10647_,
    new_n10648_, new_n10649_, new_n10650_, new_n10651_, new_n10652_,
    new_n10653_, new_n10654_, new_n10655_, new_n10656_, new_n10657_,
    new_n10658_, new_n10659_, new_n10660_, new_n10661_, new_n10662_,
    new_n10663_, new_n10664_, new_n10665_, new_n10666_, new_n10667_,
    new_n10668_, new_n10669_, new_n10670_, new_n10671_, new_n10672_,
    new_n10673_, new_n10674_, new_n10675_, new_n10676_, new_n10677_,
    new_n10678_, new_n10679_, new_n10680_, new_n10681_, new_n10682_,
    new_n10683_, new_n10684_, new_n10685_, new_n10686_, new_n10687_,
    new_n10688_, new_n10689_, new_n10690_, new_n10691_, new_n10692_,
    new_n10693_, new_n10694_, new_n10695_, new_n10696_, new_n10697_,
    new_n10698_, new_n10699_, new_n10700_, new_n10701_, new_n10702_,
    new_n10703_, new_n10704_, new_n10705_, new_n10706_, new_n10707_,
    new_n10708_, new_n10709_, new_n10710_, new_n10711_, new_n10712_,
    new_n10713_, new_n10714_, new_n10715_, new_n10716_, new_n10717_,
    new_n10718_, new_n10719_, new_n10720_, new_n10721_, new_n10722_,
    new_n10723_, new_n10724_, new_n10725_, new_n10726_, new_n10727_,
    new_n10728_, new_n10729_, new_n10730_, new_n10731_, new_n10732_,
    new_n10733_, new_n10734_, new_n10735_, new_n10736_, new_n10737_,
    new_n10738_, new_n10739_, new_n10740_, new_n10741_, new_n10742_,
    new_n10743_, new_n10744_, new_n10745_, new_n10746_, new_n10747_,
    new_n10748_, new_n10749_, new_n10750_, new_n10751_, new_n10752_,
    new_n10753_, new_n10754_, new_n10755_, new_n10756_, new_n10757_,
    new_n10758_, new_n10759_, new_n10760_, new_n10761_, new_n10762_,
    new_n10763_, new_n10764_, new_n10765_, new_n10766_, new_n10767_,
    new_n10768_, new_n10769_, new_n10770_, new_n10771_, new_n10772_,
    new_n10773_, new_n10774_, new_n10775_, new_n10776_, new_n10777_,
    new_n10778_, new_n10779_, new_n10780_, new_n10781_, new_n10782_,
    new_n10783_, new_n10784_, new_n10785_, new_n10786_, new_n10787_,
    new_n10788_, new_n10789_, new_n10790_, new_n10791_, new_n10792_,
    new_n10793_, new_n10794_, new_n10795_, new_n10796_, new_n10797_,
    new_n10798_, new_n10799_, new_n10800_, new_n10801_, new_n10802_,
    new_n10803_, new_n10804_, new_n10805_, new_n10806_, new_n10807_,
    new_n10808_, new_n10809_, new_n10810_, new_n10811_, new_n10812_,
    new_n10813_, new_n10814_, new_n10815_, new_n10816_, new_n10817_,
    new_n10818_, new_n10819_, new_n10820_, new_n10821_, new_n10822_,
    new_n10823_, new_n10824_, new_n10825_, new_n10826_, new_n10827_,
    new_n10828_, new_n10829_, new_n10830_, new_n10831_, new_n10832_,
    new_n10833_, new_n10834_, new_n10835_, new_n10836_, new_n10837_,
    new_n10838_, new_n10839_, new_n10840_, new_n10841_, new_n10842_,
    new_n10843_, new_n10844_, new_n10845_, new_n10846_, new_n10847_,
    new_n10848_, new_n10849_, new_n10850_, new_n10851_, new_n10852_,
    new_n10853_, new_n10854_, new_n10855_, new_n10856_, new_n10857_,
    new_n10858_, new_n10859_, new_n10860_, new_n10861_, new_n10862_,
    new_n10863_, new_n10864_, new_n10865_, new_n10866_, new_n10867_,
    new_n10868_, new_n10869_, new_n10870_, new_n10871_, new_n10872_,
    new_n10873_, new_n10874_, new_n10875_, new_n10876_, new_n10877_,
    new_n10878_, new_n10879_, new_n10880_, new_n10881_, new_n10882_,
    new_n10883_, new_n10884_, new_n10885_, new_n10886_, new_n10887_,
    new_n10888_, new_n10889_, new_n10890_, new_n10891_, new_n10892_,
    new_n10893_, new_n10894_, new_n10895_, new_n10896_, new_n10897_,
    new_n10898_, new_n10899_, new_n10900_, new_n10901_, new_n10902_,
    new_n10903_, new_n10904_, new_n10905_, new_n10906_, new_n10907_,
    new_n10908_, new_n10909_, new_n10910_, new_n10911_, new_n10912_,
    new_n10913_, new_n10914_, new_n10915_, new_n10916_, new_n10917_,
    new_n10918_, new_n10919_, new_n10920_, new_n10921_, new_n10922_,
    new_n10923_, new_n10924_, new_n10925_, new_n10926_, new_n10927_,
    new_n10928_, new_n10929_, new_n10930_, new_n10931_, new_n10932_,
    new_n10933_, new_n10934_, new_n10935_, new_n10936_, new_n10937_,
    new_n10938_, new_n10939_, new_n10940_, new_n10941_, new_n10942_,
    new_n10943_, new_n10944_, new_n10945_, new_n10946_, new_n10947_,
    new_n10948_, new_n10949_, new_n10950_, new_n10951_, new_n10952_,
    new_n10953_, new_n10954_, new_n10955_, new_n10956_, new_n10957_,
    new_n10958_, new_n10959_, new_n10960_, new_n10961_, new_n10962_,
    new_n10963_, new_n10964_, new_n10965_, new_n10966_, new_n10967_,
    new_n10968_, new_n10969_, new_n10970_, new_n10971_, new_n10972_,
    new_n10973_, new_n10974_, new_n10975_, new_n10976_, new_n10977_,
    new_n10978_, new_n10979_, new_n10980_, new_n10981_, new_n10982_,
    new_n10983_, new_n10984_, new_n10985_, new_n10986_, new_n10987_,
    new_n10988_, new_n10989_, new_n10990_, new_n10991_, new_n10992_,
    new_n10993_, new_n10994_, new_n10995_, new_n10996_, new_n10997_,
    new_n10998_, new_n10999_, new_n11000_, new_n11001_, new_n11002_,
    new_n11003_, new_n11004_, new_n11005_, new_n11006_, new_n11007_,
    new_n11008_, new_n11009_, new_n11010_, new_n11011_, new_n11012_,
    new_n11013_, new_n11014_, new_n11015_, new_n11016_, new_n11017_,
    new_n11018_, new_n11019_, new_n11020_, new_n11021_, new_n11022_,
    new_n11023_, new_n11024_, new_n11025_, new_n11026_, new_n11027_,
    new_n11028_, new_n11029_, new_n11030_, new_n11031_, new_n11032_,
    new_n11033_, new_n11034_, new_n11035_, new_n11036_, new_n11037_,
    new_n11038_, new_n11039_, new_n11040_, new_n11041_, new_n11042_,
    new_n11043_, new_n11044_, new_n11045_, new_n11046_, new_n11047_,
    new_n11048_, new_n11049_, new_n11050_, new_n11051_, new_n11052_,
    new_n11053_, new_n11054_, new_n11055_, new_n11056_, new_n11057_,
    new_n11058_, new_n11059_, new_n11060_, new_n11061_, new_n11062_,
    new_n11063_, new_n11064_, new_n11065_, new_n11066_, new_n11067_,
    new_n11068_, new_n11069_, new_n11070_, new_n11071_, new_n11072_,
    new_n11073_, new_n11074_, new_n11075_, new_n11076_, new_n11077_,
    new_n11078_, new_n11079_, new_n11080_, new_n11081_, new_n11082_,
    new_n11083_, new_n11084_, new_n11085_, new_n11086_, new_n11087_,
    new_n11088_, new_n11089_, new_n11090_, new_n11091_, new_n11092_,
    new_n11093_, new_n11094_, new_n11095_, new_n11096_, new_n11097_,
    new_n11098_, new_n11099_, new_n11100_, new_n11101_, new_n11102_,
    new_n11103_, new_n11104_, new_n11105_, new_n11106_, new_n11107_,
    new_n11108_, new_n11109_, new_n11110_, new_n11111_, new_n11112_,
    new_n11113_, new_n11114_, new_n11115_, new_n11116_, new_n11117_,
    new_n11118_, new_n11119_, new_n11120_, new_n11121_, new_n11122_,
    new_n11123_, new_n11124_, new_n11125_, new_n11126_, new_n11127_,
    new_n11128_, new_n11129_, new_n11130_, new_n11131_, new_n11132_,
    new_n11133_, new_n11134_, new_n11135_, new_n11136_, new_n11137_,
    new_n11138_, new_n11139_, new_n11140_, new_n11141_, new_n11142_,
    new_n11143_, new_n11144_, new_n11145_, new_n11146_, new_n11147_,
    new_n11148_, new_n11149_, new_n11150_, new_n11151_, new_n11152_,
    new_n11153_, new_n11154_, new_n11155_, new_n11156_, new_n11157_,
    new_n11158_, new_n11159_, new_n11160_, new_n11161_, new_n11162_,
    new_n11163_, new_n11164_, new_n11165_, new_n11166_, new_n11167_,
    new_n11168_, new_n11169_, new_n11170_, new_n11171_, new_n11172_,
    new_n11173_, new_n11174_, new_n11175_, new_n11176_, new_n11177_,
    new_n11178_, new_n11179_, new_n11180_, new_n11181_, new_n11182_,
    new_n11183_, new_n11184_, new_n11185_, new_n11186_, new_n11187_,
    new_n11188_, new_n11189_, new_n11190_, new_n11191_, new_n11192_,
    new_n11193_, new_n11194_, new_n11195_, new_n11196_, new_n11197_,
    new_n11198_, new_n11199_, new_n11200_, new_n11201_, new_n11202_,
    new_n11203_, new_n11204_, new_n11205_, new_n11206_, new_n11207_,
    new_n11208_, new_n11209_, new_n11210_, new_n11211_, new_n11212_,
    new_n11213_, new_n11214_, new_n11215_, new_n11216_, new_n11217_,
    new_n11218_, new_n11219_, new_n11220_, new_n11221_, new_n11222_,
    new_n11223_, new_n11224_, new_n11225_, new_n11226_, new_n11227_,
    new_n11228_, new_n11229_, new_n11230_, new_n11231_, new_n11232_,
    new_n11233_, new_n11234_, new_n11235_, new_n11236_, new_n11237_,
    new_n11238_, new_n11239_, new_n11240_, new_n11241_, new_n11242_,
    new_n11243_, new_n11244_, new_n11245_, new_n11246_, new_n11247_,
    new_n11248_, new_n11249_, new_n11250_, new_n11251_, new_n11252_,
    new_n11253_, new_n11254_, new_n11255_, new_n11256_, new_n11257_,
    new_n11258_, new_n11259_, new_n11260_, new_n11261_, new_n11262_,
    new_n11263_, new_n11264_, new_n11265_, new_n11266_, new_n11267_,
    new_n11268_, new_n11269_, new_n11270_, new_n11271_, new_n11272_,
    new_n11273_, new_n11274_, new_n11275_, new_n11276_, new_n11277_,
    new_n11278_, new_n11279_, new_n11280_, new_n11281_, new_n11282_,
    new_n11283_, new_n11284_, new_n11285_, new_n11286_, new_n11287_,
    new_n11288_, new_n11289_, new_n11290_, new_n11291_, new_n11292_,
    new_n11293_, new_n11294_, new_n11295_, new_n11296_, new_n11297_,
    new_n11298_, new_n11299_, new_n11300_, new_n11301_, new_n11302_,
    new_n11303_, new_n11304_, new_n11305_, new_n11306_, new_n11307_,
    new_n11308_, new_n11309_, new_n11310_, new_n11311_, new_n11312_,
    new_n11313_, new_n11314_, new_n11315_, new_n11316_, new_n11317_,
    new_n11318_, new_n11319_, new_n11320_, new_n11321_, new_n11322_,
    new_n11323_, new_n11324_, new_n11325_, new_n11326_, new_n11327_,
    new_n11328_, new_n11329_, new_n11330_, new_n11331_, new_n11332_,
    new_n11333_, new_n11334_, new_n11335_, new_n11336_, new_n11337_,
    new_n11338_, new_n11339_, new_n11340_, new_n11341_, new_n11342_,
    new_n11343_, new_n11344_, new_n11345_, new_n11346_, new_n11347_,
    new_n11348_, new_n11349_, new_n11350_, new_n11351_, new_n11352_,
    new_n11353_, new_n11354_, new_n11355_, new_n11356_, new_n11357_,
    new_n11358_, new_n11359_, new_n11360_, new_n11361_, new_n11362_,
    new_n11363_, new_n11364_, new_n11365_, new_n11366_, new_n11367_,
    new_n11368_, new_n11369_, new_n11370_, new_n11371_, new_n11372_,
    new_n11373_, new_n11374_, new_n11375_, new_n11376_, new_n11377_,
    new_n11378_, new_n11379_, new_n11380_, new_n11381_, new_n11382_,
    new_n11383_, new_n11384_, new_n11385_, new_n11386_, new_n11387_,
    new_n11388_, new_n11389_, new_n11390_, new_n11391_, new_n11392_,
    new_n11393_, new_n11394_, new_n11395_, new_n11396_, new_n11397_,
    new_n11398_, new_n11399_, new_n11400_, new_n11401_, new_n11402_,
    new_n11403_, new_n11404_, new_n11405_, new_n11406_, new_n11407_,
    new_n11408_, new_n11409_, new_n11410_, new_n11411_, new_n11412_,
    new_n11413_, new_n11414_, new_n11415_, new_n11416_, new_n11417_,
    new_n11418_, new_n11419_, new_n11420_, new_n11421_, new_n11422_,
    new_n11423_, new_n11424_, new_n11425_, new_n11426_, new_n11427_,
    new_n11428_, new_n11429_, new_n11430_, new_n11431_, new_n11432_,
    new_n11433_, new_n11434_, new_n11435_, new_n11436_, new_n11437_,
    new_n11438_, new_n11439_, new_n11440_, new_n11441_, new_n11442_,
    new_n11443_, new_n11444_, new_n11445_, new_n11446_, new_n11447_,
    new_n11448_, new_n11449_, new_n11450_, new_n11451_, new_n11452_,
    new_n11453_, new_n11454_, new_n11455_, new_n11456_, new_n11457_,
    new_n11458_, new_n11459_, new_n11460_, new_n11461_, new_n11462_,
    new_n11463_, new_n11464_, new_n11465_, new_n11466_, new_n11467_,
    new_n11468_, new_n11469_, new_n11470_, new_n11471_, new_n11472_,
    new_n11473_, new_n11474_, new_n11475_, new_n11476_, new_n11477_,
    new_n11478_, new_n11479_, new_n11480_, new_n11481_, new_n11482_,
    new_n11483_, new_n11484_, new_n11485_, new_n11486_, new_n11487_,
    new_n11488_, new_n11489_, new_n11490_, new_n11491_, new_n11492_,
    new_n11493_, new_n11494_, new_n11495_, new_n11496_, new_n11497_,
    new_n11498_, new_n11499_, new_n11500_, new_n11501_, new_n11502_,
    new_n11503_, new_n11504_, new_n11505_, new_n11506_, new_n11507_,
    new_n11508_, new_n11509_, new_n11510_, new_n11511_, new_n11512_,
    new_n11513_, new_n11514_, new_n11515_, new_n11516_, new_n11517_,
    new_n11518_, new_n11519_, new_n11520_, new_n11521_, new_n11522_,
    new_n11523_, new_n11524_, new_n11525_, new_n11526_, new_n11527_,
    new_n11528_, new_n11529_, new_n11530_, new_n11531_, new_n11532_,
    new_n11533_, new_n11534_, new_n11535_, new_n11536_, new_n11537_,
    new_n11538_, new_n11539_, new_n11540_, new_n11541_, new_n11542_,
    new_n11543_, new_n11544_, new_n11545_, new_n11546_, new_n11547_,
    new_n11548_, new_n11549_, new_n11550_, new_n11551_, new_n11552_,
    new_n11553_, new_n11554_, new_n11555_, new_n11556_, new_n11557_,
    new_n11558_, new_n11559_, new_n11560_, new_n11561_, new_n11562_,
    new_n11563_, new_n11564_, new_n11565_, new_n11566_, new_n11567_,
    new_n11568_, new_n11569_, new_n11570_, new_n11571_, new_n11572_,
    new_n11573_, new_n11574_, new_n11575_, new_n11576_, new_n11577_,
    new_n11578_, new_n11579_, new_n11580_, new_n11581_, new_n11582_,
    new_n11583_, new_n11584_, new_n11585_, new_n11586_, new_n11587_,
    new_n11588_, new_n11589_, new_n11590_, new_n11591_, new_n11592_,
    new_n11593_, new_n11594_, new_n11595_, new_n11596_, new_n11597_,
    new_n11598_, new_n11599_, new_n11600_, new_n11601_, new_n11602_,
    new_n11603_, new_n11604_, new_n11605_, new_n11606_, new_n11607_,
    new_n11608_, new_n11609_, new_n11610_, new_n11611_, new_n11612_,
    new_n11613_, new_n11614_, new_n11615_, new_n11616_, new_n11617_,
    new_n11618_, new_n11619_, new_n11620_, new_n11621_, new_n11622_,
    new_n11623_, new_n11624_, new_n11625_, new_n11626_, new_n11627_,
    new_n11628_, new_n11629_, new_n11630_, new_n11631_, new_n11632_,
    new_n11633_, new_n11634_, new_n11635_, new_n11636_, new_n11637_,
    new_n11638_, new_n11639_, new_n11640_, new_n11641_, new_n11642_,
    new_n11643_, new_n11644_, new_n11645_, new_n11646_, new_n11647_,
    new_n11648_, new_n11649_, new_n11650_, new_n11651_, new_n11652_,
    new_n11653_, new_n11654_, new_n11655_, new_n11656_, new_n11657_,
    new_n11658_, new_n11659_, new_n11660_, new_n11661_, new_n11662_,
    new_n11663_, new_n11664_, new_n11665_, new_n11666_, new_n11667_,
    new_n11668_, new_n11669_, new_n11670_, new_n11671_, new_n11672_,
    new_n11673_, new_n11674_, new_n11675_, new_n11676_, new_n11677_,
    new_n11678_, new_n11679_, new_n11680_, new_n11681_, new_n11682_,
    new_n11683_, new_n11684_, new_n11685_, new_n11686_, new_n11687_,
    new_n11688_, new_n11689_, new_n11690_, new_n11691_, new_n11692_,
    new_n11693_, new_n11694_, new_n11695_, new_n11696_, new_n11697_,
    new_n11698_, new_n11699_, new_n11700_, new_n11701_, new_n11702_,
    new_n11703_, new_n11704_, new_n11705_, new_n11706_, new_n11707_,
    new_n11708_, new_n11709_, new_n11710_, new_n11711_, new_n11712_,
    new_n11713_, new_n11714_, new_n11715_, new_n11716_, new_n11717_,
    new_n11718_, new_n11719_, new_n11720_, new_n11721_, new_n11722_,
    new_n11723_, new_n11724_, new_n11725_, new_n11726_, new_n11727_,
    new_n11728_, new_n11729_, new_n11730_, new_n11731_, new_n11732_,
    new_n11733_, new_n11734_, new_n11735_, new_n11736_, new_n11737_,
    new_n11738_, new_n11739_, new_n11740_, new_n11741_, new_n11742_,
    new_n11743_, new_n11744_, new_n11745_, new_n11746_, new_n11747_,
    new_n11748_, new_n11749_, new_n11750_, new_n11751_, new_n11752_,
    new_n11753_, new_n11754_, new_n11755_, new_n11756_, new_n11757_,
    new_n11758_, new_n11759_, new_n11760_, new_n11761_, new_n11762_,
    new_n11763_, new_n11764_, new_n11765_, new_n11766_, new_n11767_,
    new_n11768_, new_n11769_, new_n11770_, new_n11771_, new_n11772_,
    new_n11773_, new_n11774_, new_n11775_, new_n11776_, new_n11777_,
    new_n11778_, new_n11779_, new_n11780_, new_n11781_, new_n11782_,
    new_n11783_, new_n11784_, new_n11785_, new_n11786_, new_n11787_,
    new_n11788_, new_n11789_, new_n11790_, new_n11791_, new_n11792_,
    new_n11793_, new_n11794_, new_n11795_, new_n11796_, new_n11797_,
    new_n11798_, new_n11799_, new_n11800_, new_n11801_, new_n11802_,
    new_n11803_, new_n11804_, new_n11805_, new_n11806_, new_n11807_,
    new_n11808_, new_n11809_, new_n11810_, new_n11811_, new_n11812_,
    new_n11813_, new_n11814_, new_n11815_, new_n11816_, new_n11817_,
    new_n11818_, new_n11819_, new_n11820_, new_n11821_, new_n11822_,
    new_n11823_, new_n11824_, new_n11825_, new_n11826_, new_n11827_,
    new_n11828_, new_n11829_, new_n11830_, new_n11831_, new_n11832_,
    new_n11833_, new_n11834_, new_n11835_, new_n11836_, new_n11837_,
    new_n11838_, new_n11839_, new_n11840_, new_n11841_, new_n11842_,
    new_n11843_, new_n11844_, new_n11845_, new_n11846_, new_n11847_,
    new_n11848_, new_n11849_, new_n11850_, new_n11851_, new_n11852_,
    new_n11853_, new_n11854_, new_n11855_, new_n11856_, new_n11857_,
    new_n11858_, new_n11859_, new_n11860_, new_n11861_, new_n11862_,
    new_n11863_, new_n11864_, new_n11865_, new_n11866_, new_n11867_,
    new_n11868_, new_n11869_, new_n11870_, new_n11871_, new_n11872_,
    new_n11873_, new_n11874_, new_n11875_, new_n11876_, new_n11877_,
    new_n11878_, new_n11879_, new_n11880_, new_n11881_, new_n11882_,
    new_n11883_, new_n11884_, new_n11885_, new_n11886_, new_n11887_,
    new_n11888_, new_n11889_, new_n11890_, new_n11891_, new_n11892_,
    new_n11893_, new_n11894_, new_n11895_, new_n11896_, new_n11897_,
    new_n11898_, new_n11899_, new_n11900_, new_n11901_, new_n11902_,
    new_n11903_, new_n11904_, new_n11905_, new_n11906_, new_n11907_,
    new_n11908_, new_n11909_, new_n11910_, new_n11911_, new_n11912_,
    new_n11913_, new_n11914_, new_n11915_, new_n11916_, new_n11917_,
    new_n11918_, new_n11919_, new_n11920_, new_n11921_, new_n11922_,
    new_n11923_, new_n11924_, new_n11925_, new_n11926_, new_n11927_,
    new_n11928_, new_n11929_, new_n11930_, new_n11931_, new_n11932_,
    new_n11933_, new_n11934_, new_n11935_, new_n11936_, new_n11937_,
    new_n11938_, new_n11939_, new_n11940_, new_n11941_, new_n11942_,
    new_n11943_, new_n11944_, new_n11945_, new_n11946_, new_n11947_,
    new_n11948_, new_n11949_, new_n11950_, new_n11951_, new_n11952_,
    new_n11953_, new_n11954_, new_n11955_, new_n11956_, new_n11957_,
    new_n11958_, new_n11959_, new_n11960_, new_n11961_, new_n11962_,
    new_n11963_, new_n11964_, new_n11965_, new_n11966_, new_n11967_,
    new_n11968_, new_n11969_, new_n11970_, new_n11971_, new_n11972_,
    new_n11973_, new_n11974_, new_n11975_, new_n11976_, new_n11977_,
    new_n11978_, new_n11979_, new_n11980_, new_n11981_, new_n11982_,
    new_n11983_, new_n11984_, new_n11985_, new_n11986_, new_n11987_,
    new_n11988_, new_n11989_, new_n11990_, new_n11991_, new_n11992_,
    new_n11993_, new_n11994_, new_n11995_, new_n11996_, new_n11997_,
    new_n11998_, new_n11999_, new_n12000_, new_n12001_, new_n12002_,
    new_n12003_, new_n12004_, new_n12005_, new_n12006_, new_n12007_,
    new_n12008_, new_n12009_, new_n12010_, new_n12011_, new_n12012_,
    new_n12013_, new_n12014_, new_n12015_, new_n12016_, new_n12017_,
    new_n12018_, new_n12019_, new_n12020_, new_n12021_, new_n12022_,
    new_n12023_, new_n12024_, new_n12025_, new_n12026_, new_n12027_,
    new_n12028_, new_n12029_, new_n12030_, new_n12031_, new_n12032_,
    new_n12033_, new_n12034_, new_n12035_, new_n12036_, new_n12037_,
    new_n12038_, new_n12039_, new_n12040_, new_n12041_, new_n12042_,
    new_n12043_, new_n12044_, new_n12045_, new_n12046_, new_n12047_,
    new_n12048_, new_n12049_, new_n12050_, new_n12051_, new_n12052_,
    new_n12053_, new_n12054_, new_n12055_, new_n12056_, new_n12057_,
    new_n12058_, new_n12059_, new_n12060_, new_n12061_, new_n12062_,
    new_n12063_, new_n12064_, new_n12065_, new_n12066_, new_n12067_,
    new_n12068_, new_n12069_, new_n12070_, new_n12071_, new_n12072_,
    new_n12073_, new_n12074_, new_n12075_, new_n12076_, new_n12077_,
    new_n12078_, new_n12079_, new_n12080_, new_n12081_, new_n12082_,
    new_n12083_, new_n12084_, new_n12085_, new_n12086_, new_n12087_,
    new_n12088_, new_n12089_, new_n12090_, new_n12091_, new_n12092_,
    new_n12093_, new_n12094_, new_n12095_, new_n12096_, new_n12097_,
    new_n12098_, new_n12099_, new_n12100_, new_n12101_, new_n12102_,
    new_n12103_, new_n12104_, new_n12105_, new_n12106_, new_n12107_,
    new_n12108_, new_n12109_, new_n12110_, new_n12111_, new_n12112_,
    new_n12113_, new_n12114_, new_n12115_, new_n12116_, new_n12117_,
    new_n12118_, new_n12119_, new_n12120_, new_n12121_, new_n12122_,
    new_n12123_, new_n12124_, new_n12125_, new_n12126_, new_n12127_,
    new_n12128_, new_n12129_, new_n12130_, new_n12131_, new_n12132_,
    new_n12133_, new_n12134_, new_n12135_, new_n12136_, new_n12137_,
    new_n12138_, new_n12139_, new_n12140_, new_n12141_, new_n12142_,
    new_n12143_, new_n12144_, new_n12145_, new_n12146_, new_n12147_,
    new_n12148_, new_n12149_, new_n12150_, new_n12151_, new_n12152_,
    new_n12153_, new_n12154_, new_n12155_, new_n12156_, new_n12157_,
    new_n12158_, new_n12159_, new_n12160_, new_n12161_, new_n12162_,
    new_n12163_, new_n12164_, new_n12165_, new_n12166_, new_n12167_,
    new_n12168_, new_n12169_, new_n12170_, new_n12171_, new_n12172_,
    new_n12173_, new_n12174_, new_n12175_, new_n12176_, new_n12177_,
    new_n12178_, new_n12179_, new_n12180_, new_n12181_, new_n12182_,
    new_n12183_, new_n12184_, new_n12185_, new_n12186_, new_n12187_,
    new_n12188_, new_n12189_, new_n12190_, new_n12191_, new_n12192_,
    new_n12193_, new_n12194_, new_n12195_, new_n12196_, new_n12197_,
    new_n12198_, new_n12199_, new_n12200_, new_n12201_, new_n12202_,
    new_n12203_, new_n12204_, new_n12205_, new_n12206_, new_n12207_,
    new_n12208_, new_n12209_, new_n12210_, new_n12211_, new_n12212_,
    new_n12213_, new_n12214_, new_n12215_, new_n12216_, new_n12217_,
    new_n12218_, new_n12219_, new_n12220_, new_n12221_, new_n12222_,
    new_n12223_, new_n12224_, new_n12225_, new_n12226_, new_n12227_,
    new_n12228_, new_n12229_, new_n12230_, new_n12231_, new_n12232_,
    new_n12233_, new_n12234_, new_n12235_, new_n12236_, new_n12237_,
    new_n12238_, new_n12239_, new_n12240_, new_n12241_, new_n12242_,
    new_n12243_, new_n12244_, new_n12245_, new_n12246_, new_n12247_,
    new_n12248_, new_n12249_, new_n12250_, new_n12251_, new_n12252_,
    new_n12253_, new_n12254_, new_n12255_, new_n12256_, new_n12257_,
    new_n12258_, new_n12259_, new_n12260_, new_n12261_, new_n12262_,
    new_n12263_, new_n12264_, new_n12265_, new_n12266_, new_n12267_,
    new_n12268_, new_n12269_, new_n12270_, new_n12271_, new_n12272_,
    new_n12273_, new_n12274_, new_n12275_, new_n12276_, new_n12277_,
    new_n12278_, new_n12279_, new_n12280_, new_n12281_, new_n12282_,
    new_n12283_, new_n12284_, new_n12285_, new_n12286_, new_n12287_,
    new_n12288_, new_n12289_, new_n12290_, new_n12291_, new_n12292_,
    new_n12293_, new_n12294_, new_n12295_, new_n12296_, new_n12297_,
    new_n12298_, new_n12299_, new_n12300_, new_n12301_, new_n12302_,
    new_n12303_, new_n12304_, new_n12305_, new_n12306_, new_n12307_,
    new_n12308_, new_n12309_, new_n12310_, new_n12311_, new_n12312_,
    new_n12313_, new_n12314_, new_n12315_, new_n12316_, new_n12317_,
    new_n12318_, new_n12319_, new_n12320_, new_n12321_, new_n12322_,
    new_n12323_, new_n12324_, new_n12325_, new_n12326_, new_n12327_,
    new_n12328_, new_n12329_, new_n12330_, new_n12331_, new_n12332_,
    new_n12333_, new_n12334_, new_n12335_, new_n12336_, new_n12337_,
    new_n12338_, new_n12339_, new_n12340_, new_n12341_, new_n12342_,
    new_n12343_, new_n12344_, new_n12345_, new_n12346_, new_n12347_,
    new_n12348_, new_n12349_, new_n12350_, new_n12351_, new_n12352_,
    new_n12353_, new_n12354_, new_n12355_, new_n12356_, new_n12357_,
    new_n12358_, new_n12359_, new_n12360_, new_n12361_, new_n12362_,
    new_n12363_, new_n12364_, new_n12365_, new_n12366_, new_n12367_,
    new_n12368_, new_n12369_, new_n12370_, new_n12371_, new_n12372_,
    new_n12373_, new_n12374_, new_n12375_, new_n12376_, new_n12377_,
    new_n12378_, new_n12379_, new_n12380_, new_n12381_, new_n12382_,
    new_n12383_, new_n12384_, new_n12385_, new_n12386_, new_n12387_,
    new_n12388_, new_n12389_, new_n12390_, new_n12391_, new_n12392_,
    new_n12393_, new_n12394_, new_n12395_, new_n12396_, new_n12397_,
    new_n12398_, new_n12399_, new_n12400_, new_n12401_, new_n12402_,
    new_n12403_, new_n12404_, new_n12405_, new_n12406_, new_n12407_,
    new_n12408_, new_n12409_, new_n12410_, new_n12411_, new_n12412_,
    new_n12413_, new_n12414_, new_n12415_, new_n12416_, new_n12417_,
    new_n12418_, new_n12419_, new_n12420_, new_n12421_, new_n12422_,
    new_n12423_, new_n12424_, new_n12425_, new_n12426_, new_n12427_,
    new_n12428_, new_n12429_, new_n12430_, new_n12431_, new_n12432_,
    new_n12433_, new_n12434_, new_n12435_, new_n12436_, new_n12437_,
    new_n12438_, new_n12439_, new_n12440_, new_n12441_, new_n12442_,
    new_n12443_, new_n12444_, new_n12445_, new_n12446_, new_n12447_,
    new_n12448_, new_n12449_, new_n12450_, new_n12451_, new_n12452_,
    new_n12453_, new_n12454_, new_n12455_, new_n12456_, new_n12457_,
    new_n12458_, new_n12459_, new_n12460_, new_n12461_, new_n12462_,
    new_n12463_, new_n12464_, new_n12465_, new_n12466_, new_n12467_,
    new_n12468_, new_n12469_, new_n12470_, new_n12471_, new_n12472_,
    new_n12473_, new_n12474_, new_n12475_, new_n12476_, new_n12477_,
    new_n12478_, new_n12479_, new_n12480_, new_n12481_, new_n12482_,
    new_n12483_, new_n12484_, new_n12485_, new_n12486_, new_n12487_,
    new_n12488_, new_n12489_, new_n12490_, new_n12491_, new_n12492_,
    new_n12493_, new_n12494_, new_n12495_, new_n12496_, new_n12497_,
    new_n12498_, new_n12499_, new_n12500_, new_n12501_, new_n12502_,
    new_n12503_, new_n12504_, new_n12505_, new_n12506_, new_n12507_,
    new_n12508_, new_n12509_, new_n12510_, new_n12511_, new_n12512_,
    new_n12513_, new_n12514_, new_n12515_, new_n12516_, new_n12517_,
    new_n12518_, new_n12519_, new_n12520_, new_n12521_, new_n12522_,
    new_n12523_, new_n12524_, new_n12525_, new_n12526_, new_n12527_,
    new_n12528_, new_n12529_, new_n12530_, new_n12531_, new_n12532_,
    new_n12533_, new_n12534_, new_n12535_, new_n12536_, new_n12537_,
    new_n12538_, new_n12539_, new_n12540_, new_n12541_, new_n12542_,
    new_n12543_, new_n12544_, new_n12545_, new_n12546_, new_n12547_,
    new_n12548_, new_n12549_, new_n12550_, new_n12551_, new_n12552_,
    new_n12553_, new_n12554_, new_n12555_, new_n12556_, new_n12557_,
    new_n12558_, new_n12559_, new_n12560_, new_n12561_, new_n12562_,
    new_n12563_, new_n12564_, new_n12565_, new_n12566_, new_n12567_,
    new_n12568_, new_n12569_, new_n12570_, new_n12571_, new_n12572_,
    new_n12573_, new_n12574_, new_n12575_, new_n12576_, new_n12577_,
    new_n12578_, new_n12579_, new_n12580_, new_n12581_, new_n12582_,
    new_n12583_, new_n12584_, new_n12585_, new_n12586_, new_n12587_,
    new_n12588_, new_n12589_, new_n12590_, new_n12591_, new_n12592_,
    new_n12593_, new_n12594_, new_n12595_, new_n12596_, new_n12597_,
    new_n12598_, new_n12599_, new_n12600_, new_n12601_, new_n12602_,
    new_n12603_, new_n12604_, new_n12605_, new_n12606_, new_n12607_,
    new_n12608_, new_n12609_, new_n12610_, new_n12611_, new_n12612_,
    new_n12613_, new_n12614_, new_n12615_, new_n12616_, new_n12617_,
    new_n12618_, new_n12619_, new_n12620_, new_n12621_, new_n12622_,
    new_n12623_, new_n12624_, new_n12625_, new_n12626_, new_n12627_,
    new_n12628_, new_n12629_, new_n12630_, new_n12631_, new_n12632_,
    new_n12633_, new_n12634_, new_n12635_, new_n12636_, new_n12637_,
    new_n12638_, new_n12639_, new_n12640_, new_n12641_, new_n12642_,
    new_n12643_, new_n12644_, new_n12645_, new_n12646_, new_n12647_,
    new_n12648_, new_n12649_, new_n12650_, new_n12651_, new_n12652_,
    new_n12653_, new_n12654_, new_n12655_, new_n12656_, new_n12657_,
    new_n12658_, new_n12659_, new_n12660_, new_n12661_, new_n12662_,
    new_n12663_, new_n12664_, new_n12665_, new_n12666_, new_n12667_,
    new_n12668_, new_n12669_, new_n12670_, new_n12671_, new_n12672_,
    new_n12673_, new_n12674_, new_n12675_, new_n12676_, new_n12677_,
    new_n12678_, new_n12679_, new_n12680_, new_n12681_, new_n12682_,
    new_n12683_, new_n12684_, new_n12685_, new_n12686_, new_n12687_,
    new_n12688_, new_n12689_, new_n12690_, new_n12691_, new_n12692_,
    new_n12693_, new_n12694_, new_n12695_, new_n12696_, new_n12697_,
    new_n12698_, new_n12699_, new_n12700_, new_n12701_, new_n12702_,
    new_n12703_, new_n12704_, new_n12705_, new_n12706_, new_n12707_,
    new_n12708_, new_n12709_, new_n12710_, new_n12711_, new_n12712_,
    new_n12713_, new_n12714_, new_n12715_, new_n12716_, new_n12717_,
    new_n12718_, new_n12719_, new_n12720_, new_n12721_, new_n12722_,
    new_n12723_, new_n12724_, new_n12725_, new_n12726_, new_n12727_,
    new_n12728_, new_n12729_, new_n12730_, new_n12731_, new_n12732_,
    new_n12733_, new_n12734_, new_n12735_, new_n12736_, new_n12737_,
    new_n12738_, new_n12739_, new_n12740_, new_n12741_, new_n12742_,
    new_n12743_, new_n12744_, new_n12745_, new_n12746_, new_n12747_,
    new_n12748_, new_n12749_, new_n12750_, new_n12751_, new_n12752_,
    new_n12753_, new_n12754_, new_n12755_, new_n12756_, new_n12757_,
    new_n12758_, new_n12759_, new_n12760_, new_n12761_, new_n12762_,
    new_n12763_, new_n12764_, new_n12765_, new_n12766_, new_n12767_,
    new_n12768_, new_n12769_, new_n12770_, new_n12771_, new_n12772_,
    new_n12773_, new_n12774_, new_n12775_, new_n12776_, new_n12777_,
    new_n12778_, new_n12779_, new_n12780_, new_n12781_, new_n12782_,
    new_n12783_, new_n12784_, new_n12785_, new_n12786_, new_n12787_,
    new_n12788_, new_n12789_, new_n12790_, new_n12791_, new_n12792_,
    new_n12793_, new_n12794_, new_n12795_, new_n12796_, new_n12797_,
    new_n12798_, new_n12799_, new_n12800_, new_n12801_, new_n12802_,
    new_n12803_, new_n12804_, new_n12805_, new_n12806_, new_n12807_,
    new_n12808_, new_n12809_, new_n12810_, new_n12811_, new_n12812_,
    new_n12813_, new_n12814_, new_n12815_, new_n12816_, new_n12817_,
    new_n12818_, new_n12819_, new_n12820_, new_n12821_, new_n12822_,
    new_n12823_, new_n12824_, new_n12825_, new_n12826_, new_n12827_,
    new_n12828_, new_n12829_, new_n12830_, new_n12831_, new_n12832_,
    new_n12833_, new_n12834_, new_n12835_, new_n12836_, new_n12837_,
    new_n12838_, new_n12839_, new_n12840_, new_n12841_, new_n12842_,
    new_n12843_, new_n12844_, new_n12845_, new_n12846_, new_n12847_,
    new_n12848_, new_n12849_, new_n12850_, new_n12851_, new_n12852_,
    new_n12853_, new_n12854_, new_n12855_, new_n12856_, new_n12857_,
    new_n12858_, new_n12859_, new_n12860_, new_n12861_, new_n12862_,
    new_n12863_, new_n12864_, new_n12865_, new_n12866_, new_n12867_,
    new_n12868_, new_n12869_, new_n12870_, new_n12871_, new_n12872_,
    new_n12873_, new_n12874_, new_n12875_, new_n12876_, new_n12877_,
    new_n12878_, new_n12879_, new_n12880_, new_n12881_, new_n12882_,
    new_n12883_, new_n12884_, new_n12885_, new_n12886_, new_n12887_,
    new_n12888_, new_n12889_, new_n12890_, new_n12891_, new_n12892_,
    new_n12893_, new_n12894_, new_n12895_, new_n12896_, new_n12897_,
    new_n12898_, new_n12899_, new_n12900_, new_n12901_, new_n12902_,
    new_n12903_, new_n12904_, new_n12905_, new_n12906_, new_n12907_,
    new_n12908_, new_n12909_, new_n12910_, new_n12911_, new_n12912_,
    new_n12913_, new_n12914_, new_n12915_, new_n12916_, new_n12917_,
    new_n12918_, new_n12919_, new_n12920_, new_n12921_, new_n12922_,
    new_n12923_, new_n12924_, new_n12925_, new_n12926_, new_n12927_,
    new_n12928_, new_n12929_, new_n12930_, new_n12931_, new_n12932_,
    new_n12933_, new_n12934_, new_n12935_, new_n12936_, new_n12937_,
    new_n12938_, new_n12939_, new_n12940_, new_n12941_, new_n12942_,
    new_n12943_, new_n12944_, new_n12945_, new_n12946_, new_n12947_,
    new_n12948_, new_n12949_, new_n12950_, new_n12951_, new_n12952_,
    new_n12953_, new_n12954_, new_n12955_, new_n12956_, new_n12957_,
    new_n12958_, new_n12959_, new_n12960_, new_n12961_, new_n12962_,
    new_n12963_, new_n12964_, new_n12965_, new_n12966_, new_n12967_,
    new_n12968_, new_n12969_, new_n12970_, new_n12971_, new_n12972_,
    new_n12973_, new_n12974_, new_n12975_, new_n12976_, new_n12977_,
    new_n12978_, new_n12979_, new_n12980_, new_n12981_, new_n12982_,
    new_n12983_, new_n12984_, new_n12985_, new_n12986_, new_n12987_,
    new_n12988_, new_n12989_, new_n12990_, new_n12991_, new_n12992_,
    new_n12993_, new_n12994_, new_n12995_, new_n12996_, new_n12997_,
    new_n12998_, new_n12999_, new_n13000_, new_n13001_, new_n13002_,
    new_n13003_, new_n13004_, new_n13005_, new_n13006_, new_n13007_,
    new_n13008_, new_n13009_, new_n13010_, new_n13011_, new_n13012_,
    new_n13013_, new_n13014_, new_n13015_, new_n13016_, new_n13017_,
    new_n13018_, new_n13019_, new_n13020_, new_n13021_, new_n13022_,
    new_n13023_, new_n13024_, new_n13025_, new_n13026_, new_n13027_,
    new_n13028_, new_n13029_, new_n13030_, new_n13031_, new_n13032_,
    new_n13033_, new_n13034_, new_n13035_, new_n13036_, new_n13037_,
    new_n13038_, new_n13039_, new_n13040_, new_n13041_, new_n13042_,
    new_n13043_, new_n13044_, new_n13045_, new_n13046_, new_n13047_,
    new_n13048_, new_n13049_, new_n13050_, new_n13051_, new_n13052_,
    new_n13053_, new_n13054_, new_n13055_, new_n13056_, new_n13057_,
    new_n13058_, new_n13059_, new_n13060_, new_n13061_, new_n13062_,
    new_n13063_, new_n13064_, new_n13065_, new_n13066_, new_n13067_,
    new_n13068_, new_n13069_, new_n13070_, new_n13071_, new_n13072_,
    new_n13073_, new_n13074_, new_n13075_, new_n13076_, new_n13077_,
    new_n13078_, new_n13079_, new_n13080_, new_n13081_, new_n13082_,
    new_n13083_, new_n13084_, new_n13085_, new_n13086_, new_n13087_,
    new_n13088_, new_n13089_, new_n13090_, new_n13091_, new_n13092_,
    new_n13093_, new_n13094_, new_n13095_, new_n13096_, new_n13097_,
    new_n13098_, new_n13099_, new_n13100_, new_n13101_, new_n13102_,
    new_n13103_, new_n13104_, new_n13105_, new_n13106_, new_n13107_,
    new_n13108_, new_n13109_, new_n13110_, new_n13111_, new_n13112_,
    new_n13113_, new_n13114_, new_n13115_, new_n13116_, new_n13117_,
    new_n13118_, new_n13119_, new_n13120_, new_n13121_, new_n13122_,
    new_n13123_, new_n13124_, new_n13125_, new_n13126_, new_n13127_,
    new_n13128_, new_n13129_, new_n13130_, new_n13131_, new_n13132_,
    new_n13133_, new_n13134_, new_n13135_, new_n13136_, new_n13137_,
    new_n13138_, new_n13139_, new_n13140_, new_n13141_, new_n13142_,
    new_n13143_, new_n13144_, new_n13145_, new_n13146_, new_n13147_,
    new_n13148_, new_n13149_, new_n13150_, new_n13151_, new_n13152_,
    new_n13153_, new_n13154_, new_n13155_, new_n13156_, new_n13157_,
    new_n13158_, new_n13159_, new_n13160_, new_n13161_, new_n13162_,
    new_n13163_, new_n13164_, new_n13165_, new_n13166_, new_n13167_,
    new_n13168_, new_n13169_, new_n13170_, new_n13171_, new_n13172_,
    new_n13173_, new_n13174_, new_n13175_, new_n13176_, new_n13177_,
    new_n13178_, new_n13179_, new_n13180_, new_n13181_, new_n13182_,
    new_n13183_, new_n13184_, new_n13185_, new_n13186_, new_n13187_,
    new_n13188_, new_n13189_, new_n13190_, new_n13191_, new_n13192_,
    new_n13193_, new_n13194_, new_n13195_, new_n13196_, new_n13197_,
    new_n13198_, new_n13199_, new_n13200_, new_n13201_, new_n13202_,
    new_n13203_, new_n13204_, new_n13205_, new_n13206_, new_n13207_,
    new_n13208_, new_n13209_, new_n13210_, new_n13211_, new_n13212_,
    new_n13213_, new_n13214_, new_n13215_, new_n13216_, new_n13217_,
    new_n13218_, new_n13219_, new_n13220_, new_n13221_, new_n13222_,
    new_n13223_, new_n13224_, new_n13225_, new_n13226_, new_n13227_,
    new_n13228_, new_n13229_, new_n13230_, new_n13231_, new_n13232_,
    new_n13233_, new_n13234_, new_n13235_, new_n13236_, new_n13237_,
    new_n13238_, new_n13239_, new_n13240_, new_n13241_, new_n13242_,
    new_n13243_, new_n13244_, new_n13245_, new_n13246_, new_n13247_,
    new_n13248_, new_n13249_, new_n13250_, new_n13251_, new_n13252_,
    new_n13253_, new_n13254_, new_n13255_, new_n13256_, new_n13257_,
    new_n13258_, new_n13259_, new_n13260_, new_n13261_, new_n13262_,
    new_n13263_, new_n13264_, new_n13265_, new_n13266_, new_n13267_,
    new_n13268_, new_n13269_, new_n13270_, new_n13271_, new_n13272_,
    new_n13273_, new_n13274_, new_n13275_, new_n13276_, new_n13277_,
    new_n13278_, new_n13279_, new_n13280_, new_n13281_, new_n13282_,
    new_n13283_, new_n13284_, new_n13285_, new_n13286_, new_n13287_,
    new_n13288_, new_n13289_, new_n13290_, new_n13291_, new_n13292_,
    new_n13293_, new_n13294_, new_n13295_, new_n13296_, new_n13297_,
    new_n13298_, new_n13299_, new_n13300_, new_n13301_, new_n13302_,
    new_n13303_, new_n13304_, new_n13305_, new_n13306_, new_n13307_,
    new_n13308_, new_n13309_, new_n13310_, new_n13311_, new_n13312_,
    new_n13313_, new_n13314_, new_n13315_, new_n13316_, new_n13317_,
    new_n13318_, new_n13319_, new_n13320_, new_n13321_, new_n13322_,
    new_n13323_, new_n13324_, new_n13325_, new_n13326_, new_n13327_,
    new_n13328_, new_n13329_, new_n13330_, new_n13331_, new_n13332_,
    new_n13333_, new_n13334_, new_n13335_, new_n13336_, new_n13337_,
    new_n13338_, new_n13339_, new_n13340_, new_n13341_, new_n13342_,
    new_n13343_, new_n13344_, new_n13345_, new_n13346_, new_n13347_,
    new_n13348_, new_n13349_, new_n13350_, new_n13351_, new_n13352_,
    new_n13353_, new_n13354_, new_n13355_, new_n13356_, new_n13357_,
    new_n13358_, new_n13359_, new_n13360_, new_n13361_, new_n13362_,
    new_n13363_, new_n13364_, new_n13365_, new_n13366_, new_n13367_,
    new_n13368_, new_n13369_, new_n13370_, new_n13371_, new_n13372_,
    new_n13373_, new_n13374_, new_n13375_, new_n13376_, new_n13377_,
    new_n13378_, new_n13379_, new_n13380_, new_n13381_, new_n13382_,
    new_n13383_, new_n13384_, new_n13385_, new_n13386_, new_n13387_,
    new_n13388_, new_n13389_, new_n13390_, new_n13391_, new_n13392_,
    new_n13393_, new_n13394_, new_n13395_, new_n13396_, new_n13397_,
    new_n13398_, new_n13399_, new_n13400_, new_n13401_, new_n13402_,
    new_n13403_, new_n13404_, new_n13405_, new_n13406_, new_n13407_,
    new_n13408_, new_n13409_, new_n13410_, new_n13411_, new_n13412_,
    new_n13413_, new_n13414_, new_n13415_, new_n13416_, new_n13417_,
    new_n13418_, new_n13419_, new_n13420_, new_n13421_, new_n13422_,
    new_n13423_, new_n13424_, new_n13425_, new_n13426_, new_n13427_,
    new_n13428_, new_n13429_, new_n13430_, new_n13431_, new_n13432_,
    new_n13433_, new_n13434_, new_n13435_, new_n13436_, new_n13437_,
    new_n13438_, new_n13439_, new_n13440_, new_n13441_, new_n13442_,
    new_n13443_, new_n13444_, new_n13445_, new_n13446_, new_n13447_,
    new_n13448_, new_n13449_, new_n13450_, new_n13451_, new_n13452_,
    new_n13453_, new_n13454_, new_n13455_, new_n13456_, new_n13457_,
    new_n13458_, new_n13459_, new_n13460_, new_n13461_, new_n13462_,
    new_n13463_, new_n13464_, new_n13465_, new_n13466_, new_n13467_,
    new_n13468_, new_n13469_, new_n13470_, new_n13471_, new_n13472_,
    new_n13473_, new_n13474_, new_n13475_, new_n13476_, new_n13477_,
    new_n13478_, new_n13479_, new_n13480_, new_n13481_, new_n13482_,
    new_n13483_, new_n13484_, new_n13485_, new_n13486_, new_n13487_,
    new_n13488_, new_n13489_, new_n13490_, new_n13491_, new_n13492_,
    new_n13493_, new_n13494_, new_n13495_, new_n13496_, new_n13497_,
    new_n13498_, new_n13499_, new_n13500_, new_n13501_, new_n13502_,
    new_n13503_, new_n13504_, new_n13505_, new_n13506_, new_n13507_,
    new_n13508_, new_n13509_, new_n13510_, new_n13511_, new_n13512_,
    new_n13513_, new_n13514_, new_n13515_, new_n13516_, new_n13517_,
    new_n13518_, new_n13519_, new_n13520_, new_n13521_, new_n13522_,
    new_n13523_, new_n13524_, new_n13525_, new_n13526_, new_n13527_,
    new_n13528_, new_n13529_, new_n13530_, new_n13531_, new_n13532_,
    new_n13533_, new_n13534_, new_n13535_, new_n13536_, new_n13537_,
    new_n13538_, new_n13539_, new_n13540_, new_n13541_, new_n13542_,
    new_n13543_, new_n13544_, new_n13545_, new_n13546_, new_n13547_,
    new_n13548_, new_n13549_, new_n13550_, new_n13551_, new_n13552_,
    new_n13553_, new_n13554_, new_n13555_, new_n13556_, new_n13557_,
    new_n13558_, new_n13559_, new_n13560_, new_n13561_, new_n13562_,
    new_n13563_, new_n13564_, new_n13565_, new_n13566_, new_n13567_,
    new_n13568_, new_n13569_, new_n13570_, new_n13571_, new_n13572_,
    new_n13573_, new_n13574_, new_n13575_, new_n13576_, new_n13577_,
    new_n13578_, new_n13579_, new_n13580_, new_n13581_, new_n13582_,
    new_n13583_, new_n13584_, new_n13585_, new_n13586_, new_n13587_,
    new_n13588_, new_n13589_, new_n13590_, new_n13591_, new_n13592_,
    new_n13593_, new_n13594_, new_n13595_, new_n13596_, new_n13597_,
    new_n13598_, new_n13599_, new_n13600_, new_n13601_, new_n13602_,
    new_n13603_, new_n13604_, new_n13605_, new_n13606_, new_n13607_,
    new_n13608_, new_n13609_, new_n13610_, new_n13611_, new_n13612_,
    new_n13613_, new_n13614_, new_n13615_, new_n13616_, new_n13617_,
    new_n13618_, new_n13619_, new_n13620_, new_n13621_, new_n13622_,
    new_n13623_, new_n13624_, new_n13625_, new_n13626_, new_n13627_,
    new_n13628_, new_n13629_, new_n13630_, new_n13631_, new_n13632_,
    new_n13633_, new_n13634_, new_n13635_, new_n13636_, new_n13637_,
    new_n13638_, new_n13639_, new_n13640_, new_n13641_, new_n13642_,
    new_n13643_, new_n13644_, new_n13645_, new_n13646_, new_n13647_,
    new_n13648_, new_n13649_, new_n13650_, new_n13651_, new_n13652_,
    new_n13653_, new_n13654_, new_n13655_, new_n13656_, new_n13657_,
    new_n13658_, new_n13659_, new_n13660_, new_n13661_, new_n13662_,
    new_n13663_, new_n13664_, new_n13665_, new_n13666_, new_n13667_,
    new_n13668_, new_n13669_, new_n13670_, new_n13671_, new_n13672_,
    new_n13673_, new_n13674_, new_n13675_, new_n13676_, new_n13677_,
    new_n13678_, new_n13679_, new_n13680_, new_n13681_, new_n13682_,
    new_n13683_, new_n13684_, new_n13685_, new_n13686_, new_n13687_,
    new_n13688_, new_n13689_, new_n13690_, new_n13691_, new_n13692_,
    new_n13693_, new_n13694_, new_n13695_, new_n13696_, new_n13697_,
    new_n13698_, new_n13699_, new_n13700_, new_n13701_, new_n13702_,
    new_n13703_, new_n13704_, new_n13705_, new_n13706_, new_n13707_,
    new_n13708_, new_n13709_, new_n13710_, new_n13711_, new_n13712_,
    new_n13713_, new_n13714_, new_n13715_, new_n13716_, new_n13717_,
    new_n13718_, new_n13719_, new_n13720_, new_n13721_, new_n13722_,
    new_n13723_, new_n13724_, new_n13725_, new_n13726_, new_n13727_,
    new_n13728_, new_n13729_, new_n13730_, new_n13731_, new_n13732_,
    new_n13733_, new_n13734_, new_n13735_, new_n13736_, new_n13737_,
    new_n13738_, new_n13739_, new_n13740_, new_n13741_, new_n13742_,
    new_n13743_, new_n13744_, new_n13745_, new_n13746_, new_n13747_,
    new_n13748_, new_n13749_, new_n13750_, new_n13751_, new_n13752_,
    new_n13753_, new_n13754_, new_n13755_, new_n13756_, new_n13757_,
    new_n13758_, new_n13759_, new_n13760_, new_n13761_, new_n13762_,
    new_n13763_, new_n13764_, new_n13765_, new_n13766_, new_n13767_,
    new_n13768_, new_n13769_, new_n13770_, new_n13771_, new_n13772_,
    new_n13773_, new_n13774_, new_n13775_, new_n13776_, new_n13777_,
    new_n13778_, new_n13779_, new_n13780_, new_n13781_, new_n13782_,
    new_n13783_, new_n13784_, new_n13785_, new_n13786_, new_n13787_,
    new_n13788_, new_n13789_, new_n13790_, new_n13791_, new_n13792_,
    new_n13793_, new_n13794_, new_n13795_, new_n13796_, new_n13797_,
    new_n13798_, new_n13799_, new_n13800_, new_n13801_, new_n13802_,
    new_n13803_, new_n13804_, new_n13805_, new_n13806_, new_n13807_,
    new_n13808_, new_n13809_, new_n13810_, new_n13811_, new_n13812_,
    new_n13813_, new_n13814_, new_n13815_, new_n13816_, new_n13817_,
    new_n13818_, new_n13819_, new_n13820_, new_n13821_, new_n13822_,
    new_n13823_, new_n13824_, new_n13825_, new_n13826_, new_n13827_,
    new_n13828_, new_n13829_, new_n13830_, new_n13831_, new_n13832_,
    new_n13833_, new_n13834_, new_n13835_, new_n13836_, new_n13837_,
    new_n13838_, new_n13839_, new_n13840_, new_n13841_, new_n13842_,
    new_n13843_, new_n13844_, new_n13845_, new_n13846_, new_n13847_,
    new_n13848_, new_n13849_, new_n13850_, new_n13851_, new_n13852_,
    new_n13853_, new_n13854_, new_n13855_, new_n13856_, new_n13857_,
    new_n13858_, new_n13859_, new_n13860_, new_n13861_, new_n13862_,
    new_n13863_, new_n13864_, new_n13865_, new_n13866_, new_n13867_,
    new_n13868_, new_n13869_, new_n13870_, new_n13871_, new_n13872_,
    new_n13873_, new_n13874_, new_n13875_, new_n13876_, new_n13877_,
    new_n13878_, new_n13879_, new_n13880_, new_n13881_, new_n13882_,
    new_n13883_, new_n13884_, new_n13885_, new_n13886_, new_n13887_,
    new_n13888_, new_n13889_, new_n13890_, new_n13891_, new_n13892_,
    new_n13893_, new_n13894_, new_n13895_, new_n13896_, new_n13897_,
    new_n13898_, new_n13899_, new_n13900_, new_n13901_, new_n13902_,
    new_n13903_, new_n13904_, new_n13905_, new_n13906_, new_n13907_,
    new_n13908_, new_n13909_, new_n13910_, new_n13911_, new_n13912_,
    new_n13913_, new_n13914_, new_n13915_, new_n13916_, new_n13917_,
    new_n13918_, new_n13919_, new_n13920_, new_n13921_, new_n13922_,
    new_n13923_, new_n13924_, new_n13925_, new_n13926_, new_n13927_,
    new_n13928_, new_n13929_, new_n13930_, new_n13931_, new_n13932_,
    new_n13933_, new_n13934_, new_n13935_, new_n13936_, new_n13937_,
    new_n13938_, new_n13939_, new_n13940_, new_n13941_, new_n13942_,
    new_n13943_, new_n13944_, new_n13945_, new_n13946_, new_n13947_,
    new_n13948_, new_n13949_, new_n13950_, new_n13951_, new_n13952_,
    new_n13953_, new_n13954_, new_n13955_, new_n13956_, new_n13957_,
    new_n13958_, new_n13959_, new_n13960_, new_n13961_, new_n13962_,
    new_n13963_, new_n13964_, new_n13965_, new_n13966_, new_n13967_,
    new_n13968_, new_n13969_, new_n13970_, new_n13971_, new_n13972_,
    new_n13973_, new_n13974_, new_n13975_, new_n13976_, new_n13977_,
    new_n13978_, new_n13979_, new_n13980_, new_n13981_, new_n13982_,
    new_n13983_, new_n13984_, new_n13985_, new_n13986_, new_n13987_,
    new_n13988_, new_n13989_, new_n13990_, new_n13991_, new_n13992_,
    new_n13993_, new_n13994_, new_n13995_, new_n13996_, new_n13997_,
    new_n13998_, new_n13999_, new_n14000_, new_n14001_, new_n14002_,
    new_n14003_, new_n14004_, new_n14005_, new_n14006_, new_n14007_,
    new_n14008_, new_n14009_, new_n14010_, new_n14011_, new_n14012_,
    new_n14013_, new_n14014_, new_n14015_, new_n14016_, new_n14017_,
    new_n14018_, new_n14019_, new_n14020_, new_n14021_, new_n14022_,
    new_n14023_, new_n14024_, new_n14025_, new_n14026_, new_n14027_,
    new_n14028_, new_n14029_, new_n14030_, new_n14031_, new_n14032_,
    new_n14033_, new_n14034_, new_n14035_, new_n14036_, new_n14037_,
    new_n14038_, new_n14039_, new_n14040_, new_n14041_, new_n14042_,
    new_n14043_, new_n14044_, new_n14045_, new_n14046_, new_n14047_,
    new_n14048_, new_n14049_, new_n14050_, new_n14051_, new_n14052_,
    new_n14053_, new_n14054_, new_n14055_, new_n14056_, new_n14057_,
    new_n14058_, new_n14059_, new_n14060_, new_n14061_, new_n14062_,
    new_n14063_, new_n14064_, new_n14065_, new_n14066_, new_n14067_,
    new_n14068_, new_n14069_, new_n14070_, new_n14071_, new_n14072_,
    new_n14073_, new_n14074_, new_n14075_, new_n14076_, new_n14077_,
    new_n14078_, new_n14079_, new_n14080_, new_n14081_, new_n14082_,
    new_n14083_, new_n14084_, new_n14085_, new_n14086_, new_n14087_,
    new_n14088_, new_n14089_, new_n14090_, new_n14091_, new_n14092_,
    new_n14093_, new_n14094_, new_n14095_, new_n14096_, new_n14097_,
    new_n14098_, new_n14099_, new_n14100_, new_n14101_, new_n14102_,
    new_n14103_, new_n14104_, new_n14105_, new_n14106_, new_n14107_,
    new_n14108_, new_n14109_, new_n14110_, new_n14111_, new_n14112_,
    new_n14113_, new_n14114_, new_n14115_, new_n14116_, new_n14117_,
    new_n14118_, new_n14119_, new_n14120_, new_n14121_, new_n14122_,
    new_n14123_, new_n14124_, new_n14125_, new_n14126_, new_n14127_,
    new_n14128_, new_n14129_, new_n14130_, new_n14131_, new_n14132_,
    new_n14133_, new_n14134_, new_n14135_, new_n14136_, new_n14137_,
    new_n14138_, new_n14139_, new_n14140_, new_n14141_, new_n14142_,
    new_n14143_, new_n14144_, new_n14145_, new_n14146_, new_n14147_,
    new_n14148_, new_n14149_, new_n14150_, new_n14151_, new_n14152_,
    new_n14153_, new_n14154_, new_n14155_, new_n14156_, new_n14157_,
    new_n14158_, new_n14159_, new_n14160_, new_n14161_, new_n14162_,
    new_n14163_, new_n14164_, new_n14165_, new_n14166_, new_n14167_,
    new_n14168_, new_n14169_, new_n14170_, new_n14171_, new_n14172_,
    new_n14173_, new_n14174_, new_n14175_, new_n14176_, new_n14177_,
    new_n14178_, new_n14179_, new_n14180_, new_n14181_, new_n14182_,
    new_n14183_, new_n14184_, new_n14185_, new_n14186_, new_n14187_,
    new_n14188_, new_n14189_, new_n14190_, new_n14191_, new_n14192_,
    new_n14193_, new_n14194_, new_n14195_, new_n14196_, new_n14197_,
    new_n14198_, new_n14199_, new_n14200_, new_n14201_, new_n14202_,
    new_n14203_, new_n14204_, new_n14205_, new_n14206_, new_n14207_,
    new_n14208_, new_n14209_, new_n14210_, new_n14211_, new_n14212_,
    new_n14213_, new_n14214_, new_n14215_, new_n14216_, new_n14217_,
    new_n14218_, new_n14219_, new_n14220_, new_n14221_, new_n14222_,
    new_n14223_, new_n14224_, new_n14225_, new_n14226_, new_n14227_,
    new_n14228_, new_n14229_, new_n14230_, new_n14231_, new_n14232_,
    new_n14233_, new_n14234_, new_n14235_, new_n14236_, new_n14237_,
    new_n14238_, new_n14239_, new_n14240_, new_n14241_, new_n14242_,
    new_n14243_, new_n14244_, new_n14245_, new_n14246_, new_n14247_,
    new_n14248_, new_n14249_, new_n14250_, new_n14251_, new_n14252_,
    new_n14253_, new_n14254_, new_n14255_, new_n14256_, new_n14257_,
    new_n14258_, new_n14259_, new_n14260_, new_n14261_, new_n14262_,
    new_n14263_, new_n14264_, new_n14265_, new_n14266_, new_n14267_,
    new_n14268_, new_n14269_, new_n14270_, new_n14271_, new_n14272_,
    new_n14273_, new_n14274_, new_n14275_, new_n14276_, new_n14277_,
    new_n14278_, new_n14279_, new_n14280_, new_n14281_, new_n14282_,
    new_n14283_, new_n14284_, new_n14285_, new_n14286_, new_n14287_,
    new_n14288_, new_n14289_, new_n14290_, new_n14291_, new_n14292_,
    new_n14293_, new_n14294_, new_n14295_, new_n14296_, new_n14297_,
    new_n14298_, new_n14299_, new_n14300_, new_n14301_, new_n14302_,
    new_n14303_, new_n14304_, new_n14305_, new_n14306_, new_n14307_,
    new_n14308_, new_n14309_, new_n14310_, new_n14311_, new_n14312_,
    new_n14313_, new_n14314_, new_n14315_, new_n14316_, new_n14317_,
    new_n14318_, new_n14319_, new_n14320_, new_n14321_, new_n14322_,
    new_n14323_, new_n14324_, new_n14325_, new_n14326_, new_n14327_,
    new_n14328_, new_n14329_, new_n14330_, new_n14331_, new_n14332_,
    new_n14333_, new_n14334_, new_n14335_, new_n14336_, new_n14337_,
    new_n14338_, new_n14339_, new_n14340_, new_n14341_, new_n14342_,
    new_n14343_, new_n14344_, new_n14345_, new_n14346_, new_n14347_,
    new_n14348_, new_n14349_, new_n14350_, new_n14351_, new_n14352_,
    new_n14353_, new_n14354_, new_n14355_, new_n14356_, new_n14357_,
    new_n14358_, new_n14359_, new_n14360_, new_n14361_, new_n14362_,
    new_n14363_, new_n14364_, new_n14365_, new_n14366_, new_n14367_,
    new_n14368_, new_n14369_, new_n14370_, new_n14371_, new_n14372_,
    new_n14373_, new_n14374_, new_n14375_, new_n14376_, new_n14377_,
    new_n14378_, new_n14379_, new_n14380_, new_n14381_, new_n14382_,
    new_n14383_, new_n14384_, new_n14385_, new_n14386_, new_n14387_,
    new_n14388_, new_n14389_, new_n14390_, new_n14391_, new_n14392_,
    new_n14393_, new_n14394_, new_n14395_, new_n14396_, new_n14397_,
    new_n14398_, new_n14399_, new_n14400_, new_n14401_, new_n14402_,
    new_n14403_, new_n14404_, new_n14405_, new_n14406_, new_n14407_,
    new_n14408_, new_n14409_, new_n14410_, new_n14411_, new_n14412_,
    new_n14413_, new_n14414_, new_n14415_, new_n14416_, new_n14417_,
    new_n14418_, new_n14419_, new_n14420_, new_n14421_, new_n14422_,
    new_n14423_, new_n14424_, new_n14425_, new_n14426_, new_n14427_,
    new_n14428_, new_n14429_, new_n14430_, new_n14431_, new_n14432_,
    new_n14433_, new_n14434_, new_n14435_, new_n14436_, new_n14437_,
    new_n14438_, new_n14439_, new_n14440_, new_n14441_, new_n14442_,
    new_n14443_, new_n14444_, new_n14445_, new_n14446_, new_n14447_,
    new_n14448_, new_n14449_, new_n14450_, new_n14451_, new_n14452_,
    new_n14453_, new_n14454_, new_n14455_, new_n14456_, new_n14457_,
    new_n14458_, new_n14459_, new_n14460_, new_n14461_, new_n14462_,
    new_n14463_, new_n14464_, new_n14465_, new_n14466_, new_n14467_,
    new_n14468_, new_n14469_, new_n14470_, new_n14471_, new_n14472_,
    new_n14473_, new_n14474_, new_n14475_, new_n14476_, new_n14477_,
    new_n14478_, new_n14479_, new_n14480_, new_n14481_, new_n14482_,
    new_n14483_, new_n14484_, new_n14485_, new_n14486_, new_n14487_,
    new_n14488_, new_n14489_, new_n14490_, new_n14491_, new_n14492_,
    new_n14493_, new_n14494_, new_n14495_, new_n14496_, new_n14497_,
    new_n14498_, new_n14499_, new_n14500_, new_n14501_, new_n14502_,
    new_n14503_, new_n14504_, new_n14505_, new_n14506_, new_n14507_,
    new_n14508_, new_n14509_, new_n14510_, new_n14511_, new_n14512_,
    new_n14513_, new_n14514_, new_n14515_, new_n14516_, new_n14517_,
    new_n14518_, new_n14519_, new_n14520_, new_n14521_, new_n14522_,
    new_n14523_, new_n14524_, new_n14525_, new_n14526_, new_n14527_,
    new_n14528_, new_n14529_, new_n14530_, new_n14531_, new_n14532_,
    new_n14533_, new_n14534_, new_n14535_, new_n14536_, new_n14537_,
    new_n14538_, new_n14539_, new_n14540_, new_n14541_, new_n14542_,
    new_n14543_, new_n14544_, new_n14545_, new_n14546_, new_n14547_,
    new_n14548_, new_n14549_, new_n14550_, new_n14551_, new_n14552_,
    new_n14553_, new_n14554_, new_n14555_, new_n14556_, new_n14557_,
    new_n14558_, new_n14559_, new_n14560_, new_n14561_, new_n14562_,
    new_n14563_, new_n14564_, new_n14565_, new_n14566_, new_n14567_,
    new_n14568_, new_n14569_, new_n14570_, new_n14571_, new_n14572_,
    new_n14573_, new_n14574_, new_n14575_, new_n14576_, new_n14577_,
    new_n14578_, new_n14579_, new_n14580_, new_n14581_, new_n14582_,
    new_n14583_, new_n14584_, new_n14585_, new_n14586_, new_n14587_,
    new_n14588_, new_n14589_, new_n14590_, new_n14591_, new_n14592_,
    new_n14593_, new_n14594_, new_n14595_, new_n14596_, new_n14597_,
    new_n14598_, new_n14599_, new_n14600_, new_n14601_, new_n14602_,
    new_n14603_, new_n14604_, new_n14605_, new_n14606_, new_n14607_,
    new_n14608_, new_n14609_, new_n14610_, new_n14611_, new_n14612_,
    new_n14613_, new_n14614_, new_n14615_, new_n14616_, new_n14617_,
    new_n14618_, new_n14619_, new_n14620_, new_n14621_, new_n14622_,
    new_n14623_, new_n14624_, new_n14625_, new_n14626_, new_n14627_,
    new_n14628_, new_n14629_, new_n14630_, new_n14631_, new_n14632_,
    new_n14633_, new_n14634_, new_n14635_, new_n14636_, new_n14637_,
    new_n14638_, new_n14639_, new_n14640_, new_n14641_, new_n14642_,
    new_n14643_, new_n14644_, new_n14645_, new_n14646_, new_n14647_,
    new_n14648_, new_n14649_, new_n14650_, new_n14651_, new_n14652_,
    new_n14653_, new_n14654_, new_n14655_, new_n14656_, new_n14657_,
    new_n14658_, new_n14659_, new_n14660_, new_n14661_, new_n14662_,
    new_n14663_, new_n14664_, new_n14665_, new_n14666_, new_n14667_,
    new_n14668_, new_n14669_, new_n14670_, new_n14671_, new_n14672_,
    new_n14673_, new_n14674_, new_n14675_, new_n14676_, new_n14677_,
    new_n14678_, new_n14679_, new_n14680_, new_n14681_, new_n14682_,
    new_n14683_, new_n14684_, new_n14685_, new_n14686_, new_n14687_,
    new_n14688_, new_n14689_, new_n14690_, new_n14691_, new_n14692_,
    new_n14693_, new_n14694_, new_n14695_, new_n14696_, new_n14697_,
    new_n14698_, new_n14699_, new_n14700_, new_n14701_, new_n14702_,
    new_n14703_, new_n14704_, new_n14705_, new_n14706_, new_n14707_,
    new_n14708_, new_n14709_, new_n14710_, new_n14711_, new_n14712_,
    new_n14713_, new_n14714_, new_n14715_, new_n14716_, new_n14717_,
    new_n14718_, new_n14719_, new_n14720_, new_n14721_, new_n14722_,
    new_n14723_, new_n14724_, new_n14725_, new_n14726_, new_n14727_,
    new_n14728_, new_n14729_, new_n14730_, new_n14731_, new_n14732_,
    new_n14733_, new_n14734_, new_n14735_, new_n14736_, new_n14737_,
    new_n14738_, new_n14739_, new_n14740_, new_n14741_, new_n14742_,
    new_n14743_, new_n14744_, new_n14745_, new_n14746_, new_n14747_,
    new_n14748_, new_n14749_, new_n14750_, new_n14751_, new_n14752_,
    new_n14753_, new_n14754_, new_n14755_, new_n14756_, new_n14757_,
    new_n14758_, new_n14759_, new_n14760_, new_n14761_, new_n14762_,
    new_n14763_, new_n14764_, new_n14765_, new_n14766_, new_n14767_,
    new_n14768_, new_n14769_, new_n14770_, new_n14771_, new_n14772_,
    new_n14773_, new_n14774_, new_n14775_, new_n14776_, new_n14777_,
    new_n14778_, new_n14779_, new_n14780_, new_n14781_, new_n14782_,
    new_n14783_, new_n14784_, new_n14785_, new_n14786_, new_n14787_,
    new_n14788_, new_n14789_, new_n14790_, new_n14791_, new_n14792_,
    new_n14793_, new_n14794_, new_n14795_, new_n14796_, new_n14797_,
    new_n14798_, new_n14799_, new_n14800_, new_n14801_, new_n14802_,
    new_n14803_, new_n14804_, new_n14805_, new_n14806_, new_n14807_,
    new_n14808_, new_n14809_, new_n14810_, new_n14811_, new_n14812_,
    new_n14813_, new_n14814_, new_n14815_, new_n14816_, new_n14817_,
    new_n14818_, new_n14819_, new_n14820_, new_n14821_, new_n14822_,
    new_n14823_, new_n14824_, new_n14825_, new_n14826_, new_n14827_,
    new_n14828_, new_n14829_, new_n14830_, new_n14831_, new_n14832_,
    new_n14833_, new_n14834_, new_n14835_, new_n14836_, new_n14837_,
    new_n14838_, new_n14839_, new_n14840_, new_n14841_, new_n14842_,
    new_n14843_, new_n14844_, new_n14845_, new_n14846_, new_n14847_,
    new_n14848_, new_n14849_, new_n14850_, new_n14851_, new_n14852_,
    new_n14853_, new_n14854_, new_n14855_, new_n14856_, new_n14857_,
    new_n14858_, new_n14859_, new_n14860_, new_n14861_, new_n14862_,
    new_n14863_, new_n14864_, new_n14865_, new_n14866_, new_n14867_,
    new_n14868_, new_n14869_, new_n14870_, new_n14871_, new_n14872_,
    new_n14873_, new_n14874_, new_n14875_, new_n14876_, new_n14877_,
    new_n14878_, new_n14879_, new_n14880_, new_n14881_, new_n14882_,
    new_n14883_, new_n14884_, new_n14885_, new_n14886_, new_n14887_,
    new_n14888_, new_n14889_, new_n14890_, new_n14891_, new_n14892_,
    new_n14893_, new_n14894_, new_n14895_, new_n14896_, new_n14897_,
    new_n14898_, new_n14899_, new_n14900_, new_n14901_, new_n14902_,
    new_n14903_, new_n14904_, new_n14905_, new_n14906_, new_n14907_,
    new_n14908_, new_n14909_, new_n14910_, new_n14911_, new_n14912_,
    new_n14913_, new_n14914_, new_n14915_, new_n14916_, new_n14917_,
    new_n14918_, new_n14919_, new_n14920_, new_n14921_, new_n14922_,
    new_n14923_, new_n14924_, new_n14925_, new_n14926_, new_n14927_,
    new_n14928_, new_n14929_, new_n14930_, new_n14931_, new_n14932_,
    new_n14933_, new_n14934_, new_n14935_, new_n14936_, new_n14937_,
    new_n14938_, new_n14939_, new_n14940_, new_n14941_, new_n14942_,
    new_n14943_, new_n14944_, new_n14945_, new_n14946_, new_n14947_,
    new_n14948_, new_n14949_, new_n14950_, new_n14951_, new_n14952_,
    new_n14953_, new_n14954_, new_n14955_, new_n14956_, new_n14957_,
    new_n14958_, new_n14959_, new_n14960_, new_n14961_, new_n14962_,
    new_n14963_, new_n14964_, new_n14965_, new_n14966_, new_n14967_,
    new_n14968_, new_n14969_, new_n14970_, new_n14971_, new_n14972_,
    new_n14973_, new_n14974_, new_n14975_, new_n14976_, new_n14977_,
    new_n14978_, new_n14979_, new_n14980_, new_n14981_, new_n14982_,
    new_n14983_, new_n14984_, new_n14985_, new_n14986_, new_n14987_,
    new_n14988_, new_n14989_, new_n14990_, new_n14991_, new_n14992_,
    new_n14993_, new_n14994_, new_n14995_, new_n14996_, new_n14997_,
    new_n14998_, new_n14999_, new_n15000_, new_n15001_, new_n15002_,
    new_n15003_, new_n15004_, new_n15005_, new_n15006_, new_n15007_,
    new_n15008_, new_n15009_, new_n15010_, new_n15011_, new_n15012_,
    new_n15013_, new_n15014_, new_n15015_, new_n15016_, new_n15017_,
    new_n15018_, new_n15019_, new_n15020_, new_n15021_, new_n15022_,
    new_n15023_, new_n15024_, new_n15025_, new_n15026_, new_n15027_,
    new_n15028_, new_n15029_, new_n15030_, new_n15031_, new_n15032_,
    new_n15033_, new_n15034_, new_n15035_, new_n15036_, new_n15037_,
    new_n15038_, new_n15039_, new_n15040_, new_n15041_, new_n15042_,
    new_n15043_, new_n15044_, new_n15045_, new_n15046_, new_n15047_,
    new_n15048_, new_n15049_, new_n15050_, new_n15051_, new_n15052_,
    new_n15053_, new_n15054_, new_n15055_, new_n15056_, new_n15057_,
    new_n15058_, new_n15059_, new_n15060_, new_n15061_, new_n15062_,
    new_n15063_, new_n15064_, new_n15065_, new_n15066_, new_n15067_,
    new_n15068_, new_n15069_, new_n15070_, new_n15071_, new_n15072_,
    new_n15073_, new_n15074_, new_n15075_, new_n15076_, new_n15077_,
    new_n15078_, new_n15079_, new_n15080_, new_n15081_, new_n15082_,
    new_n15083_, new_n15084_, new_n15085_, new_n15086_, new_n15087_,
    new_n15088_, new_n15089_, new_n15090_, new_n15091_, new_n15092_,
    new_n15093_, new_n15094_, new_n15095_, new_n15096_, new_n15097_,
    new_n15098_, new_n15099_, new_n15100_, new_n15101_, new_n15102_,
    new_n15103_, new_n15104_, new_n15105_, new_n15106_, new_n15107_,
    new_n15108_, new_n15109_, new_n15110_, new_n15111_, new_n15112_,
    new_n15113_, new_n15114_, new_n15115_, new_n15116_, new_n15117_,
    new_n15118_, new_n15119_, new_n15120_, new_n15121_, new_n15122_,
    new_n15123_, new_n15124_, new_n15125_, new_n15126_, new_n15127_,
    new_n15128_, new_n15129_, new_n15130_, new_n15131_, new_n15132_,
    new_n15133_, new_n15134_, new_n15135_, new_n15136_, new_n15137_,
    new_n15138_, new_n15139_, new_n15140_, new_n15141_, new_n15142_,
    new_n15143_, new_n15144_, new_n15145_, new_n15146_, new_n15147_,
    new_n15148_, new_n15149_, new_n15150_, new_n15151_, new_n15152_,
    new_n15153_, new_n15154_, new_n15155_, new_n15156_, new_n15157_,
    new_n15158_, new_n15159_, new_n15160_, new_n15161_, new_n15162_,
    new_n15163_, new_n15164_, new_n15165_, new_n15166_, new_n15167_,
    new_n15168_, new_n15169_, new_n15170_, new_n15171_, new_n15172_,
    new_n15173_, new_n15174_, new_n15175_, new_n15176_, new_n15177_,
    new_n15178_, new_n15179_, new_n15180_, new_n15181_, new_n15182_,
    new_n15183_, new_n15184_, new_n15185_, new_n15186_, new_n15187_,
    new_n15188_, new_n15189_, new_n15190_, new_n15191_, new_n15192_,
    new_n15193_, new_n15194_, new_n15195_, new_n15196_, new_n15197_,
    new_n15198_, new_n15199_, new_n15200_, new_n15201_, new_n15202_,
    new_n15203_, new_n15204_, new_n15205_, new_n15206_, new_n15207_,
    new_n15208_, new_n15209_, new_n15210_, new_n15211_, new_n15212_,
    new_n15213_, new_n15214_, new_n15215_, new_n15216_, new_n15217_,
    new_n15218_, new_n15219_, new_n15220_, new_n15221_, new_n15222_,
    new_n15223_, new_n15224_, new_n15225_, new_n15226_, new_n15227_,
    new_n15228_, new_n15229_, new_n15230_, new_n15231_, new_n15232_,
    new_n15233_, new_n15234_, new_n15235_, new_n15236_, new_n15237_,
    new_n15238_, new_n15239_, new_n15240_, new_n15241_, new_n15242_,
    new_n15243_, new_n15244_, new_n15245_, new_n15246_, new_n15247_,
    new_n15248_, new_n15249_, new_n15250_, new_n15251_, new_n15252_,
    new_n15253_, new_n15254_, new_n15255_, new_n15256_, new_n15257_,
    new_n15258_, new_n15259_, new_n15260_, new_n15261_, new_n15262_,
    new_n15263_, new_n15264_, new_n15265_, new_n15266_, new_n15267_,
    new_n15268_, new_n15269_, new_n15270_, new_n15271_, new_n15272_,
    new_n15273_, new_n15274_, new_n15275_, new_n15276_, new_n15277_,
    new_n15278_, new_n15279_, new_n15280_, new_n15281_, new_n15282_,
    new_n15283_, new_n15284_, new_n15285_, new_n15286_, new_n15287_,
    new_n15288_, new_n15289_, new_n15290_, new_n15291_, new_n15292_,
    new_n15293_, new_n15294_, new_n15295_, new_n15296_, new_n15297_,
    new_n15298_, new_n15299_, new_n15300_, new_n15301_, new_n15302_,
    new_n15303_, new_n15304_, new_n15305_, new_n15306_, new_n15307_,
    new_n15308_, new_n15309_, new_n15310_, new_n15311_, new_n15312_,
    new_n15313_, new_n15314_, new_n15315_, new_n15316_, new_n15317_,
    new_n15318_, new_n15319_, new_n15320_, new_n15321_, new_n15322_,
    new_n15323_, new_n15324_, new_n15325_, new_n15326_, new_n15327_,
    new_n15328_, new_n15329_, new_n15330_, new_n15331_, new_n15332_,
    new_n15333_, new_n15334_, new_n15335_, new_n15336_, new_n15337_,
    new_n15338_, new_n15339_, new_n15340_, new_n15341_, new_n15342_,
    new_n15343_, new_n15344_, new_n15345_, new_n15346_, new_n15347_,
    new_n15348_, new_n15349_, new_n15350_, new_n15351_, new_n15352_,
    new_n15353_, new_n15354_, new_n15355_, new_n15356_, new_n15357_,
    new_n15358_, new_n15359_, new_n15360_, new_n15361_, new_n15362_,
    new_n15363_, new_n15364_, new_n15365_, new_n15366_, new_n15367_,
    new_n15368_, new_n15369_, new_n15370_, new_n15371_, new_n15372_,
    new_n15373_, new_n15374_, new_n15375_, new_n15376_, new_n15377_,
    new_n15378_, new_n15379_, new_n15380_, new_n15381_, new_n15382_,
    new_n15383_, new_n15384_, new_n15385_, new_n15386_, new_n15387_,
    new_n15388_, new_n15389_, new_n15390_, new_n15391_, new_n15392_,
    new_n15393_, new_n15394_, new_n15395_, new_n15396_, new_n15397_,
    new_n15398_, new_n15399_, new_n15400_, new_n15401_, new_n15402_,
    new_n15403_, new_n15404_, new_n15405_, new_n15406_, new_n15407_,
    new_n15408_, new_n15409_, new_n15410_, new_n15411_, new_n15412_,
    new_n15413_, new_n15414_, new_n15415_, new_n15416_, new_n15417_,
    new_n15418_, new_n15419_, new_n15420_, new_n15421_, new_n15422_,
    new_n15423_, new_n15424_, new_n15425_, new_n15426_, new_n15427_,
    new_n15428_, new_n15429_, new_n15430_, new_n15431_, new_n15432_,
    new_n15433_, new_n15434_, new_n15435_, new_n15436_, new_n15437_,
    new_n15438_, new_n15439_, new_n15440_, new_n15441_, new_n15442_,
    new_n15443_, new_n15444_, new_n15445_, new_n15446_, new_n15447_,
    new_n15448_, new_n15449_, new_n15450_, new_n15451_, new_n15452_,
    new_n15453_, new_n15454_, new_n15455_, new_n15456_, new_n15457_,
    new_n15458_, new_n15459_, new_n15460_, new_n15461_, new_n15462_,
    new_n15463_, new_n15464_, new_n15465_, new_n15466_, new_n15467_,
    new_n15468_, new_n15469_, new_n15470_, new_n15471_, new_n15472_,
    new_n15473_, new_n15474_, new_n15475_, new_n15476_, new_n15477_,
    new_n15478_, new_n15479_, new_n15480_, new_n15481_, new_n15482_,
    new_n15483_, new_n15484_, new_n15485_, new_n15486_, new_n15487_,
    new_n15488_, new_n15489_, new_n15490_, new_n15491_, new_n15492_,
    new_n15493_, new_n15494_, new_n15495_, new_n15496_, new_n15497_,
    new_n15498_, new_n15499_, new_n15500_, new_n15501_, new_n15502_,
    new_n15503_, new_n15504_, new_n15505_, new_n15506_, new_n15507_,
    new_n15508_, new_n15509_, new_n15510_, new_n15511_, new_n15512_,
    new_n15513_, new_n15514_, new_n15515_, new_n15516_, new_n15517_,
    new_n15518_, new_n15519_, new_n15520_, new_n15521_, new_n15522_,
    new_n15523_, new_n15524_, new_n15525_, new_n15526_, new_n15527_,
    new_n15528_, new_n15529_, new_n15530_, new_n15531_, new_n15532_,
    new_n15533_, new_n15534_, new_n15535_, new_n15536_, new_n15537_,
    new_n15538_, new_n15539_, new_n15540_, new_n15541_, new_n15542_,
    new_n15543_, new_n15544_, new_n15545_, new_n15546_, new_n15547_,
    new_n15548_, new_n15549_, new_n15550_, new_n15551_, new_n15552_,
    new_n15553_, new_n15554_, new_n15555_, new_n15556_, new_n15557_,
    new_n15558_, new_n15559_, new_n15560_, new_n15561_, new_n15562_,
    new_n15563_, new_n15564_, new_n15565_, new_n15566_, new_n15567_,
    new_n15568_, new_n15569_, new_n15570_, new_n15571_, new_n15572_,
    new_n15573_, new_n15574_, new_n15575_, new_n15576_, new_n15577_,
    new_n15578_, new_n15579_, new_n15580_, new_n15581_, new_n15582_,
    new_n15583_, new_n15584_, new_n15585_, new_n15586_, new_n15587_,
    new_n15588_, new_n15589_, new_n15590_, new_n15591_, new_n15592_,
    new_n15593_, new_n15594_, new_n15595_, new_n15596_, new_n15597_,
    new_n15598_, new_n15599_, new_n15600_, new_n15601_, new_n15602_,
    new_n15603_, new_n15604_, new_n15605_, new_n15606_, new_n15607_,
    new_n15608_, new_n15609_, new_n15610_, new_n15611_, new_n15612_,
    new_n15613_, new_n15614_, new_n15615_, new_n15616_, new_n15617_,
    new_n15618_, new_n15619_, new_n15620_, new_n15621_, new_n15622_,
    new_n15623_, new_n15624_, new_n15625_, new_n15626_, new_n15627_,
    new_n15628_, new_n15629_, new_n15630_, new_n15631_, new_n15632_,
    new_n15633_, new_n15634_, new_n15635_, new_n15636_, new_n15637_,
    new_n15638_, new_n15639_, new_n15640_, new_n15641_, new_n15642_,
    new_n15643_, new_n15644_, new_n15645_, new_n15646_, new_n15647_,
    new_n15648_, new_n15649_, new_n15650_, new_n15651_, new_n15652_,
    new_n15653_, new_n15654_, new_n15655_, new_n15656_, new_n15657_,
    new_n15658_, new_n15659_, new_n15660_, new_n15661_, new_n15662_,
    new_n15663_, new_n15664_, new_n15665_, new_n15666_, new_n15667_,
    new_n15668_, new_n15669_, new_n15670_, new_n15671_, new_n15672_,
    new_n15673_, new_n15674_, new_n15675_, new_n15676_, new_n15677_,
    new_n15678_, new_n15679_, new_n15680_, new_n15681_, new_n15682_,
    new_n15683_, new_n15684_, new_n15685_, new_n15686_, new_n15687_,
    new_n15688_, new_n15689_, new_n15690_, new_n15691_, new_n15692_,
    new_n15693_, new_n15694_, new_n15695_, new_n15696_, new_n15697_,
    new_n15698_, new_n15699_, new_n15700_, new_n15701_, new_n15702_,
    new_n15703_, new_n15704_, new_n15705_, new_n15706_, new_n15707_,
    new_n15708_, new_n15709_, new_n15710_, new_n15711_, new_n15712_,
    new_n15713_, new_n15714_, new_n15715_, new_n15716_, new_n15717_,
    new_n15718_, new_n15719_, new_n15720_, new_n15721_, new_n15722_,
    new_n15723_, new_n15724_, new_n15725_, new_n15726_, new_n15727_,
    new_n15728_, new_n15729_, new_n15730_, new_n15731_, new_n15732_,
    new_n15733_, new_n15734_, new_n15735_, new_n15736_, new_n15737_,
    new_n15738_, new_n15739_, new_n15740_, new_n15741_, new_n15742_,
    new_n15743_, new_n15744_, new_n15745_, new_n15746_, new_n15747_,
    new_n15748_, new_n15749_, new_n15750_, new_n15751_, new_n15752_,
    new_n15753_, new_n15754_, new_n15755_, new_n15756_, new_n15757_,
    new_n15758_, new_n15759_, new_n15760_, new_n15761_, new_n15762_,
    new_n15763_, new_n15764_, new_n15765_, new_n15766_, new_n15767_,
    new_n15768_, new_n15769_, new_n15770_, new_n15771_, new_n15772_,
    new_n15773_, new_n15774_, new_n15775_, new_n15776_, new_n15777_,
    new_n15778_, new_n15779_, new_n15780_, new_n15781_, new_n15782_,
    new_n15783_, new_n15784_, new_n15785_, new_n15786_, new_n15787_,
    new_n15788_, new_n15789_, new_n15790_, new_n15791_, new_n15792_,
    new_n15793_, new_n15794_, new_n15795_, new_n15796_, new_n15797_,
    new_n15798_, new_n15799_, new_n15800_, new_n15801_, new_n15802_,
    new_n15803_, new_n15804_, new_n15805_, new_n15806_, new_n15807_,
    new_n15808_, new_n15809_, new_n15810_, new_n15811_, new_n15812_,
    new_n15813_, new_n15814_, new_n15815_, new_n15816_, new_n15817_,
    new_n15818_, new_n15819_, new_n15820_, new_n15821_, new_n15822_,
    new_n15823_, new_n15824_, new_n15825_, new_n15826_, new_n15827_,
    new_n15828_, new_n15829_, new_n15830_, new_n15831_, new_n15832_,
    new_n15833_, new_n15834_, new_n15835_, new_n15836_, new_n15837_,
    new_n15838_, new_n15839_, new_n15840_, new_n15841_, new_n15842_,
    new_n15843_, new_n15844_, new_n15845_, new_n15846_, new_n15847_,
    new_n15848_, new_n15849_, new_n15850_, new_n15851_, new_n15852_,
    new_n15853_, new_n15854_, new_n15855_, new_n15856_, new_n15857_,
    new_n15858_, new_n15859_, new_n15860_, new_n15861_, new_n15862_,
    new_n15863_, new_n15864_, new_n15865_, new_n15866_, new_n15867_,
    new_n15868_, new_n15869_, new_n15870_, new_n15871_, new_n15872_,
    new_n15873_, new_n15874_, new_n15875_, new_n15876_, new_n15877_,
    new_n15878_, new_n15879_, new_n15880_, new_n15881_, new_n15882_,
    new_n15883_, new_n15884_, new_n15885_, new_n15886_, new_n15887_,
    new_n15888_, new_n15889_, new_n15890_, new_n15891_, new_n15892_,
    new_n15893_, new_n15894_, new_n15895_, new_n15896_, new_n15897_,
    new_n15898_, new_n15899_, new_n15900_, new_n15901_, new_n15902_,
    new_n15903_, new_n15904_, new_n15905_, new_n15906_, new_n15907_,
    new_n15908_, new_n15909_, new_n15910_, new_n15911_, new_n15912_,
    new_n15913_, new_n15914_, new_n15915_, new_n15916_, new_n15917_,
    new_n15918_, new_n15919_, new_n15920_, new_n15921_, new_n15922_,
    new_n15923_, new_n15924_, new_n15925_, new_n15926_, new_n15927_,
    new_n15928_, new_n15929_, new_n15930_, new_n15931_, new_n15932_,
    new_n15933_, new_n15934_, new_n15935_, new_n15936_, new_n15937_,
    new_n15938_, new_n15939_, new_n15940_, new_n15941_, new_n15942_,
    new_n15943_, new_n15944_, new_n15945_, new_n15946_, new_n15947_,
    new_n15948_, new_n15949_, new_n15950_, new_n15951_, new_n15952_,
    new_n15953_, new_n15954_, new_n15955_, new_n15956_, new_n15957_,
    new_n15958_, new_n15959_, new_n15960_, new_n15961_, new_n15962_,
    new_n15963_, new_n15964_, new_n15965_, new_n15966_, new_n15967_,
    new_n15968_, new_n15969_, new_n15970_, new_n15971_, new_n15972_,
    new_n15973_, new_n15974_, new_n15975_, new_n15976_, new_n15977_,
    new_n15978_, new_n15979_, new_n15980_, new_n15981_, new_n15982_,
    new_n15983_, new_n15984_, new_n15985_, new_n15986_, new_n15987_,
    new_n15988_, new_n15989_, new_n15990_, new_n15991_, new_n15992_,
    new_n15993_, new_n15994_, new_n15995_, new_n15996_, new_n15997_,
    new_n15998_, new_n15999_, new_n16000_, new_n16001_, new_n16002_,
    new_n16003_, new_n16004_, new_n16005_, new_n16006_, new_n16007_,
    new_n16008_, new_n16009_, new_n16010_, new_n16011_, new_n16012_,
    new_n16013_, new_n16014_, new_n16015_, new_n16016_, new_n16017_,
    new_n16018_, new_n16019_, new_n16020_, new_n16021_, new_n16022_,
    new_n16023_, new_n16024_, new_n16025_, new_n16026_, new_n16027_,
    new_n16028_, new_n16029_, new_n16030_, new_n16031_, new_n16032_,
    new_n16033_, new_n16034_, new_n16035_, new_n16036_, new_n16037_,
    new_n16038_, new_n16039_, new_n16040_, new_n16041_, new_n16042_,
    new_n16043_, new_n16044_, new_n16045_, new_n16046_, new_n16047_,
    new_n16048_, new_n16049_, new_n16050_, new_n16051_, new_n16052_,
    new_n16053_, new_n16054_, new_n16055_, new_n16056_, new_n16057_,
    new_n16058_, new_n16059_, new_n16060_, new_n16061_, new_n16062_,
    new_n16063_, new_n16064_, new_n16065_, new_n16066_, new_n16067_,
    new_n16068_, new_n16069_, new_n16070_, new_n16071_, new_n16072_,
    new_n16073_, new_n16074_, new_n16075_, new_n16076_, new_n16077_,
    new_n16078_, new_n16079_, new_n16080_, new_n16081_, new_n16082_,
    new_n16083_, new_n16084_, new_n16085_, new_n16086_, new_n16087_,
    new_n16088_, new_n16089_, new_n16090_, new_n16091_, new_n16092_,
    new_n16093_, new_n16094_, new_n16095_, new_n16096_, new_n16097_,
    new_n16098_, new_n16099_, new_n16100_, new_n16101_, new_n16102_,
    new_n16103_, new_n16104_, new_n16105_, new_n16106_, new_n16107_,
    new_n16108_, new_n16109_, new_n16110_, new_n16111_, new_n16112_,
    new_n16113_, new_n16114_, new_n16115_, new_n16116_, new_n16117_,
    new_n16118_, new_n16119_, new_n16120_, new_n16121_, new_n16122_,
    new_n16123_, new_n16124_, new_n16125_, new_n16126_, new_n16127_,
    new_n16128_, new_n16129_, new_n16130_, new_n16131_, new_n16132_,
    new_n16133_, new_n16134_, new_n16135_, new_n16136_, new_n16137_,
    new_n16138_, new_n16139_, new_n16140_, new_n16141_, new_n16142_,
    new_n16143_, new_n16144_, new_n16145_, new_n16146_, new_n16147_,
    new_n16148_, new_n16149_, new_n16150_, new_n16151_, new_n16152_,
    new_n16153_, new_n16154_, new_n16155_, new_n16156_, new_n16157_,
    new_n16158_, new_n16159_, new_n16160_, new_n16161_, new_n16162_,
    new_n16163_, new_n16164_, new_n16165_, new_n16166_, new_n16167_,
    new_n16168_, new_n16169_, new_n16170_, new_n16171_, new_n16172_,
    new_n16173_, new_n16174_, new_n16175_, new_n16176_, new_n16177_,
    new_n16178_, new_n16179_, new_n16180_, new_n16181_, new_n16182_,
    new_n16183_, new_n16184_, new_n16185_, new_n16186_, new_n16187_,
    new_n16188_, new_n16189_, new_n16190_, new_n16191_, new_n16192_,
    new_n16193_, new_n16194_, new_n16195_, new_n16196_, new_n16197_,
    new_n16198_, new_n16199_, new_n16200_, new_n16201_, new_n16202_,
    new_n16203_, new_n16204_, new_n16205_, new_n16206_, new_n16207_,
    new_n16208_, new_n16209_, new_n16210_, new_n16211_, new_n16212_,
    new_n16213_, new_n16214_, new_n16215_, new_n16216_, new_n16217_,
    new_n16218_, new_n16219_, new_n16220_, new_n16221_, new_n16222_,
    new_n16223_, new_n16224_, new_n16225_, new_n16226_, new_n16227_,
    new_n16228_, new_n16229_, new_n16230_, new_n16231_, new_n16232_,
    new_n16233_, new_n16234_, new_n16235_, new_n16236_, new_n16237_,
    new_n16238_, new_n16239_, new_n16240_, new_n16241_, new_n16242_,
    new_n16243_, new_n16244_, new_n16245_, new_n16246_, new_n16247_,
    new_n16248_, new_n16249_, new_n16250_, new_n16251_, new_n16252_,
    new_n16253_, new_n16254_, new_n16255_, new_n16256_, new_n16257_,
    new_n16258_, new_n16259_, new_n16260_, new_n16261_, new_n16262_,
    new_n16263_, new_n16264_, new_n16265_, new_n16266_, new_n16267_,
    new_n16268_, new_n16269_, new_n16270_, new_n16271_, new_n16272_,
    new_n16273_, new_n16274_, new_n16275_, new_n16276_, new_n16277_,
    new_n16278_, new_n16279_, new_n16280_, new_n16281_, new_n16282_,
    new_n16283_, new_n16284_, new_n16285_, new_n16286_, new_n16287_,
    new_n16288_, new_n16289_, new_n16290_, new_n16291_, new_n16292_,
    new_n16293_, new_n16294_, new_n16295_, new_n16296_, new_n16297_,
    new_n16298_, new_n16299_, new_n16300_, new_n16301_, new_n16302_,
    new_n16303_, new_n16304_, new_n16305_, new_n16306_, new_n16307_,
    new_n16308_, new_n16309_, new_n16310_, new_n16311_, new_n16312_,
    new_n16313_, new_n16314_, new_n16315_, new_n16316_, new_n16317_,
    new_n16318_, new_n16319_, new_n16320_, new_n16321_, new_n16322_,
    new_n16323_, new_n16324_, new_n16325_, new_n16326_, new_n16327_,
    new_n16328_, new_n16329_, new_n16330_, new_n16331_, new_n16332_,
    new_n16333_, new_n16334_, new_n16335_, new_n16336_, new_n16337_,
    new_n16338_, new_n16339_, new_n16340_, new_n16341_, new_n16342_,
    new_n16343_, new_n16344_, new_n16345_, new_n16346_, new_n16347_,
    new_n16348_, new_n16349_, new_n16350_, new_n16351_, new_n16352_,
    new_n16353_, new_n16354_, new_n16355_, new_n16356_, new_n16357_,
    new_n16358_, new_n16359_, new_n16360_, new_n16361_, new_n16362_,
    new_n16363_, new_n16364_, new_n16365_, new_n16366_, new_n16367_,
    new_n16368_, new_n16369_, new_n16370_, new_n16371_, new_n16372_,
    new_n16373_, new_n16374_, new_n16375_, new_n16376_, new_n16377_,
    new_n16378_, new_n16379_, new_n16380_, new_n16381_, new_n16382_,
    new_n16383_, new_n16384_, new_n16385_, new_n16386_, new_n16387_,
    new_n16388_, new_n16389_, new_n16390_, new_n16391_, new_n16392_,
    new_n16393_, new_n16394_, new_n16395_, new_n16396_, new_n16397_,
    new_n16398_, new_n16399_, new_n16400_, new_n16401_, new_n16402_,
    new_n16403_, new_n16404_, new_n16405_, new_n16406_, new_n16407_,
    new_n16408_, new_n16409_, new_n16410_, new_n16411_, new_n16412_,
    new_n16413_, new_n16414_, new_n16415_, new_n16416_, new_n16417_,
    new_n16418_, new_n16419_, new_n16420_, new_n16421_, new_n16422_,
    new_n16423_, new_n16424_, new_n16425_, new_n16426_, new_n16427_,
    new_n16428_, new_n16429_, new_n16430_, new_n16431_, new_n16432_,
    new_n16433_, new_n16434_, new_n16435_, new_n16436_, new_n16437_,
    new_n16438_, new_n16439_, new_n16440_, new_n16441_, new_n16442_,
    new_n16443_, new_n16444_, new_n16445_, new_n16446_, new_n16447_,
    new_n16448_, new_n16449_, new_n16450_, new_n16451_, new_n16452_,
    new_n16453_, new_n16454_, new_n16455_, new_n16456_, new_n16457_,
    new_n16458_, new_n16459_, new_n16460_, new_n16461_, new_n16462_,
    new_n16463_, new_n16464_, new_n16465_, new_n16466_, new_n16467_,
    new_n16468_, new_n16469_, new_n16470_, new_n16471_, new_n16472_,
    new_n16473_, new_n16474_, new_n16475_, new_n16476_, new_n16477_,
    new_n16478_, new_n16479_, new_n16480_, new_n16481_, new_n16482_,
    new_n16483_, new_n16484_, new_n16485_, new_n16486_, new_n16487_,
    new_n16488_, new_n16489_, new_n16490_, new_n16491_, new_n16492_,
    new_n16493_, new_n16494_, new_n16495_, new_n16496_, new_n16497_,
    new_n16498_, new_n16499_, new_n16500_, new_n16501_, new_n16502_,
    new_n16503_, new_n16504_, new_n16505_, new_n16506_, new_n16507_,
    new_n16508_, new_n16509_, new_n16510_, new_n16511_, new_n16512_,
    new_n16513_, new_n16514_, new_n16515_, new_n16516_, new_n16517_,
    new_n16518_, new_n16519_, new_n16520_, new_n16521_, new_n16522_,
    new_n16523_, new_n16524_, new_n16525_, new_n16526_, new_n16527_,
    new_n16528_, new_n16529_, new_n16530_, new_n16531_, new_n16532_,
    new_n16533_, new_n16534_, new_n16535_, new_n16536_, new_n16537_,
    new_n16538_, new_n16539_, new_n16540_, new_n16541_, new_n16542_,
    new_n16543_, new_n16544_, new_n16545_, new_n16546_, new_n16547_,
    new_n16548_, new_n16549_, new_n16550_, new_n16551_, new_n16552_,
    new_n16553_, new_n16554_, new_n16555_, new_n16556_, new_n16557_,
    new_n16558_, new_n16559_, new_n16560_, new_n16561_, new_n16562_,
    new_n16563_, new_n16564_, new_n16565_, new_n16566_, new_n16567_,
    new_n16568_, new_n16569_, new_n16570_, new_n16571_, new_n16572_,
    new_n16573_, new_n16574_, new_n16575_, new_n16576_, new_n16577_,
    new_n16578_, new_n16579_, new_n16580_, new_n16581_, new_n16582_,
    new_n16583_, new_n16584_, new_n16585_, new_n16586_, new_n16587_,
    new_n16588_, new_n16589_, new_n16590_, new_n16591_, new_n16592_,
    new_n16593_, new_n16594_, new_n16595_, new_n16596_, new_n16597_,
    new_n16598_, new_n16599_, new_n16600_, new_n16601_, new_n16602_,
    new_n16603_, new_n16604_, new_n16605_, new_n16606_, new_n16607_,
    new_n16608_, new_n16609_, new_n16610_, new_n16611_, new_n16612_,
    new_n16613_, new_n16614_, new_n16615_, new_n16616_, new_n16617_,
    new_n16618_, new_n16619_, new_n16620_, new_n16621_, new_n16622_,
    new_n16623_, new_n16624_, new_n16625_, new_n16626_, new_n16627_,
    new_n16628_, new_n16629_, new_n16630_, new_n16631_, new_n16632_,
    new_n16633_, new_n16634_, new_n16635_, new_n16636_, new_n16637_,
    new_n16638_, new_n16639_, new_n16640_, new_n16641_, new_n16642_,
    new_n16643_, new_n16644_, new_n16645_, new_n16646_, new_n16647_,
    new_n16648_, new_n16649_, new_n16650_, new_n16651_, new_n16652_,
    new_n16653_, new_n16654_, new_n16655_, new_n16656_, new_n16657_,
    new_n16658_, new_n16659_, new_n16660_, new_n16661_, new_n16662_,
    new_n16663_, new_n16664_, new_n16665_, new_n16666_, new_n16667_,
    new_n16668_, new_n16669_, new_n16670_, new_n16671_, new_n16672_,
    new_n16673_, new_n16674_, new_n16675_, new_n16676_, new_n16677_,
    new_n16678_, new_n16679_, new_n16680_, new_n16681_, new_n16682_,
    new_n16683_, new_n16684_, new_n16685_, new_n16686_, new_n16687_,
    new_n16688_, new_n16689_, new_n16690_, new_n16691_, new_n16692_,
    new_n16693_, new_n16694_, new_n16695_, new_n16696_, new_n16697_,
    new_n16698_, new_n16699_, new_n16700_, new_n16701_, new_n16702_,
    new_n16703_, new_n16704_, new_n16705_, new_n16706_, new_n16707_,
    new_n16708_, new_n16709_, new_n16710_, new_n16711_, new_n16712_,
    new_n16713_, new_n16714_, new_n16715_, new_n16716_, new_n16717_,
    new_n16718_, new_n16719_, new_n16720_, new_n16721_, new_n16722_,
    new_n16723_, new_n16724_, new_n16725_, new_n16726_, new_n16727_,
    new_n16728_, new_n16729_, new_n16730_, new_n16731_, new_n16732_,
    new_n16733_, new_n16734_, new_n16735_, new_n16736_, new_n16737_,
    new_n16738_, new_n16739_, new_n16740_, new_n16741_, new_n16742_,
    new_n16743_, new_n16744_, new_n16745_, new_n16746_, new_n16747_,
    new_n16748_, new_n16749_, new_n16750_, new_n16751_, new_n16752_,
    new_n16753_, new_n16754_, new_n16755_, new_n16756_, new_n16757_,
    new_n16758_, new_n16759_, new_n16760_, new_n16761_, new_n16762_,
    new_n16763_, new_n16764_, new_n16765_, new_n16766_, new_n16767_,
    new_n16768_, new_n16769_, new_n16770_, new_n16771_, new_n16772_,
    new_n16773_, new_n16774_, new_n16775_, new_n16776_, new_n16777_,
    new_n16778_, new_n16779_, new_n16780_, new_n16781_, new_n16782_,
    new_n16783_, new_n16784_, new_n16785_, new_n16786_, new_n16787_,
    new_n16788_, new_n16789_, new_n16790_, new_n16791_, new_n16792_,
    new_n16793_, new_n16794_, new_n16795_, new_n16796_, new_n16797_,
    new_n16798_, new_n16799_, new_n16800_, new_n16801_, new_n16802_,
    new_n16803_, new_n16804_, new_n16805_, new_n16806_, new_n16807_,
    new_n16808_, new_n16809_, new_n16810_, new_n16811_, new_n16812_,
    new_n16813_, new_n16814_, new_n16815_, new_n16816_, new_n16817_,
    new_n16818_, new_n16819_, new_n16820_, new_n16821_, new_n16822_,
    new_n16823_, new_n16824_, new_n16825_, new_n16826_, new_n16827_,
    new_n16828_, new_n16829_, new_n16830_, new_n16831_, new_n16832_,
    new_n16833_, new_n16834_, new_n16835_, new_n16836_, new_n16837_,
    new_n16838_, new_n16839_, new_n16840_, new_n16841_, new_n16842_,
    new_n16843_, new_n16844_, new_n16845_, new_n16846_, new_n16847_,
    new_n16848_, new_n16849_, new_n16850_, new_n16851_, new_n16852_,
    new_n16853_, new_n16854_, new_n16855_, new_n16856_, new_n16857_,
    new_n16858_, new_n16859_, new_n16860_, new_n16861_, new_n16862_,
    new_n16863_, new_n16864_, new_n16865_, new_n16866_, new_n16867_,
    new_n16868_, new_n16869_, new_n16870_, new_n16871_, new_n16872_,
    new_n16873_, new_n16874_, new_n16875_, new_n16876_, new_n16877_,
    new_n16878_, new_n16879_, new_n16880_, new_n16881_, new_n16882_,
    new_n16883_, new_n16884_, new_n16885_, new_n16886_, new_n16887_,
    new_n16888_, new_n16889_, new_n16890_, new_n16891_, new_n16892_,
    new_n16893_, new_n16894_, new_n16895_, new_n16896_, new_n16897_,
    new_n16898_, new_n16899_, new_n16900_, new_n16901_, new_n16902_,
    new_n16903_, new_n16904_, new_n16905_, new_n16906_, new_n16907_,
    new_n16908_, new_n16909_, new_n16910_, new_n16911_, new_n16912_,
    new_n16913_, new_n16914_, new_n16915_, new_n16916_, new_n16917_,
    new_n16918_, new_n16919_, new_n16920_, new_n16921_, new_n16922_,
    new_n16923_, new_n16924_, new_n16925_, new_n16926_, new_n16927_,
    new_n16928_, new_n16929_, new_n16930_, new_n16931_, new_n16932_,
    new_n16933_, new_n16934_, new_n16935_, new_n16936_, new_n16937_,
    new_n16938_, new_n16939_, new_n16940_, new_n16941_, new_n16942_,
    new_n16943_, new_n16944_, new_n16945_, new_n16946_, new_n16947_,
    new_n16948_, new_n16949_, new_n16950_, new_n16951_, new_n16952_,
    new_n16953_, new_n16954_, new_n16955_, new_n16956_, new_n16957_,
    new_n16958_, new_n16959_, new_n16960_, new_n16961_, new_n16962_,
    new_n16963_, new_n16964_, new_n16965_, new_n16966_, new_n16967_,
    new_n16968_, new_n16969_, new_n16970_, new_n16971_, new_n16972_,
    new_n16973_, new_n16974_, new_n16975_, new_n16976_, new_n16977_,
    new_n16978_, new_n16979_, new_n16980_, new_n16981_, new_n16982_,
    new_n16983_, new_n16984_, new_n16985_, new_n16986_, new_n16987_,
    new_n16988_, new_n16989_, new_n16990_, new_n16991_, new_n16992_,
    new_n16993_, new_n16994_, new_n16995_, new_n16996_, new_n16997_,
    new_n16998_, new_n16999_, new_n17000_, new_n17001_, new_n17002_,
    new_n17003_, new_n17004_, new_n17005_, new_n17006_, new_n17007_,
    new_n17008_, new_n17009_, new_n17010_, new_n17011_, new_n17012_,
    new_n17013_, new_n17014_, new_n17015_, new_n17016_, new_n17017_,
    new_n17018_, new_n17019_, new_n17020_, new_n17021_, new_n17022_,
    new_n17023_, new_n17024_, new_n17025_, new_n17026_, new_n17027_,
    new_n17028_, new_n17029_, new_n17030_, new_n17031_, new_n17032_,
    new_n17033_, new_n17034_, new_n17035_, new_n17036_, new_n17037_,
    new_n17038_, new_n17039_, new_n17040_, new_n17041_, new_n17042_,
    new_n17043_, new_n17044_, new_n17045_, new_n17046_, new_n17047_,
    new_n17048_, new_n17049_, new_n17050_, new_n17051_, new_n17052_,
    new_n17053_, new_n17054_, new_n17055_, new_n17056_, new_n17057_,
    new_n17058_, new_n17059_, new_n17060_, new_n17061_, new_n17062_,
    new_n17063_, new_n17064_, new_n17065_, new_n17066_, new_n17067_,
    new_n17068_, new_n17069_, new_n17070_, new_n17071_, new_n17072_,
    new_n17073_, new_n17074_, new_n17075_, new_n17076_, new_n17077_,
    new_n17078_, new_n17079_, new_n17080_, new_n17081_, new_n17082_,
    new_n17083_, new_n17084_, new_n17085_, new_n17086_, new_n17087_,
    new_n17088_, new_n17089_, new_n17090_, new_n17091_, new_n17092_,
    new_n17093_, new_n17094_, new_n17095_, new_n17096_, new_n17097_,
    new_n17098_, new_n17099_, new_n17100_, new_n17101_, new_n17102_,
    new_n17103_, new_n17104_, new_n17105_, new_n17106_, new_n17107_,
    new_n17108_, new_n17109_, new_n17110_, new_n17111_, new_n17112_,
    new_n17113_, new_n17114_, new_n17115_, new_n17116_, new_n17117_,
    new_n17118_, new_n17119_, new_n17120_, new_n17121_, new_n17122_,
    new_n17123_, new_n17124_, new_n17125_, new_n17126_, new_n17127_,
    new_n17128_, new_n17129_, new_n17130_, new_n17131_, new_n17132_,
    new_n17133_, new_n17134_, new_n17135_, new_n17136_, new_n17137_,
    new_n17138_, new_n17139_, new_n17140_, new_n17141_, new_n17142_,
    new_n17143_, new_n17144_, new_n17145_, new_n17146_, new_n17147_,
    new_n17148_, new_n17149_, new_n17150_, new_n17151_, new_n17152_,
    new_n17153_, new_n17154_, new_n17155_, new_n17156_, new_n17157_,
    new_n17158_, new_n17159_, new_n17160_, new_n17161_, new_n17162_,
    new_n17163_, new_n17164_, new_n17165_, new_n17166_, new_n17167_,
    new_n17168_, new_n17169_, new_n17170_, new_n17171_, new_n17172_,
    new_n17173_, new_n17174_, new_n17175_, new_n17176_, new_n17177_,
    new_n17178_, new_n17179_, new_n17180_, new_n17181_, new_n17182_,
    new_n17183_, new_n17184_, new_n17185_, new_n17186_, new_n17187_,
    new_n17188_, new_n17189_, new_n17190_, new_n17191_, new_n17192_,
    new_n17193_, new_n17194_, new_n17195_, new_n17196_, new_n17197_,
    new_n17198_, new_n17199_, new_n17200_, new_n17201_, new_n17202_,
    new_n17203_, new_n17204_, new_n17205_, new_n17206_, new_n17207_,
    new_n17208_, new_n17209_, new_n17210_, new_n17211_, new_n17212_,
    new_n17213_, new_n17214_, new_n17215_, new_n17216_, new_n17217_,
    new_n17218_, new_n17219_, new_n17220_, new_n17221_, new_n17222_,
    new_n17223_, new_n17224_, new_n17225_, new_n17226_, new_n17227_,
    new_n17228_, new_n17229_, new_n17230_, new_n17231_, new_n17232_,
    new_n17233_, new_n17234_, new_n17235_, new_n17236_, new_n17237_,
    new_n17238_, new_n17239_, new_n17240_, new_n17241_, new_n17242_,
    new_n17243_, new_n17244_, new_n17245_, new_n17246_, new_n17247_,
    new_n17248_, new_n17249_, new_n17250_, new_n17251_, new_n17252_,
    new_n17253_, new_n17254_, new_n17255_, new_n17256_, new_n17257_,
    new_n17258_, new_n17259_, new_n17260_, new_n17261_, new_n17262_,
    new_n17263_, new_n17264_, new_n17265_, new_n17266_, new_n17267_,
    new_n17268_, new_n17269_, new_n17270_, new_n17271_, new_n17272_,
    new_n17273_, new_n17274_, new_n17275_, new_n17276_, new_n17277_,
    new_n17278_, new_n17279_, new_n17280_, new_n17281_, new_n17282_,
    new_n17283_, new_n17284_, new_n17285_, new_n17286_, new_n17287_,
    new_n17288_, new_n17289_, new_n17290_, new_n17291_, new_n17292_,
    new_n17293_, new_n17294_, new_n17295_, new_n17296_, new_n17297_,
    new_n17298_, new_n17299_, new_n17300_, new_n17301_, new_n17302_,
    new_n17303_, new_n17304_, new_n17305_, new_n17306_, new_n17307_,
    new_n17308_, new_n17309_, new_n17310_, new_n17311_, new_n17312_,
    new_n17313_, new_n17314_, new_n17315_, new_n17316_, new_n17317_,
    new_n17318_, new_n17319_, new_n17320_, new_n17321_, new_n17322_,
    new_n17323_, new_n17324_, new_n17325_, new_n17326_, new_n17327_,
    new_n17328_, new_n17329_, new_n17330_, new_n17331_, new_n17332_,
    new_n17333_, new_n17334_, new_n17335_, new_n17336_, new_n17337_,
    new_n17338_, new_n17339_, new_n17340_, new_n17341_, new_n17342_,
    new_n17343_, new_n17344_, new_n17345_, new_n17346_, new_n17347_,
    new_n17348_, new_n17349_, new_n17350_, new_n17351_, new_n17352_,
    new_n17353_, new_n17354_, new_n17355_, new_n17356_, new_n17357_,
    new_n17358_, new_n17359_, new_n17360_, new_n17361_, new_n17362_,
    new_n17363_, new_n17364_, new_n17365_, new_n17366_, new_n17367_,
    new_n17368_, new_n17369_, new_n17370_, new_n17371_, new_n17372_,
    new_n17373_, new_n17374_, new_n17375_, new_n17376_, new_n17377_,
    new_n17378_, new_n17379_, new_n17380_, new_n17381_, new_n17382_,
    new_n17383_, new_n17384_, new_n17385_, new_n17386_, new_n17387_,
    new_n17388_, new_n17389_, new_n17390_, new_n17391_, new_n17392_,
    new_n17393_, new_n17394_, new_n17395_, new_n17396_, new_n17397_,
    new_n17398_, new_n17399_, new_n17400_, new_n17401_, new_n17402_,
    new_n17403_, new_n17404_, new_n17405_, new_n17406_, new_n17407_,
    new_n17408_, new_n17409_, new_n17410_, new_n17411_, new_n17412_,
    new_n17413_, new_n17414_, new_n17415_, new_n17416_, new_n17417_,
    new_n17418_, new_n17419_, new_n17420_, new_n17421_, new_n17422_,
    new_n17423_, new_n17424_, new_n17425_, new_n17426_, new_n17427_,
    new_n17428_, new_n17429_, new_n17430_, new_n17431_, new_n17432_,
    new_n17433_, new_n17434_, new_n17435_, new_n17436_, new_n17437_,
    new_n17438_, new_n17439_, new_n17440_, new_n17441_, new_n17442_,
    new_n17443_, new_n17444_, new_n17445_, new_n17446_, new_n17447_,
    new_n17448_, new_n17449_, new_n17450_, new_n17451_, new_n17452_,
    new_n17453_, new_n17454_, new_n17455_, new_n17456_, new_n17457_,
    new_n17458_, new_n17459_, new_n17460_, new_n17461_, new_n17462_,
    new_n17463_, new_n17464_, new_n17465_, new_n17466_, new_n17467_,
    new_n17468_, new_n17469_, new_n17470_, new_n17471_, new_n17472_,
    new_n17473_, new_n17474_, new_n17475_, new_n17476_, new_n17477_,
    new_n17478_, new_n17479_, new_n17480_, new_n17481_, new_n17482_,
    new_n17483_, new_n17484_, new_n17485_, new_n17486_, new_n17487_,
    new_n17488_, new_n17489_, new_n17490_, new_n17491_, new_n17492_,
    new_n17493_, new_n17494_, new_n17495_, new_n17496_, new_n17497_,
    new_n17498_, new_n17499_, new_n17500_, new_n17501_, new_n17502_,
    new_n17503_, new_n17504_, new_n17505_, new_n17506_, new_n17507_,
    new_n17508_, new_n17509_, new_n17510_, new_n17511_, new_n17512_,
    new_n17513_, new_n17514_, new_n17515_, new_n17516_, new_n17517_,
    new_n17518_, new_n17519_, new_n17520_, new_n17521_, new_n17522_,
    new_n17523_, new_n17524_, new_n17525_, new_n17526_, new_n17527_,
    new_n17528_, new_n17529_, new_n17530_, new_n17531_, new_n17532_,
    new_n17533_, new_n17534_, new_n17535_, new_n17536_, new_n17537_,
    new_n17538_, new_n17539_, new_n17540_, new_n17541_, new_n17542_,
    new_n17543_, new_n17544_, new_n17545_, new_n17546_, new_n17547_,
    new_n17548_, new_n17549_, new_n17550_, new_n17551_, new_n17552_,
    new_n17553_, new_n17554_, new_n17555_, new_n17556_, new_n17557_,
    new_n17558_, new_n17559_, new_n17560_, new_n17561_, new_n17562_,
    new_n17563_, new_n17564_, new_n17565_, new_n17566_, new_n17567_,
    new_n17568_, new_n17569_, new_n17570_, new_n17571_, new_n17572_,
    new_n17573_, new_n17574_, new_n17575_, new_n17576_, new_n17577_,
    new_n17578_, new_n17579_, new_n17580_, new_n17581_, new_n17582_,
    new_n17583_, new_n17584_, new_n17585_, new_n17586_, new_n17587_,
    new_n17588_, new_n17589_, new_n17590_, new_n17591_, new_n17592_,
    new_n17593_, new_n17594_, new_n17595_, new_n17596_, new_n17597_,
    new_n17598_, new_n17599_, new_n17600_, new_n17601_, new_n17602_,
    new_n17603_, new_n17604_, new_n17605_, new_n17606_, new_n17607_,
    new_n17608_, new_n17609_, new_n17610_, new_n17611_, new_n17612_,
    new_n17613_, new_n17614_, new_n17615_, new_n17616_, new_n17617_,
    new_n17618_, new_n17619_, new_n17620_, new_n17621_, new_n17622_,
    new_n17623_, new_n17624_, new_n17625_, new_n17626_, new_n17627_,
    new_n17628_, new_n17629_, new_n17630_, new_n17631_, new_n17632_,
    new_n17633_, new_n17634_, new_n17635_, new_n17636_, new_n17637_,
    new_n17638_, new_n17639_, new_n17640_, new_n17641_, new_n17642_,
    new_n17643_, new_n17644_, new_n17645_, new_n17646_, new_n17647_,
    new_n17648_, new_n17649_, new_n17650_, new_n17651_, new_n17652_,
    new_n17653_, new_n17654_, new_n17655_, new_n17656_, new_n17657_,
    new_n17658_, new_n17659_, new_n17660_, new_n17661_, new_n17662_,
    new_n17663_, new_n17664_, new_n17665_, new_n17666_, new_n17667_,
    new_n17668_, new_n17669_, new_n17670_, new_n17671_, new_n17672_,
    new_n17673_, new_n17674_, new_n17675_, new_n17676_, new_n17677_,
    new_n17678_, new_n17679_, new_n17680_, new_n17681_, new_n17682_,
    new_n17683_, new_n17684_, new_n17685_, new_n17686_, new_n17687_,
    new_n17688_, new_n17689_, new_n17690_, new_n17691_, new_n17692_,
    new_n17693_, new_n17694_, new_n17695_, new_n17696_, new_n17697_,
    new_n17698_, new_n17699_, new_n17700_, new_n17701_, new_n17702_,
    new_n17703_, new_n17704_, new_n17705_, new_n17706_, new_n17707_,
    new_n17708_, new_n17709_, new_n17710_, new_n17711_, new_n17712_,
    new_n17713_, new_n17714_, new_n17715_, new_n17716_, new_n17717_,
    new_n17718_, new_n17719_, new_n17720_, new_n17721_, new_n17722_,
    new_n17723_, new_n17724_, new_n17725_, new_n17726_, new_n17727_,
    new_n17728_, new_n17729_, new_n17730_, new_n17731_, new_n17732_,
    new_n17733_, new_n17734_, new_n17735_, new_n17736_, new_n17737_,
    new_n17738_, new_n17739_, new_n17740_, new_n17741_, new_n17742_,
    new_n17743_, new_n17744_, new_n17745_, new_n17746_, new_n17747_,
    new_n17748_, new_n17749_, new_n17750_, new_n17751_, new_n17752_,
    new_n17753_, new_n17754_, new_n17755_, new_n17756_, new_n17757_,
    new_n17758_, new_n17759_, new_n17760_, new_n17761_, new_n17762_,
    new_n17763_, new_n17764_, new_n17765_, new_n17766_, new_n17767_,
    new_n17768_, new_n17769_, new_n17770_, new_n17771_, new_n17772_,
    new_n17773_, new_n17774_, new_n17775_, new_n17776_, new_n17777_,
    new_n17778_, new_n17779_, new_n17780_, new_n17781_, new_n17782_,
    new_n17783_, new_n17784_, new_n17785_, new_n17786_, new_n17787_,
    new_n17788_, new_n17789_, new_n17790_, new_n17791_, new_n17792_,
    new_n17793_, new_n17794_, new_n17795_, new_n17796_, new_n17797_,
    new_n17798_, new_n17799_, new_n17800_, new_n17801_, new_n17802_,
    new_n17803_, new_n17804_, new_n17805_, new_n17806_, new_n17807_,
    new_n17808_, new_n17809_, new_n17810_, new_n17811_, new_n17812_,
    new_n17813_, new_n17814_, new_n17815_, new_n17816_, new_n17817_,
    new_n17818_, new_n17819_, new_n17820_, new_n17821_, new_n17822_,
    new_n17823_, new_n17824_, new_n17825_, new_n17826_, new_n17827_,
    new_n17828_, new_n17829_, new_n17830_, new_n17831_, new_n17832_,
    new_n17833_, new_n17834_, new_n17835_, new_n17836_, new_n17837_,
    new_n17838_, new_n17839_, new_n17840_, new_n17841_, new_n17842_,
    new_n17843_, new_n17844_, new_n17845_, new_n17846_, new_n17847_,
    new_n17848_, new_n17849_, new_n17850_, new_n17851_, new_n17852_,
    new_n17853_, new_n17854_, new_n17855_, new_n17856_, new_n17857_,
    new_n17858_, new_n17859_, new_n17860_, new_n17861_, new_n17862_,
    new_n17863_, new_n17864_, new_n17865_, new_n17866_, new_n17867_,
    new_n17868_, new_n17869_, new_n17870_, new_n17871_, new_n17872_,
    new_n17873_, new_n17874_, new_n17875_, new_n17876_, new_n17877_,
    new_n17878_, new_n17879_, new_n17880_, new_n17881_, new_n17882_,
    new_n17883_, new_n17884_, new_n17885_, new_n17886_, new_n17887_,
    new_n17888_, new_n17889_, new_n17890_, new_n17891_, new_n17892_,
    new_n17893_, new_n17894_, new_n17895_, new_n17896_, new_n17897_,
    new_n17898_, new_n17899_, new_n17900_, new_n17901_, new_n17902_,
    new_n17903_, new_n17904_, new_n17905_, new_n17906_, new_n17907_,
    new_n17908_, new_n17909_, new_n17910_, new_n17911_, new_n17912_,
    new_n17913_, new_n17914_, new_n17915_, new_n17916_, new_n17917_,
    new_n17918_, new_n17919_, new_n17920_, new_n17921_, new_n17922_,
    new_n17923_, new_n17924_, new_n17925_, new_n17926_, new_n17927_,
    new_n17928_, new_n17929_, new_n17930_, new_n17931_, new_n17932_,
    new_n17933_, new_n17934_, new_n17935_, new_n17936_, new_n17937_,
    new_n17938_, new_n17939_, new_n17940_, new_n17941_, new_n17942_,
    new_n17943_, new_n17944_, new_n17945_, new_n17946_, new_n17947_,
    new_n17948_, new_n17949_, new_n17950_, new_n17951_, new_n17952_,
    new_n17953_, new_n17954_, new_n17955_, new_n17956_, new_n17957_,
    new_n17958_, new_n17959_, new_n17960_, new_n17961_, new_n17962_,
    new_n17963_, new_n17964_, new_n17965_, new_n17966_, new_n17967_,
    new_n17968_, new_n17969_, new_n17970_, new_n17971_, new_n17972_,
    new_n17973_, new_n17974_, new_n17975_, new_n17976_, new_n17977_,
    new_n17978_, new_n17979_, new_n17980_, new_n17981_, new_n17982_,
    new_n17983_, new_n17984_, new_n17985_, new_n17986_, new_n17987_,
    new_n17988_, new_n17989_, new_n17990_, new_n17991_, new_n17992_,
    new_n17993_, new_n17994_, new_n17995_, new_n17996_, new_n17997_,
    new_n17998_, new_n17999_, new_n18000_, new_n18001_, new_n18002_,
    new_n18003_, new_n18004_, new_n18005_, new_n18006_, new_n18007_,
    new_n18008_, new_n18009_, new_n18010_, new_n18011_, new_n18012_,
    new_n18013_, new_n18014_, new_n18015_, new_n18016_, new_n18017_,
    new_n18018_, new_n18019_, new_n18020_, new_n18021_, new_n18022_,
    new_n18023_, new_n18024_, new_n18025_, new_n18026_, new_n18027_,
    new_n18028_, new_n18029_, new_n18030_, new_n18031_, new_n18032_,
    new_n18033_, new_n18034_, new_n18035_, new_n18036_, new_n18037_,
    new_n18038_, new_n18039_, new_n18040_, new_n18041_, new_n18042_,
    new_n18043_, new_n18044_, new_n18045_, new_n18046_, new_n18047_,
    new_n18048_, new_n18049_, new_n18050_, new_n18051_, new_n18052_,
    new_n18053_, new_n18054_, new_n18055_, new_n18056_, new_n18057_,
    new_n18058_, new_n18059_, new_n18060_, new_n18061_, new_n18062_,
    new_n18063_, new_n18064_, new_n18065_, new_n18066_, new_n18067_,
    new_n18068_, new_n18069_, new_n18070_, new_n18071_, new_n18072_,
    new_n18073_, new_n18074_, new_n18075_, new_n18076_, new_n18077_,
    new_n18078_, new_n18079_, new_n18080_, new_n18081_, new_n18082_,
    new_n18083_, new_n18084_, new_n18085_, new_n18086_, new_n18087_,
    new_n18088_, new_n18089_, new_n18090_, new_n18091_, new_n18092_,
    new_n18093_, new_n18094_, new_n18095_, new_n18096_, new_n18097_,
    new_n18098_, new_n18099_, new_n18100_, new_n18101_, new_n18102_,
    new_n18103_, new_n18104_, new_n18105_, new_n18106_, new_n18107_,
    new_n18108_, new_n18109_, new_n18110_, new_n18111_, new_n18112_,
    new_n18113_, new_n18114_, new_n18115_, new_n18116_, new_n18117_,
    new_n18118_, new_n18119_, new_n18120_, new_n18121_, new_n18122_,
    new_n18123_, new_n18124_, new_n18125_, new_n18126_, new_n18127_,
    new_n18128_, new_n18129_, new_n18130_, new_n18131_, new_n18132_,
    new_n18133_, new_n18134_, new_n18135_, new_n18136_, new_n18137_,
    new_n18138_, new_n18139_, new_n18140_, new_n18141_, new_n18142_,
    new_n18143_, new_n18144_, new_n18145_, new_n18146_, new_n18147_,
    new_n18148_, new_n18149_, new_n18150_, new_n18151_, new_n18152_,
    new_n18153_, new_n18154_, new_n18155_, new_n18156_, new_n18157_,
    new_n18158_, new_n18159_, new_n18160_, new_n18161_, new_n18162_,
    new_n18163_, new_n18164_, new_n18165_, new_n18166_, new_n18167_,
    new_n18168_, new_n18169_, new_n18170_, new_n18171_, new_n18172_,
    new_n18173_, new_n18174_, new_n18175_, new_n18176_, new_n18177_,
    new_n18178_, new_n18179_, new_n18180_, new_n18181_, new_n18182_,
    new_n18183_, new_n18184_, new_n18185_, new_n18186_, new_n18187_,
    new_n18188_, new_n18189_, new_n18190_, new_n18191_, new_n18192_,
    new_n18193_, new_n18194_, new_n18195_, new_n18196_, new_n18197_,
    new_n18198_, new_n18199_, new_n18200_, new_n18201_, new_n18202_,
    new_n18203_, new_n18204_, new_n18205_, new_n18206_, new_n18207_,
    new_n18208_, new_n18209_, new_n18210_, new_n18211_, new_n18212_,
    new_n18213_, new_n18214_, new_n18215_, new_n18216_, new_n18217_,
    new_n18218_, new_n18219_, new_n18220_, new_n18221_, new_n18222_,
    new_n18223_, new_n18224_, new_n18225_, new_n18226_, new_n18227_,
    new_n18228_, new_n18229_, new_n18230_, new_n18231_, new_n18232_,
    new_n18233_, new_n18234_, new_n18235_, new_n18236_, new_n18237_,
    new_n18238_, new_n18239_, new_n18240_, new_n18241_, new_n18242_,
    new_n18243_, new_n18244_, new_n18245_, new_n18246_, new_n18247_,
    new_n18248_, new_n18249_, new_n18250_, new_n18251_, new_n18252_,
    new_n18253_, new_n18254_, new_n18255_, new_n18256_, new_n18257_,
    new_n18258_, new_n18259_, new_n18260_, new_n18261_, new_n18262_,
    new_n18263_, new_n18264_, new_n18265_, new_n18266_, new_n18267_,
    new_n18268_, new_n18269_, new_n18270_, new_n18271_, new_n18272_,
    new_n18273_, new_n18274_, new_n18275_, new_n18276_, new_n18277_,
    new_n18278_, new_n18279_, new_n18280_, new_n18281_, new_n18282_,
    new_n18283_, new_n18284_, new_n18285_, new_n18286_, new_n18287_,
    new_n18288_, new_n18289_, new_n18290_, new_n18291_, new_n18292_,
    new_n18293_, new_n18294_, new_n18295_, new_n18296_, new_n18297_,
    new_n18298_, new_n18299_, new_n18300_, new_n18301_, new_n18302_,
    new_n18303_, new_n18304_, new_n18305_, new_n18306_, new_n18307_,
    new_n18308_, new_n18309_, new_n18310_, new_n18311_, new_n18312_,
    new_n18313_, new_n18314_, new_n18315_, new_n18316_, new_n18317_,
    new_n18318_, new_n18319_, new_n18320_, new_n18321_, new_n18322_,
    new_n18323_, new_n18324_, new_n18325_, new_n18326_, new_n18327_,
    new_n18328_, new_n18329_, new_n18330_, new_n18331_, new_n18332_,
    new_n18333_, new_n18334_, new_n18335_, new_n18336_, new_n18337_,
    new_n18338_, new_n18339_, new_n18340_, new_n18341_, new_n18342_,
    new_n18343_, new_n18344_, new_n18345_, new_n18346_, new_n18347_,
    new_n18348_, new_n18349_, new_n18350_, new_n18351_, new_n18352_,
    new_n18353_, new_n18354_, new_n18355_, new_n18356_, new_n18357_,
    new_n18358_, new_n18359_, new_n18360_, new_n18361_, new_n18362_,
    new_n18363_, new_n18364_, new_n18365_, new_n18366_, new_n18367_,
    new_n18368_, new_n18369_, new_n18370_, new_n18371_, new_n18372_,
    new_n18373_, new_n18374_, new_n18375_, new_n18376_, new_n18377_,
    new_n18378_, new_n18379_, new_n18380_, new_n18381_, new_n18382_,
    new_n18383_, new_n18384_, new_n18385_, new_n18386_, new_n18387_,
    new_n18388_, new_n18389_, new_n18390_, new_n18391_, new_n18392_,
    new_n18393_, new_n18394_, new_n18395_, new_n18396_, new_n18397_,
    new_n18398_, new_n18399_, new_n18400_, new_n18401_, new_n18402_,
    new_n18403_, new_n18404_, new_n18405_, new_n18406_, new_n18407_,
    new_n18408_, new_n18409_, new_n18410_, new_n18411_, new_n18412_,
    new_n18413_, new_n18414_, new_n18415_, new_n18416_, new_n18417_,
    new_n18418_, new_n18419_, new_n18420_, new_n18421_, new_n18422_,
    new_n18423_, new_n18424_, new_n18425_, new_n18426_, new_n18427_,
    new_n18428_, new_n18429_, new_n18430_, new_n18431_, new_n18432_,
    new_n18433_, new_n18434_, new_n18435_, new_n18436_, new_n18437_,
    new_n18438_, new_n18439_, new_n18440_, new_n18441_, new_n18442_,
    new_n18443_, new_n18444_, new_n18445_, new_n18446_, new_n18447_,
    new_n18448_, new_n18449_, new_n18450_, new_n18451_, new_n18452_,
    new_n18453_, new_n18454_, new_n18455_, new_n18456_, new_n18457_,
    new_n18458_, new_n18459_, new_n18460_, new_n18461_, new_n18462_,
    new_n18463_, new_n18464_, new_n18465_, new_n18466_, new_n18467_,
    new_n18468_, new_n18469_, new_n18470_, new_n18471_, new_n18472_,
    new_n18473_, new_n18474_, new_n18475_, new_n18476_, new_n18477_,
    new_n18478_, new_n18479_, new_n18480_, new_n18481_, new_n18482_,
    new_n18483_, new_n18484_, new_n18485_, new_n18486_, new_n18487_,
    new_n18488_, new_n18489_, new_n18490_, new_n18491_, new_n18492_,
    new_n18493_, new_n18494_, new_n18495_, new_n18496_, new_n18497_,
    new_n18498_, new_n18499_, new_n18500_, new_n18501_, new_n18502_,
    new_n18503_, new_n18504_, new_n18505_, new_n18506_, new_n18507_,
    new_n18508_, new_n18509_, new_n18510_, new_n18511_, new_n18512_,
    new_n18513_, new_n18514_, new_n18515_, new_n18516_, new_n18517_,
    new_n18518_, new_n18519_, new_n18520_, new_n18521_, new_n18522_,
    new_n18523_, new_n18524_, new_n18525_, new_n18526_, new_n18527_,
    new_n18528_, new_n18529_, new_n18530_, new_n18531_, new_n18532_,
    new_n18533_, new_n18534_, new_n18535_, new_n18536_, new_n18537_,
    new_n18538_, new_n18539_, new_n18540_, new_n18541_, new_n18542_,
    new_n18543_, new_n18544_, new_n18545_, new_n18546_, new_n18547_,
    new_n18548_, new_n18549_, new_n18550_, new_n18551_, new_n18552_,
    new_n18553_, new_n18554_, new_n18555_, new_n18556_, new_n18557_,
    new_n18558_, new_n18559_, new_n18560_, new_n18561_, new_n18562_,
    new_n18563_, new_n18564_, new_n18565_, new_n18566_, new_n18567_,
    new_n18568_, new_n18569_, new_n18570_, new_n18571_, new_n18572_,
    new_n18573_, new_n18574_, new_n18575_, new_n18576_, new_n18577_,
    new_n18578_, new_n18579_, new_n18580_, new_n18581_, new_n18582_,
    new_n18583_, new_n18584_, new_n18585_, new_n18586_, new_n18587_,
    new_n18588_, new_n18589_, new_n18590_, new_n18591_, new_n18592_,
    new_n18593_, new_n18594_, new_n18595_, new_n18596_, new_n18597_,
    new_n18598_, new_n18599_, new_n18600_, new_n18601_, new_n18602_,
    new_n18603_, new_n18604_, new_n18605_, new_n18606_, new_n18607_,
    new_n18608_, new_n18609_, new_n18610_, new_n18611_, new_n18612_,
    new_n18613_, new_n18614_, new_n18615_, new_n18616_, new_n18617_,
    new_n18618_, new_n18619_, new_n18620_, new_n18621_, new_n18622_,
    new_n18623_, new_n18624_, new_n18625_, new_n18626_, new_n18627_,
    new_n18628_, new_n18629_, new_n18630_, new_n18631_, new_n18632_,
    new_n18633_, new_n18634_, new_n18635_, new_n18636_, new_n18637_,
    new_n18638_, new_n18639_, new_n18640_, new_n18641_, new_n18642_,
    new_n18643_, new_n18644_, new_n18645_, new_n18646_, new_n18647_,
    new_n18648_, new_n18649_, new_n18650_, new_n18651_, new_n18652_,
    new_n18653_, new_n18654_, new_n18655_, new_n18656_, new_n18657_,
    new_n18658_, new_n18659_, new_n18660_, new_n18661_, new_n18662_,
    new_n18663_, new_n18664_, new_n18665_, new_n18666_, new_n18667_,
    new_n18668_, new_n18669_, new_n18670_, new_n18671_, new_n18672_,
    new_n18673_, new_n18674_, new_n18675_, new_n18676_, new_n18677_,
    new_n18678_, new_n18679_, new_n18680_, new_n18681_, new_n18682_,
    new_n18683_, new_n18684_, new_n18685_, new_n18686_, new_n18687_,
    new_n18688_, new_n18689_, new_n18690_, new_n18691_, new_n18692_,
    new_n18693_, new_n18694_, new_n18695_, new_n18696_, new_n18697_,
    new_n18698_, new_n18699_, new_n18700_, new_n18701_, new_n18702_,
    new_n18703_, new_n18704_, new_n18705_, new_n18706_, new_n18707_,
    new_n18708_, new_n18709_, new_n18710_, new_n18711_, new_n18712_,
    new_n18713_, new_n18714_, new_n18715_, new_n18716_, new_n18717_,
    new_n18718_, new_n18719_, new_n18720_, new_n18721_, new_n18722_,
    new_n18723_, new_n18724_, new_n18725_, new_n18726_, new_n18727_,
    new_n18728_, new_n18729_, new_n18730_, new_n18731_, new_n18732_,
    new_n18733_, new_n18734_, new_n18735_, new_n18736_, new_n18737_,
    new_n18738_, new_n18739_, new_n18740_, new_n18741_, new_n18742_,
    new_n18743_, new_n18744_, new_n18745_, new_n18746_, new_n18747_,
    new_n18748_, new_n18749_, new_n18750_, new_n18751_, new_n18752_,
    new_n18753_, new_n18754_, new_n18755_, new_n18756_, new_n18757_,
    new_n18758_, new_n18759_, new_n18760_, new_n18761_, new_n18762_,
    new_n18763_, new_n18764_, new_n18765_, new_n18766_, new_n18767_,
    new_n18768_, new_n18769_, new_n18770_, new_n18771_, new_n18772_,
    new_n18773_, new_n18774_, new_n18775_, new_n18776_, new_n18777_,
    new_n18778_, new_n18779_, new_n18780_, new_n18781_, new_n18782_,
    new_n18783_, new_n18784_, new_n18785_, new_n18786_, new_n18787_,
    new_n18788_, new_n18789_, new_n18790_, new_n18791_, new_n18792_,
    new_n18793_, new_n18794_, new_n18795_, new_n18796_, new_n18797_,
    new_n18798_, new_n18799_, new_n18800_, new_n18801_, new_n18802_,
    new_n18803_, new_n18804_, new_n18805_, new_n18806_, new_n18807_,
    new_n18808_, new_n18809_, new_n18810_, new_n18811_, new_n18812_,
    new_n18813_, new_n18814_, new_n18815_, new_n18816_, new_n18817_,
    new_n18818_, new_n18819_, new_n18820_, new_n18821_, new_n18822_,
    new_n18823_, new_n18824_, new_n18825_, new_n18826_, new_n18827_,
    new_n18828_, new_n18829_, new_n18830_, new_n18831_, new_n18832_,
    new_n18833_, new_n18834_, new_n18835_, new_n18836_, new_n18837_,
    new_n18838_, new_n18839_, new_n18840_, new_n18841_, new_n18842_,
    new_n18843_, new_n18844_, new_n18845_, new_n18846_, new_n18847_,
    new_n18848_, new_n18849_, new_n18850_, new_n18851_, new_n18852_,
    new_n18853_, new_n18854_, new_n18855_, new_n18856_, new_n18857_,
    new_n18858_, new_n18859_, new_n18860_, new_n18861_, new_n18862_,
    new_n18863_, new_n18864_, new_n18865_, new_n18866_, new_n18867_,
    new_n18868_, new_n18869_, new_n18870_, new_n18871_, new_n18872_,
    new_n18873_, new_n18874_, new_n18875_, new_n18876_, new_n18877_,
    new_n18878_, new_n18879_, new_n18880_, new_n18881_, new_n18882_,
    new_n18883_, new_n18884_, new_n18885_, new_n18886_, new_n18887_,
    new_n18888_, new_n18889_, new_n18890_, new_n18891_, new_n18892_,
    new_n18893_, new_n18894_, new_n18895_, new_n18896_, new_n18897_,
    new_n18898_, new_n18899_, new_n18900_, new_n18901_, new_n18902_,
    new_n18903_, new_n18904_, new_n18905_, new_n18906_, new_n18907_,
    new_n18908_, new_n18909_, new_n18910_, new_n18911_, new_n18912_,
    new_n18913_, new_n18914_, new_n18915_, new_n18916_, new_n18917_,
    new_n18918_, new_n18919_, new_n18920_, new_n18921_, new_n18922_,
    new_n18923_, new_n18924_, new_n18925_, new_n18926_, new_n18927_,
    new_n18928_, new_n18929_, new_n18930_, new_n18931_, new_n18932_,
    new_n18933_, new_n18934_, new_n18935_, new_n18936_, new_n18937_,
    new_n18938_, new_n18939_, new_n18940_, new_n18941_, new_n18942_,
    new_n18943_, new_n18944_, new_n18945_, new_n18946_, new_n18947_,
    new_n18948_, new_n18949_, new_n18950_, new_n18951_, new_n18952_,
    new_n18953_, new_n18954_, new_n18955_, new_n18956_, new_n18957_,
    new_n18958_, new_n18959_, new_n18960_, new_n18961_, new_n18962_,
    new_n18963_, new_n18964_, new_n18965_, new_n18966_, new_n18967_,
    new_n18968_, new_n18969_, new_n18970_, new_n18971_, new_n18972_,
    new_n18973_, new_n18974_, new_n18975_, new_n18976_, new_n18977_,
    new_n18978_, new_n18979_, new_n18980_, new_n18981_, new_n18982_,
    new_n18983_, new_n18984_, new_n18985_, new_n18986_, new_n18987_,
    new_n18988_, new_n18989_, new_n18990_, new_n18991_, new_n18992_,
    new_n18993_, new_n18994_, new_n18995_, new_n18996_, new_n18997_,
    new_n18998_, new_n18999_, new_n19000_, new_n19001_, new_n19002_,
    new_n19003_, new_n19004_, new_n19005_, new_n19006_, new_n19007_,
    new_n19008_, new_n19009_, new_n19010_, new_n19011_, new_n19012_,
    new_n19013_, new_n19014_, new_n19015_, new_n19016_, new_n19017_,
    new_n19018_, new_n19019_, new_n19020_, new_n19021_, new_n19022_,
    new_n19023_, new_n19024_, new_n19025_, new_n19026_, new_n19027_,
    new_n19028_, new_n19029_, new_n19030_, new_n19031_, new_n19032_,
    new_n19033_, new_n19034_, new_n19035_, new_n19036_, new_n19037_,
    new_n19038_, new_n19039_, new_n19040_, new_n19041_, new_n19042_,
    new_n19043_, new_n19044_, new_n19045_, new_n19046_, new_n19047_,
    new_n19048_, new_n19049_, new_n19050_, new_n19051_, new_n19052_,
    new_n19053_, new_n19054_, new_n19055_, new_n19056_, new_n19057_,
    new_n19058_, new_n19059_, new_n19060_, new_n19061_, new_n19062_,
    new_n19063_, new_n19064_, new_n19065_, new_n19066_, new_n19067_,
    new_n19068_, new_n19069_, new_n19070_, new_n19071_, new_n19072_,
    new_n19073_, new_n19074_, new_n19075_, new_n19076_, new_n19077_,
    new_n19078_, new_n19079_, new_n19080_, new_n19081_, new_n19082_,
    new_n19083_, new_n19084_, new_n19085_, new_n19086_, new_n19087_,
    new_n19088_, new_n19089_, new_n19090_, new_n19091_, new_n19092_,
    new_n19093_, new_n19094_, new_n19095_, new_n19096_, new_n19097_,
    new_n19098_, new_n19099_, new_n19100_, new_n19101_, new_n19102_,
    new_n19103_, new_n19104_, new_n19105_, new_n19106_, new_n19107_,
    new_n19108_, new_n19109_, new_n19110_, new_n19111_, new_n19112_,
    new_n19113_, new_n19114_, new_n19115_, new_n19116_, new_n19117_,
    new_n19118_, new_n19119_, new_n19120_, new_n19121_, new_n19122_,
    new_n19123_, new_n19124_, new_n19125_, new_n19126_, new_n19127_,
    new_n19128_, new_n19129_, new_n19130_, new_n19131_, new_n19132_,
    new_n19133_, new_n19134_, new_n19135_, new_n19136_, new_n19137_,
    new_n19138_, new_n19139_, new_n19140_, new_n19141_, new_n19142_,
    new_n19143_, new_n19144_, new_n19145_, new_n19146_, new_n19147_,
    new_n19148_, new_n19149_, new_n19150_, new_n19151_, new_n19152_,
    new_n19153_, new_n19154_, new_n19155_, new_n19156_, new_n19157_,
    new_n19158_, new_n19159_, new_n19160_, new_n19161_, new_n19162_,
    new_n19163_, new_n19164_, new_n19165_, new_n19166_, new_n19167_,
    new_n19168_, new_n19169_, new_n19170_, new_n19171_, new_n19172_,
    new_n19173_, new_n19174_, new_n19175_, new_n19176_, new_n19177_,
    new_n19178_, new_n19179_, new_n19180_, new_n19181_, new_n19182_,
    new_n19183_, new_n19184_, new_n19185_, new_n19186_, new_n19187_,
    new_n19188_, new_n19189_, new_n19190_, new_n19191_, new_n19192_,
    new_n19193_, new_n19194_, new_n19195_, new_n19196_, new_n19197_,
    new_n19198_, new_n19199_, new_n19200_, new_n19201_, new_n19202_,
    new_n19203_, new_n19204_, new_n19205_, new_n19206_, new_n19207_,
    new_n19208_, new_n19209_, new_n19210_, new_n19211_, new_n19212_,
    new_n19213_, new_n19214_, new_n19215_, new_n19216_, new_n19217_,
    new_n19218_, new_n19219_, new_n19220_, new_n19221_, new_n19222_,
    new_n19223_, new_n19224_, new_n19225_, new_n19226_, new_n19227_,
    new_n19228_, new_n19229_, new_n19230_, new_n19231_, new_n19232_,
    new_n19233_, new_n19234_, new_n19235_, new_n19236_, new_n19237_,
    new_n19238_, new_n19239_, new_n19240_, new_n19241_, new_n19242_,
    new_n19243_, new_n19244_, new_n19245_, new_n19246_, new_n19247_,
    new_n19248_, new_n19249_, new_n19250_, new_n19251_, new_n19252_,
    new_n19253_, new_n19254_, new_n19255_, new_n19256_, new_n19257_,
    new_n19258_, new_n19259_, new_n19260_, new_n19261_, new_n19262_,
    new_n19263_, new_n19264_, new_n19265_, new_n19266_, new_n19267_,
    new_n19268_, new_n19269_, new_n19270_, new_n19271_, new_n19272_,
    new_n19273_, new_n19274_, new_n19275_, new_n19276_, new_n19277_,
    new_n19278_, new_n19279_, new_n19280_, new_n19281_, new_n19282_,
    new_n19283_, new_n19284_, new_n19285_, new_n19286_, new_n19287_,
    new_n19288_, new_n19289_, new_n19290_, new_n19291_, new_n19292_,
    new_n19293_, new_n19294_, new_n19295_, new_n19296_, new_n19297_,
    new_n19298_, new_n19299_, new_n19300_, new_n19301_, new_n19302_,
    new_n19303_, new_n19304_, new_n19305_, new_n19306_, new_n19307_,
    new_n19308_, new_n19309_, new_n19310_, new_n19311_, new_n19312_,
    new_n19313_, new_n19314_, new_n19315_, new_n19316_, new_n19317_,
    new_n19318_, new_n19319_, new_n19320_, new_n19321_, new_n19322_,
    new_n19323_, new_n19324_, new_n19325_, new_n19326_, new_n19327_,
    new_n19328_, new_n19329_, new_n19330_, new_n19331_, new_n19332_,
    new_n19333_, new_n19334_, new_n19335_, new_n19336_, new_n19337_,
    new_n19338_, new_n19339_, new_n19340_, new_n19341_, new_n19342_,
    new_n19343_, new_n19344_, new_n19345_, new_n19346_, new_n19347_,
    new_n19348_, new_n19349_, new_n19350_, new_n19351_, new_n19352_,
    new_n19353_, new_n19354_, new_n19355_, new_n19356_, new_n19357_,
    new_n19358_, new_n19359_, new_n19360_, new_n19361_, new_n19362_,
    new_n19363_, new_n19364_, new_n19365_, new_n19366_, new_n19367_,
    new_n19368_, new_n19369_, new_n19370_, new_n19371_, new_n19372_,
    new_n19373_, new_n19374_, new_n19375_, new_n19376_, new_n19377_,
    new_n19378_, new_n19379_, new_n19380_, new_n19381_, new_n19382_,
    new_n19383_, new_n19384_, new_n19385_, new_n19386_, new_n19387_,
    new_n19388_, new_n19389_, new_n19390_, new_n19391_, new_n19392_,
    new_n19393_, new_n19394_, new_n19395_, new_n19396_, new_n19397_,
    new_n19398_, new_n19399_, new_n19400_, new_n19401_, new_n19402_,
    new_n19403_, new_n19404_, new_n19405_, new_n19406_, new_n19407_,
    new_n19408_, new_n19409_, new_n19410_, new_n19411_, new_n19412_,
    new_n19413_, new_n19414_, new_n19415_, new_n19416_, new_n19417_,
    new_n19418_, new_n19419_, new_n19420_, new_n19421_, new_n19422_,
    new_n19423_, new_n19424_, new_n19425_, new_n19426_, new_n19427_,
    new_n19428_, new_n19429_, new_n19430_, new_n19431_, new_n19432_,
    new_n19433_, new_n19434_, new_n19435_, new_n19436_, new_n19437_,
    new_n19438_, new_n19439_, new_n19440_, new_n19441_, new_n19442_,
    new_n19443_, new_n19444_, new_n19445_, new_n19446_, new_n19447_,
    new_n19448_, new_n19449_, new_n19450_, new_n19451_, new_n19452_,
    new_n19453_, new_n19454_, new_n19455_, new_n19456_, new_n19457_,
    new_n19458_, new_n19459_, new_n19460_, new_n19461_, new_n19462_,
    new_n19463_, new_n19464_, new_n19465_, new_n19466_, new_n19467_,
    new_n19468_, new_n19469_, new_n19470_, new_n19471_, new_n19472_,
    new_n19473_, new_n19474_, new_n19475_, new_n19476_, new_n19477_,
    new_n19478_, new_n19479_, new_n19480_, new_n19481_, new_n19482_,
    new_n19483_, new_n19484_, new_n19485_, new_n19486_, new_n19487_,
    new_n19488_, new_n19489_, new_n19490_, new_n19491_, new_n19492_,
    new_n19493_, new_n19494_, new_n19495_, new_n19496_, new_n19497_,
    new_n19498_, new_n19499_, new_n19500_, new_n19501_, new_n19502_,
    new_n19503_, new_n19504_, new_n19505_, new_n19506_, new_n19507_,
    new_n19508_, new_n19509_, new_n19510_, new_n19511_, new_n19512_,
    new_n19513_, new_n19514_, new_n19515_, new_n19516_, new_n19517_,
    new_n19518_, new_n19519_, new_n19520_, new_n19521_, new_n19522_,
    new_n19523_, new_n19524_, new_n19525_, new_n19526_, new_n19527_,
    new_n19528_, new_n19529_, new_n19530_, new_n19531_, new_n19532_,
    new_n19533_, new_n19534_, new_n19535_, new_n19536_, new_n19537_,
    new_n19538_, new_n19539_, new_n19540_, new_n19541_, new_n19542_,
    new_n19543_, new_n19544_, new_n19545_, new_n19546_, new_n19547_,
    new_n19548_, new_n19549_, new_n19550_, new_n19551_, new_n19552_,
    new_n19553_, new_n19554_, new_n19555_, new_n19556_, new_n19557_,
    new_n19558_, new_n19559_, new_n19560_, new_n19561_, new_n19562_,
    new_n19563_, new_n19564_, new_n19565_, new_n19566_, new_n19567_,
    new_n19568_, new_n19569_, new_n19570_, new_n19571_, new_n19572_,
    new_n19573_, new_n19574_, new_n19575_, new_n19576_, new_n19577_,
    new_n19578_, new_n19579_, new_n19580_, new_n19581_, new_n19582_,
    new_n19583_, new_n19584_, new_n19585_, new_n19586_, new_n19587_,
    new_n19588_, new_n19589_, new_n19590_, new_n19591_, new_n19592_,
    new_n19593_, new_n19594_, new_n19595_, new_n19596_, new_n19597_,
    new_n19598_, new_n19599_, new_n19600_, new_n19601_, new_n19602_,
    new_n19603_, new_n19604_, new_n19605_, new_n19606_, new_n19607_,
    new_n19608_, new_n19609_, new_n19610_, new_n19611_, new_n19612_,
    new_n19613_, new_n19614_, new_n19615_, new_n19616_, new_n19617_,
    new_n19618_, new_n19619_, new_n19620_, new_n19621_, new_n19622_,
    new_n19623_, new_n19624_, new_n19625_, new_n19626_, new_n19627_,
    new_n19628_, new_n19629_, new_n19630_, new_n19631_, new_n19632_,
    new_n19633_, new_n19634_, new_n19635_, new_n19636_, new_n19637_,
    new_n19638_, new_n19639_, new_n19640_, new_n19641_, new_n19642_,
    new_n19643_, new_n19644_, new_n19645_, new_n19646_, new_n19647_,
    new_n19648_, new_n19649_, new_n19650_, new_n19651_, new_n19652_,
    new_n19653_, new_n19654_, new_n19655_, new_n19656_, new_n19657_,
    new_n19658_, new_n19659_, new_n19660_, new_n19661_, new_n19662_,
    new_n19663_, new_n19664_, new_n19665_, new_n19666_, new_n19667_,
    new_n19668_, new_n19669_, new_n19670_, new_n19671_, new_n19672_,
    new_n19673_, new_n19674_, new_n19675_, new_n19676_, new_n19677_,
    new_n19678_, new_n19679_, new_n19680_, new_n19681_, new_n19682_,
    new_n19683_, new_n19684_, new_n19685_, new_n19686_, new_n19687_,
    new_n19688_, new_n19689_, new_n19690_, new_n19691_, new_n19692_,
    new_n19693_, new_n19694_, new_n19695_, new_n19696_, new_n19697_,
    new_n19698_, new_n19699_, new_n19700_, new_n19701_, new_n19702_,
    new_n19703_, new_n19704_, new_n19705_, new_n19706_, new_n19707_,
    new_n19708_, new_n19709_, new_n19710_, new_n19711_, new_n19712_,
    new_n19713_, new_n19714_, new_n19715_, new_n19716_, new_n19717_,
    new_n19718_, new_n19719_, new_n19720_, new_n19721_, new_n19722_,
    new_n19723_, new_n19724_, new_n19725_, new_n19726_, new_n19727_,
    new_n19728_, new_n19729_, new_n19730_, new_n19731_, new_n19732_,
    new_n19733_, new_n19734_, new_n19735_, new_n19736_, new_n19737_,
    new_n19738_, new_n19739_, new_n19740_, new_n19741_, new_n19742_,
    new_n19743_, new_n19744_, new_n19745_, new_n19746_, new_n19747_,
    new_n19748_, new_n19749_, new_n19750_, new_n19751_, new_n19752_,
    new_n19753_, new_n19754_, new_n19755_, new_n19756_, new_n19757_,
    new_n19758_, new_n19759_, new_n19760_, new_n19761_, new_n19762_,
    new_n19763_, new_n19764_, new_n19765_, new_n19766_, new_n19767_,
    new_n19768_, new_n19769_, new_n19770_, new_n19771_, new_n19772_,
    new_n19773_, new_n19774_, new_n19775_, new_n19776_, new_n19777_,
    new_n19778_, new_n19779_, new_n19780_, new_n19781_, new_n19782_,
    new_n19783_, new_n19784_, new_n19785_, new_n19786_, new_n19787_,
    new_n19788_, new_n19789_, new_n19790_, new_n19791_, new_n19792_,
    new_n19793_, new_n19794_, new_n19795_, new_n19796_, new_n19797_,
    new_n19798_, new_n19799_, new_n19800_, new_n19801_, new_n19802_,
    new_n19803_, new_n19804_, new_n19805_, new_n19806_, new_n19807_,
    new_n19808_, new_n19809_, new_n19810_, new_n19811_, new_n19812_,
    new_n19813_, new_n19814_, new_n19815_, new_n19816_, new_n19817_,
    new_n19818_, new_n19819_, new_n19820_, new_n19821_, new_n19822_,
    new_n19823_, new_n19824_, new_n19825_, new_n19826_, new_n19827_,
    new_n19828_, new_n19829_, new_n19830_, new_n19831_, new_n19832_,
    new_n19833_, new_n19834_, new_n19835_, new_n19836_, new_n19837_,
    new_n19838_, new_n19839_, new_n19840_, new_n19841_, new_n19842_,
    new_n19843_, new_n19844_, new_n19845_, new_n19846_, new_n19847_,
    new_n19848_, new_n19849_, new_n19850_, new_n19851_, new_n19852_,
    new_n19853_, new_n19854_, new_n19855_, new_n19856_, new_n19857_,
    new_n19858_, new_n19859_, new_n19860_, new_n19861_, new_n19862_,
    new_n19863_, new_n19864_, new_n19865_, new_n19866_, new_n19867_,
    new_n19868_, new_n19869_, new_n19870_, new_n19871_, new_n19872_,
    new_n19873_, new_n19874_, new_n19875_, new_n19876_, new_n19877_,
    new_n19878_, new_n19879_, new_n19880_, new_n19881_, new_n19882_,
    new_n19883_, new_n19884_, new_n19885_, new_n19886_, new_n19887_,
    new_n19888_, new_n19889_, new_n19890_, new_n19891_, new_n19892_,
    new_n19893_, new_n19894_, new_n19895_, new_n19896_, new_n19897_,
    new_n19898_, new_n19899_, new_n19900_, new_n19901_, new_n19902_,
    new_n19903_, new_n19904_, new_n19905_, new_n19906_, new_n19907_,
    new_n19908_, new_n19909_, new_n19910_, new_n19911_, new_n19912_,
    new_n19913_, new_n19914_, new_n19915_, new_n19916_, new_n19917_,
    new_n19918_, new_n19919_, new_n19920_, new_n19921_, new_n19922_,
    new_n19923_, new_n19924_, new_n19925_, new_n19926_, new_n19927_,
    new_n19928_, new_n19929_, new_n19930_, new_n19931_, new_n19932_,
    new_n19933_, new_n19934_, new_n19935_, new_n19936_, new_n19937_,
    new_n19938_, new_n19939_, new_n19940_, new_n19941_, new_n19942_,
    new_n19943_, new_n19944_, new_n19945_, new_n19946_, new_n19947_,
    new_n19948_, new_n19949_, new_n19950_, new_n19951_, new_n19952_,
    new_n19953_, new_n19954_, new_n19955_, new_n19956_, new_n19957_,
    new_n19958_, new_n19959_, new_n19960_, new_n19961_, new_n19962_,
    new_n19963_, new_n19964_, new_n19965_, new_n19966_, new_n19967_,
    new_n19968_, new_n19969_, new_n19970_, new_n19971_, new_n19972_,
    new_n19973_, new_n19974_, new_n19975_, new_n19976_, new_n19977_,
    new_n19978_, new_n19979_, new_n19980_, new_n19981_, new_n19982_,
    new_n19983_, new_n19984_, new_n19985_, new_n19986_, new_n19987_,
    new_n19988_, new_n19989_, new_n19990_, new_n19991_, new_n19992_,
    new_n19993_, new_n19994_, new_n19995_, new_n19996_, new_n19997_,
    new_n19998_, new_n19999_, new_n20000_, new_n20001_, new_n20002_,
    new_n20003_, new_n20004_, new_n20005_, new_n20006_, new_n20007_,
    new_n20008_, new_n20009_, new_n20010_, new_n20011_, new_n20012_,
    new_n20013_, new_n20014_, new_n20015_, new_n20016_, new_n20017_,
    new_n20018_, new_n20019_, new_n20020_, new_n20021_, new_n20022_,
    new_n20023_, new_n20024_, new_n20025_, new_n20026_, new_n20027_,
    new_n20028_, new_n20029_, new_n20030_, new_n20031_, new_n20032_,
    new_n20033_, new_n20034_, new_n20035_, new_n20036_, new_n20037_,
    new_n20038_, new_n20039_, new_n20040_, new_n20041_, new_n20042_,
    new_n20043_, new_n20044_, new_n20045_, new_n20046_, new_n20047_,
    new_n20048_, new_n20049_, new_n20050_, new_n20051_, new_n20052_,
    new_n20053_, new_n20054_, new_n20055_, new_n20056_, new_n20057_,
    new_n20058_, new_n20059_, new_n20060_, new_n20061_, new_n20062_,
    new_n20063_, new_n20064_, new_n20065_, new_n20066_, new_n20067_,
    new_n20068_, new_n20069_, new_n20070_, new_n20071_, new_n20072_,
    new_n20073_, new_n20074_, new_n20075_, new_n20076_, new_n20077_,
    new_n20078_, new_n20079_, new_n20080_, new_n20081_, new_n20082_,
    new_n20083_, new_n20084_, new_n20085_, new_n20086_, new_n20087_,
    new_n20088_, new_n20089_, new_n20090_, new_n20091_, new_n20092_,
    new_n20093_, new_n20094_, new_n20095_, new_n20096_, new_n20097_,
    new_n20098_, new_n20099_, new_n20100_, new_n20101_, new_n20102_,
    new_n20103_, new_n20104_, new_n20105_, new_n20106_, new_n20107_,
    new_n20108_, new_n20109_, new_n20110_, new_n20111_, new_n20112_,
    new_n20113_, new_n20114_, new_n20115_, new_n20116_, new_n20117_,
    new_n20118_, new_n20119_, new_n20120_, new_n20121_, new_n20122_,
    new_n20123_, new_n20124_, new_n20125_, new_n20126_, new_n20127_,
    new_n20128_, new_n20129_, new_n20130_, new_n20131_, new_n20132_,
    new_n20133_, new_n20134_, new_n20135_, new_n20136_, new_n20137_,
    new_n20138_, new_n20139_, new_n20140_, new_n20141_, new_n20142_,
    new_n20143_, new_n20144_, new_n20145_, new_n20146_, new_n20147_,
    new_n20148_, new_n20149_, new_n20150_, new_n20151_, new_n20152_,
    new_n20153_, new_n20154_, new_n20155_, new_n20156_, new_n20157_,
    new_n20158_, new_n20159_, new_n20160_, new_n20161_, new_n20162_,
    new_n20163_, new_n20164_, new_n20165_, new_n20166_, new_n20167_,
    new_n20168_, new_n20169_, new_n20170_, new_n20171_, new_n20172_,
    new_n20173_, new_n20174_, new_n20175_, new_n20176_, new_n20177_,
    new_n20178_, new_n20179_, new_n20180_, new_n20181_, new_n20182_,
    new_n20183_, new_n20184_, new_n20185_, new_n20186_, new_n20187_,
    new_n20188_, new_n20189_, new_n20190_, new_n20191_, new_n20192_,
    new_n20193_, new_n20194_, new_n20195_, new_n20196_, new_n20197_,
    new_n20198_, new_n20199_, new_n20200_, new_n20201_, new_n20202_,
    new_n20203_, new_n20204_, new_n20205_, new_n20206_, new_n20207_,
    new_n20208_, new_n20209_, new_n20210_, new_n20211_, new_n20212_,
    new_n20213_, new_n20214_, new_n20215_, new_n20216_, new_n20217_,
    new_n20218_, new_n20219_, new_n20220_, new_n20221_, new_n20222_,
    new_n20223_, new_n20224_, new_n20225_, new_n20226_, new_n20227_,
    new_n20228_, new_n20229_, new_n20230_, new_n20231_, new_n20232_,
    new_n20233_, new_n20234_, new_n20235_, new_n20236_, new_n20237_,
    new_n20238_, new_n20239_, new_n20240_, new_n20241_, new_n20242_,
    new_n20243_, new_n20244_, new_n20245_, new_n20246_, new_n20247_,
    new_n20248_, new_n20249_, new_n20250_, new_n20251_, new_n20252_,
    new_n20253_, new_n20254_, new_n20255_, new_n20256_, new_n20257_,
    new_n20258_, new_n20259_, new_n20260_, new_n20261_, new_n20262_,
    new_n20263_, new_n20264_, new_n20265_, new_n20266_, new_n20267_,
    new_n20268_, new_n20269_, new_n20270_, new_n20271_, new_n20272_,
    new_n20273_, new_n20274_, new_n20275_, new_n20276_, new_n20277_,
    new_n20278_, new_n20279_, new_n20280_, new_n20281_, new_n20282_,
    new_n20283_, new_n20284_, new_n20285_, new_n20286_, new_n20287_,
    new_n20288_, new_n20289_, new_n20290_, new_n20291_, new_n20292_,
    new_n20293_, new_n20294_, new_n20295_, new_n20296_, new_n20297_,
    new_n20298_, new_n20299_, new_n20300_, new_n20301_, new_n20302_,
    new_n20303_, new_n20304_, new_n20305_, new_n20306_, new_n20307_,
    new_n20308_, new_n20309_, new_n20310_, new_n20311_, new_n20312_,
    new_n20313_, new_n20314_, new_n20315_, new_n20316_, new_n20317_,
    new_n20318_, new_n20319_, new_n20320_, new_n20321_, new_n20322_,
    new_n20323_, new_n20324_, new_n20325_, new_n20326_, new_n20327_,
    new_n20328_, new_n20329_, new_n20330_, new_n20331_, new_n20332_,
    new_n20333_, new_n20334_, new_n20335_, new_n20336_, new_n20337_,
    new_n20338_, new_n20339_, new_n20340_, new_n20341_, new_n20342_,
    new_n20343_, new_n20344_, new_n20345_, new_n20346_, new_n20347_,
    new_n20348_, new_n20349_, new_n20350_, new_n20351_, new_n20352_,
    new_n20353_, new_n20354_, new_n20355_, new_n20356_, new_n20357_,
    new_n20358_, new_n20359_, new_n20360_, new_n20361_, new_n20362_,
    new_n20363_, new_n20364_, new_n20365_, new_n20366_, new_n20367_,
    new_n20368_, new_n20369_, new_n20370_, new_n20371_, new_n20372_,
    new_n20373_, new_n20374_, new_n20375_, new_n20376_, new_n20377_,
    new_n20378_, new_n20379_, new_n20380_, new_n20381_, new_n20382_,
    new_n20383_, new_n20384_, new_n20385_, new_n20386_, new_n20387_,
    new_n20388_, new_n20389_, new_n20390_, new_n20391_, new_n20392_,
    new_n20393_, new_n20394_, new_n20395_, new_n20396_, new_n20397_,
    new_n20398_, new_n20399_, new_n20400_, new_n20401_, new_n20402_,
    new_n20403_, new_n20404_, new_n20405_, new_n20406_, new_n20407_,
    new_n20408_, new_n20409_, new_n20410_, new_n20411_, new_n20412_,
    new_n20413_, new_n20414_, new_n20415_, new_n20416_, new_n20417_,
    new_n20418_, new_n20419_, new_n20420_, new_n20421_, new_n20422_,
    new_n20423_, new_n20424_, new_n20425_, new_n20426_, new_n20427_,
    new_n20428_, new_n20429_, new_n20430_, new_n20431_, new_n20432_,
    new_n20433_, new_n20434_, new_n20435_, new_n20436_, new_n20437_,
    new_n20438_, new_n20439_, new_n20440_, new_n20441_, new_n20442_,
    new_n20443_, new_n20444_, new_n20445_, new_n20446_, new_n20447_,
    new_n20448_, new_n20449_, new_n20450_, new_n20451_, new_n20452_,
    new_n20453_, new_n20454_, new_n20455_, new_n20456_, new_n20457_,
    new_n20458_, new_n20459_, new_n20460_, new_n20461_, new_n20462_,
    new_n20463_, new_n20464_, new_n20465_, new_n20466_, new_n20467_,
    new_n20468_, new_n20469_, new_n20470_, new_n20471_, new_n20472_,
    new_n20473_, new_n20474_, new_n20475_, new_n20476_, new_n20477_,
    new_n20478_, new_n20479_, new_n20480_, new_n20481_, new_n20482_,
    new_n20483_, new_n20484_, new_n20485_, new_n20486_, new_n20487_,
    new_n20488_, new_n20489_, new_n20490_, new_n20491_, new_n20492_,
    new_n20493_, new_n20494_, new_n20495_, new_n20496_, new_n20497_,
    new_n20498_, new_n20499_, new_n20500_, new_n20501_, new_n20502_,
    new_n20503_, new_n20504_, new_n20505_, new_n20506_, new_n20507_,
    new_n20508_, new_n20509_, new_n20510_, new_n20511_, new_n20512_,
    new_n20513_, new_n20514_, new_n20515_, new_n20516_, new_n20517_,
    new_n20518_, new_n20519_, new_n20520_, new_n20521_, new_n20522_,
    new_n20523_, new_n20524_, new_n20525_, new_n20526_, new_n20527_,
    new_n20528_, new_n20529_, new_n20530_, new_n20531_, new_n20532_,
    new_n20533_, new_n20534_, new_n20535_, new_n20536_, new_n20537_,
    new_n20538_, new_n20539_, new_n20540_, new_n20541_, new_n20542_,
    new_n20543_, new_n20544_, new_n20545_, new_n20546_, new_n20547_,
    new_n20548_, new_n20549_, new_n20550_, new_n20551_, new_n20552_,
    new_n20553_, new_n20554_, new_n20555_, new_n20556_, new_n20557_,
    new_n20558_, new_n20559_, new_n20560_, new_n20561_, new_n20562_,
    new_n20563_, new_n20564_, new_n20565_, new_n20566_, new_n20567_,
    new_n20568_, new_n20569_, new_n20570_, new_n20571_, new_n20572_,
    new_n20573_, new_n20574_, new_n20575_, new_n20576_, new_n20577_,
    new_n20578_, new_n20579_, new_n20580_, new_n20581_, new_n20582_,
    new_n20583_, new_n20584_, new_n20585_, new_n20586_, new_n20587_,
    new_n20588_, new_n20589_, new_n20590_, new_n20591_, new_n20592_,
    new_n20593_, new_n20594_, new_n20595_, new_n20596_, new_n20597_,
    new_n20598_, new_n20599_, new_n20600_, new_n20601_, new_n20602_,
    new_n20603_, new_n20604_, new_n20605_, new_n20606_, new_n20607_,
    new_n20608_, new_n20609_, new_n20610_, new_n20611_, new_n20612_,
    new_n20613_, new_n20614_, new_n20615_, new_n20616_, new_n20617_,
    new_n20618_, new_n20619_, new_n20620_, new_n20621_, new_n20622_,
    new_n20623_, new_n20624_, new_n20625_, new_n20626_, new_n20627_,
    new_n20628_, new_n20629_, new_n20630_, new_n20631_, new_n20632_,
    new_n20633_, new_n20634_, new_n20635_, new_n20636_, new_n20637_,
    new_n20638_, new_n20639_, new_n20640_, new_n20641_, new_n20642_,
    new_n20643_, new_n20644_, new_n20645_, new_n20646_, new_n20647_,
    new_n20648_, new_n20649_, new_n20650_, new_n20651_, new_n20652_,
    new_n20653_, new_n20654_, new_n20655_, new_n20656_, new_n20657_,
    new_n20658_, new_n20659_, new_n20660_, new_n20661_, new_n20662_,
    new_n20663_, new_n20664_, new_n20665_, new_n20666_, new_n20667_,
    new_n20668_, new_n20669_, new_n20670_, new_n20671_, new_n20672_,
    new_n20673_, new_n20674_, new_n20675_, new_n20676_, new_n20677_,
    new_n20678_, new_n20679_, new_n20680_, new_n20681_, new_n20682_,
    new_n20683_, new_n20684_, new_n20685_, new_n20686_, new_n20687_,
    new_n20688_, new_n20689_, new_n20690_, new_n20691_, new_n20692_,
    new_n20693_, new_n20694_, new_n20695_, new_n20696_, new_n20697_,
    new_n20698_, new_n20699_, new_n20700_, new_n20701_, new_n20702_,
    new_n20703_, new_n20704_, new_n20705_, new_n20706_, new_n20707_,
    new_n20708_, new_n20709_, new_n20710_, new_n20711_, new_n20712_,
    new_n20713_, new_n20714_, new_n20715_, new_n20716_, new_n20717_,
    new_n20718_, new_n20719_, new_n20720_, new_n20721_, new_n20722_,
    new_n20723_, new_n20724_, new_n20725_, new_n20726_, new_n20727_,
    new_n20728_, new_n20729_, new_n20730_, new_n20731_, new_n20732_,
    new_n20733_, new_n20734_, new_n20735_, new_n20736_, new_n20737_,
    new_n20738_, new_n20739_, new_n20740_, new_n20741_, new_n20742_,
    new_n20743_, new_n20744_, new_n20745_, new_n20746_, new_n20747_,
    new_n20748_, new_n20749_, new_n20750_, new_n20751_, new_n20752_,
    new_n20753_, new_n20754_, new_n20755_, new_n20756_, new_n20757_,
    new_n20758_, new_n20759_, new_n20760_, new_n20761_, new_n20762_,
    new_n20763_, new_n20764_, new_n20765_, new_n20766_, new_n20767_,
    new_n20768_, new_n20769_, new_n20770_, new_n20771_, new_n20772_,
    new_n20773_, new_n20774_, new_n20775_, new_n20776_, new_n20777_,
    new_n20778_, new_n20779_, new_n20780_, new_n20781_, new_n20782_,
    new_n20783_, new_n20784_, new_n20785_, new_n20786_, new_n20787_,
    new_n20788_, new_n20789_, new_n20790_, new_n20791_, new_n20792_,
    new_n20793_, new_n20794_, new_n20795_, new_n20796_, new_n20797_,
    new_n20798_, new_n20799_, new_n20800_, new_n20801_, new_n20802_,
    new_n20803_, new_n20804_, new_n20805_, new_n20806_, new_n20807_,
    new_n20808_, new_n20809_, new_n20810_, new_n20811_, new_n20812_,
    new_n20813_, new_n20814_, new_n20815_, new_n20816_, new_n20817_,
    new_n20818_, new_n20819_, new_n20820_, new_n20821_, new_n20822_,
    new_n20823_, new_n20824_, new_n20825_, new_n20826_, new_n20827_,
    new_n20828_, new_n20829_, new_n20830_, new_n20831_, new_n20832_,
    new_n20833_, new_n20834_, new_n20835_, new_n20836_, new_n20837_,
    new_n20838_, new_n20839_, new_n20840_, new_n20841_, new_n20842_,
    new_n20843_, new_n20844_, new_n20845_, new_n20846_, new_n20847_,
    new_n20848_, new_n20849_, new_n20850_, new_n20851_, new_n20852_,
    new_n20853_, new_n20854_, new_n20855_, new_n20856_, new_n20857_,
    new_n20858_, new_n20859_, new_n20860_, new_n20861_, new_n20862_,
    new_n20863_, new_n20864_, new_n20865_, new_n20866_, new_n20867_,
    new_n20868_, new_n20869_, new_n20870_, new_n20871_, new_n20872_,
    new_n20873_, new_n20874_, new_n20875_, new_n20876_, new_n20877_,
    new_n20878_, new_n20879_, new_n20880_, new_n20881_, new_n20882_,
    new_n20883_, new_n20884_, new_n20885_, new_n20886_, new_n20887_,
    new_n20888_, new_n20889_, new_n20890_, new_n20891_, new_n20892_,
    new_n20893_, new_n20894_, new_n20895_, new_n20896_, new_n20897_,
    new_n20898_, new_n20899_, new_n20900_, new_n20901_, new_n20902_,
    new_n20903_, new_n20904_, new_n20905_, new_n20906_, new_n20907_,
    new_n20908_, new_n20909_, new_n20910_, new_n20911_, new_n20912_,
    new_n20913_, new_n20914_, new_n20915_, new_n20916_, new_n20917_,
    new_n20918_, new_n20919_, new_n20920_, new_n20921_, new_n20922_,
    new_n20923_, new_n20924_, new_n20925_, new_n20926_, new_n20927_,
    new_n20928_, new_n20929_, new_n20930_, new_n20931_, new_n20932_,
    new_n20933_, new_n20934_, new_n20935_, new_n20936_, new_n20937_,
    new_n20938_, new_n20939_, new_n20940_, new_n20941_, new_n20942_,
    new_n20943_, new_n20944_, new_n20945_, new_n20946_, new_n20947_,
    new_n20948_, new_n20949_, new_n20950_, new_n20951_, new_n20952_,
    new_n20953_, new_n20954_, new_n20955_, new_n20956_, new_n20957_,
    new_n20958_, new_n20959_, new_n20960_, new_n20961_, new_n20962_,
    new_n20963_, new_n20964_, new_n20965_, new_n20966_, new_n20967_,
    new_n20968_, new_n20969_, new_n20970_, new_n20971_, new_n20972_,
    new_n20973_, new_n20974_, new_n20975_, new_n20976_, new_n20977_,
    new_n20978_, new_n20979_, new_n20980_, new_n20981_, new_n20982_,
    new_n20983_, new_n20984_, new_n20985_, new_n20986_, new_n20987_,
    new_n20988_, new_n20989_, new_n20990_, new_n20991_, new_n20992_,
    new_n20993_, new_n20994_, new_n20995_, new_n20996_, new_n20997_,
    new_n20998_, new_n20999_, new_n21000_, new_n21001_, new_n21002_,
    new_n21003_, new_n21004_, new_n21005_, new_n21006_, new_n21007_,
    new_n21008_, new_n21009_, new_n21010_, new_n21011_, new_n21012_,
    new_n21013_, new_n21014_, new_n21015_, new_n21016_, new_n21017_,
    new_n21018_, new_n21019_, new_n21020_, new_n21021_, new_n21022_,
    new_n21023_, new_n21024_, new_n21025_, new_n21026_, new_n21027_,
    new_n21028_, new_n21029_, new_n21030_, new_n21031_, new_n21032_,
    new_n21033_, new_n21034_, new_n21035_, new_n21036_, new_n21037_,
    new_n21038_, new_n21039_, new_n21040_, new_n21041_, new_n21042_,
    new_n21043_, new_n21044_, new_n21045_, new_n21046_, new_n21047_,
    new_n21048_, new_n21049_, new_n21050_, new_n21051_, new_n21052_,
    new_n21053_, new_n21054_, new_n21055_, new_n21056_, new_n21057_,
    new_n21058_, new_n21059_, new_n21060_, new_n21061_, new_n21062_,
    new_n21063_, new_n21064_, new_n21065_, new_n21066_, new_n21067_,
    new_n21068_, new_n21069_, new_n21070_, new_n21071_, new_n21072_,
    new_n21073_, new_n21074_, new_n21075_, new_n21076_, new_n21077_,
    new_n21078_, new_n21079_, new_n21080_, new_n21081_, new_n21082_,
    new_n21083_, new_n21084_, new_n21085_, new_n21086_, new_n21087_,
    new_n21088_, new_n21089_, new_n21090_, new_n21091_, new_n21092_,
    new_n21093_, new_n21094_, new_n21095_, new_n21096_, new_n21097_,
    new_n21098_, new_n21099_, new_n21100_, new_n21101_, new_n21102_,
    new_n21103_, new_n21104_, new_n21105_, new_n21106_, new_n21107_,
    new_n21108_, new_n21109_, new_n21110_, new_n21111_, new_n21112_,
    new_n21113_, new_n21114_, new_n21115_, new_n21116_, new_n21117_,
    new_n21118_, new_n21119_, new_n21120_, new_n21121_, new_n21122_,
    new_n21123_, new_n21124_, new_n21125_, new_n21126_, new_n21127_,
    new_n21128_, new_n21129_, new_n21130_, new_n21131_, new_n21132_,
    new_n21133_, new_n21134_, new_n21135_, new_n21136_, new_n21137_,
    new_n21138_, new_n21139_, new_n21140_, new_n21141_, new_n21142_,
    new_n21143_, new_n21144_, new_n21145_, new_n21146_, new_n21147_,
    new_n21148_, new_n21149_, new_n21150_, new_n21151_, new_n21152_,
    new_n21153_, new_n21154_, new_n21155_, new_n21156_, new_n21157_,
    new_n21158_, new_n21159_, new_n21160_, new_n21161_, new_n21162_,
    new_n21163_, new_n21164_, new_n21165_, new_n21166_, new_n21167_,
    new_n21168_, new_n21169_, new_n21170_, new_n21171_, new_n21172_,
    new_n21173_, new_n21174_, new_n21175_, new_n21176_, new_n21177_,
    new_n21178_, new_n21179_, new_n21180_, new_n21181_, new_n21182_,
    new_n21183_, new_n21184_, new_n21185_, new_n21186_, new_n21187_,
    new_n21188_, new_n21189_, new_n21190_, new_n21191_, new_n21192_,
    new_n21193_, new_n21194_, new_n21195_, new_n21196_, new_n21197_,
    new_n21198_, new_n21199_, new_n21200_, new_n21201_, new_n21202_,
    new_n21203_, new_n21204_, new_n21205_, new_n21206_, new_n21207_,
    new_n21208_, new_n21209_, new_n21210_, new_n21211_, new_n21212_,
    new_n21213_, new_n21214_, new_n21215_, new_n21216_, new_n21217_,
    new_n21218_, new_n21219_, new_n21220_, new_n21221_, new_n21222_,
    new_n21223_, new_n21224_, new_n21225_, new_n21226_, new_n21227_,
    new_n21228_, new_n21229_, new_n21230_, new_n21231_, new_n21232_,
    new_n21233_, new_n21234_, new_n21235_, new_n21236_, new_n21237_,
    new_n21238_, new_n21239_, new_n21240_, new_n21241_, new_n21242_,
    new_n21243_, new_n21244_, new_n21245_, new_n21246_, new_n21247_,
    new_n21248_, new_n21249_, new_n21250_, new_n21251_, new_n21252_,
    new_n21253_, new_n21254_, new_n21255_, new_n21256_, new_n21257_,
    new_n21258_, new_n21259_, new_n21260_, new_n21261_, new_n21262_,
    new_n21263_, new_n21264_, new_n21265_, new_n21266_, new_n21267_,
    new_n21268_, new_n21269_, new_n21270_, new_n21271_, new_n21272_,
    new_n21273_, new_n21274_, new_n21275_, new_n21276_, new_n21277_,
    new_n21278_, new_n21279_, new_n21280_, new_n21281_, new_n21282_,
    new_n21283_, new_n21284_, new_n21285_, new_n21286_, new_n21287_,
    new_n21288_, new_n21289_, new_n21290_, new_n21291_, new_n21292_,
    new_n21293_, new_n21294_, new_n21295_, new_n21296_, new_n21297_,
    new_n21298_, new_n21299_, new_n21300_, new_n21301_, new_n21302_,
    new_n21303_, new_n21304_, new_n21305_, new_n21306_, new_n21307_,
    new_n21308_, new_n21309_, new_n21310_, new_n21311_, new_n21312_,
    new_n21313_, new_n21314_, new_n21315_, new_n21316_, new_n21317_,
    new_n21318_, new_n21319_, new_n21320_, new_n21321_, new_n21322_,
    new_n21323_, new_n21324_, new_n21325_, new_n21326_, new_n21327_,
    new_n21328_, new_n21329_, new_n21330_, new_n21331_, new_n21332_,
    new_n21333_, new_n21334_, new_n21335_, new_n21336_, new_n21337_,
    new_n21338_, new_n21339_, new_n21340_, new_n21341_, new_n21342_,
    new_n21343_, new_n21344_, new_n21345_, new_n21346_, new_n21347_,
    new_n21348_, new_n21349_, new_n21350_, new_n21351_, new_n21352_,
    new_n21353_, new_n21354_, new_n21355_, new_n21356_, new_n21357_,
    new_n21358_, new_n21359_, new_n21360_, new_n21361_, new_n21362_,
    new_n21363_, new_n21364_, new_n21365_, new_n21366_, new_n21367_,
    new_n21368_, new_n21369_, new_n21370_, new_n21371_, new_n21372_,
    new_n21373_, new_n21374_, new_n21375_, new_n21376_, new_n21377_,
    new_n21378_, new_n21379_, new_n21380_, new_n21381_, new_n21382_,
    new_n21383_, new_n21384_, new_n21385_, new_n21386_, new_n21387_,
    new_n21388_, new_n21389_, new_n21390_, new_n21391_, new_n21392_,
    new_n21393_, new_n21394_, new_n21395_, new_n21396_, new_n21397_,
    new_n21398_, new_n21399_, new_n21400_, new_n21401_, new_n21402_,
    new_n21403_, new_n21404_, new_n21405_, new_n21406_, new_n21407_,
    new_n21408_, new_n21409_, new_n21410_, new_n21411_, new_n21412_,
    new_n21413_, new_n21414_, new_n21415_, new_n21416_, new_n21417_,
    new_n21418_, new_n21419_, new_n21420_, new_n21421_, new_n21422_,
    new_n21423_, new_n21424_, new_n21425_, new_n21426_, new_n21427_,
    new_n21428_, new_n21429_, new_n21430_, new_n21431_, new_n21432_,
    new_n21433_, new_n21434_, new_n21435_, new_n21436_, new_n21437_,
    new_n21438_, new_n21439_, new_n21440_, new_n21441_, new_n21442_,
    new_n21443_, new_n21444_, new_n21445_, new_n21446_, new_n21447_,
    new_n21448_, new_n21449_, new_n21450_, new_n21451_, new_n21452_,
    new_n21453_, new_n21454_, new_n21455_, new_n21456_, new_n21457_,
    new_n21458_, new_n21459_, new_n21460_, new_n21461_, new_n21462_,
    new_n21463_, new_n21464_, new_n21465_, new_n21466_, new_n21467_,
    new_n21468_, new_n21469_, new_n21470_, new_n21471_, new_n21472_,
    new_n21473_, new_n21474_, new_n21475_, new_n21476_, new_n21477_,
    new_n21478_, new_n21479_, new_n21480_, new_n21481_, new_n21482_,
    new_n21483_, new_n21484_, new_n21485_, new_n21486_, new_n21487_,
    new_n21488_, new_n21489_, new_n21490_, new_n21491_, new_n21492_,
    new_n21493_, new_n21494_, new_n21495_, new_n21496_, new_n21497_,
    new_n21498_, new_n21499_, new_n21500_, new_n21501_, new_n21502_,
    new_n21503_, new_n21504_, new_n21505_, new_n21506_, new_n21507_,
    new_n21508_, new_n21509_, new_n21510_, new_n21511_, new_n21512_,
    new_n21513_, new_n21514_, new_n21515_, new_n21516_, new_n21517_,
    new_n21518_, new_n21519_, new_n21520_, new_n21521_, new_n21522_,
    new_n21523_, new_n21524_, new_n21525_, new_n21526_, new_n21527_,
    new_n21528_, new_n21529_, new_n21530_, new_n21531_, new_n21532_,
    new_n21533_, new_n21534_, new_n21535_, new_n21536_, new_n21537_,
    new_n21538_, new_n21539_, new_n21540_, new_n21541_, new_n21542_,
    new_n21543_, new_n21544_, new_n21545_, new_n21546_, new_n21547_,
    new_n21548_, new_n21549_, new_n21550_, new_n21551_, new_n21552_,
    new_n21553_, new_n21554_, new_n21555_, new_n21556_, new_n21557_,
    new_n21558_, new_n21559_, new_n21560_, new_n21561_, new_n21562_,
    new_n21563_, new_n21564_, new_n21565_, new_n21566_, new_n21567_,
    new_n21568_, new_n21569_, new_n21570_, new_n21571_, new_n21572_,
    new_n21573_, new_n21574_, new_n21575_, new_n21576_, new_n21577_,
    new_n21578_, new_n21579_, new_n21580_, new_n21581_, new_n21582_,
    new_n21583_, new_n21584_, new_n21585_, new_n21586_, new_n21587_,
    new_n21588_, new_n21589_, new_n21590_, new_n21591_, new_n21592_,
    new_n21593_, new_n21594_, new_n21595_, new_n21596_, new_n21597_,
    new_n21598_, new_n21599_, new_n21600_, new_n21601_, new_n21602_,
    new_n21603_, new_n21604_, new_n21605_, new_n21606_, new_n21607_,
    new_n21608_, new_n21609_, new_n21610_, new_n21611_, new_n21612_,
    new_n21613_, new_n21614_, new_n21615_, new_n21616_, new_n21617_,
    new_n21618_, new_n21619_, new_n21620_, new_n21621_, new_n21622_,
    new_n21623_, new_n21624_, new_n21625_, new_n21626_, new_n21627_,
    new_n21628_, new_n21629_, new_n21630_, new_n21631_, new_n21632_,
    new_n21633_, new_n21634_, new_n21635_, new_n21636_, new_n21637_,
    new_n21638_, new_n21639_, new_n21640_, new_n21641_, new_n21642_,
    new_n21643_, new_n21644_, new_n21645_, new_n21646_, new_n21647_,
    new_n21648_, new_n21649_, new_n21650_, new_n21651_, new_n21652_,
    new_n21653_, new_n21654_, new_n21655_, new_n21656_, new_n21657_,
    new_n21658_, new_n21659_, new_n21660_, new_n21661_, new_n21662_,
    new_n21663_, new_n21664_, new_n21665_, new_n21666_, new_n21667_,
    new_n21668_, new_n21669_, new_n21670_, new_n21671_, new_n21672_,
    new_n21673_, new_n21674_, new_n21675_, new_n21676_, new_n21677_,
    new_n21678_, new_n21679_, new_n21680_, new_n21681_, new_n21682_,
    new_n21683_, new_n21684_, new_n21685_, new_n21686_, new_n21687_,
    new_n21688_, new_n21689_, new_n21690_, new_n21691_, new_n21692_,
    new_n21693_, new_n21694_, new_n21695_, new_n21696_, new_n21697_,
    new_n21698_, new_n21699_, new_n21700_, new_n21701_, new_n21702_,
    new_n21703_, new_n21704_, new_n21705_, new_n21706_, new_n21707_,
    new_n21708_, new_n21709_, new_n21710_, new_n21711_, new_n21712_,
    new_n21713_, new_n21714_, new_n21715_, new_n21716_, new_n21717_,
    new_n21718_, new_n21719_, new_n21720_, new_n21721_, new_n21722_,
    new_n21723_, new_n21724_, new_n21725_, new_n21726_, new_n21727_,
    new_n21728_, new_n21729_, new_n21730_, new_n21731_, new_n21732_,
    new_n21733_, new_n21734_, new_n21735_, new_n21736_, new_n21737_,
    new_n21738_, new_n21739_, new_n21740_, new_n21741_, new_n21742_,
    new_n21743_, new_n21744_, new_n21745_, new_n21746_, new_n21747_,
    new_n21748_, new_n21749_, new_n21750_, new_n21751_, new_n21752_,
    new_n21753_, new_n21754_, new_n21755_, new_n21756_, new_n21757_,
    new_n21758_, new_n21759_, new_n21760_, new_n21761_, new_n21762_,
    new_n21763_, new_n21764_, new_n21765_, new_n21766_, new_n21767_,
    new_n21768_, new_n21769_, new_n21770_, new_n21771_, new_n21772_,
    new_n21773_, new_n21774_, new_n21775_, new_n21776_, new_n21777_,
    new_n21778_, new_n21779_, new_n21780_, new_n21781_, new_n21782_,
    new_n21783_, new_n21784_, new_n21785_, new_n21786_, new_n21787_,
    new_n21788_, new_n21789_, new_n21790_, new_n21791_, new_n21792_,
    new_n21793_, new_n21794_, new_n21795_, new_n21796_, new_n21797_,
    new_n21798_, new_n21799_, new_n21800_, new_n21801_, new_n21802_,
    new_n21803_, new_n21804_, new_n21805_, new_n21806_, new_n21807_,
    new_n21808_, new_n21809_, new_n21810_, new_n21811_, new_n21812_,
    new_n21813_, new_n21814_, new_n21815_, new_n21816_, new_n21817_,
    new_n21818_, new_n21819_, new_n21820_, new_n21821_, new_n21822_,
    new_n21823_, new_n21824_, new_n21825_, new_n21826_, new_n21827_,
    new_n21828_, new_n21829_, new_n21830_, new_n21831_, new_n21832_,
    new_n21833_, new_n21834_, new_n21835_, new_n21836_, new_n21837_,
    new_n21838_, new_n21839_, new_n21840_, new_n21841_, new_n21842_,
    new_n21843_, new_n21844_, new_n21845_, new_n21846_, new_n21847_,
    new_n21848_, new_n21849_, new_n21850_, new_n21851_, new_n21852_,
    new_n21853_, new_n21854_, new_n21855_, new_n21856_, new_n21857_,
    new_n21858_, new_n21859_, new_n21860_, new_n21861_, new_n21862_,
    new_n21863_, new_n21864_, new_n21865_, new_n21866_, new_n21867_,
    new_n21868_, new_n21869_, new_n21870_, new_n21871_, new_n21872_,
    new_n21873_, new_n21874_, new_n21875_, new_n21876_, new_n21877_,
    new_n21878_, new_n21879_, new_n21880_, new_n21881_, new_n21882_,
    new_n21883_, new_n21884_, new_n21885_, new_n21886_, new_n21887_,
    new_n21888_, new_n21889_, new_n21890_, new_n21891_, new_n21892_,
    new_n21893_, new_n21894_, new_n21895_, new_n21896_, new_n21897_,
    new_n21898_, new_n21899_, new_n21900_, new_n21901_, new_n21902_,
    new_n21903_, new_n21904_, new_n21905_, new_n21906_, new_n21907_,
    new_n21908_, new_n21909_, new_n21910_, new_n21911_, new_n21912_,
    new_n21913_, new_n21914_, new_n21915_, new_n21916_, new_n21917_,
    new_n21918_, new_n21919_, new_n21920_, new_n21921_, new_n21922_,
    new_n21923_, new_n21924_, new_n21925_, new_n21926_, new_n21927_,
    new_n21928_, new_n21929_, new_n21930_, new_n21931_, new_n21932_,
    new_n21933_, new_n21934_, new_n21935_, new_n21936_, new_n21937_,
    new_n21938_, new_n21939_, new_n21940_, new_n21941_, new_n21942_,
    new_n21943_, new_n21944_, new_n21945_, new_n21946_, new_n21947_,
    new_n21948_, new_n21949_, new_n21950_, new_n21951_, new_n21952_,
    new_n21953_, new_n21954_, new_n21955_, new_n21956_, new_n21957_,
    new_n21958_, new_n21959_, new_n21960_, new_n21961_, new_n21962_,
    new_n21963_, new_n21964_, new_n21965_, new_n21966_, new_n21967_,
    new_n21968_, new_n21969_, new_n21970_, new_n21971_, new_n21972_,
    new_n21973_, new_n21974_, new_n21975_, new_n21976_, new_n21977_,
    new_n21978_, new_n21979_, new_n21980_, new_n21981_, new_n21982_,
    new_n21983_, new_n21984_, new_n21985_, new_n21986_, new_n21987_,
    new_n21988_, new_n21989_, new_n21990_, new_n21991_, new_n21992_,
    new_n21993_, new_n21994_, new_n21995_, new_n21996_, new_n21997_,
    new_n21998_, new_n21999_, new_n22000_, new_n22001_, new_n22002_,
    new_n22003_, new_n22004_, new_n22005_, new_n22006_, new_n22007_,
    new_n22008_, new_n22009_, new_n22010_, new_n22011_, new_n22012_,
    new_n22013_, new_n22014_, new_n22015_, new_n22016_, new_n22017_,
    new_n22018_, new_n22019_, new_n22020_, new_n22021_, new_n22022_,
    new_n22023_, new_n22024_, new_n22025_, new_n22026_, new_n22027_,
    new_n22028_, new_n22029_, new_n22030_, new_n22031_, new_n22032_,
    new_n22033_, new_n22034_, new_n22035_, new_n22036_, new_n22037_,
    new_n22038_, new_n22039_, new_n22040_, new_n22041_, new_n22042_,
    new_n22043_, new_n22044_, new_n22045_, new_n22046_, new_n22047_,
    new_n22048_, new_n22049_, new_n22050_, new_n22051_, new_n22052_,
    new_n22053_, new_n22054_, new_n22055_, new_n22056_, new_n22057_,
    new_n22058_, new_n22059_, new_n22060_, new_n22061_, new_n22062_,
    new_n22063_, new_n22064_, new_n22065_, new_n22066_, new_n22067_,
    new_n22068_, new_n22069_, new_n22070_, new_n22071_, new_n22072_,
    new_n22073_, new_n22074_, new_n22075_, new_n22076_, new_n22077_,
    new_n22078_, new_n22079_, new_n22080_, new_n22081_, new_n22082_,
    new_n22083_, new_n22084_, new_n22085_, new_n22086_, new_n22087_,
    new_n22088_, new_n22089_, new_n22090_, new_n22091_, new_n22092_,
    new_n22093_, new_n22094_, new_n22095_, new_n22096_, new_n22097_,
    new_n22098_, new_n22099_, new_n22100_, new_n22101_, new_n22102_,
    new_n22103_, new_n22104_, new_n22105_, new_n22106_, new_n22107_,
    new_n22108_, new_n22109_, new_n22110_, new_n22111_, new_n22112_,
    new_n22113_, new_n22114_, new_n22115_, new_n22116_, new_n22117_,
    new_n22118_, new_n22119_, new_n22120_, new_n22121_, new_n22122_,
    new_n22123_, new_n22124_, new_n22125_, new_n22126_, new_n22127_,
    new_n22128_, new_n22129_, new_n22130_, new_n22131_, new_n22132_,
    new_n22133_, new_n22134_, new_n22135_, new_n22136_, new_n22137_,
    new_n22138_, new_n22139_, new_n22140_, new_n22141_, new_n22142_,
    new_n22143_, new_n22144_, new_n22145_, new_n22146_, new_n22147_,
    new_n22148_, new_n22149_, new_n22150_, new_n22151_, new_n22152_,
    new_n22153_, new_n22154_, new_n22155_, new_n22156_, new_n22157_,
    new_n22158_, new_n22159_, new_n22160_, new_n22161_, new_n22162_,
    new_n22163_, new_n22164_, new_n22165_, new_n22166_, new_n22167_,
    new_n22168_, new_n22169_, new_n22170_, new_n22171_, new_n22172_,
    new_n22173_, new_n22174_, new_n22175_, new_n22176_, new_n22177_,
    new_n22178_, new_n22179_, new_n22180_, new_n22181_, new_n22182_,
    new_n22183_, new_n22184_, new_n22185_, new_n22186_, new_n22187_,
    new_n22188_, new_n22189_, new_n22190_, new_n22191_, new_n22192_,
    new_n22193_, new_n22194_, new_n22195_, new_n22196_, new_n22197_,
    new_n22198_, new_n22199_, new_n22200_, new_n22201_, new_n22202_,
    new_n22203_, new_n22204_, new_n22205_, new_n22206_, new_n22207_,
    new_n22208_, new_n22209_, new_n22210_, new_n22211_, new_n22212_,
    new_n22213_, new_n22214_, new_n22215_, new_n22216_, new_n22217_,
    new_n22218_, new_n22219_, new_n22220_, new_n22221_, new_n22222_,
    new_n22223_, new_n22224_, new_n22225_, new_n22226_, new_n22227_,
    new_n22228_, new_n22229_, new_n22230_, new_n22231_, new_n22232_,
    new_n22233_, new_n22234_, new_n22235_, new_n22236_, new_n22237_,
    new_n22238_, new_n22239_, new_n22240_, new_n22241_, new_n22242_,
    new_n22243_, new_n22244_, new_n22245_, new_n22246_, new_n22247_,
    new_n22248_, new_n22249_, new_n22250_, new_n22251_, new_n22252_,
    new_n22253_, new_n22254_, new_n22255_, new_n22256_, new_n22257_,
    new_n22258_, new_n22259_, new_n22260_, new_n22261_, new_n22262_,
    new_n22263_, new_n22264_, new_n22265_, new_n22266_, new_n22267_,
    new_n22268_, new_n22269_, new_n22270_, new_n22271_, new_n22272_,
    new_n22273_, new_n22274_, new_n22275_, new_n22276_, new_n22277_,
    new_n22278_, new_n22279_, new_n22280_, new_n22281_, new_n22282_,
    new_n22283_, new_n22284_, new_n22285_, new_n22286_, new_n22287_,
    new_n22288_, new_n22289_, new_n22290_, new_n22291_, new_n22292_,
    new_n22293_, new_n22294_, new_n22295_, new_n22296_, new_n22297_,
    new_n22298_, new_n22299_, new_n22300_, new_n22301_, new_n22302_,
    new_n22303_, new_n22304_, new_n22305_, new_n22306_, new_n22307_,
    new_n22308_, new_n22309_, new_n22310_, new_n22311_, new_n22312_,
    new_n22313_, new_n22314_, new_n22315_, new_n22316_, new_n22317_,
    new_n22318_, new_n22319_, new_n22320_, new_n22321_, new_n22322_,
    new_n22323_, new_n22324_, new_n22325_, new_n22326_, new_n22327_,
    new_n22328_, new_n22329_, new_n22330_, new_n22331_, new_n22332_,
    new_n22333_, new_n22334_, new_n22335_, new_n22336_, new_n22337_,
    new_n22338_, new_n22339_, new_n22340_, new_n22341_, new_n22342_,
    new_n22343_, new_n22344_, new_n22345_, new_n22346_, new_n22347_,
    new_n22348_, new_n22349_, new_n22350_, new_n22351_, new_n22352_,
    new_n22353_, new_n22354_, new_n22355_, new_n22356_, new_n22357_,
    new_n22358_, new_n22359_, new_n22360_, new_n22361_, new_n22362_,
    new_n22363_, new_n22364_, new_n22365_, new_n22366_, new_n22367_,
    new_n22368_, new_n22369_, new_n22370_, new_n22371_, new_n22372_,
    new_n22373_, new_n22374_, new_n22375_, new_n22376_, new_n22377_,
    new_n22378_, new_n22379_, new_n22380_, new_n22381_, new_n22382_,
    new_n22383_, new_n22384_, new_n22385_, new_n22386_, new_n22387_,
    new_n22388_, new_n22389_, new_n22390_, new_n22391_, new_n22392_,
    new_n22393_, new_n22394_, new_n22395_, new_n22396_, new_n22397_,
    new_n22398_, new_n22399_, new_n22400_, new_n22401_, new_n22402_,
    new_n22403_, new_n22404_, new_n22405_, new_n22406_, new_n22407_,
    new_n22408_, new_n22409_, new_n22410_, new_n22411_, new_n22412_,
    new_n22413_, new_n22414_, new_n22415_, new_n22416_, new_n22417_,
    new_n22418_, new_n22419_, new_n22420_, new_n22421_, new_n22422_,
    new_n22423_, new_n22424_, new_n22425_, new_n22426_, new_n22427_,
    new_n22428_, new_n22429_, new_n22430_, new_n22431_, new_n22432_,
    new_n22433_, new_n22434_, new_n22435_, new_n22436_, new_n22437_,
    new_n22438_, new_n22439_, new_n22440_, new_n22441_, new_n22442_,
    new_n22443_, new_n22444_, new_n22445_, new_n22446_, new_n22447_,
    new_n22448_, new_n22449_, new_n22450_, new_n22451_, new_n22452_,
    new_n22453_, new_n22454_, new_n22455_, new_n22456_, new_n22457_,
    new_n22458_, new_n22459_, new_n22460_, new_n22461_, new_n22462_,
    new_n22463_, new_n22464_, new_n22465_, new_n22466_, new_n22467_,
    new_n22468_, new_n22469_, new_n22470_, new_n22471_, new_n22472_,
    new_n22473_, new_n22474_, new_n22475_, new_n22476_, new_n22477_,
    new_n22478_, new_n22479_, new_n22480_, new_n22481_, new_n22482_,
    new_n22483_, new_n22484_, new_n22485_, new_n22486_, new_n22487_,
    new_n22488_, new_n22489_, new_n22490_, new_n22491_, new_n22492_,
    new_n22493_, new_n22494_, new_n22495_, new_n22496_, new_n22497_,
    new_n22498_, new_n22499_, new_n22500_, new_n22501_, new_n22502_,
    new_n22503_, new_n22504_, new_n22505_, new_n22506_, new_n22507_,
    new_n22508_, new_n22509_, new_n22510_, new_n22511_, new_n22512_,
    new_n22513_, new_n22514_, new_n22515_, new_n22516_, new_n22517_,
    new_n22518_, new_n22519_, new_n22520_, new_n22521_, new_n22522_,
    new_n22523_, new_n22524_, new_n22525_, new_n22526_, new_n22527_,
    new_n22528_, new_n22529_, new_n22530_, new_n22531_, new_n22532_,
    new_n22533_, new_n22534_, new_n22535_, new_n22536_, new_n22537_,
    new_n22538_, new_n22539_, new_n22540_, new_n22541_, new_n22542_,
    new_n22543_, new_n22544_, new_n22545_, new_n22546_, new_n22547_,
    new_n22548_, new_n22549_, new_n22550_, new_n22551_, new_n22552_,
    new_n22553_, new_n22554_, new_n22555_, new_n22556_, new_n22557_,
    new_n22558_, new_n22559_, new_n22560_, new_n22561_, new_n22562_,
    new_n22563_, new_n22564_, new_n22565_, new_n22566_, new_n22567_,
    new_n22568_, new_n22569_, new_n22570_, new_n22571_, new_n22572_,
    new_n22573_, new_n22574_, new_n22575_, new_n22576_, new_n22577_,
    new_n22578_, new_n22579_, new_n22580_, new_n22581_, new_n22582_,
    new_n22583_, new_n22584_, new_n22585_, new_n22586_, new_n22587_,
    new_n22588_, new_n22589_, new_n22590_, new_n22591_, new_n22592_,
    new_n22593_, new_n22594_, new_n22595_, new_n22596_, new_n22597_,
    new_n22598_, new_n22599_, new_n22600_, new_n22601_, new_n22602_,
    new_n22603_, new_n22604_, new_n22605_, new_n22606_, new_n22607_,
    new_n22608_, new_n22609_, new_n22610_, new_n22611_, new_n22612_,
    new_n22613_, new_n22614_, new_n22615_, new_n22616_, new_n22617_,
    new_n22618_, new_n22619_, new_n22620_, new_n22621_, new_n22622_,
    new_n22623_, new_n22624_, new_n22625_, new_n22626_, new_n22627_,
    new_n22628_, new_n22629_, new_n22630_, new_n22631_, new_n22632_,
    new_n22633_, new_n22634_, new_n22635_, new_n22636_, new_n22637_,
    new_n22638_, new_n22639_, new_n22640_, new_n22641_, new_n22642_,
    new_n22643_, new_n22644_, new_n22645_, new_n22646_, new_n22647_,
    new_n22648_, new_n22649_, new_n22650_, new_n22651_, new_n22652_,
    new_n22653_, new_n22654_, new_n22655_, new_n22656_, new_n22657_,
    new_n22658_, new_n22659_, new_n22660_, new_n22661_, new_n22662_,
    new_n22663_, new_n22664_, new_n22665_, new_n22666_, new_n22667_,
    new_n22668_, new_n22669_, new_n22670_, new_n22671_, new_n22672_,
    new_n22673_, new_n22674_, new_n22675_, new_n22676_, new_n22677_,
    new_n22678_, new_n22679_, new_n22680_, new_n22681_, new_n22682_,
    new_n22683_, new_n22684_, new_n22685_, new_n22686_, new_n22687_,
    new_n22688_, new_n22689_, new_n22690_, new_n22691_, new_n22692_,
    new_n22693_, new_n22694_, new_n22695_, new_n22696_, new_n22697_,
    new_n22698_, new_n22699_, new_n22700_, new_n22701_, new_n22702_,
    new_n22703_, new_n22704_, new_n22705_, new_n22706_, new_n22707_,
    new_n22708_, new_n22709_, new_n22710_, new_n22711_, new_n22712_,
    new_n22713_, new_n22714_, new_n22715_, new_n22716_, new_n22717_,
    new_n22718_, new_n22719_, new_n22720_, new_n22721_, new_n22722_,
    new_n22723_, new_n22724_, new_n22725_, new_n22726_, new_n22727_,
    new_n22728_, new_n22729_, new_n22730_, new_n22731_, new_n22732_,
    new_n22733_, new_n22734_, new_n22735_, new_n22736_, new_n22737_,
    new_n22738_, new_n22739_, new_n22740_, new_n22741_, new_n22742_,
    new_n22743_, new_n22744_, new_n22745_, new_n22746_, new_n22747_,
    new_n22748_, new_n22749_, new_n22750_, new_n22751_, new_n22752_,
    new_n22753_, new_n22754_, new_n22755_, new_n22756_, new_n22757_,
    new_n22758_, new_n22759_, new_n22760_, new_n22761_, new_n22762_,
    new_n22763_, new_n22764_, new_n22765_, new_n22766_, new_n22767_,
    new_n22768_, new_n22769_, new_n22770_, new_n22771_, new_n22772_,
    new_n22773_, new_n22774_, new_n22775_, new_n22776_, new_n22777_,
    new_n22778_, new_n22779_, new_n22780_, new_n22781_, new_n22782_,
    new_n22783_, new_n22784_, new_n22785_, new_n22786_, new_n22787_,
    new_n22788_, new_n22789_, new_n22790_, new_n22791_, new_n22792_,
    new_n22793_, new_n22794_, new_n22795_, new_n22796_, new_n22797_,
    new_n22798_, new_n22799_, new_n22800_, new_n22801_, new_n22802_,
    new_n22803_, new_n22804_, new_n22805_, new_n22806_, new_n22807_,
    new_n22808_, new_n22809_, new_n22810_, new_n22811_, new_n22812_,
    new_n22813_, new_n22814_, new_n22815_, new_n22816_, new_n22817_,
    new_n22818_, new_n22819_, new_n22820_, new_n22821_, new_n22822_,
    new_n22823_, new_n22824_, new_n22825_, new_n22826_, new_n22827_,
    new_n22828_, new_n22829_, new_n22830_, new_n22831_, new_n22832_,
    new_n22833_, new_n22834_, new_n22835_, new_n22836_, new_n22837_,
    new_n22838_, new_n22839_, new_n22840_, new_n22841_, new_n22842_,
    new_n22843_, new_n22844_, new_n22845_, new_n22846_, new_n22847_,
    new_n22848_, new_n22849_, new_n22850_, new_n22851_, new_n22852_,
    new_n22853_, new_n22854_, new_n22855_, new_n22856_, new_n22857_,
    new_n22858_, new_n22859_, new_n22860_, new_n22861_, new_n22862_,
    new_n22863_, new_n22864_, new_n22865_, new_n22866_, new_n22867_,
    new_n22868_, new_n22869_, new_n22870_, new_n22871_, new_n22872_,
    new_n22873_, new_n22874_, new_n22875_, new_n22876_, new_n22877_,
    new_n22878_, new_n22879_, new_n22880_, new_n22881_, new_n22882_,
    new_n22883_, new_n22884_, new_n22885_, new_n22886_, new_n22887_,
    new_n22888_, new_n22889_, new_n22890_, new_n22891_, new_n22892_,
    new_n22893_, new_n22894_, new_n22895_, new_n22896_, new_n22897_,
    new_n22898_, new_n22899_, new_n22900_, new_n22901_, new_n22902_,
    new_n22903_, new_n22904_, new_n22905_, new_n22906_, new_n22907_,
    new_n22908_, new_n22909_, new_n22910_, new_n22911_, new_n22912_,
    new_n22913_, new_n22914_, new_n22915_, new_n22916_, new_n22917_,
    new_n22918_, new_n22919_, new_n22920_, new_n22921_, new_n22922_,
    new_n22923_, new_n22924_, new_n22925_, new_n22926_, new_n22927_,
    new_n22928_, new_n22929_, new_n22930_, new_n22931_, new_n22932_,
    new_n22933_, new_n22934_, new_n22935_, new_n22936_, new_n22937_,
    new_n22938_, new_n22939_, new_n22940_, new_n22941_, new_n22942_,
    new_n22943_, new_n22944_, new_n22945_, new_n22946_, new_n22947_,
    new_n22948_, new_n22949_, new_n22950_, new_n22951_, new_n22952_,
    new_n22953_, new_n22954_, new_n22955_, new_n22956_, new_n22957_,
    new_n22958_, new_n22959_, new_n22960_, new_n22961_, new_n22962_,
    new_n22963_, new_n22964_, new_n22965_, new_n22966_, new_n22967_,
    new_n22968_, new_n22969_, new_n22970_, new_n22971_, new_n22972_,
    new_n22973_, new_n22974_, new_n22975_, new_n22976_, new_n22977_,
    new_n22978_, new_n22979_, new_n22980_, new_n22981_, new_n22982_,
    new_n22983_, new_n22984_, new_n22985_, new_n22986_, new_n22987_,
    new_n22988_, new_n22989_, new_n22990_, new_n22991_, new_n22992_,
    new_n22993_, new_n22994_, new_n22995_, new_n22996_, new_n22997_,
    new_n22998_, new_n22999_, new_n23000_, new_n23001_, new_n23002_,
    new_n23003_, new_n23004_, new_n23005_, new_n23006_, new_n23007_,
    new_n23008_, new_n23009_, new_n23010_, new_n23011_, new_n23012_,
    new_n23013_, new_n23014_, new_n23015_, new_n23016_, new_n23017_,
    new_n23018_, new_n23019_, new_n23020_, new_n23021_, new_n23022_,
    new_n23023_, new_n23024_, new_n23025_, new_n23026_, new_n23027_,
    new_n23028_, new_n23029_, new_n23030_, new_n23031_, new_n23032_,
    new_n23033_, new_n23034_, new_n23035_, new_n23036_, new_n23037_,
    new_n23038_, new_n23039_, new_n23040_, new_n23041_, new_n23042_,
    new_n23043_, new_n23044_, new_n23045_, new_n23046_, new_n23047_,
    new_n23048_, new_n23049_, new_n23050_, new_n23051_, new_n23052_,
    new_n23053_, new_n23054_, new_n23055_, new_n23056_, new_n23057_,
    new_n23058_, new_n23059_, new_n23060_, new_n23061_, new_n23062_,
    new_n23063_, new_n23064_, new_n23065_, new_n23066_, new_n23067_,
    new_n23068_, new_n23069_, new_n23070_, new_n23071_, new_n23072_,
    new_n23073_, new_n23074_, new_n23075_, new_n23076_, new_n23077_,
    new_n23078_, new_n23079_, new_n23080_, new_n23081_, new_n23082_,
    new_n23083_, new_n23084_, new_n23085_, new_n23086_, new_n23087_,
    new_n23088_, new_n23089_, new_n23090_, new_n23091_, new_n23092_,
    new_n23093_, new_n23094_, new_n23095_, new_n23096_, new_n23097_,
    new_n23098_, new_n23099_, new_n23100_, new_n23101_, new_n23102_,
    new_n23103_, new_n23104_, new_n23105_, new_n23106_, new_n23107_,
    new_n23108_, new_n23109_, new_n23110_, new_n23111_, new_n23112_,
    new_n23113_, new_n23114_, new_n23115_, new_n23116_, new_n23117_,
    new_n23118_, new_n23119_, new_n23120_, new_n23121_, new_n23122_,
    new_n23123_, new_n23124_, new_n23125_, new_n23126_, new_n23127_,
    new_n23128_, new_n23129_, new_n23130_, new_n23131_, new_n23132_,
    new_n23133_, new_n23134_, new_n23135_, new_n23136_, new_n23137_,
    new_n23138_, new_n23139_, new_n23140_, new_n23141_, new_n23142_,
    new_n23143_, new_n23144_, new_n23145_, new_n23146_, new_n23147_,
    new_n23148_, new_n23149_, new_n23150_, new_n23151_, new_n23152_,
    new_n23153_, new_n23154_, new_n23155_, new_n23156_, new_n23157_,
    new_n23158_, new_n23159_, new_n23160_, new_n23161_, new_n23162_,
    new_n23163_, new_n23164_, new_n23165_, new_n23166_, new_n23167_,
    new_n23168_, new_n23169_, new_n23170_, new_n23171_, new_n23172_,
    new_n23173_, new_n23174_, new_n23175_, new_n23176_, new_n23177_,
    new_n23178_, new_n23179_, new_n23180_, new_n23181_, new_n23182_,
    new_n23183_, new_n23184_, new_n23185_, new_n23186_, new_n23187_,
    new_n23188_, new_n23189_, new_n23190_, new_n23191_, new_n23192_,
    new_n23193_, new_n23194_, new_n23195_, new_n23196_, new_n23197_,
    new_n23198_, new_n23199_, new_n23200_, new_n23201_, new_n23202_,
    new_n23203_, new_n23204_, new_n23205_, new_n23206_, new_n23207_,
    new_n23208_, new_n23209_, new_n23210_, new_n23211_, new_n23212_,
    new_n23213_, new_n23214_, new_n23215_, new_n23216_, new_n23217_,
    new_n23218_, new_n23219_, new_n23220_, new_n23221_, new_n23222_,
    new_n23223_, new_n23224_, new_n23225_, new_n23226_, new_n23227_,
    new_n23228_, new_n23229_, new_n23230_, new_n23231_, new_n23232_,
    new_n23233_, new_n23234_, new_n23235_, new_n23236_, new_n23237_,
    new_n23238_, new_n23239_, new_n23240_, new_n23241_, new_n23242_,
    new_n23243_, new_n23244_, new_n23245_, new_n23246_, new_n23247_,
    new_n23248_, new_n23249_, new_n23250_, new_n23251_, new_n23252_,
    new_n23253_, new_n23254_, new_n23255_, new_n23256_, new_n23257_,
    new_n23258_, new_n23259_, new_n23260_, new_n23261_, new_n23262_,
    new_n23263_, new_n23264_, new_n23265_, new_n23266_, new_n23267_,
    new_n23268_, new_n23269_, new_n23270_, new_n23271_, new_n23272_,
    new_n23273_, new_n23274_, new_n23275_, new_n23276_, new_n23277_,
    new_n23278_, new_n23279_, new_n23280_, new_n23281_, new_n23282_,
    new_n23283_, new_n23284_, new_n23285_, new_n23286_, new_n23287_,
    new_n23288_, new_n23289_, new_n23290_, new_n23291_, new_n23292_,
    new_n23293_, new_n23294_, new_n23295_, new_n23296_, new_n23297_,
    new_n23298_, new_n23299_, new_n23300_, new_n23301_, new_n23302_,
    new_n23303_, new_n23304_, new_n23305_, new_n23306_, new_n23307_,
    new_n23308_, new_n23309_, new_n23310_, new_n23311_, new_n23312_,
    new_n23313_, new_n23314_, new_n23315_, new_n23316_, new_n23317_,
    new_n23318_, new_n23319_, new_n23320_, new_n23321_, new_n23322_,
    new_n23323_, new_n23324_, new_n23325_, new_n23326_, new_n23327_,
    new_n23328_, new_n23329_, new_n23330_, new_n23331_, new_n23332_,
    new_n23333_, new_n23334_, new_n23335_, new_n23336_, new_n23337_,
    new_n23338_, new_n23339_, new_n23340_, new_n23341_, new_n23342_,
    new_n23343_, new_n23344_, new_n23345_, new_n23346_, new_n23347_,
    new_n23348_, new_n23349_, new_n23350_, new_n23351_, new_n23352_,
    new_n23353_, new_n23354_, new_n23355_, new_n23356_, new_n23357_,
    new_n23358_, new_n23359_, new_n23360_, new_n23361_, new_n23362_,
    new_n23363_, new_n23364_, new_n23365_, new_n23366_, new_n23367_,
    new_n23368_, new_n23369_, new_n23370_, new_n23371_, new_n23372_,
    new_n23373_, new_n23374_, new_n23375_, new_n23376_, new_n23377_,
    new_n23378_, new_n23379_, new_n23380_, new_n23381_, new_n23382_,
    new_n23383_, new_n23384_, new_n23385_, new_n23386_, new_n23387_,
    new_n23388_, new_n23389_, new_n23390_, new_n23391_, new_n23392_,
    new_n23393_, new_n23394_, new_n23395_, new_n23396_, new_n23397_,
    new_n23398_, new_n23399_, new_n23400_, new_n23401_, new_n23402_,
    new_n23403_, new_n23404_, new_n23405_, new_n23406_, new_n23407_,
    new_n23408_, new_n23409_, new_n23410_, new_n23411_, new_n23412_,
    new_n23413_, new_n23414_, new_n23415_, new_n23416_, new_n23417_,
    new_n23418_, new_n23419_, new_n23420_, new_n23421_, new_n23422_,
    new_n23423_, new_n23424_, new_n23425_, new_n23426_, new_n23427_,
    new_n23428_, new_n23429_, new_n23430_, new_n23431_, new_n23432_,
    new_n23433_, new_n23434_, new_n23435_, new_n23436_, new_n23437_,
    new_n23438_, new_n23439_, new_n23440_, new_n23441_, new_n23442_,
    new_n23443_, new_n23444_, new_n23445_, new_n23446_, new_n23447_,
    new_n23448_, new_n23449_, new_n23450_, new_n23451_, new_n23452_,
    new_n23453_, new_n23454_, new_n23455_, new_n23456_, new_n23457_,
    new_n23458_, new_n23459_, new_n23460_, new_n23461_, new_n23462_,
    new_n23463_, new_n23464_, new_n23465_, new_n23466_, new_n23467_,
    new_n23468_, new_n23469_, new_n23470_, new_n23471_, new_n23472_,
    new_n23473_, new_n23474_, new_n23475_, new_n23476_, new_n23477_,
    new_n23478_, new_n23479_, new_n23480_, new_n23481_, new_n23482_,
    new_n23483_, new_n23484_, new_n23485_, new_n23486_, new_n23487_,
    new_n23488_, new_n23489_, new_n23490_, new_n23491_, new_n23492_,
    new_n23493_, new_n23494_, new_n23495_, new_n23496_, new_n23497_,
    new_n23498_, new_n23499_, new_n23500_, new_n23501_, new_n23502_,
    new_n23503_, new_n23504_, new_n23505_, new_n23506_, new_n23507_,
    new_n23508_, new_n23509_, new_n23510_, new_n23511_, new_n23512_,
    new_n23513_, new_n23514_, new_n23515_, new_n23516_, new_n23517_,
    new_n23518_, new_n23519_, new_n23520_, new_n23521_, new_n23522_,
    new_n23523_, new_n23524_, new_n23525_, new_n23526_, new_n23527_,
    new_n23528_, new_n23529_, new_n23530_, new_n23531_, new_n23532_,
    new_n23533_, new_n23534_, new_n23535_, new_n23536_, new_n23537_,
    new_n23538_, new_n23539_, new_n23540_, new_n23541_, new_n23542_,
    new_n23543_, new_n23544_, new_n23545_, new_n23546_, new_n23547_,
    new_n23548_, new_n23549_, new_n23550_, new_n23551_, new_n23552_,
    new_n23553_, new_n23554_, new_n23555_, new_n23556_, new_n23557_,
    new_n23558_, new_n23559_, new_n23560_, new_n23561_, new_n23562_,
    new_n23563_, new_n23564_, new_n23565_, new_n23566_, new_n23567_,
    new_n23568_, new_n23569_, new_n23570_, new_n23571_, new_n23572_,
    new_n23573_, new_n23574_, new_n23575_, new_n23576_, new_n23577_,
    new_n23578_, new_n23579_, new_n23580_, new_n23581_, new_n23582_,
    new_n23583_, new_n23584_, new_n23585_, new_n23586_, new_n23587_,
    new_n23588_, new_n23589_, new_n23590_, new_n23591_, new_n23592_,
    new_n23593_, new_n23594_, new_n23595_, new_n23596_, new_n23597_,
    new_n23598_, new_n23599_, new_n23600_, new_n23601_, new_n23602_,
    new_n23603_, new_n23604_, new_n23605_, new_n23606_, new_n23607_,
    new_n23608_, new_n23609_, new_n23610_, new_n23611_, new_n23612_,
    new_n23613_, new_n23614_, new_n23615_, new_n23616_, new_n23617_,
    new_n23618_, new_n23619_, new_n23620_, new_n23621_, new_n23622_,
    new_n23623_, new_n23624_, new_n23625_, new_n23626_, new_n23627_,
    new_n23628_, new_n23629_, new_n23630_, new_n23631_, new_n23632_,
    new_n23633_, new_n23634_, new_n23635_, new_n23636_, new_n23637_,
    new_n23638_, new_n23639_, new_n23640_, new_n23641_, new_n23642_,
    new_n23643_, new_n23644_, new_n23645_, new_n23646_, new_n23647_,
    new_n23648_, new_n23649_, new_n23650_, new_n23651_, new_n23652_,
    new_n23653_, new_n23654_, new_n23655_, new_n23656_, new_n23657_,
    new_n23658_, new_n23659_, new_n23660_, new_n23661_, new_n23662_,
    new_n23663_, new_n23664_, new_n23665_, new_n23666_, new_n23667_,
    new_n23668_, new_n23669_, new_n23670_, new_n23671_, new_n23672_,
    new_n23673_, new_n23674_, new_n23675_, new_n23676_, new_n23677_,
    new_n23678_, new_n23679_, new_n23680_, new_n23681_, new_n23682_,
    new_n23683_, new_n23684_, new_n23685_, new_n23686_, new_n23687_,
    new_n23688_, new_n23689_, new_n23690_, new_n23691_, new_n23692_,
    new_n23693_, new_n23694_, new_n23695_, new_n23696_, new_n23697_,
    new_n23698_, new_n23699_, new_n23700_, new_n23701_, new_n23702_,
    new_n23703_, new_n23704_, new_n23705_, new_n23706_, new_n23707_,
    new_n23708_, new_n23709_, new_n23710_, new_n23711_, new_n23712_,
    new_n23713_, new_n23714_, new_n23715_, new_n23716_, new_n23717_,
    new_n23718_, new_n23719_, new_n23720_, new_n23721_, new_n23722_,
    new_n23723_, new_n23724_, new_n23725_, new_n23726_, new_n23727_,
    new_n23728_, new_n23729_, new_n23730_, new_n23731_, new_n23732_,
    new_n23733_, new_n23734_, new_n23735_, new_n23736_, new_n23737_,
    new_n23738_, new_n23739_, new_n23740_, new_n23741_, new_n23742_,
    new_n23743_, new_n23744_, new_n23745_, new_n23746_, new_n23747_,
    new_n23748_, new_n23749_, new_n23750_, new_n23751_, new_n23752_,
    new_n23753_, new_n23754_, new_n23755_, new_n23756_, new_n23757_,
    new_n23758_, new_n23759_, new_n23760_, new_n23761_, new_n23762_,
    new_n23763_, new_n23764_, new_n23765_, new_n23766_, new_n23767_,
    new_n23768_, new_n23769_, new_n23770_, new_n23771_, new_n23772_,
    new_n23773_, new_n23774_, new_n23775_, new_n23776_, new_n23777_,
    new_n23778_, new_n23779_, new_n23780_, new_n23781_, new_n23782_,
    new_n23783_, new_n23784_, new_n23785_, new_n23786_, new_n23787_,
    new_n23788_, new_n23789_, new_n23790_, new_n23791_, new_n23792_,
    new_n23793_, new_n23794_, new_n23795_, new_n23796_, new_n23797_,
    new_n23798_, new_n23799_, new_n23800_, new_n23801_, new_n23802_,
    new_n23803_, new_n23804_, new_n23805_, new_n23806_, new_n23807_,
    new_n23808_, new_n23809_, new_n23810_, new_n23811_, new_n23812_,
    new_n23813_, new_n23814_, new_n23815_, new_n23816_, new_n23817_,
    new_n23818_, new_n23819_, new_n23820_, new_n23821_, new_n23822_,
    new_n23823_, new_n23824_, new_n23825_, new_n23826_, new_n23827_,
    new_n23828_, new_n23829_, new_n23830_, new_n23831_, new_n23832_,
    new_n23833_, new_n23834_, new_n23835_, new_n23836_, new_n23837_,
    new_n23838_, new_n23839_, new_n23840_, new_n23841_, new_n23842_,
    new_n23843_, new_n23844_, new_n23845_, new_n23846_, new_n23847_,
    new_n23848_, new_n23849_, new_n23850_, new_n23851_, new_n23852_,
    new_n23853_, new_n23854_, new_n23855_, new_n23856_, new_n23857_,
    new_n23858_, new_n23859_, new_n23860_, new_n23861_, new_n23862_,
    new_n23863_, new_n23864_, new_n23865_, new_n23866_, new_n23867_,
    new_n23868_, new_n23869_, new_n23870_, new_n23871_, new_n23872_,
    new_n23873_, new_n23874_, new_n23875_, new_n23876_, new_n23877_,
    new_n23878_, new_n23879_, new_n23880_, new_n23881_, new_n23882_,
    new_n23883_, new_n23884_, new_n23885_, new_n23886_, new_n23887_,
    new_n23888_, new_n23889_, new_n23890_, new_n23891_, new_n23892_,
    new_n23893_, new_n23894_, new_n23895_, new_n23896_, new_n23897_,
    new_n23898_, new_n23899_, new_n23900_, new_n23901_, new_n23902_,
    new_n23903_, new_n23904_, new_n23905_, new_n23906_, new_n23907_,
    new_n23908_, new_n23909_, new_n23910_, new_n23911_, new_n23912_,
    new_n23913_, new_n23914_, new_n23915_, new_n23916_, new_n23917_,
    new_n23918_, new_n23919_, new_n23920_, new_n23921_, new_n23922_,
    new_n23923_, new_n23924_, new_n23925_, new_n23926_, new_n23927_,
    new_n23928_, new_n23929_, new_n23930_, new_n23931_, new_n23932_,
    new_n23933_, new_n23934_, new_n23935_, new_n23936_, new_n23937_,
    new_n23938_, new_n23939_, new_n23940_, new_n23941_, new_n23942_,
    new_n23943_, new_n23944_, new_n23945_, new_n23946_, new_n23947_,
    new_n23948_, new_n23949_, new_n23950_, new_n23951_, new_n23952_,
    new_n23953_, new_n23954_, new_n23955_, new_n23956_, new_n23957_,
    new_n23958_, new_n23959_, new_n23960_, new_n23961_, new_n23962_,
    new_n23963_, new_n23964_, new_n23965_, new_n23966_, new_n23967_,
    new_n23968_, new_n23969_, new_n23970_, new_n23971_, new_n23972_,
    new_n23973_, new_n23974_, new_n23975_, new_n23976_, new_n23977_,
    new_n23978_, new_n23979_, new_n23980_, new_n23981_, new_n23982_,
    new_n23983_, new_n23984_, new_n23985_, new_n23986_, new_n23987_,
    new_n23988_, new_n23989_, new_n23990_, new_n23991_, new_n23992_,
    new_n23993_, new_n23994_, new_n23995_, new_n23996_, new_n23997_,
    new_n23998_, new_n23999_, new_n24000_, new_n24001_, new_n24002_,
    new_n24003_, new_n24004_, new_n24005_, new_n24006_, new_n24007_,
    new_n24008_, new_n24009_, new_n24010_, new_n24011_, new_n24012_,
    new_n24013_, new_n24014_, new_n24015_, new_n24016_, new_n24017_,
    new_n24018_, new_n24019_, new_n24020_, new_n24021_, new_n24022_,
    new_n24023_, new_n24024_, new_n24025_, new_n24026_, new_n24027_,
    new_n24028_, new_n24029_, new_n24030_, new_n24031_, new_n24032_,
    new_n24033_, new_n24034_, new_n24035_, new_n24036_, new_n24037_,
    new_n24038_, new_n24039_, new_n24040_, new_n24041_, new_n24042_,
    new_n24043_, new_n24044_, new_n24045_, new_n24046_, new_n24047_,
    new_n24048_, new_n24049_, new_n24050_, new_n24051_, new_n24052_,
    new_n24053_, new_n24054_, new_n24055_, new_n24056_, new_n24057_,
    new_n24058_, new_n24059_, new_n24060_, new_n24061_, new_n24062_,
    new_n24063_, new_n24064_, new_n24065_, new_n24066_, new_n24067_,
    new_n24068_, new_n24069_, new_n24070_, new_n24071_, new_n24072_,
    new_n24073_, new_n24074_, new_n24075_, new_n24076_, new_n24077_,
    new_n24078_, new_n24079_, new_n24080_, new_n24081_, new_n24082_,
    new_n24083_, new_n24084_, new_n24085_, new_n24086_, new_n24087_,
    new_n24088_, new_n24089_, new_n24090_, new_n24091_, new_n24092_,
    new_n24093_, new_n24094_, new_n24095_, new_n24096_, new_n24097_,
    new_n24098_, new_n24099_, new_n24100_, new_n24101_, new_n24102_,
    new_n24103_, new_n24104_, new_n24105_, new_n24106_, new_n24107_,
    new_n24108_, new_n24109_, new_n24110_, new_n24111_, new_n24112_,
    new_n24113_, new_n24114_, new_n24115_, new_n24116_, new_n24117_,
    new_n24118_, new_n24119_, new_n24120_, new_n24121_, new_n24122_,
    new_n24123_, new_n24124_, new_n24125_, new_n24126_, new_n24127_,
    new_n24128_, new_n24129_, new_n24130_, new_n24131_, new_n24132_,
    new_n24133_, new_n24134_, new_n24135_, new_n24136_, new_n24137_,
    new_n24138_, new_n24139_, new_n24140_, new_n24141_, new_n24142_,
    new_n24143_, new_n24144_, new_n24145_, new_n24146_, new_n24147_,
    new_n24148_, new_n24149_, new_n24150_, new_n24151_, new_n24152_,
    new_n24153_, new_n24154_, new_n24155_, new_n24156_, new_n24157_,
    new_n24158_, new_n24159_, new_n24160_, new_n24161_, new_n24162_,
    new_n24163_, new_n24164_, new_n24165_, new_n24166_, new_n24167_,
    new_n24168_, new_n24169_, new_n24170_, new_n24171_, new_n24172_,
    new_n24173_, new_n24174_, new_n24175_, new_n24176_, new_n24177_,
    new_n24178_, new_n24179_, new_n24180_, new_n24181_, new_n24182_,
    new_n24183_, new_n24184_, new_n24185_, new_n24186_, new_n24187_,
    new_n24188_, new_n24189_, new_n24190_, new_n24191_, new_n24192_,
    new_n24193_, new_n24194_, new_n24195_, new_n24196_, new_n24197_,
    new_n24198_, new_n24199_, new_n24200_, new_n24201_, new_n24202_,
    new_n24203_, new_n24204_, new_n24205_, new_n24206_, new_n24207_,
    new_n24208_, new_n24209_, new_n24210_, new_n24211_, new_n24212_,
    new_n24213_, new_n24214_, new_n24215_, new_n24216_, new_n24217_,
    new_n24218_, new_n24219_, new_n24220_, new_n24221_, new_n24222_,
    new_n24223_, new_n24224_, new_n24225_, new_n24226_, new_n24227_,
    new_n24228_, new_n24229_, new_n24230_, new_n24231_, new_n24232_,
    new_n24233_, new_n24234_, new_n24235_, new_n24236_, new_n24237_,
    new_n24238_, new_n24239_, new_n24240_, new_n24241_, new_n24242_,
    new_n24243_, new_n24244_, new_n24245_, new_n24246_, new_n24247_,
    new_n24248_, new_n24249_, new_n24250_, new_n24251_, new_n24252_,
    new_n24253_, new_n24254_, new_n24255_, new_n24256_, new_n24257_,
    new_n24258_, new_n24259_, new_n24260_, new_n24261_, new_n24262_,
    new_n24263_, new_n24264_, new_n24265_, new_n24266_, new_n24267_,
    new_n24268_, new_n24269_, new_n24270_, new_n24271_, new_n24272_,
    new_n24273_, new_n24274_, new_n24275_, new_n24276_, new_n24277_,
    new_n24278_, new_n24279_, new_n24280_, new_n24281_, new_n24282_,
    new_n24283_, new_n24284_, new_n24285_, new_n24286_, new_n24287_,
    new_n24288_, new_n24289_, new_n24290_, new_n24291_, new_n24292_,
    new_n24293_, new_n24294_, new_n24295_, new_n24296_, new_n24297_,
    new_n24298_, new_n24299_, new_n24300_, new_n24301_, new_n24302_,
    new_n24303_, new_n24304_, new_n24305_, new_n24306_, new_n24307_,
    new_n24308_, new_n24309_, new_n24310_, new_n24311_, new_n24312_,
    new_n24313_, new_n24314_, new_n24315_, new_n24316_, new_n24317_,
    new_n24318_, new_n24319_, new_n24320_, new_n24321_, new_n24322_,
    new_n24323_, new_n24324_, new_n24325_, new_n24326_, new_n24327_,
    new_n24328_, new_n24329_, new_n24330_, new_n24331_, new_n24332_,
    new_n24333_, new_n24334_, new_n24335_, new_n24336_, new_n24337_,
    new_n24338_, new_n24339_, new_n24340_, new_n24341_, new_n24342_,
    new_n24343_, new_n24344_, new_n24345_, new_n24346_, new_n24347_,
    new_n24348_, new_n24349_, new_n24350_, new_n24351_, new_n24352_,
    new_n24353_, new_n24354_, new_n24355_, new_n24356_, new_n24357_,
    new_n24358_, new_n24359_, new_n24360_, new_n24361_, new_n24362_,
    new_n24363_, new_n24364_, new_n24365_, new_n24366_, new_n24367_,
    new_n24368_, new_n24369_, new_n24370_, new_n24371_, new_n24372_,
    new_n24373_, new_n24374_, new_n24375_, new_n24376_, new_n24377_,
    new_n24378_, new_n24379_, new_n24380_, new_n24381_, new_n24382_,
    new_n24383_, new_n24384_, new_n24385_, new_n24386_, new_n24387_,
    new_n24388_, new_n24389_, new_n24390_, new_n24391_, new_n24392_,
    new_n24393_, new_n24394_, new_n24395_, new_n24396_, new_n24397_,
    new_n24398_, new_n24399_, new_n24400_, new_n24401_, new_n24402_,
    new_n24403_, new_n24404_, new_n24405_, new_n24406_, new_n24407_,
    new_n24408_, new_n24409_, new_n24410_, new_n24411_, new_n24412_,
    new_n24413_, new_n24414_, new_n24415_, new_n24416_, new_n24417_,
    new_n24418_, new_n24419_, new_n24420_, new_n24421_, new_n24422_,
    new_n24423_, new_n24424_, new_n24425_, new_n24426_, new_n24427_,
    new_n24428_, new_n24429_, new_n24430_, new_n24431_, new_n24432_,
    new_n24433_, new_n24434_, new_n24435_, new_n24436_, new_n24437_,
    new_n24438_, new_n24439_, new_n24440_, new_n24441_, new_n24442_,
    new_n24443_, new_n24444_, new_n24445_, new_n24446_, new_n24447_,
    new_n24448_, new_n24449_, new_n24450_, new_n24451_, new_n24452_,
    new_n24453_, new_n24454_, new_n24455_, new_n24456_, new_n24457_,
    new_n24458_, new_n24459_, new_n24460_, new_n24461_, new_n24462_,
    new_n24463_, new_n24464_, new_n24465_, new_n24466_, new_n24467_,
    new_n24468_, new_n24469_, new_n24470_, new_n24471_, new_n24472_,
    new_n24473_, new_n24474_, new_n24475_, new_n24476_, new_n24477_,
    new_n24478_, new_n24479_, new_n24480_, new_n24481_, new_n24482_,
    new_n24483_, new_n24484_, new_n24485_, new_n24486_, new_n24487_,
    new_n24488_, new_n24489_, new_n24490_, new_n24491_, new_n24492_,
    new_n24493_, new_n24494_, new_n24495_, new_n24496_, new_n24497_,
    new_n24498_, new_n24499_, new_n24500_, new_n24501_, new_n24502_,
    new_n24503_, new_n24504_, new_n24505_, new_n24506_, new_n24507_,
    new_n24508_, new_n24509_, new_n24510_, new_n24511_, new_n24512_,
    new_n24513_, new_n24514_, new_n24515_, new_n24516_, new_n24517_,
    new_n24518_, new_n24519_, new_n24520_, new_n24521_, new_n24522_,
    new_n24523_, new_n24524_, new_n24525_, new_n24526_, new_n24527_,
    new_n24528_, new_n24529_, new_n24530_, new_n24531_, new_n24532_,
    new_n24533_, new_n24534_, new_n24535_, new_n24536_, new_n24537_,
    new_n24538_, new_n24539_, new_n24540_, new_n24541_, new_n24542_,
    new_n24543_, new_n24544_, new_n24545_, new_n24546_, new_n24547_,
    new_n24548_, new_n24549_, new_n24550_, new_n24551_, new_n24552_,
    new_n24553_, new_n24554_, new_n24555_, new_n24556_, new_n24557_,
    new_n24558_, new_n24559_, new_n24560_, new_n24561_, new_n24562_,
    new_n24563_, new_n24564_, new_n24565_, new_n24566_, new_n24567_,
    new_n24568_, new_n24569_, new_n24570_, new_n24571_, new_n24572_,
    new_n24573_, new_n24574_, new_n24575_, new_n24576_, new_n24577_,
    new_n24578_, new_n24579_, new_n24580_, new_n24581_, new_n24582_,
    new_n24583_, new_n24584_, new_n24585_, new_n24586_, new_n24587_,
    new_n24588_, new_n24589_, new_n24590_, new_n24591_, new_n24592_,
    new_n24593_, new_n24594_, new_n24595_, new_n24596_, new_n24597_,
    new_n24598_, new_n24599_, new_n24600_, new_n24601_, new_n24602_,
    new_n24603_, new_n24604_, new_n24605_, new_n24606_, new_n24607_,
    new_n24608_, new_n24609_, new_n24610_, new_n24611_, new_n24612_,
    new_n24613_, new_n24614_, new_n24615_, new_n24616_, new_n24617_,
    new_n24618_, new_n24619_, new_n24620_, new_n24621_, new_n24622_,
    new_n24623_, new_n24624_, new_n24625_, new_n24626_, new_n24627_,
    new_n24628_, new_n24629_, new_n24630_, new_n24631_, new_n24632_,
    new_n24633_, new_n24634_, new_n24635_, new_n24636_, new_n24637_,
    new_n24638_, new_n24639_, new_n24640_, new_n24641_, new_n24642_,
    new_n24643_, new_n24644_, new_n24645_, new_n24646_, new_n24647_,
    new_n24648_, new_n24649_, new_n24650_, new_n24651_, new_n24652_,
    new_n24653_, new_n24654_, new_n24655_, new_n24656_, new_n24657_,
    new_n24658_, new_n24659_, new_n24660_, new_n24661_, new_n24662_,
    new_n24663_, new_n24664_, new_n24665_, new_n24666_, new_n24667_,
    new_n24668_, new_n24669_, new_n24670_, new_n24671_, new_n24672_,
    new_n24673_, new_n24674_, new_n24675_, new_n24676_, new_n24677_,
    new_n24678_, new_n24679_, new_n24680_, new_n24681_, new_n24682_,
    new_n24683_, new_n24684_, new_n24685_, new_n24686_, new_n24687_,
    new_n24688_, new_n24689_, new_n24690_, new_n24691_, new_n24692_,
    new_n24693_, new_n24694_, new_n24695_, new_n24696_, new_n24697_,
    new_n24698_, new_n24699_, new_n24700_, new_n24701_, new_n24702_,
    new_n24703_, new_n24704_, new_n24705_, new_n24706_, new_n24707_,
    new_n24708_, new_n24709_, new_n24710_, new_n24711_, new_n24712_,
    new_n24713_, new_n24714_, new_n24715_, new_n24716_, new_n24717_,
    new_n24718_, new_n24719_, new_n24720_, new_n24721_, new_n24722_,
    new_n24723_, new_n24724_, new_n24725_, new_n24726_, new_n24727_,
    new_n24728_, new_n24729_, new_n24730_, new_n24731_, new_n24732_,
    new_n24733_, new_n24734_, new_n24735_, new_n24736_, new_n24737_,
    new_n24738_, new_n24739_, new_n24740_, new_n24741_, new_n24742_,
    new_n24743_, new_n24744_, new_n24745_, new_n24746_, new_n24747_,
    new_n24748_, new_n24749_, new_n24750_, new_n24751_, new_n24752_,
    new_n24753_, new_n24754_, new_n24755_, new_n24756_, new_n24757_,
    new_n24758_, new_n24759_, new_n24760_, new_n24761_, new_n24762_,
    new_n24763_, new_n24764_, new_n24765_, new_n24766_, new_n24767_,
    new_n24768_, new_n24769_, new_n24770_, new_n24771_, new_n24772_,
    new_n24773_, new_n24774_, new_n24775_, new_n24776_, new_n24777_,
    new_n24778_, new_n24779_, new_n24780_, new_n24781_, new_n24782_,
    new_n24783_, new_n24784_, new_n24785_, new_n24786_, new_n24787_,
    new_n24788_, new_n24789_, new_n24790_, new_n24791_, new_n24792_,
    new_n24793_, new_n24794_, new_n24795_, new_n24796_, new_n24797_,
    new_n24798_, new_n24799_, new_n24800_, new_n24801_, new_n24802_,
    new_n24803_, new_n24804_, new_n24805_, new_n24806_, new_n24807_,
    new_n24808_, new_n24809_, new_n24810_, new_n24811_, new_n24812_,
    new_n24813_, new_n24814_, new_n24815_, new_n24816_, new_n24817_,
    new_n24818_, new_n24819_, new_n24820_, new_n24821_, new_n24822_,
    new_n24823_, new_n24824_, new_n24825_, new_n24826_, new_n24827_,
    new_n24828_, new_n24829_, new_n24830_, new_n24831_, new_n24832_,
    new_n24833_, new_n24834_, new_n24835_, new_n24836_, new_n24837_,
    new_n24838_, new_n24839_, new_n24840_, new_n24841_, new_n24842_,
    new_n24843_, new_n24844_, new_n24845_, new_n24846_, new_n24847_,
    new_n24848_, new_n24849_, new_n24850_, new_n24851_, new_n24852_,
    new_n24853_, new_n24854_, new_n24855_, new_n24856_, new_n24857_,
    new_n24858_, new_n24859_, new_n24860_, new_n24861_, new_n24862_,
    new_n24863_, new_n24864_, new_n24865_, new_n24866_, new_n24867_,
    new_n24868_, new_n24869_, new_n24870_, new_n24871_, new_n24872_,
    new_n24873_, new_n24874_, new_n24875_, new_n24876_, new_n24877_,
    new_n24878_, new_n24879_, new_n24880_, new_n24881_, new_n24882_,
    new_n24883_, new_n24884_, new_n24885_, new_n24886_, new_n24887_,
    new_n24888_, new_n24889_, new_n24890_, new_n24891_, new_n24892_,
    new_n24893_, new_n24894_, new_n24895_, new_n24896_, new_n24897_,
    new_n24898_, new_n24899_, new_n24900_, new_n24901_, new_n24902_,
    new_n24903_, new_n24904_, new_n24905_, new_n24906_, new_n24907_,
    new_n24908_, new_n24909_, new_n24910_, new_n24911_, new_n24912_,
    new_n24913_, new_n24914_, new_n24915_, new_n24916_, new_n24917_,
    new_n24918_, new_n24919_, new_n24920_, new_n24921_, new_n24922_,
    new_n24923_, new_n24924_, new_n24925_, new_n24926_, new_n24927_,
    new_n24928_, new_n24929_, new_n24930_, new_n24931_, new_n24932_,
    new_n24933_, new_n24934_, new_n24935_, new_n24936_, new_n24937_,
    new_n24938_, new_n24939_, new_n24940_, new_n24941_, new_n24942_,
    new_n24943_, new_n24944_, new_n24945_, new_n24946_, new_n24947_,
    new_n24948_, new_n24949_, new_n24950_, new_n24951_, new_n24952_,
    new_n24953_, new_n24954_, new_n24955_, new_n24956_, new_n24957_,
    new_n24958_, new_n24959_, new_n24960_, new_n24961_, new_n24962_,
    new_n24963_, new_n24964_, new_n24965_, new_n24966_, new_n24967_,
    new_n24968_, new_n24969_, new_n24970_, new_n24971_, new_n24972_,
    new_n24973_, new_n24974_, new_n24975_, new_n24976_, new_n24977_,
    new_n24978_, new_n24979_, new_n24980_, new_n24981_, new_n24982_,
    new_n24983_, new_n24984_, new_n24985_, new_n24986_, new_n24987_,
    new_n24988_, new_n24989_, new_n24990_, new_n24991_, new_n24992_,
    new_n24993_, new_n24994_, new_n24995_, new_n24996_, new_n24997_,
    new_n24998_, new_n24999_, new_n25000_, new_n25001_, new_n25002_,
    new_n25003_, new_n25004_, new_n25005_, new_n25006_, new_n25007_,
    new_n25008_, new_n25009_, new_n25010_, new_n25011_, new_n25012_,
    new_n25013_, new_n25014_, new_n25015_, new_n25016_, new_n25017_,
    new_n25018_, new_n25019_, new_n25020_, new_n25021_, new_n25022_,
    new_n25023_, new_n25024_, new_n25025_, new_n25026_, new_n25027_,
    new_n25028_, new_n25029_, new_n25030_, new_n25031_, new_n25032_,
    new_n25033_, new_n25034_, new_n25035_, new_n25036_, new_n25037_,
    new_n25038_, new_n25039_, new_n25040_, new_n25041_, new_n25042_,
    new_n25043_, new_n25044_, new_n25045_, new_n25046_, new_n25047_,
    new_n25048_, new_n25049_, new_n25050_, new_n25051_, new_n25052_,
    new_n25053_, new_n25054_, new_n25055_, new_n25056_, new_n25057_,
    new_n25058_, new_n25059_, new_n25060_, new_n25061_, new_n25062_,
    new_n25063_, new_n25064_, new_n25065_, new_n25066_, new_n25067_,
    new_n25068_, new_n25069_, new_n25070_, new_n25071_, new_n25072_,
    new_n25073_, new_n25074_, new_n25075_, new_n25076_, new_n25077_,
    new_n25078_, new_n25079_, new_n25080_, new_n25081_, new_n25082_,
    new_n25083_, new_n25084_, new_n25085_, new_n25086_, new_n25087_,
    new_n25088_, new_n25089_, new_n25090_, new_n25091_, new_n25092_,
    new_n25093_, new_n25094_, new_n25095_, new_n25096_, new_n25097_,
    new_n25098_, new_n25099_, new_n25100_, new_n25101_, new_n25102_,
    new_n25103_, new_n25104_, new_n25105_, new_n25106_, new_n25107_,
    new_n25108_, new_n25109_, new_n25110_, new_n25111_, new_n25112_,
    new_n25113_, new_n25114_, new_n25115_, new_n25116_, new_n25117_,
    new_n25118_, new_n25119_, new_n25120_, new_n25121_, new_n25122_,
    new_n25123_, new_n25124_, new_n25125_, new_n25126_, new_n25127_,
    new_n25128_, new_n25129_, new_n25130_, new_n25131_, new_n25132_,
    new_n25133_, new_n25134_, new_n25135_, new_n25136_, new_n25137_,
    new_n25138_, new_n25139_, new_n25140_, new_n25141_, new_n25142_,
    new_n25143_, new_n25144_, new_n25145_, new_n25146_, new_n25147_,
    new_n25148_, new_n25149_, new_n25150_, new_n25151_, new_n25152_,
    new_n25153_, new_n25154_, new_n25155_, new_n25156_, new_n25157_,
    new_n25158_, new_n25159_, new_n25160_, new_n25161_, new_n25162_,
    new_n25163_, new_n25164_, new_n25165_, new_n25166_, new_n25167_,
    new_n25168_, new_n25169_, new_n25170_, new_n25171_, new_n25172_,
    new_n25173_, new_n25174_, new_n25175_, new_n25176_, new_n25177_,
    new_n25178_, new_n25179_, new_n25180_, new_n25181_, new_n25182_,
    new_n25183_, new_n25184_, new_n25185_, new_n25186_, new_n25187_,
    new_n25188_, new_n25189_, new_n25190_, new_n25191_, new_n25192_,
    new_n25193_, new_n25194_, new_n25195_, new_n25196_, new_n25197_,
    new_n25198_, new_n25199_, new_n25200_, new_n25201_, new_n25202_,
    new_n25203_, new_n25204_, new_n25205_, new_n25206_, new_n25207_,
    new_n25208_, new_n25209_, new_n25210_, new_n25211_, new_n25212_,
    new_n25213_, new_n25214_, new_n25215_, new_n25216_, new_n25217_,
    new_n25218_, new_n25219_, new_n25220_, new_n25221_, new_n25222_,
    new_n25223_, new_n25224_, new_n25225_, new_n25226_, new_n25227_,
    new_n25228_, new_n25229_, new_n25230_, new_n25231_, new_n25232_,
    new_n25233_, new_n25234_, new_n25235_, new_n25236_, new_n25237_,
    new_n25238_, new_n25239_, new_n25240_, new_n25241_, new_n25242_,
    new_n25243_, new_n25244_, new_n25245_, new_n25246_, new_n25247_,
    new_n25248_, new_n25249_, new_n25250_, new_n25251_, new_n25252_,
    new_n25253_, new_n25254_, new_n25255_, new_n25256_, new_n25257_,
    new_n25258_, new_n25259_, new_n25260_, new_n25261_, new_n25262_,
    new_n25263_, new_n25264_, new_n25265_, new_n25266_, new_n25267_,
    new_n25268_, new_n25269_, new_n25270_, new_n25271_, new_n25272_,
    new_n25273_, new_n25274_, new_n25275_, new_n25276_, new_n25277_,
    new_n25278_, new_n25279_, new_n25280_, new_n25281_, new_n25282_,
    new_n25283_, new_n25284_, new_n25285_, new_n25286_, new_n25287_,
    new_n25288_, new_n25289_, new_n25290_, new_n25291_, new_n25292_,
    new_n25293_, new_n25294_, new_n25295_, new_n25296_, new_n25297_,
    new_n25298_, new_n25299_, new_n25300_, new_n25301_, new_n25302_,
    new_n25303_, new_n25304_, new_n25305_, new_n25306_, new_n25307_,
    new_n25308_, new_n25309_, new_n25310_, new_n25311_, new_n25312_,
    new_n25313_, new_n25314_, new_n25315_, new_n25316_, new_n25317_,
    new_n25318_, new_n25319_, new_n25320_, new_n25321_, new_n25322_,
    new_n25323_, new_n25324_, new_n25325_, new_n25326_, new_n25327_,
    new_n25328_, new_n25329_, new_n25330_, new_n25331_, new_n25332_,
    new_n25333_, new_n25334_, new_n25335_, new_n25336_, new_n25337_,
    new_n25338_, new_n25339_, new_n25340_, new_n25341_, new_n25342_,
    new_n25343_, new_n25344_, new_n25345_, new_n25346_, new_n25347_,
    new_n25348_, new_n25349_, new_n25350_, new_n25351_, new_n25352_,
    new_n25353_, new_n25354_, new_n25355_, new_n25356_, new_n25357_,
    new_n25358_, new_n25359_, new_n25360_, new_n25361_, new_n25362_,
    new_n25363_, new_n25364_, new_n25365_, new_n25366_, new_n25367_,
    new_n25368_, new_n25369_, new_n25370_, new_n25371_, new_n25372_,
    new_n25373_, new_n25374_, new_n25375_, new_n25376_, new_n25377_,
    new_n25378_, new_n25379_, new_n25380_, new_n25381_, new_n25382_,
    new_n25383_, new_n25384_, new_n25385_, new_n25386_, new_n25387_,
    new_n25388_, new_n25389_, new_n25390_, new_n25391_, new_n25392_,
    new_n25393_, new_n25394_, new_n25395_, new_n25396_, new_n25397_,
    new_n25398_, new_n25399_, new_n25400_, new_n25401_, new_n25402_,
    new_n25403_, new_n25404_, new_n25405_, new_n25406_, new_n25407_,
    new_n25408_, new_n25409_, new_n25410_, new_n25411_, new_n25412_,
    new_n25413_, new_n25414_, new_n25415_, new_n25416_, new_n25417_,
    new_n25418_, new_n25419_, new_n25420_, new_n25421_, new_n25422_,
    new_n25423_, new_n25424_, new_n25425_, new_n25426_, new_n25427_,
    new_n25428_, new_n25429_, new_n25430_, new_n25431_, new_n25432_,
    new_n25433_, new_n25434_, new_n25435_, new_n25436_, new_n25437_,
    new_n25438_, new_n25439_, new_n25440_, new_n25441_, new_n25442_,
    new_n25443_, new_n25444_, new_n25445_, new_n25446_, new_n25447_,
    new_n25448_, new_n25449_, new_n25450_, new_n25451_, new_n25452_,
    new_n25453_, new_n25454_, new_n25455_, new_n25456_, new_n25457_,
    new_n25458_, new_n25459_, new_n25460_, new_n25461_, new_n25462_,
    new_n25463_, new_n25464_, new_n25465_, new_n25466_, new_n25467_,
    new_n25468_, new_n25469_, new_n25470_, new_n25471_, new_n25472_,
    new_n25473_, new_n25474_, new_n25475_, new_n25476_, new_n25477_,
    new_n25478_, new_n25479_, new_n25480_, new_n25481_, new_n25482_,
    new_n25483_, new_n25484_, new_n25485_, new_n25486_, new_n25487_,
    new_n25488_, new_n25489_, new_n25490_, new_n25491_, new_n25492_,
    new_n25493_, new_n25494_, new_n25495_, new_n25496_, new_n25497_,
    new_n25498_, new_n25499_, new_n25500_, new_n25501_, new_n25502_,
    new_n25503_, new_n25504_, new_n25505_, new_n25506_, new_n25507_,
    new_n25508_, new_n25509_, new_n25510_, new_n25511_, new_n25512_,
    new_n25513_, new_n25514_, new_n25515_, new_n25516_, new_n25517_,
    new_n25518_, new_n25519_, new_n25520_, new_n25521_, new_n25522_,
    new_n25523_, new_n25524_, new_n25525_, new_n25526_, new_n25527_,
    new_n25528_, new_n25529_, new_n25530_, new_n25531_, new_n25532_,
    new_n25533_, new_n25534_, new_n25535_, new_n25536_, new_n25537_,
    new_n25538_, new_n25539_, new_n25540_, new_n25541_, new_n25542_,
    new_n25543_, new_n25544_, new_n25545_, new_n25546_, new_n25547_,
    new_n25548_, new_n25549_, new_n25550_, new_n25551_, new_n25552_,
    new_n25553_, new_n25554_, new_n25555_, new_n25556_, new_n25557_,
    new_n25558_, new_n25559_, new_n25560_, new_n25561_, new_n25562_,
    new_n25563_, new_n25564_, new_n25565_, new_n25566_, new_n25567_,
    new_n25568_, new_n25569_, new_n25570_, new_n25571_, new_n25572_,
    new_n25573_, new_n25574_, new_n25575_, new_n25576_, new_n25577_,
    new_n25578_, new_n25579_, new_n25580_, new_n25581_, new_n25582_,
    new_n25583_, new_n25584_, new_n25585_, new_n25586_, new_n25587_,
    new_n25588_, new_n25589_, new_n25590_, new_n25591_, new_n25592_,
    new_n25593_, new_n25594_, new_n25595_, new_n25596_, new_n25597_,
    new_n25598_, new_n25599_, new_n25600_, new_n25601_, new_n25602_,
    new_n25603_, new_n25604_, new_n25605_, new_n25606_, new_n25607_,
    new_n25608_, new_n25609_, new_n25610_, new_n25611_, new_n25612_,
    new_n25613_, new_n25614_, new_n25615_, new_n25616_, new_n25617_,
    new_n25618_, new_n25619_, new_n25620_, new_n25621_, new_n25622_,
    new_n25623_, new_n25624_, new_n25625_, new_n25626_, new_n25627_,
    new_n25628_, new_n25629_, new_n25630_, new_n25631_, new_n25632_,
    new_n25633_, new_n25634_, new_n25635_, new_n25636_, new_n25637_,
    new_n25638_, new_n25639_, new_n25640_, new_n25641_, new_n25642_,
    new_n25643_, new_n25644_, new_n25645_, new_n25646_, new_n25647_,
    new_n25648_, new_n25649_, new_n25650_, new_n25651_, new_n25652_,
    new_n25653_, new_n25654_, new_n25655_, new_n25656_, new_n25657_,
    new_n25658_, new_n25659_, new_n25660_, new_n25661_, new_n25662_,
    new_n25663_, new_n25664_, new_n25665_, new_n25666_, new_n25667_,
    new_n25668_, new_n25669_, new_n25670_, new_n25671_, new_n25672_,
    new_n25673_, new_n25674_, new_n25675_, new_n25676_, new_n25677_,
    new_n25678_, new_n25679_, new_n25680_, new_n25681_, new_n25682_,
    new_n25683_, new_n25684_, new_n25685_, new_n25686_, new_n25687_,
    new_n25688_, new_n25689_, new_n25690_, new_n25691_, new_n25692_,
    new_n25693_, new_n25694_, new_n25695_, new_n25696_, new_n25697_,
    new_n25698_, new_n25699_, new_n25700_, new_n25701_, new_n25702_,
    new_n25703_, new_n25704_, new_n25705_, new_n25706_, new_n25707_,
    new_n25708_, new_n25709_, new_n25710_, new_n25711_, new_n25712_,
    new_n25713_, new_n25714_, new_n25715_, new_n25716_, new_n25717_,
    new_n25718_, new_n25719_, new_n25720_, new_n25721_, new_n25722_,
    new_n25723_, new_n25724_, new_n25725_, new_n25726_, new_n25727_,
    new_n25728_, new_n25729_, new_n25730_, new_n25731_, new_n25732_,
    new_n25733_, new_n25734_, new_n25735_, new_n25736_, new_n25737_,
    new_n25738_, new_n25739_, new_n25740_, new_n25741_, new_n25742_,
    new_n25743_, new_n25744_, new_n25745_, new_n25746_, new_n25747_,
    new_n25748_, new_n25749_, new_n25750_, new_n25751_, new_n25752_,
    new_n25753_, new_n25754_, new_n25755_, new_n25756_, new_n25757_,
    new_n25758_, new_n25759_, new_n25760_, new_n25761_, new_n25762_,
    new_n25763_, new_n25764_, new_n25765_, new_n25766_, new_n25767_,
    new_n25768_, new_n25769_, new_n25770_, new_n25771_, new_n25772_,
    new_n25773_, new_n25774_, new_n25775_, new_n25776_, new_n25777_,
    new_n25778_, new_n25779_, new_n25780_, new_n25781_, new_n25782_,
    new_n25783_, new_n25784_, new_n25785_, new_n25786_, new_n25787_,
    new_n25788_, new_n25789_, new_n25790_, new_n25791_, new_n25792_,
    new_n25793_, new_n25794_, new_n25795_, new_n25796_, new_n25797_,
    new_n25798_, new_n25799_, new_n25800_, new_n25801_, new_n25802_,
    new_n25803_, new_n25804_, new_n25805_, new_n25806_, new_n25807_,
    new_n25808_, new_n25809_, new_n25810_, new_n25811_, new_n25812_,
    new_n25813_, new_n25814_, new_n25815_, new_n25816_, new_n25817_,
    new_n25818_, new_n25819_, new_n25820_, new_n25821_, new_n25822_,
    new_n25823_, new_n25824_, new_n25825_, new_n25826_, new_n25827_,
    new_n25828_, new_n25829_, new_n25830_, new_n25831_, new_n25832_,
    new_n25833_, new_n25834_, new_n25835_, new_n25836_, new_n25837_,
    new_n25838_, new_n25839_, new_n25840_, new_n25841_, new_n25842_,
    new_n25843_, new_n25844_, new_n25845_, new_n25846_, new_n25847_,
    new_n25848_, new_n25849_, new_n25850_, new_n25851_, new_n25852_,
    new_n25853_, new_n25854_, new_n25855_, new_n25856_, new_n25857_,
    new_n25858_, new_n25859_, new_n25860_, new_n25861_, new_n25862_,
    new_n25863_, new_n25864_, new_n25865_, new_n25866_, new_n25867_,
    new_n25868_, new_n25869_, new_n25870_, new_n25871_, new_n25872_,
    new_n25873_, new_n25874_, new_n25875_, new_n25876_, new_n25877_,
    new_n25878_, new_n25879_, new_n25880_, new_n25881_, new_n25882_,
    new_n25883_, new_n25884_, new_n25885_, new_n25886_, new_n25887_,
    new_n25888_, new_n25889_, new_n25890_, new_n25891_, new_n25892_,
    new_n25893_, new_n25894_, new_n25895_, new_n25896_, new_n25897_,
    new_n25898_, new_n25899_, new_n25900_, new_n25901_, new_n25902_,
    new_n25903_, new_n25904_, new_n25905_, new_n25906_, new_n25907_,
    new_n25908_, new_n25909_, new_n25910_, new_n25911_, new_n25912_,
    new_n25913_, new_n25914_, new_n25915_, new_n25916_, new_n25917_,
    new_n25918_, new_n25919_, new_n25920_, new_n25921_, new_n25922_,
    new_n25923_, new_n25924_, new_n25925_, new_n25926_, new_n25927_,
    new_n25928_, new_n25929_, new_n25930_, new_n25931_, new_n25932_,
    new_n25933_, new_n25934_, new_n25935_, new_n25936_, new_n25937_,
    new_n25938_, new_n25939_, new_n25940_, new_n25941_, new_n25942_,
    new_n25943_, new_n25944_, new_n25945_, new_n25946_, new_n25947_,
    new_n25948_, new_n25949_, new_n25950_, new_n25951_, new_n25952_,
    new_n25953_, new_n25954_, new_n25955_, new_n25956_, new_n25957_,
    new_n25958_, new_n25959_, new_n25960_, new_n25961_, new_n25962_,
    new_n25963_, new_n25964_, new_n25965_, new_n25966_, new_n25967_,
    new_n25968_, new_n25969_, new_n25970_, new_n25971_, new_n25972_,
    new_n25973_, new_n25974_, new_n25975_, new_n25976_, new_n25977_,
    new_n25978_, new_n25979_, new_n25980_, new_n25981_, new_n25982_,
    new_n25983_, new_n25984_, new_n25985_, new_n25986_, new_n25987_,
    new_n25988_, new_n25989_, new_n25990_, new_n25991_, new_n25992_,
    new_n25993_, new_n25994_, new_n25995_, new_n25996_, new_n25997_,
    new_n25998_, new_n25999_, new_n26000_, new_n26001_, new_n26002_,
    new_n26003_, new_n26004_, new_n26005_, new_n26006_, new_n26007_,
    new_n26008_, new_n26009_, new_n26010_, new_n26011_, new_n26012_,
    new_n26013_, new_n26014_, new_n26015_, new_n26016_, new_n26017_,
    new_n26018_, new_n26019_, new_n26020_, new_n26021_, new_n26022_,
    new_n26023_, new_n26024_, new_n26025_, new_n26026_, new_n26027_,
    new_n26028_, new_n26029_, new_n26030_, new_n26031_, new_n26032_,
    new_n26033_, new_n26034_, new_n26035_, new_n26036_, new_n26037_,
    new_n26038_, new_n26039_, new_n26040_, new_n26041_, new_n26042_,
    new_n26043_, new_n26044_, new_n26045_, new_n26046_, new_n26047_,
    new_n26048_, new_n26049_, new_n26050_, new_n26051_, new_n26052_,
    new_n26053_, new_n26054_, new_n26055_, new_n26056_, new_n26057_,
    new_n26058_, new_n26059_, new_n26060_, new_n26061_, new_n26062_,
    new_n26063_, new_n26064_, new_n26065_, new_n26066_, new_n26067_,
    new_n26068_, new_n26069_, new_n26070_, new_n26071_, new_n26072_,
    new_n26073_, new_n26074_, new_n26075_, new_n26076_, new_n26077_,
    new_n26078_, new_n26079_, new_n26080_, new_n26081_, new_n26082_,
    new_n26083_, new_n26084_, new_n26085_, new_n26086_, new_n26087_,
    new_n26088_, new_n26089_, new_n26090_, new_n26091_, new_n26092_,
    new_n26093_, new_n26094_, new_n26095_, new_n26096_, new_n26097_,
    new_n26098_, new_n26099_, new_n26100_, new_n26101_, new_n26102_,
    new_n26103_, new_n26104_, new_n26105_, new_n26106_, new_n26107_,
    new_n26108_, new_n26109_, new_n26110_, new_n26111_, new_n26112_,
    new_n26113_, new_n26114_, new_n26115_, new_n26116_, new_n26117_,
    new_n26118_, new_n26119_, new_n26120_, new_n26121_, new_n26122_,
    new_n26123_, new_n26124_, new_n26125_, new_n26126_, new_n26127_,
    new_n26128_, new_n26129_, new_n26130_, new_n26131_, new_n26132_,
    new_n26133_, new_n26134_, new_n26135_, new_n26136_, new_n26137_,
    new_n26138_, new_n26139_, new_n26140_, new_n26141_, new_n26142_,
    new_n26143_, new_n26144_, new_n26145_, new_n26146_, new_n26147_,
    new_n26148_, new_n26149_, new_n26150_, new_n26151_, new_n26152_,
    new_n26153_, new_n26154_, new_n26155_, new_n26156_, new_n26157_,
    new_n26158_, new_n26159_, new_n26160_, new_n26161_, new_n26162_,
    new_n26163_, new_n26164_, new_n26165_, new_n26166_, new_n26167_,
    new_n26168_, new_n26169_, new_n26170_, new_n26171_, new_n26172_,
    new_n26173_, new_n26174_, new_n26175_, new_n26176_, new_n26177_,
    new_n26178_, new_n26179_, new_n26180_, new_n26181_, new_n26182_,
    new_n26183_, new_n26184_, new_n26185_, new_n26186_, new_n26187_,
    new_n26188_, new_n26189_, new_n26190_, new_n26191_, new_n26192_,
    new_n26193_, new_n26194_, new_n26195_, new_n26196_, new_n26197_,
    new_n26198_, new_n26199_, new_n26200_, new_n26201_, new_n26202_,
    new_n26203_, new_n26204_, new_n26205_, new_n26206_, new_n26207_,
    new_n26208_, new_n26209_, new_n26210_, new_n26211_, new_n26212_,
    new_n26213_, new_n26214_, new_n26215_, new_n26216_, new_n26217_,
    new_n26218_, new_n26219_, new_n26220_, new_n26221_, new_n26222_,
    new_n26223_, new_n26224_, new_n26225_, new_n26226_, new_n26227_,
    new_n26228_, new_n26229_, new_n26230_, new_n26231_, new_n26232_,
    new_n26233_, new_n26234_, new_n26235_, new_n26236_, new_n26237_,
    new_n26238_, new_n26239_, new_n26240_, new_n26241_, new_n26242_,
    new_n26243_, new_n26244_, new_n26245_, new_n26246_, new_n26247_,
    new_n26248_, new_n26249_, new_n26250_, new_n26251_, new_n26252_,
    new_n26253_, new_n26254_, new_n26255_, new_n26256_, new_n26257_,
    new_n26258_, new_n26259_, new_n26260_, new_n26261_, new_n26262_,
    new_n26263_, new_n26264_, new_n26265_, new_n26266_, new_n26267_,
    new_n26268_, new_n26269_, new_n26270_, new_n26271_, new_n26272_,
    new_n26273_, new_n26274_, new_n26275_, new_n26276_, new_n26277_,
    new_n26278_, new_n26279_, new_n26280_, new_n26281_, new_n26282_,
    new_n26283_, new_n26284_, new_n26285_, new_n26286_, new_n26287_,
    new_n26288_, new_n26289_, new_n26290_, new_n26291_, new_n26292_,
    new_n26293_, new_n26294_, new_n26295_, new_n26296_, new_n26297_,
    new_n26298_, new_n26299_, new_n26300_, new_n26301_, new_n26302_,
    new_n26303_, new_n26304_, new_n26305_, new_n26306_, new_n26307_,
    new_n26308_, new_n26309_, new_n26310_, new_n26311_, new_n26312_,
    new_n26313_, new_n26314_, new_n26315_, new_n26316_, new_n26317_,
    new_n26318_, new_n26319_, new_n26320_, new_n26321_, new_n26322_,
    new_n26323_, new_n26324_, new_n26325_, new_n26326_, new_n26327_,
    new_n26328_, new_n26329_, new_n26330_, new_n26331_, new_n26332_,
    new_n26333_, new_n26334_, new_n26335_, new_n26336_, new_n26337_,
    new_n26338_, new_n26339_, new_n26340_, new_n26341_, new_n26342_,
    new_n26343_, new_n26344_, new_n26345_, new_n26346_, new_n26347_,
    new_n26348_, new_n26349_, new_n26350_, new_n26351_, new_n26352_,
    new_n26353_, new_n26354_, new_n26355_, new_n26356_, new_n26357_,
    new_n26358_, new_n26359_, new_n26360_, new_n26361_, new_n26362_,
    new_n26363_, new_n26364_, new_n26365_, new_n26366_, new_n26367_,
    new_n26368_, new_n26369_, new_n26370_, new_n26371_, new_n26372_,
    new_n26373_, new_n26374_, new_n26375_, new_n26376_, new_n26377_,
    new_n26378_, new_n26379_, new_n26380_, new_n26381_, new_n26382_,
    new_n26383_, new_n26384_, new_n26385_, new_n26386_, new_n26387_,
    new_n26388_, new_n26389_, new_n26390_, new_n26391_, new_n26392_,
    new_n26393_, new_n26394_, new_n26395_, new_n26396_, new_n26397_,
    new_n26398_, new_n26399_, new_n26400_, new_n26401_, new_n26402_,
    new_n26403_, new_n26404_, new_n26405_, new_n26406_, new_n26407_,
    new_n26408_, new_n26409_, new_n26410_, new_n26411_, new_n26412_,
    new_n26413_, new_n26414_, new_n26415_, new_n26416_, new_n26417_,
    new_n26418_, new_n26419_, new_n26420_, new_n26421_, new_n26422_,
    new_n26423_, new_n26424_, new_n26425_, new_n26426_, new_n26427_,
    new_n26428_, new_n26429_, new_n26430_, new_n26431_, new_n26432_,
    new_n26433_, new_n26434_, new_n26435_, new_n26436_, new_n26437_,
    new_n26438_, new_n26439_, new_n26440_, new_n26441_, new_n26442_,
    new_n26443_, new_n26444_, new_n26445_, new_n26446_, new_n26447_,
    new_n26448_, new_n26449_, new_n26450_, new_n26451_, new_n26452_,
    new_n26453_, new_n26454_, new_n26455_, new_n26456_, new_n26457_,
    new_n26458_, new_n26459_, new_n26460_, new_n26461_, new_n26462_,
    new_n26463_, new_n26464_, new_n26465_, new_n26466_, new_n26467_,
    new_n26468_, new_n26469_, new_n26470_, new_n26471_, new_n26472_,
    new_n26473_, new_n26474_, new_n26475_, new_n26476_, new_n26477_,
    new_n26478_, new_n26479_, new_n26480_, new_n26481_, new_n26482_,
    new_n26483_, new_n26484_, new_n26485_, new_n26486_, new_n26487_,
    new_n26488_, new_n26489_, new_n26490_, new_n26491_, new_n26492_,
    new_n26493_, new_n26494_, new_n26495_, new_n26496_, new_n26497_,
    new_n26498_, new_n26499_, new_n26500_, new_n26501_, new_n26502_,
    new_n26503_, new_n26504_, new_n26505_, new_n26506_, new_n26507_,
    new_n26508_, new_n26509_, new_n26510_, new_n26511_, new_n26512_,
    new_n26513_, new_n26514_, new_n26515_, new_n26516_, new_n26517_,
    new_n26518_, new_n26519_, new_n26520_, new_n26521_, new_n26522_,
    new_n26523_, new_n26524_, new_n26525_, new_n26526_, new_n26527_,
    new_n26528_, new_n26529_, new_n26530_, new_n26531_, new_n26532_,
    new_n26533_, new_n26534_, new_n26535_, new_n26536_, new_n26537_,
    new_n26538_, new_n26539_, new_n26540_, new_n26541_, new_n26542_,
    new_n26543_, new_n26544_, new_n26545_, new_n26546_, new_n26547_,
    new_n26548_, new_n26549_, new_n26550_, new_n26551_, new_n26552_,
    new_n26553_, new_n26554_, new_n26555_, new_n26556_, new_n26557_,
    new_n26558_, new_n26559_, new_n26560_, new_n26561_, new_n26562_,
    new_n26563_, new_n26564_, new_n26565_, new_n26566_, new_n26567_,
    new_n26568_, new_n26569_, new_n26570_, new_n26571_, new_n26572_,
    new_n26573_, new_n26574_, new_n26575_, new_n26576_, new_n26577_,
    new_n26578_, new_n26579_, new_n26580_, new_n26581_, new_n26582_,
    new_n26583_, new_n26584_, new_n26585_, new_n26586_, new_n26587_,
    new_n26588_, new_n26589_, new_n26590_, new_n26591_, new_n26592_,
    new_n26593_, new_n26594_, new_n26595_, new_n26596_, new_n26597_,
    new_n26598_, new_n26599_, new_n26600_, new_n26601_, new_n26602_,
    new_n26603_, new_n26604_, new_n26605_, new_n26606_, new_n26607_,
    new_n26608_, new_n26609_, new_n26610_, new_n26611_, new_n26612_,
    new_n26613_, new_n26614_, new_n26615_, new_n26616_, new_n26617_,
    new_n26618_, new_n26619_, new_n26620_, new_n26621_, new_n26622_,
    new_n26623_, new_n26624_, new_n26625_, new_n26626_, new_n26627_,
    new_n26628_, new_n26629_, new_n26630_, new_n26631_, new_n26632_,
    new_n26633_, new_n26634_, new_n26635_, new_n26636_, new_n26637_,
    new_n26638_, new_n26639_, new_n26640_, new_n26641_, new_n26642_,
    new_n26643_, new_n26644_, new_n26645_, new_n26646_, new_n26647_,
    new_n26648_, new_n26649_, new_n26650_, new_n26651_, new_n26652_,
    new_n26653_, new_n26654_, new_n26655_, new_n26656_, new_n26657_,
    new_n26658_, new_n26659_, new_n26660_, new_n26661_, new_n26662_,
    new_n26663_, new_n26664_, new_n26665_, new_n26666_, new_n26667_,
    new_n26668_, new_n26669_, new_n26670_, new_n26671_, new_n26672_,
    new_n26673_, new_n26674_, new_n26675_, new_n26676_, new_n26677_,
    new_n26678_, new_n26679_, new_n26680_, new_n26681_, new_n26682_,
    new_n26683_, new_n26684_, new_n26685_, new_n26686_, new_n26687_,
    new_n26688_, new_n26689_, new_n26690_, new_n26691_, new_n26692_,
    new_n26693_, new_n26694_, new_n26695_, new_n26696_, new_n26697_,
    new_n26698_, new_n26699_, new_n26700_, new_n26701_, new_n26702_,
    new_n26703_, new_n26704_, new_n26705_, new_n26706_, new_n26707_,
    new_n26708_, new_n26709_, new_n26710_, new_n26711_, new_n26712_,
    new_n26713_, new_n26714_, new_n26715_, new_n26716_, new_n26717_,
    new_n26718_, new_n26719_, new_n26720_, new_n26721_, new_n26722_,
    new_n26723_, new_n26724_, new_n26725_, new_n26726_, new_n26727_,
    new_n26728_, new_n26729_, new_n26730_, new_n26731_, new_n26732_,
    new_n26733_, new_n26734_, new_n26735_, new_n26736_, new_n26737_,
    new_n26738_, new_n26739_, new_n26740_, new_n26741_, new_n26742_,
    new_n26743_, new_n26744_, new_n26745_, new_n26746_, new_n26747_,
    new_n26748_, new_n26749_, new_n26750_, new_n26751_, new_n26752_,
    new_n26753_, new_n26754_, new_n26755_, new_n26756_, new_n26757_,
    new_n26758_, new_n26759_, new_n26760_, new_n26761_, new_n26762_,
    new_n26763_, new_n26764_, new_n26765_, new_n26766_, new_n26767_,
    new_n26768_, new_n26769_, new_n26770_, new_n26771_, new_n26772_,
    new_n26773_, new_n26774_, new_n26775_, new_n26776_, new_n26777_,
    new_n26778_, new_n26779_, new_n26780_, new_n26781_, new_n26782_,
    new_n26783_, new_n26784_, new_n26785_, new_n26786_, new_n26787_,
    new_n26788_, new_n26789_, new_n26790_, new_n26791_, new_n26792_,
    new_n26793_, new_n26794_, new_n26795_, new_n26796_, new_n26797_,
    new_n26798_, new_n26799_, new_n26800_, new_n26801_, new_n26802_,
    new_n26803_, new_n26804_, new_n26805_, new_n26806_, new_n26807_,
    new_n26808_, new_n26809_, new_n26810_, new_n26811_, new_n26812_,
    new_n26813_, new_n26814_, new_n26815_, new_n26816_, new_n26817_,
    new_n26818_, new_n26819_, new_n26820_, new_n26821_, new_n26822_,
    new_n26823_, new_n26824_, new_n26825_, new_n26826_, new_n26827_,
    new_n26828_, new_n26829_, new_n26830_, new_n26831_, new_n26832_,
    new_n26833_, new_n26834_, new_n26835_, new_n26836_, new_n26837_,
    new_n26838_, new_n26839_, new_n26840_, new_n26841_, new_n26842_,
    new_n26843_, new_n26844_, new_n26845_, new_n26846_, new_n26847_,
    new_n26848_, new_n26849_, new_n26850_, new_n26851_, new_n26852_,
    new_n26853_, new_n26854_, new_n26855_, new_n26856_, new_n26857_,
    new_n26858_, new_n26859_, new_n26860_, new_n26861_, new_n26862_,
    new_n26863_, new_n26864_, new_n26865_, new_n26866_, new_n26867_,
    new_n26868_, new_n26869_, new_n26870_, new_n26871_, new_n26872_,
    new_n26873_, new_n26874_, new_n26875_, new_n26876_, new_n26877_,
    new_n26878_, new_n26879_, new_n26880_, new_n26881_, new_n26882_,
    new_n26883_, new_n26884_, new_n26885_, new_n26886_, new_n26887_,
    new_n26888_, new_n26889_, new_n26890_, new_n26891_, new_n26892_,
    new_n26893_, new_n26894_, new_n26895_, new_n26896_, new_n26897_,
    new_n26898_, new_n26899_, new_n26900_, new_n26901_, new_n26902_,
    new_n26903_, new_n26904_, new_n26905_, new_n26906_, new_n26907_,
    new_n26908_, new_n26909_, new_n26910_, new_n26911_, new_n26912_,
    new_n26913_, new_n26914_, new_n26915_, new_n26916_, new_n26917_,
    new_n26918_, new_n26919_, new_n26920_, new_n26921_, new_n26922_,
    new_n26923_, new_n26924_, new_n26925_, new_n26926_, new_n26927_,
    new_n26928_, new_n26929_, new_n26930_, new_n26931_, new_n26932_,
    new_n26933_, new_n26934_, new_n26935_, new_n26936_, new_n26937_,
    new_n26938_, new_n26939_, new_n26940_, new_n26941_, new_n26942_,
    new_n26943_, new_n26944_, new_n26945_, new_n26946_, new_n26947_,
    new_n26948_, new_n26949_, new_n26950_, new_n26951_, new_n26952_,
    new_n26953_, new_n26954_, new_n26955_, new_n26956_, new_n26957_,
    new_n26958_, new_n26959_, new_n26960_, new_n26961_, new_n26962_,
    new_n26963_, new_n26964_, new_n26965_, new_n26966_, new_n26967_,
    new_n26968_, new_n26969_, new_n26970_, new_n26971_, new_n26972_,
    new_n26973_, new_n26974_, new_n26975_, new_n26976_, new_n26977_,
    new_n26978_, new_n26979_, new_n26980_, new_n26981_, new_n26982_,
    new_n26983_, new_n26984_, new_n26985_, new_n26986_, new_n26987_,
    new_n26988_, new_n26989_, new_n26990_, new_n26991_, new_n26992_,
    new_n26993_, new_n26994_, new_n26995_, new_n26996_, new_n26997_,
    new_n26998_, new_n26999_, new_n27000_, new_n27001_, new_n27002_,
    new_n27003_, new_n27004_, new_n27005_, new_n27006_, new_n27007_,
    new_n27008_, new_n27009_, new_n27010_, new_n27011_, new_n27012_,
    new_n27013_, new_n27014_, new_n27015_, new_n27016_, new_n27017_,
    new_n27018_, new_n27019_, new_n27020_, new_n27021_, new_n27022_,
    new_n27023_, new_n27024_, new_n27025_, new_n27026_, new_n27027_,
    new_n27028_, new_n27029_, new_n27030_, new_n27031_, new_n27032_,
    new_n27033_, new_n27034_, new_n27035_, new_n27036_, new_n27037_,
    new_n27038_, new_n27039_, new_n27040_, new_n27041_, new_n27042_,
    new_n27043_, new_n27044_, new_n27045_, new_n27046_, new_n27047_,
    new_n27048_, new_n27049_, new_n27050_, new_n27051_, new_n27052_,
    new_n27053_, new_n27054_, new_n27055_, new_n27056_, new_n27057_,
    new_n27058_, new_n27059_, new_n27060_, new_n27061_, new_n27062_,
    new_n27063_, new_n27064_, new_n27065_, new_n27066_, new_n27067_,
    new_n27068_, new_n27069_, new_n27070_, new_n27071_, new_n27072_,
    new_n27073_, new_n27074_, new_n27075_, new_n27076_, new_n27077_,
    new_n27078_, new_n27079_, new_n27080_, new_n27081_, new_n27082_,
    new_n27083_, new_n27084_, new_n27085_, new_n27086_, new_n27087_,
    new_n27088_, new_n27089_, new_n27090_, new_n27091_, new_n27092_,
    new_n27093_, new_n27094_, new_n27095_, new_n27096_, new_n27097_,
    new_n27098_, new_n27099_, new_n27100_, new_n27101_, new_n27102_,
    new_n27103_, new_n27104_, new_n27105_, new_n27106_, new_n27107_,
    new_n27108_, new_n27109_, new_n27110_, new_n27111_, new_n27112_,
    new_n27113_, new_n27114_, new_n27115_, new_n27116_, new_n27117_,
    new_n27118_, new_n27119_, new_n27120_, new_n27121_, new_n27122_,
    new_n27123_, new_n27124_, new_n27125_, new_n27126_, new_n27127_,
    new_n27128_, new_n27129_, new_n27130_, new_n27131_, new_n27132_,
    new_n27133_, new_n27134_, new_n27135_, new_n27136_, new_n27137_,
    new_n27138_, new_n27139_, new_n27140_, new_n27141_, new_n27142_,
    new_n27143_, new_n27144_, new_n27145_, new_n27146_, new_n27147_,
    new_n27148_, new_n27149_, new_n27150_, new_n27151_, new_n27152_,
    new_n27153_, new_n27154_, new_n27155_, new_n27156_, new_n27157_,
    new_n27158_, new_n27159_, new_n27160_, new_n27161_, new_n27162_,
    new_n27163_, new_n27164_, new_n27165_, new_n27166_, new_n27167_,
    new_n27168_, new_n27169_, new_n27170_, new_n27171_, new_n27172_,
    new_n27173_, new_n27174_, new_n27175_, new_n27176_, new_n27177_,
    new_n27178_, new_n27179_, new_n27180_, new_n27181_, new_n27182_,
    new_n27183_, new_n27184_, new_n27185_, new_n27186_, new_n27187_,
    new_n27188_, new_n27189_, new_n27190_, new_n27191_, new_n27192_,
    new_n27193_, new_n27194_, new_n27195_, new_n27196_, new_n27197_,
    new_n27198_, new_n27199_, new_n27200_, new_n27201_, new_n27202_,
    new_n27203_, new_n27204_, new_n27205_, new_n27206_, new_n27207_,
    new_n27208_, new_n27209_, new_n27210_, new_n27211_, new_n27212_,
    new_n27213_, new_n27214_, new_n27215_, new_n27216_, new_n27217_,
    new_n27218_, new_n27219_, new_n27220_, new_n27221_, new_n27222_,
    new_n27223_, new_n27224_, new_n27225_, new_n27226_, new_n27227_,
    new_n27228_, new_n27229_, new_n27230_, new_n27231_, new_n27232_,
    new_n27233_, new_n27234_, new_n27235_, new_n27236_, new_n27237_,
    new_n27238_, new_n27239_, new_n27240_, new_n27241_, new_n27242_,
    new_n27243_, new_n27244_, new_n27245_, new_n27246_, new_n27247_,
    new_n27248_, new_n27249_, new_n27250_, new_n27251_, new_n27252_,
    new_n27253_, new_n27254_, new_n27255_, new_n27256_, new_n27257_,
    new_n27258_, new_n27259_, new_n27260_, new_n27261_, new_n27262_,
    new_n27263_, new_n27264_, new_n27265_, new_n27266_, new_n27267_,
    new_n27268_, new_n27269_, new_n27270_, new_n27271_, new_n27272_,
    new_n27273_, new_n27274_, new_n27275_, new_n27276_, new_n27277_,
    new_n27278_, new_n27279_, new_n27280_, new_n27281_, new_n27282_,
    new_n27283_, new_n27284_, new_n27285_, new_n27286_, new_n27287_,
    new_n27288_, new_n27289_, new_n27290_, new_n27291_, new_n27292_,
    new_n27293_, new_n27294_, new_n27295_, new_n27296_, new_n27297_,
    new_n27298_, new_n27299_, new_n27300_, new_n27301_, new_n27302_,
    new_n27303_, new_n27304_, new_n27305_, new_n27306_, new_n27307_,
    new_n27308_, new_n27309_, new_n27310_, new_n27311_, new_n27312_,
    new_n27313_, new_n27314_, new_n27315_, new_n27316_, new_n27317_,
    new_n27318_, new_n27319_, new_n27320_, new_n27321_, new_n27322_,
    new_n27323_, new_n27324_, new_n27325_, new_n27326_, new_n27327_,
    new_n27328_, new_n27329_, new_n27330_, new_n27331_, new_n27332_,
    new_n27333_, new_n27334_, new_n27335_, new_n27336_, new_n27337_,
    new_n27338_, new_n27339_, new_n27340_, new_n27341_, new_n27342_,
    new_n27343_, new_n27344_, new_n27345_, new_n27346_, new_n27347_,
    new_n27348_, new_n27349_, new_n27350_, new_n27351_, new_n27352_,
    new_n27353_, new_n27354_, new_n27355_, new_n27356_, new_n27357_,
    new_n27358_, new_n27359_, new_n27360_, new_n27361_, new_n27362_,
    new_n27363_, new_n27364_, new_n27365_, new_n27366_, new_n27367_,
    new_n27368_, new_n27369_, new_n27370_, new_n27371_, new_n27372_,
    new_n27373_, new_n27374_, new_n27375_, new_n27376_, new_n27377_,
    new_n27378_, new_n27379_, new_n27380_, new_n27381_, new_n27382_,
    new_n27383_, new_n27384_, new_n27385_, new_n27386_, new_n27387_,
    new_n27388_, new_n27389_, new_n27390_, new_n27391_, new_n27392_,
    new_n27393_, new_n27394_, new_n27395_, new_n27396_, new_n27397_,
    new_n27398_, new_n27399_, new_n27400_, new_n27401_, new_n27402_,
    new_n27403_, new_n27404_, new_n27405_, new_n27406_, new_n27407_,
    new_n27408_, new_n27409_, new_n27410_, new_n27411_, new_n27412_,
    new_n27413_, new_n27414_, new_n27415_, new_n27416_, new_n27417_,
    new_n27418_, new_n27419_, new_n27420_, new_n27421_, new_n27422_,
    new_n27423_, new_n27424_, new_n27425_, new_n27426_, new_n27427_,
    new_n27428_, new_n27429_, new_n27430_, new_n27431_, new_n27432_,
    new_n27433_, new_n27434_, new_n27435_, new_n27436_, new_n27437_,
    new_n27438_, new_n27439_, new_n27440_, new_n27441_, new_n27442_,
    new_n27443_, new_n27444_, new_n27445_, new_n27446_, new_n27447_,
    new_n27448_, new_n27449_, new_n27450_, new_n27451_, new_n27452_,
    new_n27453_, new_n27454_, new_n27455_, new_n27456_, new_n27457_,
    new_n27458_, new_n27459_, new_n27460_, new_n27461_, new_n27462_,
    new_n27463_, new_n27464_, new_n27465_, new_n27466_, new_n27467_,
    new_n27468_, new_n27469_, new_n27470_, new_n27471_, new_n27472_,
    new_n27473_, new_n27474_, new_n27475_, new_n27476_, new_n27477_,
    new_n27478_, new_n27479_, new_n27480_, new_n27481_, new_n27482_,
    new_n27483_, new_n27484_, new_n27485_, new_n27486_, new_n27487_,
    new_n27488_, new_n27489_, new_n27490_, new_n27491_, new_n27492_,
    new_n27493_, new_n27494_, new_n27495_, new_n27496_, new_n27497_,
    new_n27498_, new_n27499_, new_n27500_, new_n27501_, new_n27502_,
    new_n27503_, new_n27504_, new_n27505_, new_n27506_, new_n27507_,
    new_n27508_, new_n27509_, new_n27510_, new_n27511_, new_n27512_,
    new_n27513_, new_n27514_, new_n27515_, new_n27516_, new_n27517_,
    new_n27518_, new_n27519_, new_n27520_, new_n27521_, new_n27522_,
    new_n27523_, new_n27524_, new_n27525_, new_n27526_, new_n27527_,
    new_n27528_, new_n27529_, new_n27530_, new_n27531_, new_n27532_,
    new_n27533_, new_n27534_, new_n27535_, new_n27536_, new_n27537_,
    new_n27538_, new_n27539_, new_n27540_, new_n27541_, new_n27542_,
    new_n27543_, new_n27544_, new_n27545_, new_n27546_, new_n27547_,
    new_n27548_, new_n27549_, new_n27550_, new_n27551_, new_n27552_,
    new_n27553_, new_n27554_, new_n27555_, new_n27556_, new_n27557_,
    new_n27558_, new_n27559_, new_n27560_, new_n27561_, new_n27562_,
    new_n27563_, new_n27564_, new_n27565_, new_n27566_, new_n27567_,
    new_n27568_, new_n27569_, new_n27570_, new_n27571_, new_n27572_,
    new_n27573_, new_n27574_, new_n27575_, new_n27576_, new_n27577_,
    new_n27578_, new_n27579_, new_n27580_, new_n27581_, new_n27582_,
    new_n27583_, new_n27584_, new_n27585_, new_n27586_, new_n27587_,
    new_n27588_, new_n27589_, new_n27590_, new_n27591_, new_n27592_,
    new_n27593_, new_n27594_, new_n27595_, new_n27596_, new_n27597_,
    new_n27598_, new_n27599_, new_n27600_, new_n27601_, new_n27602_,
    new_n27603_, new_n27604_, new_n27605_, new_n27606_, new_n27607_,
    new_n27608_, new_n27609_, new_n27610_, new_n27611_, new_n27612_,
    new_n27613_, new_n27614_, new_n27615_, new_n27616_, new_n27617_,
    new_n27618_, new_n27619_, new_n27620_, new_n27621_, new_n27622_,
    new_n27623_, new_n27624_, new_n27625_, new_n27626_, new_n27627_,
    new_n27628_, new_n27629_, new_n27630_, new_n27631_, new_n27632_,
    new_n27633_, new_n27634_, new_n27635_, new_n27636_, new_n27637_,
    new_n27638_, new_n27639_, new_n27640_, new_n27641_, new_n27642_,
    new_n27643_, new_n27644_, new_n27645_, new_n27646_, new_n27647_,
    new_n27648_, new_n27649_, new_n27650_, new_n27651_, new_n27652_,
    new_n27653_, new_n27654_, new_n27655_, new_n27656_, new_n27657_,
    new_n27658_, new_n27659_, new_n27660_, new_n27661_, new_n27662_,
    new_n27663_, new_n27664_, new_n27665_, new_n27666_, new_n27667_,
    new_n27668_, new_n27669_, new_n27670_, new_n27671_, new_n27672_,
    new_n27673_, new_n27674_, new_n27675_, new_n27676_, new_n27677_,
    new_n27678_, new_n27679_, new_n27680_, new_n27681_, new_n27682_,
    new_n27683_, new_n27684_, new_n27685_, new_n27686_, new_n27687_,
    new_n27688_, new_n27689_, new_n27690_, new_n27691_, new_n27692_,
    new_n27693_, new_n27694_, new_n27695_, new_n27696_, new_n27697_,
    new_n27698_, new_n27699_, new_n27700_, new_n27701_, new_n27702_,
    new_n27703_, new_n27704_, new_n27705_, new_n27706_, new_n27707_,
    new_n27708_, new_n27709_, new_n27710_, new_n27711_, new_n27712_,
    new_n27713_, new_n27714_, new_n27715_, new_n27716_, new_n27717_,
    new_n27718_, new_n27719_, new_n27720_, new_n27721_, new_n27722_,
    new_n27723_, new_n27724_, new_n27725_, new_n27726_, new_n27727_,
    new_n27728_, new_n27729_, new_n27730_, new_n27731_, new_n27732_,
    new_n27733_, new_n27734_, new_n27735_, new_n27736_, new_n27737_,
    new_n27738_, new_n27739_, new_n27740_, new_n27741_, new_n27742_,
    new_n27743_, new_n27744_, new_n27745_, new_n27746_, new_n27747_,
    new_n27748_, new_n27749_, new_n27750_, new_n27751_, new_n27752_,
    new_n27753_, new_n27754_, new_n27755_, new_n27756_, new_n27757_,
    new_n27758_, new_n27759_, new_n27760_, new_n27761_, new_n27762_,
    new_n27763_, new_n27764_, new_n27765_, new_n27766_, new_n27767_,
    new_n27768_, new_n27769_, new_n27770_, new_n27771_, new_n27772_,
    new_n27773_, new_n27774_, new_n27775_, new_n27776_, new_n27777_,
    new_n27778_, new_n27779_, new_n27780_, new_n27781_, new_n27782_,
    new_n27783_, new_n27784_, new_n27785_, new_n27786_, new_n27787_,
    new_n27788_, new_n27789_, new_n27790_, new_n27791_, new_n27792_,
    new_n27793_, new_n27794_, new_n27795_, new_n27796_, new_n27797_,
    new_n27798_, new_n27799_, new_n27800_, new_n27801_, new_n27802_,
    new_n27803_, new_n27804_, new_n27805_, new_n27806_, new_n27807_,
    new_n27808_, new_n27809_, new_n27810_, new_n27811_, new_n27812_,
    new_n27813_, new_n27814_, new_n27815_, new_n27816_, new_n27817_,
    new_n27818_, new_n27819_, new_n27820_, new_n27821_, new_n27822_,
    new_n27823_, new_n27824_, new_n27825_, new_n27826_, new_n27827_,
    new_n27828_, new_n27829_, new_n27830_, new_n27831_, new_n27832_,
    new_n27833_, new_n27834_, new_n27835_, new_n27836_, new_n27837_,
    new_n27838_, new_n27839_, new_n27840_, new_n27841_, new_n27842_,
    new_n27843_, new_n27844_, new_n27845_, new_n27846_, new_n27847_,
    new_n27848_, new_n27849_, new_n27850_, new_n27851_, new_n27852_,
    new_n27853_, new_n27854_, new_n27855_, new_n27856_, new_n27857_,
    new_n27858_, new_n27859_, new_n27860_, new_n27861_, new_n27862_,
    new_n27863_, new_n27864_, new_n27865_, new_n27866_, new_n27867_,
    new_n27868_, new_n27869_, new_n27870_, new_n27871_, new_n27872_,
    new_n27873_, new_n27874_, new_n27875_, new_n27876_, new_n27877_,
    new_n27878_, new_n27879_, new_n27880_, new_n27881_, new_n27882_,
    new_n27883_, new_n27884_, new_n27885_, new_n27886_, new_n27887_,
    new_n27888_, new_n27889_, new_n27890_, new_n27891_, new_n27892_,
    new_n27893_, new_n27894_, new_n27895_, new_n27896_, new_n27897_,
    new_n27898_, new_n27899_, new_n27900_, new_n27901_, new_n27902_,
    new_n27903_, new_n27904_, new_n27905_, new_n27906_, new_n27907_,
    new_n27908_, new_n27909_, new_n27910_, new_n27911_, new_n27912_,
    new_n27913_, new_n27914_, new_n27915_, new_n27916_, new_n27917_,
    new_n27918_, new_n27919_, new_n27920_, new_n27921_, new_n27922_,
    new_n27923_, new_n27924_, new_n27925_, new_n27926_, new_n27927_,
    new_n27928_, new_n27929_, new_n27930_, new_n27931_, new_n27932_,
    new_n27933_, new_n27934_, new_n27935_, new_n27936_, new_n27937_,
    new_n27938_, new_n27939_, new_n27940_, new_n27941_, new_n27942_,
    new_n27943_, new_n27944_, new_n27945_, new_n27946_, new_n27947_,
    new_n27948_, new_n27949_, new_n27950_, new_n27951_, new_n27952_,
    new_n27953_, new_n27954_, new_n27955_, new_n27956_, new_n27957_,
    new_n27958_, new_n27959_, new_n27960_, new_n27961_, new_n27962_,
    new_n27963_, new_n27964_, new_n27965_, new_n27966_, new_n27967_,
    new_n27968_, new_n27969_, new_n27970_, new_n27971_, new_n27972_,
    new_n27973_, new_n27974_, new_n27975_, new_n27976_, new_n27977_,
    new_n27978_, new_n27979_, new_n27980_, new_n27981_, new_n27982_,
    new_n27983_, new_n27984_, new_n27985_, new_n27986_, new_n27987_,
    new_n27988_, new_n27989_, new_n27990_, new_n27991_, new_n27992_,
    new_n27993_, new_n27994_, new_n27995_, new_n27996_, new_n27997_,
    new_n27998_, new_n27999_, new_n28000_, new_n28001_, new_n28002_,
    new_n28003_, new_n28004_, new_n28005_, new_n28006_, new_n28007_,
    new_n28008_, new_n28009_, new_n28010_, new_n28011_, new_n28012_,
    new_n28013_, new_n28014_, new_n28015_, new_n28016_, new_n28017_,
    new_n28018_, new_n28019_, new_n28020_, new_n28021_, new_n28022_,
    new_n28023_, new_n28024_, new_n28025_, new_n28026_, new_n28027_,
    new_n28028_, new_n28029_, new_n28030_, new_n28031_, new_n28032_,
    new_n28033_, new_n28034_, new_n28035_, new_n28036_, new_n28037_,
    new_n28038_, new_n28039_, new_n28040_, new_n28041_, new_n28042_,
    new_n28043_, new_n28044_, new_n28045_, new_n28046_, new_n28047_,
    new_n28048_, new_n28049_, new_n28050_, new_n28051_, new_n28052_,
    new_n28053_, new_n28054_, new_n28055_, new_n28056_, new_n28057_,
    new_n28058_, new_n28059_, new_n28060_, new_n28061_, new_n28062_,
    new_n28063_, new_n28064_, new_n28065_, new_n28066_, new_n28067_,
    new_n28068_, new_n28069_, new_n28070_, new_n28071_, new_n28072_,
    new_n28073_, new_n28074_, new_n28075_, new_n28076_, new_n28077_,
    new_n28078_, new_n28079_, new_n28080_, new_n28081_, new_n28082_,
    new_n28083_, new_n28084_, new_n28085_, new_n28086_, new_n28087_,
    new_n28088_, new_n28089_, new_n28090_, new_n28091_, new_n28092_,
    new_n28093_, new_n28094_, new_n28095_, new_n28096_, new_n28097_,
    new_n28098_, new_n28099_, new_n28100_, new_n28101_, new_n28102_,
    new_n28103_, new_n28104_, new_n28105_, new_n28106_, new_n28107_,
    new_n28108_, new_n28109_, new_n28110_, new_n28111_, new_n28112_,
    new_n28113_, new_n28114_, new_n28115_, new_n28116_, new_n28117_,
    new_n28118_, new_n28119_, new_n28120_, new_n28121_, new_n28122_,
    new_n28123_, new_n28124_, new_n28125_, new_n28126_, new_n28127_,
    new_n28128_, new_n28129_, new_n28130_, new_n28131_, new_n28132_,
    new_n28133_, new_n28134_, new_n28135_, new_n28136_, new_n28137_,
    new_n28138_, new_n28139_, new_n28140_, new_n28141_, new_n28142_,
    new_n28143_, new_n28144_, new_n28145_, new_n28146_, new_n28147_,
    new_n28148_, new_n28149_, new_n28150_, new_n28151_, new_n28152_,
    new_n28153_, new_n28154_, new_n28155_, new_n28156_, new_n28157_,
    new_n28158_, new_n28159_, new_n28160_, new_n28161_, new_n28162_,
    new_n28163_, new_n28164_, new_n28165_, new_n28166_, new_n28167_,
    new_n28168_, new_n28169_, new_n28170_, new_n28171_, new_n28172_,
    new_n28173_, new_n28174_, new_n28175_, new_n28176_, new_n28177_,
    new_n28178_, new_n28179_, new_n28180_, new_n28181_, new_n28182_,
    new_n28183_, new_n28184_, new_n28185_, new_n28186_, new_n28187_,
    new_n28188_, new_n28189_, new_n28190_, new_n28191_, new_n28192_,
    new_n28193_, new_n28194_, new_n28195_, new_n28196_, new_n28197_,
    new_n28198_, new_n28199_, new_n28200_, new_n28201_, new_n28202_,
    new_n28203_, new_n28204_, new_n28205_, new_n28206_, new_n28207_,
    new_n28208_, new_n28209_, new_n28210_, new_n28211_, new_n28212_,
    new_n28213_, new_n28214_, new_n28215_, new_n28216_, new_n28217_,
    new_n28218_, new_n28219_, new_n28220_, new_n28221_, new_n28222_,
    new_n28223_, new_n28224_, new_n28225_, new_n28226_, new_n28227_,
    new_n28228_, new_n28229_, new_n28230_, new_n28231_, new_n28232_,
    new_n28233_, new_n28234_, new_n28235_, new_n28236_, new_n28237_,
    new_n28238_, new_n28239_, new_n28240_, new_n28241_, new_n28242_,
    new_n28243_, new_n28244_, new_n28245_, new_n28246_, new_n28247_,
    new_n28248_, new_n28249_, new_n28250_, new_n28251_, new_n28252_,
    new_n28253_, new_n28254_, new_n28255_, new_n28256_, new_n28257_,
    new_n28258_, new_n28259_, new_n28260_, new_n28261_, new_n28262_,
    new_n28263_, new_n28264_, new_n28265_, new_n28266_, new_n28267_,
    new_n28268_, new_n28269_, new_n28270_, new_n28271_, new_n28272_,
    new_n28273_, new_n28274_, new_n28275_, new_n28276_, new_n28277_,
    new_n28278_, new_n28279_, new_n28280_, new_n28281_, new_n28282_,
    new_n28283_, new_n28284_, new_n28285_, new_n28286_, new_n28287_,
    new_n28288_, new_n28289_, new_n28290_, new_n28291_, new_n28292_,
    new_n28293_, new_n28294_, new_n28295_, new_n28296_, new_n28297_,
    new_n28298_, new_n28299_, new_n28300_, new_n28301_, new_n28302_,
    new_n28303_, new_n28304_, new_n28305_, new_n28306_, new_n28307_,
    new_n28308_, new_n28309_, new_n28310_, new_n28311_, new_n28312_,
    new_n28313_, new_n28314_, new_n28315_, new_n28316_, new_n28317_,
    new_n28318_, new_n28319_, new_n28320_, new_n28321_, new_n28322_,
    new_n28323_, new_n28324_, new_n28325_, new_n28326_, new_n28327_,
    new_n28328_, new_n28329_, new_n28330_, new_n28331_, new_n28332_,
    new_n28333_, new_n28334_, new_n28335_, new_n28336_, new_n28337_,
    new_n28338_, new_n28339_, new_n28340_, new_n28341_, new_n28342_,
    new_n28343_, new_n28344_, new_n28345_, new_n28346_, new_n28347_,
    new_n28348_, new_n28349_, new_n28350_, new_n28351_, new_n28352_,
    new_n28353_, new_n28354_, new_n28355_, new_n28356_, new_n28357_,
    new_n28358_, new_n28359_, new_n28360_, new_n28361_, new_n28362_,
    new_n28363_, new_n28364_, new_n28365_, new_n28366_, new_n28367_,
    new_n28368_, new_n28369_, new_n28370_, new_n28371_, new_n28372_,
    new_n28373_, new_n28374_, new_n28375_, new_n28376_, new_n28377_,
    new_n28378_, new_n28379_, new_n28380_, new_n28381_, new_n28382_,
    new_n28383_, new_n28384_, new_n28385_, new_n28386_, new_n28387_,
    new_n28388_, new_n28389_, new_n28390_, new_n28391_, new_n28392_,
    new_n28393_, new_n28394_, new_n28395_, new_n28396_, new_n28397_,
    new_n28398_, new_n28399_, new_n28400_, new_n28401_, new_n28402_,
    new_n28403_, new_n28404_, new_n28405_, new_n28406_, new_n28407_,
    new_n28408_, new_n28409_, new_n28410_, new_n28411_, new_n28412_,
    new_n28413_, new_n28414_, new_n28415_, new_n28416_, new_n28417_,
    new_n28418_, new_n28419_, new_n28420_, new_n28421_, new_n28422_,
    new_n28423_, new_n28424_, new_n28425_, new_n28426_, new_n28427_,
    new_n28428_, new_n28429_, new_n28430_, new_n28431_, new_n28432_,
    new_n28433_, new_n28434_, new_n28435_, new_n28436_, new_n28437_,
    new_n28438_, new_n28439_, new_n28440_, new_n28441_, new_n28442_,
    new_n28443_, new_n28444_, new_n28445_, new_n28446_, new_n28447_,
    new_n28448_, new_n28449_, new_n28450_, new_n28451_, new_n28452_,
    new_n28453_, new_n28454_, new_n28455_, new_n28456_, new_n28457_,
    new_n28458_, new_n28459_, new_n28460_, new_n28461_, new_n28462_,
    new_n28463_, new_n28464_, new_n28465_, new_n28466_, new_n28467_,
    new_n28468_, new_n28469_, new_n28470_, new_n28471_, new_n28472_,
    new_n28473_, new_n28474_, new_n28475_, new_n28476_, new_n28477_,
    new_n28478_, new_n28479_, new_n28480_, new_n28481_, new_n28482_,
    new_n28483_, new_n28484_, new_n28485_, new_n28486_, new_n28487_,
    new_n28488_, new_n28489_, new_n28490_, new_n28491_, new_n28492_,
    new_n28493_, new_n28494_, new_n28495_, new_n28496_, new_n28497_,
    new_n28498_, new_n28499_, new_n28500_, new_n28501_, new_n28502_,
    new_n28503_, new_n28504_, new_n28505_, new_n28506_, new_n28507_,
    new_n28508_, new_n28509_, new_n28510_, new_n28511_, new_n28512_,
    new_n28513_, new_n28514_, new_n28515_, new_n28516_, new_n28517_,
    new_n28518_, new_n28519_, new_n28520_, new_n28521_, new_n28522_,
    new_n28523_, new_n28524_, new_n28525_, new_n28526_, new_n28527_,
    new_n28528_, new_n28529_, new_n28530_, new_n28531_, new_n28532_,
    new_n28533_, new_n28534_, new_n28535_, new_n28536_, new_n28537_,
    new_n28538_, new_n28539_, new_n28540_, new_n28541_, new_n28542_,
    new_n28543_, new_n28544_, new_n28545_, new_n28546_, new_n28547_,
    new_n28548_, new_n28549_, new_n28550_, new_n28551_, new_n28552_,
    new_n28553_, new_n28554_, new_n28555_, new_n28556_, new_n28557_,
    new_n28558_, new_n28559_, new_n28560_, new_n28561_, new_n28562_,
    new_n28563_, new_n28564_, new_n28565_, new_n28566_, new_n28567_,
    new_n28568_, new_n28569_, new_n28570_, new_n28571_, new_n28572_,
    new_n28573_, new_n28574_, new_n28575_, new_n28576_, new_n28577_,
    new_n28578_, new_n28579_, new_n28580_, new_n28581_, new_n28582_,
    new_n28583_, new_n28584_, new_n28585_, new_n28586_, new_n28587_,
    new_n28588_, new_n28589_, new_n28590_, new_n28591_, new_n28592_,
    new_n28593_, new_n28594_, new_n28595_, new_n28596_, new_n28597_,
    new_n28598_, new_n28599_, new_n28600_, new_n28601_, new_n28602_,
    new_n28603_, new_n28604_, new_n28605_, new_n28606_, new_n28607_,
    new_n28608_, new_n28609_, new_n28610_, new_n28611_, new_n28612_,
    new_n28613_, new_n28614_, new_n28615_, new_n28616_, new_n28617_,
    new_n28618_, new_n28619_, new_n28620_, new_n28621_, new_n28622_,
    new_n28623_, new_n28624_, new_n28625_, new_n28626_, new_n28627_,
    new_n28628_, new_n28629_, new_n28630_, new_n28631_, new_n28632_,
    new_n28633_, new_n28634_, new_n28635_, new_n28636_, new_n28637_,
    new_n28638_, new_n28639_, new_n28640_, new_n28641_, new_n28642_,
    new_n28643_, new_n28644_, new_n28645_, new_n28646_, new_n28647_,
    new_n28648_, new_n28649_, new_n28650_, new_n28651_, new_n28652_,
    new_n28653_, new_n28654_, new_n28655_, new_n28656_, new_n28657_,
    new_n28658_, new_n28659_, new_n28660_, new_n28661_, new_n28662_,
    new_n28663_, new_n28664_, new_n28665_, new_n28666_, new_n28667_,
    new_n28668_, new_n28669_, new_n28670_, new_n28671_, new_n28672_,
    new_n28673_, new_n28674_, new_n28675_, new_n28676_, new_n28677_,
    new_n28678_, new_n28679_, new_n28680_, new_n28681_, new_n28682_,
    new_n28683_, new_n28684_, new_n28685_, new_n28686_, new_n28687_,
    new_n28688_, new_n28689_, new_n28690_, new_n28691_, new_n28692_,
    new_n28693_, new_n28694_, new_n28695_, new_n28696_, new_n28697_,
    new_n28698_, new_n28699_, new_n28700_, new_n28701_, new_n28702_,
    new_n28703_, new_n28704_, new_n28705_, new_n28706_, new_n28707_,
    new_n28708_, new_n28709_, new_n28710_, new_n28711_, new_n28712_,
    new_n28713_, new_n28714_, new_n28715_, new_n28716_, new_n28717_,
    new_n28718_, new_n28719_, new_n28720_, new_n28721_, new_n28722_,
    new_n28723_, new_n28724_, new_n28725_, new_n28726_, new_n28727_,
    new_n28728_, new_n28729_, new_n28730_, new_n28731_, new_n28732_,
    new_n28733_, new_n28734_, new_n28735_, new_n28736_, new_n28737_,
    new_n28738_, new_n28739_, new_n28740_, new_n28741_, new_n28742_,
    new_n28743_, new_n28744_, new_n28745_, new_n28746_, new_n28747_,
    new_n28748_, new_n28749_, new_n28750_, new_n28751_, new_n28752_,
    new_n28753_, new_n28754_, new_n28755_, new_n28756_, new_n28757_,
    new_n28758_, new_n28759_, new_n28760_, new_n28761_, new_n28762_,
    new_n28763_, new_n28764_, new_n28765_, new_n28766_, new_n28767_,
    new_n28768_, new_n28769_, new_n28770_, new_n28771_, new_n28772_,
    new_n28773_, new_n28774_, new_n28775_, new_n28776_, new_n28777_,
    new_n28778_, new_n28779_, new_n28780_, new_n28781_, new_n28782_,
    new_n28783_, new_n28784_, new_n28785_, new_n28786_, new_n28787_,
    new_n28788_, new_n28789_, new_n28790_, new_n28791_, new_n28792_,
    new_n28793_, new_n28794_, new_n28795_, new_n28796_, new_n28797_,
    new_n28798_, new_n28799_, new_n28800_, new_n28801_, new_n28802_,
    new_n28803_, new_n28804_, new_n28805_, new_n28806_, new_n28807_,
    new_n28808_, new_n28809_, new_n28810_, new_n28811_, new_n28812_,
    new_n28813_, new_n28814_, new_n28815_, new_n28816_, new_n28817_,
    new_n28818_, new_n28819_, new_n28820_, new_n28821_, new_n28822_,
    new_n28823_, new_n28824_, new_n28825_, new_n28826_, new_n28827_,
    new_n28828_, new_n28829_, new_n28830_, new_n28831_, new_n28832_,
    new_n28833_, new_n28834_, new_n28835_, new_n28836_, new_n28837_,
    new_n28838_, new_n28839_, new_n28840_, new_n28841_, new_n28842_,
    new_n28843_, new_n28844_, new_n28845_, new_n28846_, new_n28847_,
    new_n28848_, new_n28849_, new_n28850_, new_n28851_, new_n28852_,
    new_n28853_, new_n28854_, new_n28855_, new_n28856_, new_n28857_,
    new_n28858_, new_n28859_, new_n28860_, new_n28861_, new_n28862_,
    new_n28863_, new_n28864_, new_n28865_, new_n28866_, new_n28867_,
    new_n28868_, new_n28869_, new_n28870_, new_n28871_, new_n28872_,
    new_n28873_, new_n28874_, new_n28875_, new_n28876_, new_n28877_,
    new_n28878_, new_n28879_, new_n28880_, new_n28881_, new_n28882_,
    new_n28883_, new_n28884_, new_n28885_, new_n28886_, new_n28887_,
    new_n28888_, new_n28889_, new_n28890_, new_n28891_, new_n28892_,
    new_n28893_, new_n28894_, new_n28895_, new_n28896_, new_n28897_,
    new_n28898_, new_n28899_, new_n28900_, new_n28901_, new_n28902_,
    new_n28903_, new_n28904_, new_n28905_, new_n28906_, new_n28907_,
    new_n28908_, new_n28909_, new_n28910_, new_n28911_, new_n28912_,
    new_n28913_, new_n28914_, new_n28915_, new_n28916_, new_n28917_,
    new_n28918_, new_n28919_, new_n28920_, new_n28921_, new_n28922_,
    new_n28923_, new_n28924_, new_n28925_, new_n28926_, new_n28927_,
    new_n28928_, new_n28929_, new_n28930_, new_n28931_, new_n28932_,
    new_n28933_, new_n28934_, new_n28935_, new_n28936_, new_n28937_,
    new_n28938_, new_n28939_, new_n28940_, new_n28941_, new_n28942_,
    new_n28943_, new_n28944_, new_n28945_, new_n28946_, new_n28947_,
    new_n28948_, new_n28949_, new_n28950_, new_n28951_, new_n28952_,
    new_n28953_, new_n28954_, new_n28955_, new_n28956_, new_n28957_,
    new_n28958_, new_n28959_, new_n28960_, new_n28961_, new_n28962_,
    new_n28963_, new_n28964_, new_n28965_, new_n28966_, new_n28967_,
    new_n28968_, new_n28969_, new_n28970_, new_n28971_, new_n28972_,
    new_n28973_, new_n28974_, new_n28975_, new_n28976_, new_n28977_,
    new_n28978_, new_n28979_, new_n28980_, new_n28981_, new_n28982_,
    new_n28983_, new_n28984_, new_n28985_, new_n28986_, new_n28987_,
    new_n28988_, new_n28989_, new_n28990_, new_n28991_, new_n28992_,
    new_n28993_, new_n28994_, new_n28995_, new_n28996_, new_n28997_,
    new_n28998_, new_n28999_, new_n29000_, new_n29001_, new_n29002_,
    new_n29003_, new_n29004_, new_n29005_, new_n29006_, new_n29007_,
    new_n29008_, new_n29009_, new_n29010_, new_n29011_, new_n29012_,
    new_n29013_, new_n29014_, new_n29015_, new_n29016_, new_n29017_,
    new_n29018_, new_n29019_, new_n29020_, new_n29021_, new_n29022_,
    new_n29023_, new_n29024_, new_n29025_, new_n29026_, new_n29027_,
    new_n29028_, new_n29029_, new_n29030_, new_n29031_, new_n29032_,
    new_n29033_, new_n29034_, new_n29035_, new_n29036_, new_n29037_,
    new_n29038_, new_n29039_, new_n29040_, new_n29041_, new_n29042_,
    new_n29043_, new_n29044_, new_n29045_, new_n29046_, new_n29047_,
    new_n29048_, new_n29049_, new_n29050_, new_n29051_, new_n29052_,
    new_n29053_, new_n29054_, new_n29055_, new_n29056_, new_n29057_,
    new_n29058_, new_n29059_, new_n29060_, new_n29061_, new_n29062_,
    new_n29063_, new_n29064_, new_n29065_, new_n29066_, new_n29067_,
    new_n29068_, new_n29069_, new_n29070_, new_n29071_, new_n29072_,
    new_n29073_, new_n29074_, new_n29075_, new_n29076_, new_n29077_,
    new_n29078_, new_n29079_, new_n29080_, new_n29081_, new_n29082_,
    new_n29083_, new_n29084_, new_n29085_, new_n29086_, new_n29087_,
    new_n29088_, new_n29089_, new_n29090_, new_n29091_, new_n29092_,
    new_n29093_, new_n29094_, new_n29095_, new_n29096_, new_n29097_,
    new_n29098_, new_n29099_, new_n29100_, new_n29101_, new_n29102_,
    new_n29103_, new_n29104_, new_n29105_, new_n29106_, new_n29107_,
    new_n29108_, new_n29109_, new_n29110_, new_n29111_, new_n29112_,
    new_n29113_, new_n29114_, new_n29115_, new_n29116_, new_n29117_,
    new_n29118_, new_n29119_, new_n29120_, new_n29121_, new_n29122_,
    new_n29123_, new_n29124_, new_n29125_, new_n29126_, new_n29127_,
    new_n29128_, new_n29129_, new_n29130_, new_n29131_, new_n29132_,
    new_n29133_, new_n29134_, new_n29135_, new_n29136_, new_n29137_,
    new_n29138_, new_n29139_, new_n29140_, new_n29141_, new_n29142_,
    new_n29143_, new_n29144_, new_n29145_, new_n29146_, new_n29147_,
    new_n29148_, new_n29149_, new_n29150_, new_n29151_, new_n29152_,
    new_n29153_, new_n29154_, new_n29155_, new_n29156_, new_n29157_,
    new_n29158_, new_n29159_, new_n29160_, new_n29161_, new_n29162_,
    new_n29163_, new_n29164_, new_n29165_, new_n29166_, new_n29167_,
    new_n29168_, new_n29169_, new_n29170_, new_n29171_, new_n29172_,
    new_n29173_, new_n29174_, new_n29175_, new_n29176_, new_n29177_,
    new_n29178_, new_n29179_, new_n29180_, new_n29181_, new_n29182_,
    new_n29183_, new_n29184_, new_n29185_, new_n29186_, new_n29187_,
    new_n29188_, new_n29189_, new_n29190_, new_n29191_, new_n29192_,
    new_n29193_, new_n29194_, new_n29195_, new_n29196_, new_n29197_,
    new_n29198_, new_n29199_, new_n29200_, new_n29201_, new_n29202_,
    new_n29203_, new_n29204_, new_n29205_, new_n29206_, new_n29207_,
    new_n29208_, new_n29209_, new_n29210_, new_n29211_, new_n29212_,
    new_n29213_, new_n29214_, new_n29215_, new_n29216_, new_n29217_,
    new_n29218_, new_n29219_, new_n29220_, new_n29221_, new_n29222_,
    new_n29223_, new_n29224_, new_n29225_, new_n29226_, new_n29227_,
    new_n29228_, new_n29229_, new_n29230_, new_n29231_, new_n29232_,
    new_n29233_, new_n29234_, new_n29235_, new_n29236_, new_n29237_,
    new_n29238_, new_n29239_, new_n29240_, new_n29241_, new_n29242_,
    new_n29243_, new_n29244_, new_n29245_, new_n29246_, new_n29247_,
    new_n29248_, new_n29249_, new_n29250_, new_n29251_, new_n29252_,
    new_n29253_, new_n29254_, new_n29255_, new_n29256_, new_n29257_,
    new_n29258_, new_n29259_, new_n29260_, new_n29261_, new_n29262_,
    new_n29263_, new_n29264_, new_n29265_, new_n29266_, new_n29267_,
    new_n29268_, new_n29269_, new_n29270_, new_n29271_, new_n29272_,
    new_n29273_, new_n29274_, new_n29275_, new_n29276_, new_n29277_,
    new_n29278_, new_n29279_, new_n29280_, new_n29281_, new_n29282_,
    new_n29283_, new_n29284_, new_n29285_, new_n29286_, new_n29287_,
    new_n29288_, new_n29289_, new_n29290_, new_n29291_, new_n29292_,
    new_n29293_, new_n29294_, new_n29295_, new_n29296_, new_n29297_,
    new_n29298_, new_n29299_, new_n29300_, new_n29301_, new_n29302_,
    new_n29303_, new_n29304_, new_n29305_, new_n29306_, new_n29307_,
    new_n29308_, new_n29309_, new_n29310_, new_n29311_, new_n29312_,
    new_n29313_, new_n29314_, new_n29315_, new_n29316_, new_n29317_,
    new_n29318_, new_n29319_, new_n29320_, new_n29321_, new_n29322_,
    new_n29323_, new_n29324_, new_n29325_, new_n29326_, new_n29327_,
    new_n29328_, new_n29329_, new_n29330_, new_n29331_, new_n29332_,
    new_n29333_, new_n29334_, new_n29335_, new_n29336_, new_n29337_,
    new_n29338_, new_n29339_, new_n29340_, new_n29341_, new_n29342_,
    new_n29343_, new_n29344_, new_n29345_, new_n29346_, new_n29347_,
    new_n29348_, new_n29349_, new_n29350_, new_n29351_, new_n29352_,
    new_n29353_, new_n29354_, new_n29355_, new_n29356_, new_n29357_,
    new_n29358_, new_n29359_, new_n29360_, new_n29361_, new_n29362_,
    new_n29363_, new_n29364_, new_n29365_, new_n29366_, new_n29367_,
    new_n29368_, new_n29369_, new_n29370_, new_n29371_, new_n29372_,
    new_n29373_, new_n29374_, new_n29375_, new_n29376_, new_n29377_,
    new_n29378_, new_n29379_, new_n29380_, new_n29381_, new_n29382_,
    new_n29383_, new_n29384_, new_n29385_, new_n29386_, new_n29387_,
    new_n29388_, new_n29389_, new_n29390_, new_n29391_, new_n29392_,
    new_n29393_, new_n29394_, new_n29395_, new_n29396_, new_n29397_,
    new_n29398_, new_n29399_, new_n29400_, new_n29401_, new_n29402_,
    new_n29403_, new_n29404_, new_n29405_, new_n29406_, new_n29407_,
    new_n29408_, new_n29409_, new_n29410_, new_n29411_, new_n29412_,
    new_n29413_, new_n29414_, new_n29415_, new_n29416_, new_n29417_,
    new_n29418_, new_n29419_, new_n29420_, new_n29421_, new_n29422_,
    new_n29423_, new_n29424_, new_n29425_, new_n29426_, new_n29427_,
    new_n29428_, new_n29429_, new_n29430_, new_n29431_, new_n29432_,
    new_n29433_, new_n29434_, new_n29435_, new_n29436_, new_n29437_,
    new_n29438_, new_n29439_, new_n29440_, new_n29441_, new_n29442_,
    new_n29443_, new_n29444_, new_n29445_, new_n29446_, new_n29447_,
    new_n29448_, new_n29449_, new_n29450_, new_n29451_, new_n29452_,
    new_n29453_, new_n29454_, new_n29455_, new_n29456_, new_n29457_,
    new_n29458_, new_n29459_, new_n29460_, new_n29461_, new_n29462_,
    new_n29463_, new_n29464_, new_n29465_, new_n29466_, new_n29467_,
    new_n29468_, new_n29469_, new_n29470_, new_n29471_, new_n29472_,
    new_n29473_, new_n29474_, new_n29475_, new_n29476_, new_n29477_,
    new_n29478_, new_n29479_, new_n29480_, new_n29481_, new_n29482_,
    new_n29483_, new_n29484_, new_n29485_, new_n29486_, new_n29487_,
    new_n29488_, new_n29489_, new_n29490_, new_n29491_, new_n29492_,
    new_n29493_, new_n29494_, new_n29495_, new_n29496_, new_n29497_,
    new_n29498_, new_n29499_, new_n29500_, new_n29501_, new_n29502_,
    new_n29503_, new_n29504_, new_n29505_, new_n29506_, new_n29507_,
    new_n29508_, new_n29509_, new_n29510_, new_n29511_, new_n29512_,
    new_n29513_, new_n29514_, new_n29515_, new_n29516_, new_n29517_,
    new_n29518_, new_n29519_, new_n29520_, new_n29521_, new_n29522_,
    new_n29523_, new_n29524_, new_n29525_, new_n29526_, new_n29527_,
    new_n29528_, new_n29529_, new_n29530_, new_n29531_, new_n29532_,
    new_n29533_, new_n29534_, new_n29535_, new_n29536_, new_n29537_,
    new_n29538_, new_n29539_, new_n29540_, new_n29541_, new_n29542_,
    new_n29543_, new_n29544_, new_n29545_, new_n29546_, new_n29547_,
    new_n29548_, new_n29549_, new_n29550_, new_n29551_, new_n29552_,
    new_n29553_, new_n29554_, new_n29555_, new_n29556_, new_n29557_,
    new_n29558_, new_n29559_, new_n29560_, new_n29561_, new_n29562_,
    new_n29563_, new_n29564_, new_n29565_, new_n29566_, new_n29567_,
    new_n29568_, new_n29569_, new_n29570_, new_n29571_, new_n29572_,
    new_n29573_, new_n29574_, new_n29575_, new_n29576_, new_n29577_,
    new_n29578_, new_n29579_, new_n29580_, new_n29581_, new_n29582_,
    new_n29583_, new_n29584_, new_n29585_, new_n29586_, new_n29587_,
    new_n29588_, new_n29589_, new_n29590_, new_n29591_, new_n29592_,
    new_n29593_, new_n29594_, new_n29595_, new_n29596_, new_n29597_,
    new_n29598_, new_n29599_, new_n29600_, new_n29601_, new_n29602_,
    new_n29603_, new_n29604_, new_n29605_, new_n29606_, new_n29607_,
    new_n29608_, new_n29609_, new_n29610_, new_n29611_, new_n29612_,
    new_n29613_, new_n29614_, new_n29615_, new_n29616_, new_n29617_,
    new_n29618_, new_n29619_, new_n29620_, new_n29621_, new_n29622_,
    new_n29623_, new_n29624_, new_n29625_, new_n29626_, new_n29627_,
    new_n29628_, new_n29629_, new_n29630_, new_n29631_, new_n29632_,
    new_n29633_, new_n29634_, new_n29635_, new_n29636_, new_n29637_,
    new_n29638_, new_n29639_, new_n29640_, new_n29641_, new_n29642_,
    new_n29643_, new_n29644_, new_n29645_, new_n29646_, new_n29647_,
    new_n29648_, new_n29649_, new_n29650_, new_n29651_, new_n29652_,
    new_n29653_, new_n29654_, new_n29655_, new_n29656_, new_n29657_,
    new_n29658_, new_n29659_, new_n29660_, new_n29661_, new_n29662_,
    new_n29663_, new_n29664_, new_n29665_, new_n29666_, new_n29667_,
    new_n29668_, new_n29669_, new_n29670_, new_n29671_, new_n29672_,
    new_n29673_, new_n29674_, new_n29675_, new_n29676_, new_n29677_,
    new_n29678_, new_n29679_, new_n29680_, new_n29681_, new_n29682_,
    new_n29683_, new_n29684_, new_n29685_, new_n29686_, new_n29687_,
    new_n29688_, new_n29689_, new_n29690_, new_n29691_, new_n29692_,
    new_n29693_, new_n29694_, new_n29695_, new_n29696_, new_n29697_,
    new_n29698_, new_n29699_, new_n29700_, new_n29701_, new_n29702_,
    new_n29703_, new_n29704_, new_n29705_, new_n29706_, new_n29707_,
    new_n29708_, new_n29709_, new_n29710_, new_n29711_, new_n29712_,
    new_n29713_, new_n29714_, new_n29715_, new_n29716_, new_n29717_,
    new_n29718_, new_n29719_, new_n29720_, new_n29721_, new_n29722_,
    new_n29723_, new_n29724_, new_n29725_, new_n29726_, new_n29727_,
    new_n29728_, new_n29729_, new_n29730_, new_n29731_, new_n29732_,
    new_n29733_, new_n29734_, new_n29735_, new_n29736_, new_n29737_,
    new_n29738_, new_n29739_, new_n29740_, new_n29741_, new_n29742_,
    new_n29743_, new_n29744_, new_n29745_, new_n29746_, new_n29747_,
    new_n29748_, new_n29749_, new_n29750_, new_n29751_, new_n29752_,
    new_n29753_, new_n29754_, new_n29755_, new_n29756_, new_n29757_,
    new_n29758_, new_n29759_, new_n29760_, new_n29761_, new_n29762_,
    new_n29763_, new_n29764_, new_n29765_, new_n29766_, new_n29767_,
    new_n29768_, new_n29769_, new_n29770_, new_n29771_, new_n29772_,
    new_n29773_, new_n29774_, new_n29775_, new_n29776_, new_n29777_,
    new_n29778_, new_n29779_, new_n29780_, new_n29781_, new_n29782_,
    new_n29783_, new_n29784_, new_n29785_, new_n29786_, new_n29787_,
    new_n29788_, new_n29789_, new_n29790_, new_n29791_, new_n29792_,
    new_n29793_, new_n29794_, new_n29795_, new_n29796_, new_n29797_,
    new_n29798_, new_n29799_, new_n29800_, new_n29801_, new_n29802_,
    new_n29803_, new_n29804_, new_n29805_, new_n29806_, new_n29807_,
    new_n29808_, new_n29809_, new_n29810_, new_n29811_, new_n29812_,
    new_n29813_, new_n29814_, new_n29815_, new_n29816_, new_n29817_,
    new_n29818_, new_n29819_, new_n29820_, new_n29821_, new_n29822_,
    new_n29823_, new_n29824_, new_n29825_, new_n29826_, new_n29827_,
    new_n29828_, new_n29829_, new_n29830_, new_n29831_, new_n29832_,
    new_n29833_, new_n29834_, new_n29835_, new_n29836_, new_n29837_,
    new_n29838_, new_n29839_, new_n29840_, new_n29841_, new_n29842_,
    new_n29843_, new_n29844_, new_n29845_, new_n29846_, new_n29847_,
    new_n29848_, new_n29849_, new_n29850_, new_n29851_, new_n29852_,
    new_n29853_, new_n29854_, new_n29855_, new_n29856_, new_n29857_,
    new_n29858_, new_n29859_, new_n29860_, new_n29861_, new_n29862_,
    new_n29863_, new_n29864_, new_n29865_, new_n29866_, new_n29867_,
    new_n29868_, new_n29869_, new_n29870_, new_n29871_, new_n29872_,
    new_n29873_, new_n29874_, new_n29875_, new_n29876_, new_n29877_,
    new_n29878_, new_n29879_, new_n29880_, new_n29881_, new_n29882_,
    new_n29883_, new_n29884_, new_n29885_, new_n29886_, new_n29887_,
    new_n29888_, new_n29889_, new_n29890_, new_n29891_, new_n29892_,
    new_n29893_, new_n29894_, new_n29895_, new_n29896_, new_n29897_,
    new_n29898_, new_n29899_, new_n29900_, new_n29901_, new_n29902_,
    new_n29903_, new_n29904_, new_n29905_, new_n29906_, new_n29907_,
    new_n29908_, new_n29909_, new_n29910_, new_n29911_, new_n29912_,
    new_n29913_, new_n29914_, new_n29915_, new_n29916_, new_n29917_,
    new_n29918_, new_n29919_, new_n29920_, new_n29921_, new_n29922_,
    new_n29923_, new_n29924_, new_n29925_, new_n29926_, new_n29927_,
    new_n29928_, new_n29929_, new_n29930_, new_n29931_, new_n29932_,
    new_n29933_, new_n29934_, new_n29935_, new_n29936_, new_n29937_,
    new_n29938_, new_n29939_, new_n29940_, new_n29941_, new_n29942_,
    new_n29943_, new_n29944_, new_n29945_, new_n29946_, new_n29947_,
    new_n29948_, new_n29949_, new_n29950_, new_n29951_, new_n29952_,
    new_n29953_, new_n29954_, new_n29955_, new_n29956_, new_n29957_,
    new_n29958_, new_n29959_, new_n29960_, new_n29961_, new_n29962_,
    new_n29963_, new_n29964_, new_n29965_, new_n29966_, new_n29967_,
    new_n29968_, new_n29969_, new_n29970_, new_n29971_, new_n29972_,
    new_n29973_, new_n29974_, new_n29975_, new_n29976_, new_n29977_,
    new_n29978_, new_n29979_, new_n29980_, new_n29981_, new_n29982_,
    new_n29983_, new_n29984_, new_n29985_, new_n29986_, new_n29987_,
    new_n29988_, new_n29989_, new_n29990_, new_n29991_, new_n29992_,
    new_n29993_, new_n29994_, new_n29995_, new_n29996_, new_n29997_,
    new_n29998_, new_n29999_, new_n30000_, new_n30001_, new_n30002_,
    new_n30003_, new_n30004_, new_n30005_, new_n30006_, new_n30007_,
    new_n30008_, new_n30009_, new_n30010_, new_n30011_, new_n30012_,
    new_n30013_, new_n30014_, new_n30015_, new_n30016_, new_n30017_,
    new_n30018_, new_n30019_, new_n30020_, new_n30021_, new_n30022_,
    new_n30023_, new_n30024_, new_n30025_, new_n30026_, new_n30027_,
    new_n30028_, new_n30029_, new_n30030_, new_n30031_, new_n30032_,
    new_n30033_, new_n30034_, new_n30035_, new_n30036_, new_n30037_,
    new_n30038_, new_n30039_, new_n30040_, new_n30041_, new_n30042_,
    new_n30043_, new_n30044_, new_n30045_, new_n30046_, new_n30047_,
    new_n30048_, new_n30049_, new_n30050_, new_n30051_, new_n30052_,
    new_n30053_, new_n30054_, new_n30055_, new_n30056_, new_n30057_,
    new_n30058_, new_n30059_, new_n30060_, new_n30061_, new_n30062_,
    new_n30063_, new_n30064_, new_n30065_, new_n30066_, new_n30067_,
    new_n30068_, new_n30069_, new_n30070_, new_n30071_, new_n30072_,
    new_n30073_, new_n30074_, new_n30075_, new_n30076_, new_n30077_,
    new_n30078_, new_n30079_, new_n30080_, new_n30081_, new_n30082_,
    new_n30083_, new_n30084_, new_n30085_, new_n30086_, new_n30087_,
    new_n30088_, new_n30089_, new_n30090_, new_n30091_, new_n30092_,
    new_n30093_, new_n30094_, new_n30095_, new_n30096_, new_n30097_,
    new_n30098_, new_n30099_, new_n30100_, new_n30101_, new_n30102_,
    new_n30103_, new_n30104_, new_n30105_, new_n30106_, new_n30107_,
    new_n30108_, new_n30109_, new_n30110_, new_n30111_, new_n30112_,
    new_n30113_, new_n30114_, new_n30115_, new_n30116_, new_n30117_,
    new_n30118_, new_n30119_, new_n30120_, new_n30121_, new_n30122_,
    new_n30123_, new_n30124_, new_n30125_, new_n30126_, new_n30127_,
    new_n30128_, new_n30129_, new_n30130_, new_n30131_, new_n30132_,
    new_n30133_, new_n30134_, new_n30135_, new_n30136_, new_n30137_,
    new_n30138_, new_n30139_, new_n30140_, new_n30141_, new_n30142_,
    new_n30143_, new_n30144_, new_n30145_, new_n30146_, new_n30147_,
    new_n30148_, new_n30149_, new_n30150_, new_n30151_, new_n30152_,
    new_n30153_, new_n30154_, new_n30155_, new_n30156_, new_n30157_,
    new_n30158_, new_n30159_, new_n30160_, new_n30161_, new_n30162_,
    new_n30163_, new_n30164_, new_n30165_, new_n30166_, new_n30167_,
    new_n30168_, new_n30169_, new_n30170_, new_n30171_, new_n30172_,
    new_n30173_, new_n30174_, new_n30175_, new_n30176_, new_n30177_,
    new_n30178_, new_n30179_, new_n30180_, new_n30181_, new_n30182_,
    new_n30183_, new_n30184_, new_n30185_, new_n30186_, new_n30187_,
    new_n30188_, new_n30189_, new_n30190_, new_n30191_, new_n30192_,
    new_n30193_, new_n30194_, new_n30195_, new_n30196_, new_n30197_,
    new_n30198_, new_n30199_, new_n30200_, new_n30201_, new_n30202_,
    new_n30203_, new_n30204_, new_n30205_, new_n30206_, new_n30207_,
    new_n30208_, new_n30209_, new_n30210_, new_n30211_, new_n30212_,
    new_n30213_, new_n30214_, new_n30215_, new_n30216_, new_n30217_,
    new_n30218_, new_n30219_, new_n30220_, new_n30221_, new_n30222_,
    new_n30223_, new_n30224_, new_n30225_, new_n30226_, new_n30227_,
    new_n30228_, new_n30229_, new_n30230_, new_n30231_, new_n30232_,
    new_n30233_, new_n30234_, new_n30235_, new_n30236_, new_n30237_,
    new_n30238_, new_n30239_, new_n30240_, new_n30241_, new_n30242_,
    new_n30243_, new_n30244_, new_n30245_, new_n30246_, new_n30247_,
    new_n30248_, new_n30249_, new_n30250_, new_n30251_, new_n30252_,
    new_n30253_, new_n30254_, new_n30255_, new_n30256_, new_n30257_,
    new_n30258_, new_n30259_, new_n30260_, new_n30261_, new_n30262_,
    new_n30263_, new_n30264_, new_n30265_, new_n30266_, new_n30267_,
    new_n30268_, new_n30269_, new_n30270_, new_n30271_, new_n30272_,
    new_n30273_, new_n30274_, new_n30275_, new_n30276_, new_n30277_,
    new_n30278_, new_n30279_, new_n30280_, new_n30281_, new_n30282_,
    new_n30283_, new_n30284_, new_n30285_, new_n30286_, new_n30287_,
    new_n30288_, new_n30289_, new_n30290_, new_n30291_, new_n30292_,
    new_n30293_, new_n30294_, new_n30295_, new_n30296_, new_n30297_,
    new_n30298_, new_n30299_, new_n30300_, new_n30301_, new_n30302_,
    new_n30303_, new_n30304_, new_n30305_, new_n30306_, new_n30307_,
    new_n30308_, new_n30309_, new_n30310_, new_n30311_, new_n30312_,
    new_n30313_, new_n30314_, new_n30315_, new_n30316_, new_n30317_,
    new_n30318_, new_n30319_, new_n30320_, new_n30321_, new_n30322_,
    new_n30323_, new_n30324_, new_n30325_, new_n30326_, new_n30327_,
    new_n30328_, new_n30329_, new_n30330_, new_n30331_, new_n30332_,
    new_n30333_, new_n30334_, new_n30335_, new_n30336_, new_n30337_,
    new_n30338_, new_n30339_, new_n30340_, new_n30341_, new_n30342_,
    new_n30343_, new_n30344_, new_n30345_, new_n30346_, new_n30347_,
    new_n30348_, new_n30349_, new_n30350_, new_n30351_, new_n30352_,
    new_n30353_, new_n30354_, new_n30355_, new_n30356_, new_n30357_,
    new_n30358_, new_n30359_, new_n30360_, new_n30361_, new_n30362_,
    new_n30363_, new_n30364_, new_n30365_, new_n30366_, new_n30367_,
    new_n30368_, new_n30369_, new_n30370_, new_n30371_, new_n30372_,
    new_n30373_, new_n30374_, new_n30375_, new_n30376_, new_n30377_,
    new_n30378_, new_n30379_, new_n30380_, new_n30381_, new_n30382_,
    new_n30383_, new_n30384_, new_n30385_, new_n30386_, new_n30387_,
    new_n30388_, new_n30389_, new_n30390_, new_n30391_, new_n30392_,
    new_n30393_, new_n30394_, new_n30395_, new_n30396_, new_n30397_,
    new_n30398_, new_n30399_, new_n30400_, new_n30401_, new_n30402_,
    new_n30403_, new_n30404_, new_n30405_, new_n30406_, new_n30407_,
    new_n30408_, new_n30409_, new_n30410_, new_n30411_, new_n30412_,
    new_n30413_, new_n30414_, new_n30415_, new_n30416_, new_n30417_,
    new_n30418_, new_n30419_, new_n30420_, new_n30421_, new_n30422_,
    new_n30423_, new_n30424_, new_n30425_, new_n30426_, new_n30427_,
    new_n30428_, new_n30429_, new_n30430_, new_n30431_, new_n30432_,
    new_n30433_, new_n30434_, new_n30435_, new_n30436_, new_n30437_,
    new_n30438_, new_n30439_, new_n30440_, new_n30441_, new_n30442_,
    new_n30443_, new_n30444_, new_n30445_, new_n30446_, new_n30447_,
    new_n30448_, new_n30449_, new_n30450_, new_n30451_, new_n30452_,
    new_n30453_, new_n30454_, new_n30455_, new_n30456_, new_n30457_,
    new_n30458_, new_n30459_, new_n30460_, new_n30461_, new_n30462_,
    new_n30463_, new_n30464_, new_n30465_, new_n30466_, new_n30467_,
    new_n30468_, new_n30469_, new_n30470_, new_n30471_, new_n30472_,
    new_n30473_, new_n30474_, new_n30475_, new_n30476_, new_n30477_,
    new_n30478_, new_n30479_, new_n30480_, new_n30481_, new_n30482_,
    new_n30483_, new_n30484_, new_n30485_, new_n30486_, new_n30487_,
    new_n30488_, new_n30489_, new_n30490_, new_n30491_, new_n30492_,
    new_n30493_, new_n30494_, new_n30495_, new_n30496_, new_n30497_,
    new_n30498_, new_n30499_, new_n30500_, new_n30501_, new_n30502_,
    new_n30503_, new_n30504_, new_n30505_, new_n30506_, new_n30507_,
    new_n30508_, new_n30509_, new_n30510_, new_n30511_, new_n30512_,
    new_n30513_, new_n30514_, new_n30515_, new_n30516_, new_n30517_,
    new_n30518_, new_n30519_, new_n30520_, new_n30521_, new_n30522_,
    new_n30523_, new_n30524_, new_n30525_, new_n30526_, new_n30527_,
    new_n30528_, new_n30529_, new_n30530_, new_n30531_, new_n30532_,
    new_n30533_, new_n30534_, new_n30535_, new_n30536_, new_n30537_,
    new_n30538_, new_n30539_, new_n30540_, new_n30541_, new_n30542_,
    new_n30543_, new_n30544_, new_n30545_, new_n30546_, new_n30547_,
    new_n30548_, new_n30549_, new_n30550_, new_n30551_, new_n30552_,
    new_n30553_, new_n30554_, new_n30555_, new_n30556_, new_n30557_,
    new_n30558_, new_n30559_, new_n30560_, new_n30561_, new_n30562_,
    new_n30563_, new_n30564_, new_n30565_, new_n30566_, new_n30567_,
    new_n30568_, new_n30569_, new_n30570_, new_n30571_, new_n30572_,
    new_n30573_, new_n30574_, new_n30575_, new_n30576_, new_n30577_,
    new_n30578_, new_n30579_, new_n30580_, new_n30581_, new_n30582_,
    new_n30583_, new_n30584_, new_n30585_, new_n30586_, new_n30587_,
    new_n30588_, new_n30589_, new_n30590_, new_n30591_, new_n30592_,
    new_n30593_, new_n30594_, new_n30595_, new_n30596_, new_n30597_,
    new_n30598_, new_n30599_, new_n30600_, new_n30601_, new_n30602_,
    new_n30603_, new_n30604_, new_n30605_, new_n30606_, new_n30607_,
    new_n30608_, new_n30609_, new_n30610_, new_n30611_, new_n30612_,
    new_n30613_, new_n30614_, new_n30615_, new_n30616_, new_n30617_,
    new_n30618_, new_n30619_, new_n30620_, new_n30621_, new_n30622_,
    new_n30623_, new_n30624_, new_n30625_, new_n30626_, new_n30627_,
    new_n30628_, new_n30629_, new_n30630_, new_n30631_, new_n30632_,
    new_n30633_, new_n30634_, new_n30635_, new_n30636_, new_n30637_,
    new_n30638_, new_n30639_, new_n30640_, new_n30641_, new_n30642_,
    new_n30643_, new_n30644_, new_n30645_, new_n30646_, new_n30647_,
    new_n30648_, new_n30649_, new_n30650_, new_n30651_, new_n30652_,
    new_n30653_, new_n30654_, new_n30655_, new_n30656_, new_n30657_,
    new_n30658_, new_n30659_, new_n30660_, new_n30661_, new_n30662_,
    new_n30663_, new_n30664_, new_n30665_, new_n30666_, new_n30667_,
    new_n30668_, new_n30669_, new_n30670_, new_n30671_, new_n30672_,
    new_n30673_, new_n30674_, new_n30675_, new_n30676_, new_n30677_,
    new_n30678_, new_n30679_, new_n30680_, new_n30681_, new_n30682_,
    new_n30683_, new_n30684_, new_n30685_, new_n30686_, new_n30687_,
    new_n30688_, new_n30689_, new_n30690_, new_n30691_, new_n30692_,
    new_n30693_, new_n30694_, new_n30695_, new_n30696_, new_n30697_,
    new_n30698_, new_n30699_, new_n30700_, new_n30701_, new_n30702_,
    new_n30703_, new_n30704_, new_n30705_, new_n30706_, new_n30707_,
    new_n30708_, new_n30709_, new_n30710_, new_n30711_, new_n30712_,
    new_n30713_, new_n30714_, new_n30715_, new_n30716_, new_n30717_,
    new_n30718_, new_n30719_, new_n30720_, new_n30721_, new_n30722_,
    new_n30723_, new_n30724_, new_n30725_, new_n30726_, new_n30727_,
    new_n30728_, new_n30729_, new_n30730_, new_n30731_, new_n30732_,
    new_n30733_, new_n30734_, new_n30735_, new_n30736_, new_n30737_,
    new_n30738_, new_n30739_, new_n30740_, new_n30741_, new_n30742_,
    new_n30743_, new_n30744_, new_n30745_, new_n30746_, new_n30747_,
    new_n30748_, new_n30749_, new_n30750_, new_n30751_, new_n30752_,
    new_n30753_, new_n30754_, new_n30755_, new_n30756_, new_n30757_,
    new_n30758_, new_n30759_, new_n30760_, new_n30761_, new_n30762_,
    new_n30763_, new_n30764_, new_n30765_, new_n30766_, new_n30767_,
    new_n30768_, new_n30769_, new_n30770_, new_n30771_, new_n30772_,
    new_n30773_, new_n30774_, new_n30775_, new_n30776_, new_n30777_,
    new_n30778_, new_n30779_, new_n30780_, new_n30781_, new_n30782_,
    new_n30783_, new_n30784_, new_n30785_, new_n30786_, new_n30787_,
    new_n30788_, new_n30789_, new_n30790_, new_n30791_, new_n30792_,
    new_n30793_, new_n30794_, new_n30795_, new_n30796_, new_n30797_,
    new_n30798_, new_n30799_, new_n30800_, new_n30801_, new_n30802_,
    new_n30803_, new_n30804_, new_n30805_, new_n30806_, new_n30807_,
    new_n30808_, new_n30809_, new_n30810_, new_n30811_, new_n30812_,
    new_n30813_, new_n30814_, new_n30815_, new_n30816_, new_n30817_,
    new_n30818_, new_n30819_, new_n30820_, new_n30821_, new_n30822_,
    new_n30823_, new_n30824_, new_n30825_, new_n30826_, new_n30827_,
    new_n30828_, new_n30829_, new_n30830_, new_n30831_, new_n30832_,
    new_n30833_, new_n30834_, new_n30835_, new_n30836_, new_n30837_,
    new_n30838_, new_n30839_, new_n30840_, new_n30841_, new_n30842_,
    new_n30843_, new_n30844_, new_n30845_, new_n30846_, new_n30847_,
    new_n30848_, new_n30849_, new_n30850_, new_n30851_, new_n30852_,
    new_n30853_, new_n30854_, new_n30855_, new_n30856_, new_n30857_,
    new_n30858_, new_n30859_, new_n30860_, new_n30861_, new_n30862_,
    new_n30863_, new_n30864_, new_n30865_, new_n30866_, new_n30867_,
    new_n30868_, new_n30869_, new_n30870_, new_n30871_, new_n30872_,
    new_n30873_, new_n30874_, new_n30875_, new_n30876_, new_n30877_,
    new_n30878_, new_n30879_, new_n30880_, new_n30881_, new_n30882_,
    new_n30883_, new_n30884_, new_n30885_, new_n30886_, new_n30887_,
    new_n30888_, new_n30889_, new_n30890_, new_n30891_, new_n30892_,
    new_n30893_, new_n30894_, new_n30895_, new_n30896_, new_n30897_,
    new_n30898_, new_n30899_, new_n30900_, new_n30901_, new_n30902_,
    new_n30903_, new_n30904_, new_n30905_, new_n30906_, new_n30907_,
    new_n30908_, new_n30909_, new_n30910_, new_n30911_, new_n30912_,
    new_n30913_, new_n30914_, new_n30915_, new_n30916_, new_n30917_,
    new_n30918_, new_n30919_, new_n30920_, new_n30921_, new_n30922_,
    new_n30923_, new_n30924_, new_n30925_, new_n30926_, new_n30927_,
    new_n30928_, new_n30929_, new_n30930_, new_n30931_, new_n30932_,
    new_n30933_, new_n30934_, new_n30935_, new_n30936_, new_n30937_,
    new_n30938_, new_n30939_, new_n30940_, new_n30941_, new_n30942_,
    new_n30943_, new_n30944_, new_n30945_, new_n30946_, new_n30947_,
    new_n30948_, new_n30949_, new_n30950_, new_n30951_, new_n30952_,
    new_n30953_, new_n30954_, new_n30955_, new_n30956_, new_n30957_,
    new_n30958_, new_n30959_, new_n30960_, new_n30961_, new_n30962_,
    new_n30963_, new_n30964_, new_n30965_, new_n30966_, new_n30967_,
    new_n30968_, new_n30969_, new_n30970_, new_n30971_, new_n30972_,
    new_n30973_, new_n30974_, new_n30975_, new_n30976_, new_n30977_,
    new_n30978_, new_n30979_, new_n30980_, new_n30981_, new_n30982_,
    new_n30983_, new_n30984_, new_n30985_, new_n30986_, new_n30987_,
    new_n30988_, new_n30989_, new_n30990_, new_n30991_, new_n30992_,
    new_n30993_, new_n30994_, new_n30995_, new_n30996_, new_n30997_,
    new_n30998_, new_n30999_, new_n31000_, new_n31001_, new_n31002_,
    new_n31003_, new_n31004_, new_n31005_, new_n31006_, new_n31007_,
    new_n31008_, new_n31009_, new_n31010_, new_n31011_, new_n31012_,
    new_n31013_, new_n31014_, new_n31015_, new_n31016_, new_n31017_,
    new_n31018_, new_n31019_, new_n31020_, new_n31021_, new_n31022_,
    new_n31023_, new_n31024_, new_n31025_, new_n31026_, new_n31027_,
    new_n31028_, new_n31029_, new_n31030_, new_n31031_, new_n31032_,
    new_n31033_, new_n31034_, new_n31035_, new_n31036_, new_n31037_,
    new_n31038_, new_n31039_, new_n31040_, new_n31041_, new_n31042_,
    new_n31043_, new_n31044_, new_n31045_, new_n31046_, new_n31047_,
    new_n31048_, new_n31049_, new_n31050_, new_n31051_, new_n31052_,
    new_n31053_, new_n31054_, new_n31055_, new_n31056_, new_n31057_,
    new_n31058_, new_n31059_, new_n31060_, new_n31061_, new_n31062_,
    new_n31063_, new_n31064_, new_n31065_, new_n31066_, new_n31067_,
    new_n31068_, new_n31069_, new_n31070_, new_n31071_, new_n31072_,
    new_n31073_, new_n31074_, new_n31075_, new_n31076_, new_n31077_,
    new_n31078_, new_n31079_, new_n31080_, new_n31081_, new_n31082_,
    new_n31083_, new_n31084_, new_n31085_, new_n31086_, new_n31087_,
    new_n31088_, new_n31089_, new_n31090_, new_n31091_, new_n31092_,
    new_n31093_, new_n31094_, new_n31095_, new_n31096_, new_n31097_,
    new_n31098_, new_n31099_, new_n31100_, new_n31101_, new_n31102_,
    new_n31103_, new_n31104_, new_n31105_, new_n31106_, new_n31107_,
    new_n31108_, new_n31109_, new_n31110_, new_n31111_, new_n31112_,
    new_n31113_, new_n31114_, new_n31115_, new_n31116_, new_n31117_,
    new_n31118_, new_n31119_, new_n31120_, new_n31121_, new_n31122_,
    new_n31123_, new_n31124_, new_n31125_, new_n31126_, new_n31127_,
    new_n31128_, new_n31129_, new_n31130_, new_n31131_, new_n31132_,
    new_n31133_, new_n31134_, new_n31135_, new_n31136_, new_n31137_,
    new_n31138_, new_n31139_, new_n31140_, new_n31141_, new_n31142_,
    new_n31143_, new_n31144_, new_n31145_, new_n31146_, new_n31147_,
    new_n31148_, new_n31149_, new_n31150_, new_n31151_, new_n31152_,
    new_n31153_, new_n31154_, new_n31155_, new_n31156_, new_n31157_,
    new_n31158_, new_n31159_, new_n31160_, new_n31161_, new_n31162_,
    new_n31163_, new_n31164_, new_n31165_, new_n31166_, new_n31167_,
    new_n31168_, new_n31169_, new_n31170_, new_n31171_, new_n31172_,
    new_n31173_, new_n31174_, new_n31175_, new_n31176_, new_n31177_,
    new_n31178_, new_n31179_, new_n31180_, new_n31181_, new_n31182_,
    new_n31183_, new_n31184_, new_n31185_, new_n31186_, new_n31187_,
    new_n31188_, new_n31189_, new_n31190_, new_n31191_, new_n31192_,
    new_n31193_, new_n31194_, new_n31195_, new_n31196_, new_n31197_,
    new_n31198_, new_n31199_, new_n31200_, new_n31201_, new_n31202_,
    new_n31203_, new_n31204_, new_n31205_, new_n31206_, new_n31207_,
    new_n31208_, new_n31209_, new_n31210_, new_n31211_, new_n31212_,
    new_n31213_, new_n31214_, new_n31215_, new_n31216_, new_n31217_,
    new_n31218_, new_n31219_, new_n31220_, new_n31221_, new_n31222_,
    new_n31223_, new_n31224_, new_n31225_, new_n31226_, new_n31227_,
    new_n31228_, new_n31229_, new_n31230_, new_n31231_, new_n31232_,
    new_n31233_, new_n31234_, new_n31235_, new_n31236_, new_n31237_,
    new_n31238_, new_n31239_, new_n31240_, new_n31241_, new_n31242_,
    new_n31243_, new_n31244_, new_n31245_, new_n31246_, new_n31247_,
    new_n31248_, new_n31249_, new_n31250_, new_n31251_, new_n31252_,
    new_n31253_, new_n31254_, new_n31255_, new_n31256_, new_n31257_,
    new_n31258_, new_n31259_, new_n31260_, new_n31261_, new_n31262_,
    new_n31263_, new_n31264_, new_n31265_, new_n31266_, new_n31267_,
    new_n31268_, new_n31269_, new_n31270_, new_n31271_, new_n31272_,
    new_n31273_, new_n31274_, new_n31275_, new_n31276_, new_n31277_,
    new_n31278_, new_n31279_, new_n31280_, new_n31281_, new_n31282_,
    new_n31283_, new_n31284_, new_n31285_, new_n31286_, new_n31287_,
    new_n31288_, new_n31289_, new_n31290_, new_n31291_, new_n31292_,
    new_n31293_, new_n31294_, new_n31295_, new_n31296_, new_n31297_,
    new_n31298_, new_n31299_, new_n31300_, new_n31301_, new_n31302_,
    new_n31303_, new_n31304_, new_n31305_, new_n31306_, new_n31307_,
    new_n31308_, new_n31309_, new_n31310_, new_n31311_, new_n31312_,
    new_n31313_, new_n31314_, new_n31315_, new_n31316_, new_n31317_,
    new_n31318_, new_n31319_, new_n31320_, new_n31321_, new_n31322_,
    new_n31323_, new_n31324_, new_n31325_, new_n31326_, new_n31327_,
    new_n31328_, new_n31329_, new_n31330_, new_n31331_, new_n31332_,
    new_n31333_, new_n31334_, new_n31335_, new_n31336_, new_n31337_,
    new_n31338_, new_n31339_, new_n31340_, new_n31341_, new_n31342_,
    new_n31343_, new_n31344_, new_n31345_, new_n31346_, new_n31347_,
    new_n31348_, new_n31349_, new_n31350_, new_n31351_, new_n31352_,
    new_n31353_, new_n31354_, new_n31355_, new_n31356_, new_n31357_,
    new_n31358_, new_n31359_, new_n31360_, new_n31361_, new_n31362_,
    new_n31363_, new_n31364_, new_n31365_, new_n31366_, new_n31367_,
    new_n31368_, new_n31369_, new_n31370_, new_n31371_, new_n31372_,
    new_n31373_, new_n31374_, new_n31375_, new_n31376_, new_n31377_,
    new_n31378_, new_n31379_, new_n31380_, new_n31381_, new_n31382_,
    new_n31383_, new_n31384_, new_n31385_, new_n31386_, new_n31387_,
    new_n31388_, new_n31389_, new_n31390_, new_n31391_, new_n31392_,
    new_n31393_, new_n31394_, new_n31395_, new_n31396_, new_n31397_,
    new_n31398_, new_n31399_, new_n31400_, new_n31401_, new_n31402_,
    new_n31403_, new_n31404_, new_n31405_, new_n31406_, new_n31407_,
    new_n31408_, new_n31409_, new_n31410_, new_n31411_, new_n31412_,
    new_n31413_, new_n31414_, new_n31415_, new_n31416_, new_n31417_,
    new_n31418_, new_n31419_, new_n31420_, new_n31421_, new_n31422_,
    new_n31423_, new_n31424_, new_n31425_, new_n31426_, new_n31427_,
    new_n31428_, new_n31429_, new_n31430_, new_n31431_, new_n31432_,
    new_n31433_, new_n31434_, new_n31435_, new_n31436_, new_n31437_,
    new_n31438_, new_n31439_, new_n31440_, new_n31441_, new_n31442_,
    new_n31443_, new_n31444_, new_n31445_, new_n31446_, new_n31447_,
    new_n31448_, new_n31449_, new_n31450_, new_n31451_, new_n31452_,
    new_n31453_, new_n31454_, new_n31455_, new_n31456_, new_n31457_,
    new_n31458_, new_n31459_, new_n31460_, new_n31461_, new_n31462_,
    new_n31463_, new_n31464_, new_n31465_, new_n31466_, new_n31467_,
    new_n31468_, new_n31469_, new_n31470_, new_n31471_, new_n31472_,
    new_n31473_, new_n31474_, new_n31475_, new_n31476_, new_n31477_,
    new_n31478_, new_n31479_, new_n31480_, new_n31481_, new_n31482_,
    new_n31483_, new_n31484_, new_n31485_, new_n31486_, new_n31487_,
    new_n31488_, new_n31489_, new_n31490_, new_n31491_, new_n31492_,
    new_n31493_, new_n31494_, new_n31495_, new_n31496_, new_n31497_,
    new_n31498_, new_n31499_, new_n31500_, new_n31501_, new_n31502_,
    new_n31503_, new_n31504_, new_n31505_, new_n31506_, new_n31507_,
    new_n31508_, new_n31509_, new_n31510_, new_n31511_, new_n31512_,
    new_n31513_, new_n31514_, new_n31515_, new_n31516_, new_n31517_,
    new_n31518_, new_n31519_, new_n31520_, new_n31521_, new_n31522_,
    new_n31523_, new_n31524_, new_n31525_, new_n31526_, new_n31527_,
    new_n31528_, new_n31529_, new_n31530_, new_n31531_, new_n31532_,
    new_n31533_, new_n31534_, new_n31535_, new_n31536_, new_n31537_,
    new_n31538_, new_n31539_, new_n31540_, new_n31541_, new_n31542_,
    new_n31543_, new_n31544_, new_n31545_, new_n31546_, new_n31547_,
    new_n31548_, new_n31549_, new_n31550_, new_n31551_, new_n31552_,
    new_n31553_, new_n31554_, new_n31555_, new_n31556_, new_n31557_,
    new_n31558_, new_n31559_, new_n31560_, new_n31561_, new_n31562_,
    new_n31563_, new_n31564_, new_n31565_, new_n31566_, new_n31567_,
    new_n31568_, new_n31569_, new_n31570_, new_n31571_, new_n31572_,
    new_n31573_, new_n31574_, new_n31575_, new_n31576_, new_n31577_,
    new_n31578_, new_n31579_, new_n31580_, new_n31581_, new_n31582_,
    new_n31583_, new_n31584_, new_n31585_, new_n31586_, new_n31587_,
    new_n31588_, new_n31589_, new_n31590_, new_n31591_, new_n31592_,
    new_n31593_, new_n31594_, new_n31595_, new_n31596_, new_n31597_,
    new_n31598_, new_n31599_, new_n31600_, new_n31601_, new_n31602_,
    new_n31603_, new_n31604_, new_n31605_, new_n31606_, new_n31607_,
    new_n31608_, new_n31609_, new_n31610_, new_n31611_, new_n31612_,
    new_n31613_, new_n31614_, new_n31615_, new_n31616_, new_n31617_,
    new_n31618_, new_n31619_, new_n31620_, new_n31621_, new_n31622_,
    new_n31623_, new_n31624_, new_n31625_, new_n31626_, new_n31627_,
    new_n31628_, new_n31629_, new_n31630_, new_n31631_, new_n31632_,
    new_n31633_, new_n31634_, new_n31635_, new_n31636_, new_n31637_,
    new_n31638_, new_n31639_, new_n31640_, new_n31641_, new_n31642_,
    new_n31643_, new_n31644_, new_n31645_, new_n31646_, new_n31647_,
    new_n31648_, new_n31649_, new_n31650_, new_n31651_, new_n31652_,
    new_n31653_, new_n31654_, new_n31655_, new_n31656_, new_n31657_,
    new_n31658_, new_n31659_, new_n31660_, new_n31661_, new_n31662_,
    new_n31663_, new_n31664_, new_n31665_, new_n31666_, new_n31667_,
    new_n31668_, new_n31669_, new_n31670_, new_n31671_, new_n31672_,
    new_n31673_, new_n31674_, new_n31675_, new_n31676_, new_n31677_,
    new_n31678_, new_n31679_, new_n31680_, new_n31681_, new_n31682_,
    new_n31683_, new_n31684_, new_n31685_, new_n31686_, new_n31687_,
    new_n31688_, new_n31689_, new_n31690_, new_n31691_, new_n31692_,
    new_n31693_, new_n31694_, new_n31695_, new_n31696_, new_n31697_,
    new_n31698_, new_n31699_, new_n31700_, new_n31701_, new_n31702_,
    new_n31703_, new_n31704_, new_n31705_, new_n31706_, new_n31707_,
    new_n31708_, new_n31709_, new_n31710_, new_n31711_, new_n31712_,
    new_n31713_, new_n31714_, new_n31715_, new_n31716_, new_n31717_,
    new_n31718_, new_n31719_, new_n31720_, new_n31721_, new_n31722_,
    new_n31723_, new_n31724_, new_n31725_, new_n31726_, new_n31727_,
    new_n31728_, new_n31729_, new_n31730_, new_n31731_, new_n31732_,
    new_n31733_, new_n31734_, new_n31735_, new_n31736_, new_n31737_,
    new_n31738_, new_n31739_, new_n31740_, new_n31741_, new_n31742_,
    new_n31743_, new_n31744_, new_n31745_, new_n31746_, new_n31747_,
    new_n31748_, new_n31749_, new_n31750_, new_n31751_, new_n31752_,
    new_n31753_, new_n31754_, new_n31755_, new_n31756_, new_n31757_,
    new_n31758_, new_n31759_, new_n31760_, new_n31761_, new_n31762_,
    new_n31763_, new_n31764_, new_n31765_, new_n31766_, new_n31767_,
    new_n31768_, new_n31769_, new_n31770_, new_n31771_, new_n31772_,
    new_n31773_, new_n31774_, new_n31775_, new_n31776_, new_n31777_,
    new_n31778_, new_n31779_, new_n31780_, new_n31781_, new_n31782_,
    new_n31783_, new_n31784_, new_n31785_, new_n31786_, new_n31787_,
    new_n31788_, new_n31789_, new_n31790_, new_n31791_, new_n31792_,
    new_n31793_, new_n31794_, new_n31795_, new_n31796_, new_n31797_,
    new_n31798_, new_n31799_, new_n31800_, new_n31801_, new_n31802_,
    new_n31803_, new_n31804_, new_n31805_, new_n31806_, new_n31807_,
    new_n31808_, new_n31809_, new_n31810_, new_n31811_, new_n31812_,
    new_n31813_, new_n31814_, new_n31815_, new_n31816_, new_n31817_,
    new_n31818_, new_n31819_, new_n31820_, new_n31821_, new_n31822_,
    new_n31823_, new_n31824_, new_n31825_, new_n31826_, new_n31827_,
    new_n31828_, new_n31829_, new_n31830_, new_n31831_, new_n31832_,
    new_n31833_, new_n31834_, new_n31835_, new_n31836_, new_n31837_,
    new_n31838_, new_n31839_, new_n31840_, new_n31841_, new_n31842_,
    new_n31843_, new_n31844_, new_n31845_, new_n31846_, new_n31847_,
    new_n31848_, new_n31849_, new_n31850_, new_n31851_, new_n31852_,
    new_n31853_, new_n31854_, new_n31855_, new_n31856_, new_n31857_,
    new_n31858_, new_n31859_, new_n31860_, new_n31861_, new_n31862_,
    new_n31863_, new_n31864_, new_n31865_, new_n31866_, new_n31867_,
    new_n31868_, new_n31869_, new_n31870_, new_n31871_, new_n31872_,
    new_n31873_, new_n31874_, new_n31875_, new_n31876_, new_n31877_,
    new_n31878_, new_n31879_, new_n31880_, new_n31881_, new_n31882_,
    new_n31883_, new_n31884_, new_n31885_, new_n31886_, new_n31887_,
    new_n31888_, new_n31889_, new_n31890_, new_n31891_, new_n31892_,
    new_n31893_, new_n31894_, new_n31895_, new_n31896_, new_n31897_,
    new_n31898_, new_n31899_, new_n31900_, new_n31901_, new_n31902_,
    new_n31903_, new_n31904_, new_n31905_, new_n31906_, new_n31907_,
    new_n31908_, new_n31909_, new_n31910_, new_n31911_, new_n31912_,
    new_n31913_, new_n31914_, new_n31915_, new_n31916_, new_n31917_,
    new_n31918_, new_n31919_, new_n31920_, new_n31921_, new_n31922_,
    new_n31923_, new_n31924_, new_n31925_, new_n31926_, new_n31927_,
    new_n31928_, new_n31929_, new_n31930_, new_n31931_, new_n31932_,
    new_n31933_, new_n31934_, new_n31935_, new_n31936_, new_n31937_,
    new_n31938_, new_n31939_, new_n31940_, new_n31941_, new_n31942_,
    new_n31943_, new_n31944_, new_n31945_, new_n31946_, new_n31947_,
    new_n31948_, new_n31949_, new_n31950_, new_n31951_, new_n31952_,
    new_n31953_, new_n31954_, new_n31955_, new_n31956_, new_n31957_,
    new_n31958_, new_n31959_, new_n31960_, new_n31961_, new_n31962_,
    new_n31963_, new_n31964_, new_n31965_, new_n31966_, new_n31967_,
    new_n31968_, new_n31969_, new_n31970_, new_n31971_, new_n31972_,
    new_n31973_, new_n31974_, new_n31975_, new_n31976_, new_n31977_,
    new_n31978_, new_n31979_, new_n31980_, new_n31981_, new_n31982_,
    new_n31983_, new_n31984_, new_n31985_, new_n31986_, new_n31987_,
    new_n31988_, new_n31989_, new_n31990_, new_n31991_, new_n31992_,
    new_n31993_, new_n31994_, new_n31995_, new_n31996_, new_n31997_,
    new_n31998_, new_n31999_, new_n32000_, new_n32001_, new_n32002_,
    new_n32003_, new_n32004_, new_n32005_, new_n32006_, new_n32007_,
    new_n32008_, new_n32009_, new_n32010_, new_n32011_, new_n32012_,
    new_n32013_, new_n32014_, new_n32015_, new_n32016_, new_n32017_,
    new_n32018_, new_n32019_, new_n32020_, new_n32021_, new_n32022_,
    new_n32023_, new_n32024_, new_n32025_, new_n32026_, new_n32027_,
    new_n32028_, new_n32029_, new_n32030_, new_n32031_, new_n32032_,
    new_n32033_, new_n32034_, new_n32035_, new_n32036_, new_n32037_,
    new_n32038_, new_n32039_, new_n32040_, new_n32041_, new_n32042_,
    new_n32043_, new_n32044_, new_n32045_, new_n32046_, new_n32047_,
    new_n32048_, new_n32049_, new_n32050_, new_n32051_, new_n32052_,
    new_n32053_, new_n32054_, new_n32055_, new_n32056_, new_n32057_,
    new_n32058_, new_n32059_, new_n32060_, new_n32061_, new_n32062_,
    new_n32063_, new_n32064_, new_n32065_, new_n32066_, new_n32067_,
    new_n32068_, new_n32069_, new_n32070_, new_n32071_, new_n32072_,
    new_n32073_, new_n32074_, new_n32075_, new_n32076_, new_n32077_,
    new_n32078_, new_n32079_, new_n32080_, new_n32081_, new_n32082_,
    new_n32083_, new_n32084_, new_n32085_, new_n32086_, new_n32087_,
    new_n32088_, new_n32089_, new_n32090_, new_n32091_, new_n32092_,
    new_n32093_, new_n32094_, new_n32095_, new_n32096_, new_n32097_,
    new_n32098_, new_n32099_, new_n32100_, new_n32101_, new_n32102_,
    new_n32103_, new_n32104_, new_n32105_, new_n32106_, new_n32107_,
    new_n32108_, new_n32109_, new_n32110_, new_n32111_, new_n32112_,
    new_n32113_, new_n32114_, new_n32115_, new_n32116_, new_n32117_,
    new_n32118_, new_n32119_, new_n32120_, new_n32121_, new_n32122_,
    new_n32123_, new_n32124_, new_n32125_, new_n32126_, new_n32127_,
    new_n32128_, new_n32129_, new_n32130_, new_n32131_, new_n32132_,
    new_n32133_, new_n32134_, new_n32135_, new_n32136_, new_n32137_,
    new_n32138_, new_n32139_, new_n32140_, new_n32141_, new_n32142_,
    new_n32143_, new_n32144_, new_n32145_, new_n32146_, new_n32147_,
    new_n32148_, new_n32149_, new_n32150_, new_n32151_, new_n32152_,
    new_n32153_, new_n32154_, new_n32155_, new_n32156_, new_n32157_,
    new_n32158_, new_n32159_, new_n32160_, new_n32161_, new_n32162_,
    new_n32163_, new_n32164_, new_n32165_, new_n32166_, new_n32167_,
    new_n32168_, new_n32169_, new_n32170_, new_n32171_, new_n32172_,
    new_n32173_, new_n32174_, new_n32175_, new_n32176_, new_n32177_,
    new_n32178_, new_n32179_, new_n32180_, new_n32181_, new_n32182_,
    new_n32183_, new_n32184_, new_n32185_, new_n32186_, new_n32187_,
    new_n32188_, new_n32189_, new_n32190_, new_n32191_, new_n32192_,
    new_n32193_, new_n32194_, new_n32195_, new_n32196_, new_n32197_,
    new_n32198_, new_n32199_, new_n32200_, new_n32201_, new_n32202_,
    new_n32203_, new_n32204_, new_n32205_, new_n32206_, new_n32207_,
    new_n32208_, new_n32209_, new_n32210_, new_n32211_, new_n32212_,
    new_n32213_, new_n32214_, new_n32215_, new_n32216_, new_n32217_,
    new_n32218_, new_n32219_, new_n32220_, new_n32221_, new_n32222_,
    new_n32223_, new_n32224_, new_n32225_, new_n32226_, new_n32227_,
    new_n32228_, new_n32229_, new_n32230_, new_n32231_, new_n32232_,
    new_n32233_, new_n32234_, new_n32235_, new_n32236_, new_n32237_,
    new_n32238_, new_n32239_, new_n32240_, new_n32241_, new_n32242_,
    new_n32243_, new_n32244_, new_n32245_, new_n32246_, new_n32247_,
    new_n32248_, new_n32249_, new_n32250_, new_n32251_, new_n32252_,
    new_n32253_, new_n32254_, new_n32255_, new_n32256_, new_n32257_,
    new_n32258_, new_n32259_, new_n32260_, new_n32261_, new_n32262_,
    new_n32263_, new_n32264_, new_n32265_, new_n32266_, new_n32267_,
    new_n32268_, new_n32269_, new_n32270_, new_n32271_, new_n32272_,
    new_n32273_, new_n32274_, new_n32275_, new_n32276_, new_n32277_,
    new_n32278_, new_n32279_, new_n32280_, new_n32281_, new_n32282_,
    new_n32283_, new_n32284_, new_n32285_, new_n32286_, new_n32287_,
    new_n32288_, new_n32289_, new_n32290_, new_n32291_, new_n32292_,
    new_n32293_, new_n32294_, new_n32295_, new_n32296_, new_n32297_,
    new_n32298_, new_n32299_, new_n32300_, new_n32301_, new_n32302_,
    new_n32303_, new_n32304_, new_n32305_, new_n32306_, new_n32307_,
    new_n32308_, new_n32309_, new_n32310_, new_n32311_, new_n32312_,
    new_n32313_, new_n32314_, new_n32315_, new_n32316_, new_n32317_,
    new_n32318_, new_n32319_, new_n32320_, new_n32321_, new_n32322_,
    new_n32323_, new_n32324_, new_n32325_, new_n32326_, new_n32327_,
    new_n32328_, new_n32329_, new_n32330_, new_n32331_, new_n32332_,
    new_n32333_, new_n32334_, new_n32335_, new_n32336_, new_n32337_,
    new_n32338_, new_n32339_, new_n32340_, new_n32341_, new_n32342_,
    new_n32343_, new_n32344_, new_n32345_, new_n32346_, new_n32347_,
    new_n32348_, new_n32349_, new_n32350_, new_n32351_, new_n32352_,
    new_n32353_, new_n32354_, new_n32355_, new_n32356_, new_n32357_,
    new_n32358_, new_n32359_, new_n32360_, new_n32361_, new_n32362_,
    new_n32363_, new_n32364_, new_n32365_, new_n32366_, new_n32367_,
    new_n32368_, new_n32369_, new_n32370_, new_n32371_, new_n32372_,
    new_n32373_, new_n32374_, new_n32375_, new_n32376_, new_n32377_,
    new_n32378_, new_n32379_, new_n32380_, new_n32381_, new_n32382_,
    new_n32383_, new_n32384_, new_n32385_, new_n32386_, new_n32387_,
    new_n32388_, new_n32389_, new_n32390_, new_n32391_, new_n32392_,
    new_n32393_, new_n32394_, new_n32395_, new_n32396_, new_n32397_,
    new_n32398_, new_n32399_, new_n32400_, new_n32401_, new_n32402_,
    new_n32403_, new_n32404_, new_n32405_, new_n32406_, new_n32407_,
    new_n32408_, new_n32409_, new_n32410_, new_n32411_, new_n32412_,
    new_n32413_, new_n32414_, new_n32415_, new_n32416_, new_n32417_,
    new_n32418_, new_n32419_, new_n32420_, new_n32421_, new_n32422_,
    new_n32423_, new_n32424_, new_n32425_, new_n32426_, new_n32427_,
    new_n32428_, new_n32429_, new_n32430_, new_n32431_, new_n32432_,
    new_n32433_, new_n32434_, new_n32435_, new_n32436_, new_n32437_,
    new_n32438_, new_n32439_, new_n32440_, new_n32441_, new_n32442_,
    new_n32443_, new_n32444_, new_n32445_, new_n32446_, new_n32447_,
    new_n32448_, new_n32449_, new_n32450_, new_n32451_, new_n32452_,
    new_n32453_, new_n32454_, new_n32455_, new_n32456_, new_n32457_,
    new_n32458_, new_n32459_, new_n32460_, new_n32461_, new_n32462_,
    new_n32463_, new_n32464_, new_n32465_, new_n32466_, new_n32467_,
    new_n32468_, new_n32469_, new_n32470_, new_n32471_, new_n32472_,
    new_n32473_, new_n32474_, new_n32475_, new_n32476_, new_n32477_,
    new_n32478_, new_n32479_, new_n32480_, new_n32481_, new_n32482_,
    new_n32483_, new_n32484_, new_n32485_, new_n32486_, new_n32487_,
    new_n32488_, new_n32489_, new_n32490_, new_n32491_, new_n32492_,
    new_n32493_, new_n32494_, new_n32495_, new_n32496_, new_n32497_,
    new_n32498_, new_n32499_, new_n32500_, new_n32501_, new_n32502_,
    new_n32503_, new_n32504_, new_n32505_, new_n32506_, new_n32507_,
    new_n32508_, new_n32509_, new_n32510_, new_n32511_, new_n32512_,
    new_n32513_, new_n32514_, new_n32515_, new_n32516_, new_n32517_,
    new_n32518_, new_n32519_, new_n32520_, new_n32521_, new_n32522_,
    new_n32523_, new_n32524_, new_n32525_, new_n32526_, new_n32527_,
    new_n32528_, new_n32529_, new_n32530_, new_n32531_, new_n32532_,
    new_n32533_, new_n32534_, new_n32535_, new_n32536_, new_n32537_,
    new_n32538_, new_n32539_, new_n32540_, new_n32541_, new_n32542_,
    new_n32543_, new_n32544_, new_n32545_, new_n32546_, new_n32547_,
    new_n32548_, new_n32549_, new_n32550_, new_n32551_, new_n32552_,
    new_n32553_, new_n32554_, new_n32555_, new_n32556_, new_n32557_,
    new_n32558_, new_n32559_, new_n32560_, new_n32561_, new_n32562_,
    new_n32563_, new_n32564_, new_n32565_, new_n32566_, new_n32567_,
    new_n32568_, new_n32569_, new_n32570_, new_n32571_, new_n32572_,
    new_n32573_, new_n32574_, new_n32575_, new_n32576_, new_n32577_,
    new_n32578_, new_n32579_, new_n32580_, new_n32581_, new_n32582_,
    new_n32583_, new_n32584_, new_n32585_, new_n32586_, new_n32587_,
    new_n32588_, new_n32589_, new_n32590_, new_n32591_, new_n32592_,
    new_n32593_, new_n32594_, new_n32595_, new_n32596_, new_n32597_,
    new_n32598_, new_n32599_, new_n32600_, new_n32601_, new_n32602_,
    new_n32603_, new_n32604_, new_n32605_, new_n32606_, new_n32607_,
    new_n32608_, new_n32609_, new_n32610_, new_n32611_, new_n32612_,
    new_n32613_, new_n32614_, new_n32615_, new_n32616_, new_n32617_,
    new_n32618_, new_n32619_, new_n32620_, new_n32621_, new_n32622_,
    new_n32623_, new_n32624_, new_n32625_, new_n32626_, new_n32627_,
    new_n32628_, new_n32629_, new_n32630_, new_n32631_, new_n32632_,
    new_n32633_, new_n32634_, new_n32635_, new_n32636_, new_n32637_,
    new_n32638_, new_n32639_, new_n32640_, new_n32641_, new_n32642_,
    new_n32643_, new_n32644_, new_n32645_, new_n32646_, new_n32647_,
    new_n32648_, new_n32649_, new_n32650_, new_n32651_, new_n32652_,
    new_n32653_, new_n32654_, new_n32655_, new_n32656_, new_n32657_,
    new_n32658_, new_n32659_, new_n32660_, new_n32661_, new_n32662_,
    new_n32663_, new_n32664_, new_n32665_, new_n32666_, new_n32667_,
    new_n32668_, new_n32669_, new_n32670_, new_n32671_, new_n32672_,
    new_n32673_, new_n32674_, new_n32675_, new_n32676_, new_n32677_,
    new_n32678_, new_n32679_, new_n32680_, new_n32681_, new_n32682_,
    new_n32683_, new_n32684_, new_n32685_, new_n32686_, new_n32687_,
    new_n32688_, new_n32689_, new_n32690_, new_n32691_, new_n32692_,
    new_n32693_, new_n32694_, new_n32695_, new_n32696_, new_n32697_,
    new_n32698_, new_n32699_, new_n32700_, new_n32701_, new_n32702_,
    new_n32703_, new_n32704_, new_n32705_, new_n32706_, new_n32707_,
    new_n32708_, new_n32709_, new_n32710_, new_n32711_, new_n32712_,
    new_n32713_, new_n32714_, new_n32715_, new_n32716_, new_n32717_,
    new_n32718_, new_n32719_, new_n32720_, new_n32721_, new_n32722_,
    new_n32723_, new_n32724_, new_n32725_, new_n32726_, new_n32727_,
    new_n32728_, new_n32729_, new_n32730_, new_n32731_, new_n32732_,
    new_n32733_, new_n32734_, new_n32735_, new_n32736_, new_n32737_,
    new_n32738_, new_n32739_, new_n32740_, new_n32741_, new_n32742_,
    new_n32743_, new_n32744_, new_n32745_, new_n32746_, new_n32747_,
    new_n32748_, new_n32749_, new_n32750_, new_n32751_, new_n32752_,
    new_n32753_, new_n32754_, new_n32755_, new_n32756_, new_n32757_,
    new_n32758_, new_n32759_, new_n32760_, new_n32761_, new_n32762_,
    new_n32763_, new_n32764_, new_n32765_, new_n32766_, new_n32767_,
    new_n32768_, new_n32769_, new_n32770_, new_n32771_, new_n32772_,
    new_n32773_, new_n32774_, new_n32775_, new_n32776_, new_n32777_,
    new_n32778_, new_n32779_, new_n32780_, new_n32781_, new_n32782_,
    new_n32783_, new_n32784_, new_n32785_, new_n32786_, new_n32787_,
    new_n32788_, new_n32789_, new_n32790_, new_n32791_, new_n32792_,
    new_n32793_, new_n32794_, new_n32795_, new_n32796_, new_n32797_,
    new_n32798_, new_n32799_, new_n32800_, new_n32801_, new_n32802_,
    new_n32803_, new_n32804_, new_n32805_, new_n32806_, new_n32807_,
    new_n32808_, new_n32809_, new_n32810_, new_n32811_, new_n32812_,
    new_n32813_, new_n32814_, new_n32815_, new_n32816_, new_n32817_,
    new_n32818_, new_n32819_, new_n32820_, new_n32821_, new_n32822_,
    new_n32823_, new_n32824_, new_n32825_, new_n32826_, new_n32827_,
    new_n32828_, new_n32829_, new_n32830_, new_n32831_, new_n32832_,
    new_n32833_, new_n32834_, new_n32835_, new_n32836_, new_n32837_,
    new_n32838_, new_n32839_, new_n32840_, new_n32841_, new_n32842_,
    new_n32843_, new_n32844_, new_n32845_, new_n32846_, new_n32847_,
    new_n32848_, new_n32849_, new_n32850_, new_n32851_, new_n32852_,
    new_n32853_, new_n32854_, new_n32855_, new_n32856_, new_n32857_,
    new_n32858_, new_n32859_, new_n32860_, new_n32861_, new_n32862_,
    new_n32863_, new_n32864_, new_n32865_, new_n32866_, new_n32867_,
    new_n32868_, new_n32869_, new_n32870_, new_n32871_, new_n32872_,
    new_n32873_, new_n32874_, new_n32875_, new_n32876_, new_n32877_,
    new_n32878_, new_n32879_, new_n32880_, new_n32881_, new_n32882_,
    new_n32883_, new_n32884_, new_n32885_, new_n32886_, new_n32887_,
    new_n32888_, new_n32889_, new_n32890_, new_n32891_, new_n32892_,
    new_n32893_, new_n32894_, new_n32895_, new_n32896_, new_n32897_,
    new_n32898_, new_n32899_, new_n32900_, new_n32901_, new_n32902_,
    new_n32903_, new_n32904_, new_n32905_, new_n32906_, new_n32907_,
    new_n32908_, new_n32909_, new_n32910_, new_n32911_, new_n32912_,
    new_n32913_, new_n32914_, new_n32915_, new_n32916_, new_n32917_,
    new_n32918_, new_n32919_, new_n32920_, new_n32921_, new_n32922_,
    new_n32923_, new_n32924_, new_n32925_, new_n32926_, new_n32927_,
    new_n32928_, new_n32929_, new_n32930_, new_n32931_, new_n32932_,
    new_n32933_, new_n32934_, new_n32935_, new_n32936_, new_n32937_,
    new_n32938_, new_n32939_, new_n32940_, new_n32941_, new_n32942_,
    new_n32943_, new_n32944_, new_n32945_, new_n32946_, new_n32947_,
    new_n32948_, new_n32949_, new_n32950_, new_n32951_, new_n32952_,
    new_n32953_, new_n32954_, new_n32955_, new_n32956_, new_n32957_,
    new_n32958_, new_n32959_, new_n32960_, new_n32961_, new_n32962_,
    new_n32963_, new_n32964_, new_n32965_, new_n32966_, new_n32967_,
    new_n32968_, new_n32969_, new_n32970_, new_n32971_, new_n32972_,
    new_n32973_, new_n32974_, new_n32975_, new_n32976_, new_n32977_,
    new_n32978_, new_n32979_, new_n32980_, new_n32981_, new_n32982_,
    new_n32983_, new_n32984_, new_n32985_, new_n32986_, new_n32987_,
    new_n32988_, new_n32989_, new_n32990_, new_n32991_, new_n32992_,
    new_n32993_, new_n32994_, new_n32995_, new_n32996_, new_n32997_,
    new_n32998_, new_n32999_, new_n33000_, new_n33001_, new_n33002_,
    new_n33003_, new_n33004_, new_n33005_, new_n33006_, new_n33007_,
    new_n33008_, new_n33009_, new_n33010_, new_n33011_, new_n33012_,
    new_n33013_, new_n33014_, new_n33015_, new_n33016_, new_n33017_,
    new_n33018_, new_n33019_, new_n33020_, new_n33021_, new_n33022_,
    new_n33023_, new_n33024_, new_n33025_, new_n33026_, new_n33027_,
    new_n33028_, new_n33029_, new_n33030_, new_n33031_, new_n33032_,
    new_n33033_, new_n33034_, new_n33035_, new_n33036_, new_n33037_,
    new_n33038_, new_n33039_, new_n33040_, new_n33041_, new_n33042_,
    new_n33043_, new_n33044_, new_n33045_, new_n33046_, new_n33047_,
    new_n33048_, new_n33049_, new_n33050_, new_n33051_, new_n33052_,
    new_n33053_, new_n33054_, new_n33055_, new_n33056_, new_n33057_,
    new_n33058_, new_n33059_, new_n33060_, new_n33061_, new_n33062_,
    new_n33063_, new_n33064_, new_n33065_, new_n33066_, new_n33067_,
    new_n33068_, new_n33069_, new_n33070_, new_n33071_, new_n33072_,
    new_n33073_, new_n33074_, new_n33075_, new_n33076_, new_n33077_,
    new_n33078_, new_n33079_, new_n33080_, new_n33081_, new_n33082_,
    new_n33083_, new_n33084_, new_n33085_, new_n33086_, new_n33087_,
    new_n33088_, new_n33089_, new_n33090_, new_n33091_, new_n33092_,
    new_n33093_, new_n33094_, new_n33095_, new_n33096_, new_n33097_,
    new_n33098_, new_n33099_, new_n33100_, new_n33101_, new_n33102_,
    new_n33103_, new_n33104_, new_n33105_, new_n33106_, new_n33107_,
    new_n33108_, new_n33109_, new_n33110_, new_n33111_, new_n33112_,
    new_n33113_, new_n33114_, new_n33115_, new_n33116_, new_n33117_,
    new_n33118_, new_n33119_, new_n33120_, new_n33121_, new_n33122_,
    new_n33123_, new_n33124_, new_n33125_, new_n33126_, new_n33127_,
    new_n33128_, new_n33129_, new_n33130_, new_n33131_, new_n33132_,
    new_n33133_, new_n33134_, new_n33135_, new_n33136_, new_n33137_,
    new_n33138_, new_n33139_, new_n33140_, new_n33141_, new_n33142_,
    new_n33143_, new_n33144_, new_n33145_, new_n33146_, new_n33147_,
    new_n33148_, new_n33149_, new_n33150_, new_n33151_, new_n33152_,
    new_n33153_, new_n33154_, new_n33155_, new_n33156_, new_n33157_,
    new_n33158_, new_n33159_, new_n33160_, new_n33161_, new_n33162_,
    new_n33163_, new_n33164_, new_n33165_, new_n33166_, new_n33167_,
    new_n33168_, new_n33169_, new_n33170_, new_n33171_, new_n33172_,
    new_n33173_, new_n33174_, new_n33175_, new_n33176_, new_n33177_,
    new_n33178_, new_n33179_, new_n33180_, new_n33181_, new_n33182_,
    new_n33183_, new_n33184_, new_n33185_, new_n33186_, new_n33187_,
    new_n33188_, new_n33189_, new_n33190_, new_n33191_, new_n33192_,
    new_n33193_, new_n33194_, new_n33195_, new_n33196_, new_n33197_,
    new_n33198_, new_n33199_, new_n33200_, new_n33201_, new_n33202_,
    new_n33203_, new_n33204_, new_n33205_, new_n33206_, new_n33207_,
    new_n33208_, new_n33209_, new_n33210_, new_n33211_, new_n33212_,
    new_n33213_, new_n33214_, new_n33215_, new_n33216_, new_n33217_,
    new_n33218_, new_n33219_, new_n33220_, new_n33221_, new_n33222_,
    new_n33223_, new_n33224_, new_n33225_, new_n33226_, new_n33227_,
    new_n33228_, new_n33229_, new_n33230_, new_n33231_, new_n33232_,
    new_n33233_, new_n33234_, new_n33235_, new_n33236_, new_n33237_,
    new_n33238_, new_n33239_, new_n33240_, new_n33241_, new_n33242_,
    new_n33243_, new_n33244_, new_n33245_, new_n33246_, new_n33247_,
    new_n33248_, new_n33249_, new_n33250_, new_n33251_, new_n33252_,
    new_n33253_, new_n33254_, new_n33255_, new_n33256_, new_n33257_,
    new_n33258_, new_n33259_, new_n33260_, new_n33261_, new_n33262_,
    new_n33263_, new_n33264_, new_n33265_, new_n33266_, new_n33267_,
    new_n33268_, new_n33269_, new_n33270_, new_n33271_, new_n33272_,
    new_n33273_, new_n33274_, new_n33275_, new_n33276_, new_n33277_,
    new_n33278_, new_n33279_, new_n33280_, new_n33281_, new_n33282_,
    new_n33283_, new_n33284_, new_n33285_, new_n33286_, new_n33287_,
    new_n33288_, new_n33289_, new_n33290_, new_n33291_, new_n33292_,
    new_n33293_, new_n33294_, new_n33295_, new_n33296_, new_n33297_,
    new_n33298_, new_n33299_, new_n33300_, new_n33301_, new_n33302_,
    new_n33303_, new_n33304_, new_n33305_, new_n33306_, new_n33307_,
    new_n33308_, new_n33309_, new_n33310_, new_n33311_, new_n33312_,
    new_n33313_, new_n33314_, new_n33315_, new_n33316_, new_n33317_,
    new_n33318_, new_n33319_, new_n33320_, new_n33321_, new_n33322_,
    new_n33323_, new_n33324_, new_n33325_, new_n33326_, new_n33327_,
    new_n33328_, new_n33329_, new_n33330_, new_n33331_, new_n33332_,
    new_n33333_, new_n33334_, new_n33335_, new_n33336_, new_n33337_,
    new_n33338_, new_n33339_, new_n33340_, new_n33341_, new_n33342_,
    new_n33343_, new_n33344_, new_n33345_, new_n33346_, new_n33347_,
    new_n33348_, new_n33349_, new_n33350_, new_n33351_, new_n33352_,
    new_n33353_, new_n33354_, new_n33355_, new_n33356_, new_n33357_,
    new_n33358_, new_n33359_, new_n33360_, new_n33361_, new_n33362_,
    new_n33363_, new_n33364_, new_n33365_, new_n33366_, new_n33367_,
    new_n33368_, new_n33369_, new_n33370_, new_n33371_, new_n33372_,
    new_n33373_, new_n33374_, new_n33375_, new_n33376_, new_n33377_,
    new_n33378_, new_n33379_, new_n33380_, new_n33381_, new_n33382_,
    new_n33383_, new_n33384_, new_n33385_, new_n33386_, new_n33387_,
    new_n33388_, new_n33389_, new_n33390_, new_n33391_, new_n33392_,
    new_n33393_, new_n33394_, new_n33395_, new_n33396_, new_n33397_,
    new_n33398_, new_n33399_, new_n33400_, new_n33401_, new_n33402_,
    new_n33403_, new_n33404_, new_n33405_, new_n33406_, new_n33407_,
    new_n33408_, new_n33409_, new_n33410_, new_n33411_, new_n33412_,
    new_n33413_, new_n33414_, new_n33415_, new_n33416_, new_n33417_,
    new_n33418_, new_n33419_, new_n33420_, new_n33421_, new_n33422_,
    new_n33423_, new_n33424_, new_n33425_, new_n33426_, new_n33427_,
    new_n33428_, new_n33429_, new_n33430_, new_n33431_, new_n33432_,
    new_n33433_, new_n33434_, new_n33435_, new_n33436_, new_n33437_,
    new_n33438_, new_n33439_, new_n33440_, new_n33441_, new_n33442_,
    new_n33443_, new_n33444_, new_n33445_, new_n33446_, new_n33447_,
    new_n33448_, new_n33449_, new_n33450_, new_n33451_, new_n33452_,
    new_n33453_, new_n33454_, new_n33455_, new_n33456_, new_n33457_,
    new_n33458_, new_n33459_, new_n33460_, new_n33461_, new_n33462_,
    new_n33463_, new_n33464_, new_n33465_, new_n33466_, new_n33467_,
    new_n33468_, new_n33469_, new_n33470_, new_n33471_, new_n33472_,
    new_n33473_, new_n33474_, new_n33475_, new_n33476_, new_n33477_,
    new_n33478_, new_n33479_, new_n33480_, new_n33481_, new_n33482_,
    new_n33483_, new_n33484_, new_n33485_, new_n33486_, new_n33487_,
    new_n33488_, new_n33489_, new_n33490_, new_n33491_, new_n33492_,
    new_n33493_, new_n33494_, new_n33495_, new_n33496_, new_n33497_,
    new_n33498_, new_n33499_, new_n33500_, new_n33501_, new_n33502_,
    new_n33503_, new_n33504_, new_n33505_, new_n33506_, new_n33507_,
    new_n33508_, new_n33509_, new_n33510_, new_n33511_, new_n33512_,
    new_n33513_, new_n33514_, new_n33515_, new_n33516_, new_n33517_,
    new_n33518_, new_n33519_, new_n33520_, new_n33521_, new_n33522_,
    new_n33523_, new_n33524_, new_n33525_, new_n33526_, new_n33527_,
    new_n33528_, new_n33529_, new_n33530_, new_n33531_, new_n33532_,
    new_n33533_, new_n33534_, new_n33535_, new_n33536_, new_n33537_,
    new_n33538_, new_n33539_, new_n33540_, new_n33541_, new_n33542_,
    new_n33543_, new_n33544_, new_n33545_, new_n33546_, new_n33547_,
    new_n33548_, new_n33549_, new_n33550_, new_n33551_, new_n33552_,
    new_n33553_, new_n33554_, new_n33555_, new_n33556_, new_n33557_,
    new_n33558_, new_n33559_, new_n33560_, new_n33561_, new_n33562_,
    new_n33563_, new_n33564_, new_n33565_, new_n33566_, new_n33567_,
    new_n33568_, new_n33569_, new_n33570_, new_n33571_, new_n33572_,
    new_n33573_, new_n33574_, new_n33575_, new_n33576_, new_n33577_,
    new_n33578_, new_n33579_, new_n33580_, new_n33581_, new_n33582_,
    new_n33583_, new_n33584_, new_n33585_, new_n33586_, new_n33587_,
    new_n33588_, new_n33589_, new_n33590_, new_n33591_, new_n33592_,
    new_n33593_, new_n33594_, new_n33595_, new_n33596_, new_n33597_,
    new_n33598_, new_n33599_, new_n33600_, new_n33601_, new_n33602_,
    new_n33603_, new_n33604_, new_n33605_, new_n33606_, new_n33607_,
    new_n33608_, new_n33609_, new_n33610_, new_n33611_, new_n33612_,
    new_n33613_, new_n33614_, new_n33615_, new_n33616_, new_n33617_,
    new_n33618_, new_n33619_, new_n33620_, new_n33621_, new_n33622_,
    new_n33623_, new_n33624_, new_n33625_, new_n33626_, new_n33627_,
    new_n33628_, new_n33629_, new_n33630_, new_n33631_, new_n33632_,
    new_n33633_, new_n33634_, new_n33635_, new_n33636_, new_n33637_,
    new_n33638_, new_n33639_, new_n33640_, new_n33641_, new_n33642_,
    new_n33643_, new_n33644_, new_n33645_, new_n33646_, new_n33647_,
    new_n33648_, new_n33649_, new_n33650_, new_n33651_, new_n33652_,
    new_n33653_, new_n33654_, new_n33655_, new_n33656_, new_n33657_,
    new_n33658_, new_n33659_, new_n33660_, new_n33661_, new_n33662_,
    new_n33663_, new_n33664_, new_n33665_, new_n33666_, new_n33667_,
    new_n33668_, new_n33669_, new_n33670_, new_n33671_, new_n33672_,
    new_n33673_, new_n33674_, new_n33675_, new_n33676_, new_n33677_,
    new_n33678_, new_n33679_, new_n33680_, new_n33681_, new_n33682_,
    new_n33683_, new_n33684_, new_n33685_, new_n33686_, new_n33687_,
    new_n33688_, new_n33689_, new_n33690_, new_n33691_, new_n33692_,
    new_n33693_, new_n33694_, new_n33695_, new_n33696_, new_n33697_,
    new_n33698_, new_n33699_, new_n33700_, new_n33701_, new_n33702_,
    new_n33703_, new_n33704_, new_n33705_, new_n33706_, new_n33707_,
    new_n33708_, new_n33709_, new_n33710_, new_n33711_, new_n33712_,
    new_n33713_, new_n33714_, new_n33715_, new_n33716_, new_n33717_,
    new_n33718_, new_n33719_, new_n33720_, new_n33721_, new_n33722_,
    new_n33723_, new_n33724_, new_n33725_, new_n33726_, new_n33727_,
    new_n33728_, new_n33729_, new_n33730_, new_n33731_, new_n33732_,
    new_n33733_, new_n33734_, new_n33735_, new_n33736_, new_n33737_,
    new_n33738_, new_n33739_, new_n33740_, new_n33741_, new_n33742_,
    new_n33743_, new_n33744_, new_n33745_, new_n33746_, new_n33747_,
    new_n33748_, new_n33749_, new_n33750_, new_n33751_, new_n33752_,
    new_n33753_, new_n33754_, new_n33755_, new_n33756_, new_n33757_,
    new_n33758_, new_n33759_, new_n33760_, new_n33761_, new_n33762_,
    new_n33763_, new_n33764_, new_n33765_, new_n33766_, new_n33767_,
    new_n33768_, new_n33769_, new_n33770_, new_n33771_, new_n33772_,
    new_n33773_, new_n33774_, new_n33775_, new_n33776_, new_n33777_,
    new_n33778_, new_n33779_, new_n33780_, new_n33781_, new_n33782_,
    new_n33783_, new_n33784_, new_n33785_, new_n33786_, new_n33787_,
    new_n33788_, new_n33789_, new_n33790_, new_n33791_, new_n33792_,
    new_n33793_, new_n33794_, new_n33795_, new_n33796_, new_n33797_,
    new_n33798_, new_n33799_, new_n33800_, new_n33801_, new_n33802_,
    new_n33803_, new_n33804_, new_n33805_, new_n33806_, new_n33807_,
    new_n33808_, new_n33809_, new_n33810_, new_n33811_, new_n33812_,
    new_n33813_, new_n33814_, new_n33815_, new_n33816_, new_n33817_,
    new_n33818_, new_n33819_, new_n33820_, new_n33821_, new_n33822_,
    new_n33823_, new_n33824_, new_n33825_, new_n33826_, new_n33827_,
    new_n33828_, new_n33829_, new_n33830_, new_n33831_, new_n33832_,
    new_n33833_, new_n33834_, new_n33835_, new_n33836_, new_n33837_,
    new_n33838_, new_n33839_, new_n33840_, new_n33841_, new_n33842_,
    new_n33843_, new_n33844_, new_n33845_, new_n33846_, new_n33847_,
    new_n33848_, new_n33849_, new_n33850_, new_n33851_, new_n33852_,
    new_n33853_, new_n33854_, new_n33855_, new_n33856_, new_n33857_,
    new_n33858_, new_n33859_, new_n33860_, new_n33861_, new_n33862_,
    new_n33863_, new_n33864_, new_n33865_, new_n33866_, new_n33867_,
    new_n33868_, new_n33869_, new_n33870_, new_n33871_, new_n33872_,
    new_n33873_, new_n33874_, new_n33875_, new_n33876_, new_n33877_,
    new_n33878_, new_n33879_, new_n33880_, new_n33881_, new_n33882_,
    new_n33883_, new_n33884_, new_n33885_, new_n33886_, new_n33887_,
    new_n33888_, new_n33889_, new_n33890_, new_n33891_, new_n33892_,
    new_n33893_, new_n33894_, new_n33895_, new_n33896_, new_n33897_,
    new_n33898_, new_n33899_, new_n33900_, new_n33901_, new_n33902_,
    new_n33903_, new_n33904_, new_n33905_, new_n33906_, new_n33907_,
    new_n33908_, new_n33909_, new_n33910_, new_n33911_, new_n33912_,
    new_n33913_, new_n33914_, new_n33915_, new_n33916_, new_n33917_,
    new_n33918_, new_n33919_, new_n33920_, new_n33921_, new_n33922_,
    new_n33923_, new_n33924_, new_n33925_, new_n33926_, new_n33927_,
    new_n33928_, new_n33929_, new_n33930_, new_n33931_, new_n33932_,
    new_n33933_, new_n33934_, new_n33935_, new_n33936_, new_n33937_,
    new_n33938_, new_n33939_, new_n33940_, new_n33941_, new_n33942_,
    new_n33943_, new_n33944_, new_n33945_, new_n33946_, new_n33947_,
    new_n33948_, new_n33949_, new_n33950_, new_n33951_, new_n33952_,
    new_n33953_, new_n33954_, new_n33955_, new_n33956_, new_n33957_,
    new_n33958_, new_n33959_, new_n33960_, new_n33961_, new_n33962_,
    new_n33963_, new_n33964_, new_n33965_, new_n33966_, new_n33967_,
    new_n33968_, new_n33969_, new_n33970_, new_n33971_, new_n33972_,
    new_n33973_, new_n33974_, new_n33975_, new_n33976_, new_n33977_,
    new_n33978_, new_n33979_, new_n33980_, new_n33981_, new_n33982_,
    new_n33983_, new_n33984_, new_n33985_, new_n33986_, new_n33987_,
    new_n33988_, new_n33989_, new_n33990_, new_n33991_, new_n33992_,
    new_n33993_, new_n33994_, new_n33995_, new_n33996_, new_n33997_,
    new_n33998_, new_n33999_, new_n34000_, new_n34001_, new_n34002_,
    new_n34003_, new_n34004_, new_n34005_, new_n34006_, new_n34007_,
    new_n34008_, new_n34009_, new_n34010_, new_n34011_, new_n34012_,
    new_n34013_, new_n34014_, new_n34015_, new_n34016_, new_n34017_,
    new_n34018_, new_n34019_, new_n34020_, new_n34021_, new_n34022_,
    new_n34023_, new_n34024_, new_n34025_, new_n34026_, new_n34027_,
    new_n34028_, new_n34029_, new_n34030_, new_n34031_, new_n34032_,
    new_n34033_, new_n34034_, new_n34035_, new_n34036_, new_n34037_,
    new_n34038_, new_n34039_, new_n34040_, new_n34041_, new_n34042_,
    new_n34043_, new_n34044_, new_n34045_, new_n34046_, new_n34047_,
    new_n34048_, new_n34049_, new_n34050_, new_n34051_, new_n34052_,
    new_n34053_, new_n34054_, new_n34055_, new_n34056_, new_n34057_,
    new_n34058_, new_n34059_, new_n34060_, new_n34061_, new_n34062_,
    new_n34063_, new_n34064_, new_n34065_, new_n34066_, new_n34067_,
    new_n34068_, new_n34069_, new_n34070_, new_n34071_, new_n34072_,
    new_n34073_, new_n34074_, new_n34075_, new_n34076_, new_n34077_,
    new_n34078_, new_n34079_, new_n34080_, new_n34081_, new_n34082_,
    new_n34083_, new_n34084_, new_n34085_, new_n34086_, new_n34087_,
    new_n34088_, new_n34089_, new_n34090_, new_n34091_, new_n34092_,
    new_n34093_, new_n34094_, new_n34095_, new_n34096_, new_n34097_,
    new_n34098_, new_n34099_, new_n34100_, new_n34101_, new_n34102_,
    new_n34103_, new_n34104_, new_n34105_, new_n34106_, new_n34107_,
    new_n34108_, new_n34109_, new_n34110_, new_n34111_, new_n34112_,
    new_n34113_, new_n34114_, new_n34115_, new_n34116_, new_n34117_,
    new_n34118_, new_n34119_, new_n34120_, new_n34121_, new_n34122_,
    new_n34123_, new_n34124_, new_n34125_, new_n34126_, new_n34127_,
    new_n34128_, new_n34129_, new_n34130_, new_n34131_, new_n34132_,
    new_n34133_, new_n34134_, new_n34135_, new_n34136_, new_n34137_,
    new_n34138_, new_n34139_, new_n34140_, new_n34141_, new_n34142_,
    new_n34143_, new_n34144_, new_n34145_, new_n34146_, new_n34147_,
    new_n34148_, new_n34149_, new_n34150_, new_n34151_, new_n34152_,
    new_n34153_, new_n34154_, new_n34155_, new_n34156_, new_n34157_,
    new_n34158_, new_n34159_, new_n34160_, new_n34161_, new_n34162_,
    new_n34163_, new_n34164_, new_n34165_, new_n34166_, new_n34167_,
    new_n34168_, new_n34169_, new_n34170_, new_n34171_, new_n34172_,
    new_n34173_, new_n34174_, new_n34175_, new_n34176_, new_n34177_,
    new_n34178_, new_n34179_, new_n34180_, new_n34181_, new_n34182_,
    new_n34183_, new_n34184_, new_n34185_, new_n34186_, new_n34187_,
    new_n34188_, new_n34189_, new_n34190_, new_n34191_, new_n34192_,
    new_n34193_, new_n34194_, new_n34195_, new_n34196_, new_n34197_,
    new_n34198_, new_n34199_, new_n34200_, new_n34201_, new_n34202_,
    new_n34203_, new_n34204_, new_n34205_, new_n34206_, new_n34207_,
    new_n34208_, new_n34209_, new_n34210_, new_n34211_, new_n34212_,
    new_n34213_, new_n34214_, new_n34215_, new_n34216_, new_n34217_,
    new_n34218_, new_n34219_, new_n34220_, new_n34221_, new_n34222_,
    new_n34223_, new_n34224_, new_n34225_, new_n34226_, new_n34227_,
    new_n34228_, new_n34229_, new_n34230_, new_n34231_, new_n34232_,
    new_n34233_, new_n34234_, new_n34235_, new_n34236_, new_n34237_,
    new_n34238_, new_n34239_, new_n34240_, new_n34241_, new_n34242_,
    new_n34243_, new_n34244_, new_n34245_, new_n34246_, new_n34247_,
    new_n34248_, new_n34249_, new_n34250_, new_n34251_, new_n34252_,
    new_n34253_, new_n34254_, new_n34255_, new_n34256_, new_n34257_,
    new_n34258_, new_n34259_, new_n34260_, new_n34261_, new_n34262_,
    new_n34263_, new_n34264_, new_n34265_, new_n34266_, new_n34267_,
    new_n34268_, new_n34269_, new_n34270_, new_n34271_, new_n34272_,
    new_n34273_, new_n34274_, new_n34275_, new_n34276_, new_n34277_,
    new_n34278_, new_n34279_, new_n34280_, new_n34281_, new_n34282_,
    new_n34283_, new_n34284_, new_n34285_, new_n34286_, new_n34287_,
    new_n34288_, new_n34289_, new_n34290_, new_n34291_, new_n34292_,
    new_n34293_, new_n34294_, new_n34295_, new_n34296_, new_n34297_,
    new_n34298_, new_n34299_, new_n34300_, new_n34301_, new_n34302_,
    new_n34303_, new_n34304_, new_n34305_, new_n34306_, new_n34307_,
    new_n34308_, new_n34309_, new_n34310_, new_n34311_, new_n34312_,
    new_n34313_, new_n34314_, new_n34315_, new_n34316_, new_n34317_,
    new_n34318_, new_n34319_, new_n34320_, new_n34321_, new_n34322_,
    new_n34323_, new_n34324_, new_n34325_, new_n34326_, new_n34327_,
    new_n34328_, new_n34329_, new_n34330_, new_n34331_, new_n34332_,
    new_n34333_, new_n34334_, new_n34335_, new_n34336_, new_n34337_,
    new_n34338_, new_n34339_, new_n34340_, new_n34341_, new_n34342_,
    new_n34343_, new_n34344_, new_n34345_, new_n34346_, new_n34347_,
    new_n34348_, new_n34349_, new_n34350_, new_n34351_, new_n34352_,
    new_n34353_, new_n34354_, new_n34355_, new_n34356_, new_n34357_,
    new_n34358_, new_n34359_, new_n34360_, new_n34361_, new_n34362_,
    new_n34363_, new_n34364_, new_n34365_, new_n34366_, new_n34367_,
    new_n34368_, new_n34369_, new_n34370_, new_n34371_, new_n34372_,
    new_n34373_, new_n34374_, new_n34375_, new_n34376_, new_n34377_,
    new_n34378_, new_n34379_, new_n34380_, new_n34381_, new_n34382_,
    new_n34383_, new_n34384_, new_n34385_, new_n34386_, new_n34387_,
    new_n34388_, new_n34389_, new_n34390_, new_n34391_, new_n34392_,
    new_n34393_, new_n34394_, new_n34395_, new_n34396_, new_n34397_,
    new_n34398_, new_n34399_, new_n34400_, new_n34401_, new_n34402_,
    new_n34403_, new_n34404_, new_n34405_, new_n34406_, new_n34407_,
    new_n34408_, new_n34409_, new_n34410_, new_n34411_, new_n34412_,
    new_n34413_, new_n34414_, new_n34415_, new_n34416_, new_n34417_,
    new_n34418_, new_n34419_, new_n34420_, new_n34421_, new_n34422_,
    new_n34423_, new_n34424_, new_n34425_, new_n34426_, new_n34427_,
    new_n34428_, new_n34429_, new_n34430_, new_n34431_, new_n34432_,
    new_n34433_, new_n34434_, new_n34435_, new_n34436_, new_n34437_,
    new_n34438_, new_n34439_, new_n34440_, new_n34441_, new_n34442_,
    new_n34443_, new_n34444_, new_n34445_, new_n34446_, new_n34447_,
    new_n34448_, new_n34449_, new_n34450_, new_n34451_, new_n34452_,
    new_n34453_, new_n34454_, new_n34455_, new_n34456_, new_n34457_,
    new_n34458_, new_n34459_, new_n34460_, new_n34461_, new_n34462_,
    new_n34463_, new_n34464_, new_n34465_, new_n34466_, new_n34467_,
    new_n34468_, new_n34469_, new_n34470_, new_n34471_, new_n34472_,
    new_n34473_, new_n34474_, new_n34475_, new_n34476_, new_n34477_,
    new_n34478_, new_n34479_, new_n34480_, new_n34481_, new_n34482_,
    new_n34483_, new_n34484_, new_n34485_, new_n34486_, new_n34487_,
    new_n34488_, new_n34489_, new_n34490_, new_n34491_, new_n34492_,
    new_n34493_, new_n34494_, new_n34495_, new_n34496_, new_n34497_,
    new_n34498_, new_n34499_, new_n34500_, new_n34501_, new_n34502_,
    new_n34503_, new_n34504_, new_n34505_, new_n34506_, new_n34507_,
    new_n34508_, new_n34509_, new_n34510_, new_n34511_, new_n34512_,
    new_n34513_, new_n34514_, new_n34515_, new_n34516_, new_n34517_,
    new_n34518_, new_n34519_, new_n34520_, new_n34521_, new_n34522_,
    new_n34523_, new_n34524_, new_n34525_, new_n34526_, new_n34527_,
    new_n34528_, new_n34529_, new_n34530_, new_n34531_, new_n34532_,
    new_n34533_, new_n34534_, new_n34535_, new_n34536_, new_n34537_,
    new_n34538_, new_n34539_, new_n34540_, new_n34541_, new_n34542_,
    new_n34543_, new_n34544_, new_n34545_, new_n34546_, new_n34547_,
    new_n34548_, new_n34549_, new_n34550_, new_n34551_, new_n34552_,
    new_n34553_, new_n34554_, new_n34555_, new_n34556_, new_n34557_,
    new_n34558_, new_n34559_, new_n34560_, new_n34561_, new_n34562_,
    new_n34563_, new_n34564_, new_n34565_, new_n34566_, new_n34567_,
    new_n34568_, new_n34569_, new_n34570_, new_n34571_, new_n34572_,
    new_n34573_, new_n34574_, new_n34575_, new_n34576_, new_n34577_,
    new_n34578_, new_n34579_, new_n34580_, new_n34581_, new_n34582_,
    new_n34583_, new_n34584_, new_n34585_, new_n34586_, new_n34587_,
    new_n34588_, new_n34589_, new_n34590_, new_n34591_, new_n34592_,
    new_n34593_, new_n34594_, new_n34595_, new_n34596_, new_n34597_,
    new_n34598_, new_n34599_, new_n34600_, new_n34601_, new_n34602_,
    new_n34603_, new_n34604_, new_n34605_, new_n34606_, new_n34607_,
    new_n34608_, new_n34609_, new_n34610_, new_n34611_, new_n34612_,
    new_n34613_, new_n34614_, new_n34615_, new_n34616_, new_n34617_,
    new_n34618_, new_n34619_, new_n34620_, new_n34621_, new_n34622_,
    new_n34623_, new_n34624_, new_n34625_, new_n34626_, new_n34627_,
    new_n34628_, new_n34629_, new_n34630_, new_n34631_, new_n34632_,
    new_n34633_, new_n34634_, new_n34635_, new_n34636_, new_n34637_,
    new_n34638_, new_n34639_, new_n34640_, new_n34641_, new_n34642_,
    new_n34643_, new_n34644_, new_n34645_, new_n34646_, new_n34647_,
    new_n34648_, new_n34649_, new_n34650_, new_n34651_, new_n34652_,
    new_n34653_, new_n34654_, new_n34655_, new_n34656_, new_n34657_,
    new_n34658_, new_n34659_, new_n34660_, new_n34661_, new_n34662_,
    new_n34663_, new_n34664_, new_n34665_, new_n34666_, new_n34667_,
    new_n34668_, new_n34669_, new_n34670_, new_n34671_, new_n34672_,
    new_n34673_, new_n34674_, new_n34675_, new_n34676_, new_n34677_,
    new_n34678_, new_n34679_, new_n34680_, new_n34681_, new_n34682_,
    new_n34683_, new_n34684_, new_n34685_, new_n34686_, new_n34687_,
    new_n34688_, new_n34689_, new_n34690_, new_n34691_, new_n34692_,
    new_n34693_, new_n34694_, new_n34695_, new_n34696_, new_n34697_,
    new_n34698_, new_n34699_, new_n34700_, new_n34701_, new_n34702_,
    new_n34703_, new_n34704_, new_n34705_, new_n34706_, new_n34707_,
    new_n34708_, new_n34709_, new_n34710_, new_n34711_, new_n34712_,
    new_n34713_, new_n34714_, new_n34715_, new_n34716_, new_n34717_,
    new_n34718_, new_n34719_, new_n34720_, new_n34721_, new_n34722_,
    new_n34723_, new_n34724_, new_n34725_, new_n34726_, new_n34727_,
    new_n34728_, new_n34729_, new_n34730_, new_n34731_, new_n34732_,
    new_n34733_, new_n34734_, new_n34735_, new_n34736_, new_n34737_,
    new_n34738_, new_n34739_, new_n34740_, new_n34741_, new_n34742_,
    new_n34743_, new_n34744_, new_n34745_, new_n34746_, new_n34747_,
    new_n34748_, new_n34749_, new_n34750_, new_n34751_, new_n34752_,
    new_n34753_, new_n34754_, new_n34755_, new_n34756_, new_n34757_,
    new_n34758_, new_n34759_, new_n34760_, new_n34761_, new_n34762_,
    new_n34763_, new_n34764_, new_n34765_, new_n34766_, new_n34767_,
    new_n34768_, new_n34769_, new_n34770_, new_n34771_, new_n34772_,
    new_n34773_, new_n34774_, new_n34775_, new_n34776_, new_n34777_,
    new_n34778_, new_n34779_, new_n34780_, new_n34781_, new_n34782_,
    new_n34783_, new_n34784_, new_n34785_, new_n34786_, new_n34787_,
    new_n34788_, new_n34789_, new_n34790_, new_n34791_, new_n34792_,
    new_n34793_, new_n34794_, new_n34795_, new_n34796_, new_n34797_,
    new_n34798_, new_n34799_, new_n34800_, new_n34801_, new_n34802_,
    new_n34803_, new_n34804_, new_n34805_, new_n34806_, new_n34807_,
    new_n34808_, new_n34809_, new_n34810_, new_n34811_, new_n34812_,
    new_n34813_, new_n34814_, new_n34815_, new_n34816_, new_n34817_,
    new_n34818_, new_n34819_, new_n34820_, new_n34821_, new_n34822_,
    new_n34823_, new_n34824_, new_n34825_, new_n34826_, new_n34827_,
    new_n34828_, new_n34829_, new_n34830_, new_n34831_, new_n34832_,
    new_n34833_, new_n34834_, new_n34835_, new_n34836_, new_n34837_,
    new_n34838_, new_n34839_, new_n34840_, new_n34841_, new_n34842_,
    new_n34843_, new_n34844_, new_n34845_, new_n34846_, new_n34847_,
    new_n34848_, new_n34849_, new_n34850_, new_n34851_, new_n34852_,
    new_n34853_, new_n34854_, new_n34855_, new_n34856_, new_n34857_,
    new_n34858_, new_n34859_, new_n34860_, new_n34861_, new_n34862_,
    new_n34863_, new_n34864_, new_n34865_, new_n34866_, new_n34867_,
    new_n34868_, new_n34869_, new_n34870_, new_n34871_, new_n34872_,
    new_n34873_, new_n34874_, new_n34875_, new_n34876_, new_n34877_,
    new_n34878_, new_n34879_, new_n34880_, new_n34881_, new_n34882_,
    new_n34883_, new_n34884_, new_n34885_, new_n34886_, new_n34887_,
    new_n34888_, new_n34889_, new_n34890_, new_n34891_, new_n34892_,
    new_n34893_, new_n34894_, new_n34895_, new_n34896_, new_n34897_,
    new_n34898_, new_n34899_, new_n34900_, new_n34901_, new_n34902_,
    new_n34903_, new_n34904_, new_n34905_, new_n34906_, new_n34907_,
    new_n34908_, new_n34909_, new_n34910_, new_n34911_, new_n34912_,
    new_n34913_, new_n34914_, new_n34915_, new_n34916_, new_n34917_,
    new_n34918_, new_n34919_, new_n34920_, new_n34921_, new_n34922_,
    new_n34923_, new_n34924_, new_n34925_, new_n34926_, new_n34927_,
    new_n34928_, new_n34929_, new_n34930_, new_n34931_, new_n34932_,
    new_n34933_, new_n34934_, new_n34935_, new_n34936_, new_n34937_,
    new_n34938_, new_n34939_, new_n34940_, new_n34941_, new_n34942_,
    new_n34943_, new_n34944_, new_n34945_, new_n34946_, new_n34947_,
    new_n34948_, new_n34949_, new_n34950_, new_n34951_, new_n34952_,
    new_n34953_, new_n34954_, new_n34955_, new_n34956_, new_n34957_,
    new_n34958_, new_n34959_, new_n34960_, new_n34961_, new_n34962_,
    new_n34963_, new_n34964_, new_n34965_, new_n34966_, new_n34967_,
    new_n34968_, new_n34969_, new_n34970_, new_n34971_, new_n34972_,
    new_n34973_, new_n34974_, new_n34975_, new_n34976_, new_n34977_,
    new_n34978_, new_n34979_, new_n34980_, new_n34981_, new_n34982_,
    new_n34983_, new_n34984_, new_n34985_, new_n34986_, new_n34987_,
    new_n34988_, new_n34989_, new_n34990_, new_n34991_, new_n34992_,
    new_n34993_, new_n34994_, new_n34995_, new_n34996_, new_n34997_,
    new_n34998_, new_n34999_, new_n35000_, new_n35001_, new_n35002_,
    new_n35003_, new_n35004_, new_n35005_, new_n35006_, new_n35007_,
    new_n35008_, new_n35009_, new_n35010_, new_n35011_, new_n35012_,
    new_n35013_, new_n35014_, new_n35015_, new_n35016_, new_n35017_,
    new_n35018_, new_n35019_, new_n35020_, new_n35021_, new_n35022_,
    new_n35023_, new_n35024_, new_n35025_, new_n35026_, new_n35027_,
    new_n35028_, new_n35029_, new_n35030_, new_n35031_, new_n35032_,
    new_n35033_, new_n35034_, new_n35035_, new_n35036_, new_n35037_,
    new_n35038_, new_n35039_, new_n35040_, new_n35041_, new_n35042_,
    new_n35043_, new_n35044_, new_n35045_, new_n35046_, new_n35047_,
    new_n35048_, new_n35049_, new_n35050_, new_n35051_, new_n35052_,
    new_n35053_, new_n35054_, new_n35055_, new_n35056_, new_n35057_,
    new_n35058_, new_n35059_, new_n35060_, new_n35061_, new_n35062_,
    new_n35063_, new_n35064_, new_n35065_, new_n35066_, new_n35067_,
    new_n35068_, new_n35069_, new_n35070_, new_n35071_, new_n35072_,
    new_n35073_, new_n35074_, new_n35075_, new_n35076_, new_n35077_,
    new_n35078_, new_n35079_, new_n35080_, new_n35081_, new_n35082_,
    new_n35083_, new_n35084_, new_n35085_, new_n35086_, new_n35087_,
    new_n35088_, new_n35089_, new_n35090_, new_n35091_, new_n35092_,
    new_n35093_, new_n35094_, new_n35095_, new_n35096_, new_n35097_,
    new_n35098_, new_n35099_, new_n35100_, new_n35101_, new_n35102_,
    new_n35103_, new_n35104_, new_n35105_, new_n35106_, new_n35107_,
    new_n35108_, new_n35109_, new_n35110_, new_n35111_, new_n35112_,
    new_n35113_, new_n35114_, new_n35115_, new_n35116_, new_n35117_,
    new_n35118_, new_n35119_, new_n35120_, new_n35121_, new_n35122_,
    new_n35123_, new_n35124_, new_n35125_, new_n35126_, new_n35127_,
    new_n35128_, new_n35129_, new_n35130_, new_n35131_, new_n35132_,
    new_n35133_, new_n35134_, new_n35135_, new_n35136_, new_n35137_,
    new_n35138_, new_n35139_, new_n35140_, new_n35141_, new_n35142_,
    new_n35143_, new_n35144_, new_n35145_, new_n35146_, new_n35147_,
    new_n35148_, new_n35149_, new_n35150_, new_n35151_, new_n35152_,
    new_n35153_, new_n35154_, new_n35155_, new_n35156_, new_n35157_,
    new_n35158_, new_n35159_, new_n35160_, new_n35161_, new_n35162_,
    new_n35163_, new_n35164_, new_n35165_, new_n35166_, new_n35167_,
    new_n35168_, new_n35169_, new_n35170_, new_n35171_, new_n35172_,
    new_n35173_, new_n35174_, new_n35175_, new_n35176_, new_n35177_,
    new_n35178_, new_n35179_, new_n35180_, new_n35181_, new_n35182_,
    new_n35183_, new_n35184_, new_n35185_, new_n35186_, new_n35187_,
    new_n35188_, new_n35189_, new_n35190_, new_n35191_, new_n35192_,
    new_n35193_, new_n35194_, new_n35195_, new_n35196_, new_n35197_,
    new_n35198_, new_n35199_, new_n35200_, new_n35201_, new_n35202_,
    new_n35203_, new_n35204_, new_n35205_, new_n35206_, new_n35207_,
    new_n35208_, new_n35209_, new_n35210_, new_n35211_, new_n35212_,
    new_n35213_, new_n35214_, new_n35215_, new_n35216_, new_n35217_,
    new_n35218_, new_n35219_, new_n35220_, new_n35221_, new_n35222_,
    new_n35223_, new_n35224_, new_n35225_, new_n35226_, new_n35227_,
    new_n35228_, new_n35229_, new_n35230_, new_n35231_, new_n35232_,
    new_n35233_, new_n35234_, new_n35235_, new_n35236_, new_n35237_,
    new_n35238_, new_n35239_, new_n35240_, new_n35241_, new_n35242_,
    new_n35243_, new_n35244_, new_n35245_, new_n35246_, new_n35247_,
    new_n35248_, new_n35249_, new_n35250_, new_n35251_, new_n35252_,
    new_n35253_, new_n35254_, new_n35255_, new_n35256_, new_n35257_,
    new_n35258_, new_n35259_, new_n35260_, new_n35261_, new_n35262_,
    new_n35263_, new_n35264_, new_n35265_, new_n35266_, new_n35267_,
    new_n35268_, new_n35269_, new_n35270_, new_n35271_, new_n35272_,
    new_n35273_, new_n35274_, new_n35275_, new_n35276_, new_n35277_,
    new_n35278_, new_n35279_, new_n35280_, new_n35281_, new_n35282_,
    new_n35283_, new_n35284_, new_n35285_, new_n35286_, new_n35287_,
    new_n35288_, new_n35289_, new_n35290_, new_n35291_, new_n35292_,
    new_n35293_, new_n35294_, new_n35295_, new_n35296_, new_n35297_,
    new_n35298_, new_n35299_, new_n35300_, new_n35301_, new_n35302_,
    new_n35303_, new_n35304_, new_n35305_, new_n35306_, new_n35307_,
    new_n35308_, new_n35309_, new_n35310_, new_n35311_, new_n35312_,
    new_n35313_, new_n35314_, new_n35315_, new_n35316_, new_n35317_,
    new_n35318_, new_n35319_, new_n35320_, new_n35321_, new_n35322_,
    new_n35323_, new_n35324_, new_n35325_, new_n35326_, new_n35327_,
    new_n35328_, new_n35329_, new_n35330_, new_n35331_, new_n35332_,
    new_n35333_, new_n35334_, new_n35335_, new_n35336_, new_n35337_,
    new_n35338_, new_n35339_, new_n35340_, new_n35341_, new_n35342_,
    new_n35343_, new_n35344_, new_n35345_, new_n35346_, new_n35347_,
    new_n35348_, new_n35349_, new_n35350_, new_n35351_, new_n35352_,
    new_n35353_, new_n35354_, new_n35355_, new_n35356_, new_n35357_,
    new_n35358_, new_n35359_, new_n35360_, new_n35361_, new_n35362_,
    new_n35363_, new_n35364_, new_n35365_, new_n35366_, new_n35367_,
    new_n35368_, new_n35369_, new_n35370_, new_n35371_, new_n35372_,
    new_n35373_, new_n35374_, new_n35375_, new_n35376_, new_n35377_,
    new_n35378_, new_n35379_, new_n35380_, new_n35381_, new_n35382_,
    new_n35383_, new_n35384_, new_n35385_, new_n35386_, new_n35387_,
    new_n35388_, new_n35389_, new_n35390_, new_n35391_, new_n35392_,
    new_n35393_, new_n35394_, new_n35395_, new_n35396_, new_n35397_,
    new_n35398_, new_n35399_, new_n35400_, new_n35401_, new_n35402_,
    new_n35403_, new_n35404_, new_n35405_, new_n35406_, new_n35407_,
    new_n35408_, new_n35409_, new_n35410_, new_n35411_, new_n35412_,
    new_n35413_, new_n35414_, new_n35415_, new_n35416_, new_n35417_,
    new_n35418_, new_n35419_, new_n35420_, new_n35421_, new_n35422_,
    new_n35423_, new_n35424_, new_n35425_, new_n35426_, new_n35427_,
    new_n35428_, new_n35429_, new_n35430_, new_n35431_, new_n35432_,
    new_n35433_, new_n35434_, new_n35435_, new_n35436_, new_n35437_,
    new_n35438_, new_n35439_, new_n35440_, new_n35441_, new_n35442_,
    new_n35443_, new_n35444_, new_n35445_, new_n35446_, new_n35447_,
    new_n35448_, new_n35449_, new_n35450_, new_n35451_, new_n35452_,
    new_n35453_, new_n35454_, new_n35455_, new_n35456_, new_n35457_,
    new_n35458_, new_n35459_, new_n35460_, new_n35461_, new_n35462_,
    new_n35463_, new_n35464_, new_n35465_, new_n35466_, new_n35467_,
    new_n35468_, new_n35469_, new_n35470_, new_n35471_, new_n35472_,
    new_n35473_, new_n35474_, new_n35475_, new_n35476_, new_n35477_,
    new_n35478_, new_n35479_, new_n35480_, new_n35481_, new_n35482_,
    new_n35483_, new_n35484_, new_n35485_, new_n35486_, new_n35487_,
    new_n35488_, new_n35489_, new_n35490_, new_n35491_, new_n35492_,
    new_n35493_, new_n35494_, new_n35495_, new_n35496_, new_n35497_,
    new_n35498_, new_n35499_, new_n35500_, new_n35501_, new_n35502_,
    new_n35503_, new_n35504_, new_n35505_, new_n35506_, new_n35507_,
    new_n35508_, new_n35509_, new_n35510_, new_n35511_, new_n35512_,
    new_n35513_, new_n35514_, new_n35515_, new_n35516_, new_n35517_,
    new_n35518_, new_n35519_, new_n35520_, new_n35521_, new_n35522_,
    new_n35523_, new_n35524_, new_n35525_, new_n35526_, new_n35527_,
    new_n35528_, new_n35529_, new_n35530_, new_n35531_, new_n35532_,
    new_n35533_, new_n35534_, new_n35535_, new_n35536_, new_n35537_,
    new_n35538_, new_n35539_, new_n35540_, new_n35541_, new_n35542_,
    new_n35543_, new_n35544_, new_n35545_, new_n35546_, new_n35547_,
    new_n35548_, new_n35549_, new_n35550_, new_n35551_, new_n35552_,
    new_n35553_, new_n35554_, new_n35555_, new_n35556_, new_n35557_,
    new_n35558_, new_n35559_, new_n35560_, new_n35561_, new_n35562_,
    new_n35563_, new_n35564_, new_n35565_, new_n35566_, new_n35567_,
    new_n35568_, new_n35569_, new_n35570_, new_n35571_, new_n35572_,
    new_n35573_, new_n35574_, new_n35575_, new_n35576_, new_n35577_,
    new_n35578_, new_n35579_, new_n35580_, new_n35581_, new_n35582_,
    new_n35583_, new_n35584_, new_n35585_, new_n35586_, new_n35587_,
    new_n35588_, new_n35589_, new_n35590_, new_n35591_, new_n35592_,
    new_n35593_, new_n35594_, new_n35595_, new_n35596_, new_n35597_,
    new_n35598_, new_n35599_, new_n35600_, new_n35601_, new_n35602_,
    new_n35603_, new_n35604_, new_n35605_, new_n35606_, new_n35607_,
    new_n35608_, new_n35609_, new_n35610_, new_n35611_, new_n35612_,
    new_n35613_, new_n35614_, new_n35615_, new_n35616_, new_n35617_,
    new_n35618_, new_n35619_, new_n35620_, new_n35621_, new_n35622_,
    new_n35623_, new_n35624_, new_n35625_, new_n35626_, new_n35627_,
    new_n35628_, new_n35629_, new_n35630_, new_n35631_, new_n35632_,
    new_n35633_, new_n35634_, new_n35635_, new_n35636_, new_n35637_,
    new_n35638_, new_n35639_, new_n35640_, new_n35641_, new_n35642_,
    new_n35643_, new_n35644_, new_n35645_, new_n35646_, new_n35647_,
    new_n35648_, new_n35649_, new_n35650_, new_n35651_, new_n35652_,
    new_n35653_, new_n35654_, new_n35655_, new_n35656_, new_n35657_,
    new_n35658_, new_n35659_, new_n35660_, new_n35661_, new_n35662_,
    new_n35663_, new_n35664_, new_n35665_, new_n35666_, new_n35667_,
    new_n35668_, new_n35669_, new_n35670_, new_n35671_, new_n35672_,
    new_n35673_, new_n35674_, new_n35675_, new_n35676_, new_n35677_,
    new_n35678_, new_n35679_, new_n35680_, new_n35681_, new_n35682_,
    new_n35683_, new_n35684_, new_n35685_, new_n35686_, new_n35687_,
    new_n35688_, new_n35689_, new_n35690_, new_n35691_, new_n35692_,
    new_n35693_, new_n35694_, new_n35695_, new_n35696_, new_n35697_,
    new_n35698_, new_n35699_, new_n35700_, new_n35701_, new_n35702_,
    new_n35703_, new_n35704_, new_n35705_, new_n35706_, new_n35707_,
    new_n35708_, new_n35709_, new_n35710_, new_n35711_, new_n35712_,
    new_n35713_, new_n35714_, new_n35715_, new_n35716_, new_n35717_,
    new_n35718_, new_n35719_, new_n35720_, new_n35721_, new_n35722_,
    new_n35723_, new_n35724_, new_n35725_, new_n35726_, new_n35727_,
    new_n35728_, new_n35729_, new_n35730_, new_n35731_, new_n35732_,
    new_n35733_, new_n35734_, new_n35735_, new_n35736_, new_n35737_,
    new_n35738_, new_n35739_, new_n35740_, new_n35741_, new_n35742_,
    new_n35743_, new_n35744_, new_n35745_, new_n35746_, new_n35747_,
    new_n35748_, new_n35749_, new_n35750_, new_n35751_, new_n35752_,
    new_n35753_, new_n35754_, new_n35755_, new_n35756_, new_n35757_,
    new_n35758_, new_n35759_, new_n35760_, new_n35761_, new_n35762_,
    new_n35763_, new_n35764_, new_n35765_, new_n35766_, new_n35767_,
    new_n35768_, new_n35769_, new_n35770_, new_n35771_, new_n35772_,
    new_n35773_, new_n35774_, new_n35775_, new_n35776_, new_n35777_,
    new_n35778_, new_n35779_, new_n35780_, new_n35781_, new_n35782_,
    new_n35783_, new_n35784_, new_n35785_, new_n35786_, new_n35787_,
    new_n35788_, new_n35789_, new_n35790_, new_n35791_, new_n35792_,
    new_n35793_, new_n35794_, new_n35795_, new_n35796_, new_n35797_,
    new_n35798_, new_n35799_, new_n35800_, new_n35801_, new_n35802_,
    new_n35803_, new_n35804_, new_n35805_, new_n35806_, new_n35807_,
    new_n35808_, new_n35809_, new_n35810_, new_n35811_, new_n35812_,
    new_n35813_, new_n35814_, new_n35815_, new_n35816_, new_n35817_,
    new_n35818_, new_n35819_, new_n35820_, new_n35821_, new_n35822_,
    new_n35823_, new_n35824_, new_n35825_, new_n35826_, new_n35827_,
    new_n35828_, new_n35829_, new_n35830_, new_n35831_, new_n35832_,
    new_n35833_, new_n35834_, new_n35835_, new_n35836_, new_n35837_,
    new_n35838_, new_n35839_, new_n35840_, new_n35841_, new_n35842_,
    new_n35843_, new_n35844_, new_n35845_, new_n35846_, new_n35847_,
    new_n35848_, new_n35849_, new_n35850_, new_n35851_, new_n35852_,
    new_n35853_, new_n35854_, new_n35855_, new_n35856_, new_n35857_,
    new_n35858_, new_n35859_, new_n35860_, new_n35861_, new_n35862_,
    new_n35863_, new_n35864_, new_n35865_, new_n35866_, new_n35867_,
    new_n35868_, new_n35869_;
xor  ( new_n98_, RI2b1c4342dbe8_80, RI2b1c4342db70_79 );
not  ( new_n99_, RI2b1c4342d4e0_65 );
xor  ( new_n100_, RI2b1c4342d558_66, new_n99_ );
xor  ( new_n101_, RI2b1c4342d738_70, RI2b1c4342d6c0_69 );
xor  ( new_n102_, new_n101_, new_n100_ );
xnor ( new_n103_, new_n102_, new_n98_ );
xor  ( new_n104_, RI2b1c4342da08_76, RI2b1c4342d990_75 );
not  ( new_n105_, RI2b1c4342d8a0_73 );
xor  ( new_n106_, RI2b1c4342d918_74, new_n105_ );
xor  ( new_n107_, RI2b1c4342daf8_78, RI2b1c4342da80_77 );
xor  ( new_n108_, new_n107_, new_n106_ );
xor  ( new_n109_, new_n108_, new_n104_ );
not  ( new_n110_, RI2b1c4342d7b0_71 );
xor  ( new_n111_, RI2b1c4342d828_72, new_n110_ );
not  ( new_n112_, RI2b1c4342d5d0_67 );
xor  ( new_n113_, RI2b1c4342d648_68, new_n112_ );
xor  ( new_n114_, new_n113_, new_n111_ );
xor  ( new_n115_, new_n114_, new_n109_ );
xor  ( new_n116_, new_n115_, new_n103_ );
not  ( new_n117_, RI2b1c4342e110_91 );
xor  ( new_n118_, RI2b1c4342e188_92, new_n117_ );
xnor ( new_n119_, new_n118_, new_n116_ );
xor  ( new_n120_, RI2b1c4342dfa8_88, RI2b1c4342df30_87 );
not  ( new_n121_, RI2b1c4342dd50_83 );
xor  ( new_n122_, RI2b1c4342ddc8_84, new_n121_ );
xor  ( new_n123_, new_n122_, new_n120_ );
not  ( new_n124_, RI2b1c4342e2f0_95 );
xor  ( new_n125_, RI2b1c4342e368_96, new_n124_ );
not  ( new_n126_, RI2b1c4342dc60_81 );
xor  ( new_n127_, RI2b1c4342dcd8_82, new_n126_ );
xor  ( new_n128_, RI2b1c4342deb8_86, RI2b1c4342de40_85 );
xor  ( new_n129_, new_n128_, new_n127_ );
xor  ( new_n130_, new_n129_, new_n125_ );
xor  ( new_n131_, new_n130_, new_n123_ );
not  ( new_n132_, RI2b1c4342e020_89 );
xor  ( new_n133_, RI2b1c4342e098_90, new_n132_ );
xor  ( new_n134_, RI2b1c4342e278_94, RI2b1c4342e200_93 );
xor  ( new_n135_, new_n134_, new_n133_ );
xor  ( new_n136_, new_n135_, new_n131_ );
xor  ( new_n137_, new_n136_, new_n119_ );
not  ( new_n138_, new_n137_ );
and  ( new_n139_, new_n138_, RI2b1c4342bc80_13 );
and  ( new_n140_, RI2b1c4342bcf8_14, RI2b1c4342cbf8_46 );
not  ( new_n141_, RI2b1c4342cbf8_46 );
not  ( new_n142_, RI2b1c4342bcf8_14 );
and  ( new_n143_, new_n142_, new_n141_ );
and  ( new_n144_, RI2b1c4342bd70_15, RI2b1c4342cc70_47 );
and  ( new_n145_, RI2b1c4342bde8_16, RI2b1c4342cce8_48 );
not  ( new_n146_, RI2b1c4342cce8_48 );
not  ( new_n147_, RI2b1c4342bde8_16 );
and  ( new_n148_, new_n147_, new_n146_ );
and  ( new_n149_, RI2b1c4342be60_17, RI2b1c4342cd60_49 );
not  ( new_n150_, RI2b1c4342cd60_49 );
not  ( new_n151_, RI2b1c4342be60_17 );
and  ( new_n152_, new_n151_, new_n150_ );
not  ( new_n153_, RI2b1c4342cdd8_50 );
not  ( new_n154_, RI2b1c4342bed8_18 );
and  ( new_n155_, new_n154_, new_n153_ );
and  ( new_n156_, RI2b1c4342bed8_18, RI2b1c4342cdd8_50 );
not  ( new_n157_, RI2b1c4342ce50_51 );
not  ( new_n158_, RI2b1c4342bf50_19 );
and  ( new_n159_, new_n158_, new_n157_ );
and  ( new_n160_, RI2b1c4342bf50_19, RI2b1c4342ce50_51 );
not  ( new_n161_, RI2b1c4342cec8_52 );
not  ( new_n162_, RI2b1c4342bfc8_20 );
and  ( new_n163_, new_n162_, new_n161_ );
and  ( new_n164_, RI2b1c4342bfc8_20, RI2b1c4342cec8_52 );
not  ( new_n165_, RI2b1c4342cf40_53 );
not  ( new_n166_, RI2b1c4342c040_21 );
and  ( new_n167_, new_n166_, new_n165_ );
and  ( new_n168_, RI2b1c4342c040_21, RI2b1c4342cf40_53 );
not  ( new_n169_, RI2b1c4342cfb8_54 );
not  ( new_n170_, RI2b1c4342c0b8_22 );
and  ( new_n171_, new_n170_, new_n169_ );
and  ( new_n172_, RI2b1c4342c0b8_22, RI2b1c4342cfb8_54 );
not  ( new_n173_, RI2b1c4342d030_55 );
not  ( new_n174_, RI2b1c4342c130_23 );
and  ( new_n175_, new_n174_, new_n173_ );
and  ( new_n176_, RI2b1c4342c130_23, RI2b1c4342d030_55 );
not  ( new_n177_, RI2b1c4342d0a8_56 );
not  ( new_n178_, RI2b1c4342c1a8_24 );
and  ( new_n179_, new_n178_, new_n177_ );
and  ( new_n180_, RI2b1c4342c1a8_24, RI2b1c4342d0a8_56 );
not  ( new_n181_, new_n180_ );
not  ( new_n182_, RI2b1c4342d120_57 );
not  ( new_n183_, RI2b1c4342c220_25 );
and  ( new_n184_, new_n183_, new_n182_ );
and  ( new_n185_, RI2b1c4342c220_25, RI2b1c4342d120_57 );
not  ( new_n186_, RI2b1c4342d198_58 );
not  ( new_n187_, RI2b1c4342c298_26 );
and  ( new_n188_, new_n187_, new_n186_ );
and  ( new_n189_, RI2b1c4342c298_26, RI2b1c4342d198_58 );
not  ( new_n190_, new_n189_ );
not  ( new_n191_, RI2b1c4342d210_59 );
not  ( new_n192_, RI2b1c4342c310_27 );
and  ( new_n193_, new_n192_, new_n191_ );
and  ( new_n194_, RI2b1c4342c310_27, RI2b1c4342d210_59 );
not  ( new_n195_, RI2b1c4342d288_60 );
not  ( new_n196_, RI2b1c4342c388_28 );
and  ( new_n197_, new_n196_, new_n195_ );
and  ( new_n198_, RI2b1c4342c388_28, RI2b1c4342d288_60 );
not  ( new_n199_, new_n198_ );
not  ( new_n200_, RI2b1c4342d300_61 );
not  ( new_n201_, RI2b1c4342c400_29 );
and  ( new_n202_, new_n201_, new_n200_ );
and  ( new_n203_, RI2b1c4342c400_29, RI2b1c4342d300_61 );
not  ( new_n204_, RI2b1c4342d378_62 );
not  ( new_n205_, RI2b1c4342c478_30 );
and  ( new_n206_, new_n205_, new_n204_ );
and  ( new_n207_, RI2b1c4342c478_30, RI2b1c4342d378_62 );
not  ( new_n208_, RI2b1c4342d3f0_63 );
not  ( new_n209_, RI2b1c4342c4f0_31 );
and  ( new_n210_, new_n209_, new_n208_ );
and  ( new_n211_, RI2b1c4342c4f0_31, RI2b1c4342d3f0_63 );
not  ( new_n212_, new_n211_ );
and  ( new_n213_, RI2b1c4342c568_32, RI2b1c4342d468_64 );
not  ( new_n214_, new_n213_ );
and  ( new_n215_, new_n214_, new_n212_ );
nor  ( new_n216_, new_n215_, new_n210_ );
nor  ( new_n217_, new_n216_, new_n207_ );
nor  ( new_n218_, new_n217_, new_n206_ );
nor  ( new_n219_, new_n218_, new_n203_ );
nor  ( new_n220_, new_n219_, new_n202_ );
not  ( new_n221_, new_n220_ );
and  ( new_n222_, new_n221_, new_n199_ );
nor  ( new_n223_, new_n222_, new_n197_ );
nor  ( new_n224_, new_n223_, new_n194_ );
nor  ( new_n225_, new_n224_, new_n193_ );
not  ( new_n226_, new_n225_ );
and  ( new_n227_, new_n226_, new_n190_ );
nor  ( new_n228_, new_n227_, new_n188_ );
nor  ( new_n229_, new_n228_, new_n185_ );
nor  ( new_n230_, new_n229_, new_n184_ );
not  ( new_n231_, new_n230_ );
and  ( new_n232_, new_n231_, new_n181_ );
nor  ( new_n233_, new_n232_, new_n179_ );
nor  ( new_n234_, new_n233_, new_n176_ );
nor  ( new_n235_, new_n234_, new_n175_ );
nor  ( new_n236_, new_n235_, new_n172_ );
nor  ( new_n237_, new_n236_, new_n171_ );
nor  ( new_n238_, new_n237_, new_n168_ );
nor  ( new_n239_, new_n238_, new_n167_ );
nor  ( new_n240_, new_n239_, new_n164_ );
nor  ( new_n241_, new_n240_, new_n163_ );
nor  ( new_n242_, new_n241_, new_n160_ );
nor  ( new_n243_, new_n242_, new_n159_ );
nor  ( new_n244_, new_n243_, new_n156_ );
nor  ( new_n245_, new_n244_, new_n155_ );
not  ( new_n246_, new_n245_ );
nor  ( new_n247_, new_n246_, new_n152_ );
nor  ( new_n248_, new_n247_, new_n149_ );
nor  ( new_n249_, new_n248_, new_n148_ );
nor  ( new_n250_, new_n249_, new_n145_ );
not  ( new_n251_, RI2b1c4342cc70_47 );
not  ( new_n252_, RI2b1c4342bd70_15 );
and  ( new_n253_, new_n252_, new_n251_ );
nor  ( new_n254_, new_n253_, new_n250_ );
nor  ( new_n255_, new_n254_, new_n144_ );
nor  ( new_n256_, new_n255_, new_n143_ );
nor  ( new_n257_, new_n256_, new_n140_ );
xor  ( new_n258_, RI2b1c4342bc80_13, RI2b1c4342cb80_45 );
nor  ( new_n259_, new_n258_, new_n257_ );
and  ( new_n260_, new_n138_, new_n142_ );
or   ( new_n261_, new_n260_, new_n141_ );
and  ( new_n262_, new_n138_, RI2b1c4342bcf8_14 );
not  ( new_n263_, new_n262_ );
and  ( new_n264_, new_n263_, new_n141_ );
and  ( new_n265_, new_n138_, RI2b1c4342bd70_15 );
not  ( new_n266_, new_n265_ );
and  ( new_n267_, new_n266_, new_n251_ );
and  ( new_n268_, new_n138_, new_n147_ );
or   ( new_n269_, new_n268_, new_n146_ );
and  ( new_n270_, new_n138_, RI2b1c4342bde8_16 );
not  ( new_n271_, new_n270_ );
and  ( new_n272_, new_n271_, new_n146_ );
and  ( new_n273_, new_n138_, RI2b1c4342be60_17 );
not  ( new_n274_, new_n273_ );
and  ( new_n275_, new_n274_, new_n150_ );
and  ( new_n276_, new_n138_, new_n154_ );
or   ( new_n277_, new_n276_, new_n153_ );
and  ( new_n278_, new_n138_, RI2b1c4342bed8_18 );
not  ( new_n279_, new_n278_ );
and  ( new_n280_, new_n279_, new_n153_ );
and  ( new_n281_, new_n138_, RI2b1c4342bf50_19 );
not  ( new_n282_, new_n281_ );
and  ( new_n283_, new_n282_, new_n157_ );
and  ( new_n284_, new_n138_, new_n158_ );
or   ( new_n285_, new_n284_, new_n157_ );
and  ( new_n286_, new_n138_, new_n162_ );
or   ( new_n287_, new_n286_, new_n161_ );
and  ( new_n288_, new_n138_, RI2b1c4342bfc8_20 );
not  ( new_n289_, new_n288_ );
and  ( new_n290_, new_n289_, new_n161_ );
and  ( new_n291_, new_n138_, RI2b1c4342c040_21 );
not  ( new_n292_, new_n291_ );
and  ( new_n293_, new_n292_, new_n165_ );
and  ( new_n294_, new_n138_, new_n166_ );
or   ( new_n295_, new_n294_, new_n165_ );
and  ( new_n296_, new_n138_, new_n170_ );
or   ( new_n297_, new_n296_, new_n169_ );
and  ( new_n298_, new_n138_, RI2b1c4342c0b8_22 );
not  ( new_n299_, new_n298_ );
and  ( new_n300_, new_n299_, new_n169_ );
and  ( new_n301_, new_n138_, RI2b1c4342c130_23 );
not  ( new_n302_, new_n301_ );
and  ( new_n303_, new_n302_, new_n173_ );
and  ( new_n304_, new_n138_, new_n174_ );
or   ( new_n305_, new_n304_, new_n173_ );
and  ( new_n306_, new_n138_, RI2b1c4342c1a8_24 );
not  ( new_n307_, new_n306_ );
and  ( new_n308_, new_n307_, new_n177_ );
and  ( new_n309_, new_n138_, RI2b1c4342c220_25 );
not  ( new_n310_, new_n309_ );
and  ( new_n311_, new_n310_, new_n182_ );
and  ( new_n312_, new_n138_, new_n183_ );
or   ( new_n313_, new_n312_, new_n182_ );
and  ( new_n314_, new_n138_, RI2b1c4342c298_26 );
not  ( new_n315_, new_n314_ );
and  ( new_n316_, new_n315_, new_n186_ );
and  ( new_n317_, new_n138_, RI2b1c4342c310_27 );
not  ( new_n318_, new_n317_ );
and  ( new_n319_, new_n318_, new_n191_ );
and  ( new_n320_, new_n138_, new_n192_ );
or   ( new_n321_, new_n320_, new_n191_ );
and  ( new_n322_, new_n138_, RI2b1c4342c388_28 );
not  ( new_n323_, new_n322_ );
and  ( new_n324_, new_n323_, new_n195_ );
and  ( new_n325_, new_n138_, RI2b1c4342c400_29 );
not  ( new_n326_, new_n325_ );
and  ( new_n327_, new_n326_, new_n200_ );
and  ( new_n328_, new_n138_, new_n201_ );
or   ( new_n329_, new_n328_, new_n200_ );
and  ( new_n330_, new_n138_, new_n205_ );
or   ( new_n331_, new_n330_, new_n204_ );
and  ( new_n332_, new_n138_, RI2b1c4342c478_30 );
not  ( new_n333_, new_n332_ );
and  ( new_n334_, new_n333_, new_n204_ );
and  ( new_n335_, new_n138_, RI2b1c4342c4f0_31 );
not  ( new_n336_, new_n335_ );
and  ( new_n337_, new_n336_, new_n208_ );
and  ( new_n338_, new_n214_, new_n138_ );
and  ( new_n339_, new_n338_, new_n212_ );
or   ( new_n340_, new_n339_, new_n337_ );
or   ( new_n341_, new_n340_, new_n334_ );
and  ( new_n342_, new_n341_, new_n331_ );
and  ( new_n343_, new_n342_, new_n329_ );
or   ( new_n344_, new_n343_, new_n327_ );
and  ( new_n345_, new_n344_, new_n138_ );
or   ( new_n346_, new_n345_, new_n324_ );
and  ( new_n347_, new_n346_, new_n199_ );
and  ( new_n348_, new_n347_, new_n321_ );
or   ( new_n349_, new_n348_, new_n319_ );
and  ( new_n350_, new_n349_, new_n138_ );
or   ( new_n351_, new_n350_, new_n316_ );
and  ( new_n352_, new_n351_, new_n190_ );
and  ( new_n353_, new_n352_, new_n313_ );
or   ( new_n354_, new_n353_, new_n311_ );
and  ( new_n355_, new_n354_, new_n138_ );
or   ( new_n356_, new_n355_, new_n308_ );
and  ( new_n357_, new_n356_, new_n181_ );
and  ( new_n358_, new_n357_, new_n305_ );
or   ( new_n359_, new_n358_, new_n303_ );
or   ( new_n360_, new_n359_, new_n300_ );
and  ( new_n361_, new_n360_, new_n297_ );
and  ( new_n362_, new_n361_, new_n295_ );
or   ( new_n363_, new_n362_, new_n293_ );
or   ( new_n364_, new_n363_, new_n290_ );
and  ( new_n365_, new_n364_, new_n287_ );
and  ( new_n366_, new_n365_, new_n285_ );
or   ( new_n367_, new_n366_, new_n283_ );
or   ( new_n368_, new_n367_, new_n280_ );
and  ( new_n369_, new_n368_, new_n277_ );
and  ( new_n370_, new_n138_, new_n151_ );
or   ( new_n371_, new_n370_, new_n150_ );
and  ( new_n372_, new_n371_, new_n369_ );
or   ( new_n373_, new_n372_, new_n275_ );
or   ( new_n374_, new_n373_, new_n272_ );
and  ( new_n375_, new_n374_, new_n269_ );
and  ( new_n376_, new_n138_, new_n252_ );
or   ( new_n377_, new_n376_, new_n251_ );
and  ( new_n378_, new_n377_, new_n375_ );
or   ( new_n379_, new_n378_, new_n267_ );
or   ( new_n380_, new_n379_, new_n264_ );
and  ( new_n381_, new_n380_, new_n261_ );
and  ( new_n382_, new_n381_, new_n258_ );
or   ( new_n383_, new_n382_, new_n259_ );
and  ( new_n384_, new_n383_, new_n139_ );
and  ( new_n385_, new_n138_, RI2b1c4342bc08_12 );
and  ( new_n386_, RI2b1c4342bc80_13, RI2b1c4342cb80_45 );
not  ( new_n387_, RI2b1c4342cb80_45 );
not  ( new_n388_, RI2b1c4342bc80_13 );
and  ( new_n389_, new_n388_, new_n387_ );
nor  ( new_n390_, new_n389_, new_n257_ );
nor  ( new_n391_, new_n390_, new_n386_ );
xor  ( new_n392_, RI2b1c4342bc08_12, RI2b1c4342cb08_44 );
nor  ( new_n393_, new_n392_, new_n391_ );
not  ( new_n394_, new_n139_ );
and  ( new_n395_, new_n394_, new_n387_ );
and  ( new_n396_, new_n138_, new_n388_ );
or   ( new_n397_, new_n396_, new_n387_ );
and  ( new_n398_, new_n397_, new_n381_ );
or   ( new_n399_, new_n398_, new_n395_ );
and  ( new_n400_, new_n399_, new_n392_ );
or   ( new_n401_, new_n400_, new_n393_ );
and  ( new_n402_, new_n401_, new_n385_ );
and  ( new_n403_, new_n402_, new_n384_ );
not  ( new_n404_, RI2b1c4342cb08_44 );
not  ( new_n405_, RI2b1c4342bc08_12 );
and  ( new_n406_, new_n138_, new_n405_ );
or   ( new_n407_, new_n406_, new_n404_ );
not  ( new_n408_, new_n385_ );
and  ( new_n409_, new_n408_, new_n404_ );
or   ( new_n410_, new_n409_, new_n399_ );
and  ( new_n411_, new_n410_, new_n407_ );
not  ( new_n412_, RI2b1c4342ca90_43 );
and  ( new_n413_, new_n138_, RI2b1c4342bb90_11 );
xor  ( new_n414_, new_n413_, new_n412_ );
and  ( new_n415_, new_n414_, new_n411_ );
not  ( new_n416_, RI2b1c4342bb90_11 );
and  ( new_n417_, RI2b1c4342bc08_12, RI2b1c4342cb08_44 );
and  ( new_n418_, new_n405_, new_n404_ );
nor  ( new_n419_, new_n418_, new_n391_ );
nor  ( new_n420_, new_n419_, new_n417_ );
and  ( new_n421_, new_n416_, new_n412_ );
nor  ( new_n422_, new_n421_, new_n420_ );
and  ( new_n423_, RI2b1c4342bb90_11, RI2b1c4342ca90_43 );
nor  ( new_n424_, new_n423_, new_n137_ );
and  ( new_n425_, new_n424_, new_n422_ );
or   ( new_n426_, new_n425_, new_n416_ );
or   ( new_n427_, new_n426_, new_n415_ );
or   ( new_n428_, new_n427_, new_n403_ );
xor  ( new_n429_, RI2b1c4342bb90_11, RI2b1c4342ca90_43 );
nor  ( new_n430_, new_n429_, new_n420_ );
and  ( new_n431_, new_n429_, new_n411_ );
or   ( new_n432_, new_n431_, new_n430_ );
and  ( new_n433_, new_n432_, new_n413_ );
and  ( new_n434_, new_n433_, new_n402_ );
and  ( new_n435_, new_n417_, new_n138_ );
or   ( new_n436_, new_n435_, new_n409_ );
and  ( new_n437_, new_n436_, new_n399_ );
nand ( new_n438_, new_n392_, new_n138_ );
nor  ( new_n439_, new_n438_, new_n391_ );
or   ( new_n440_, new_n439_, new_n405_ );
or   ( new_n441_, new_n440_, new_n437_ );
and  ( new_n442_, new_n441_, new_n427_ );
xor  ( new_n443_, new_n139_, new_n387_ );
and  ( new_n444_, new_n443_, new_n381_ );
nand ( new_n445_, new_n258_, new_n138_ );
nor  ( new_n446_, new_n445_, new_n257_ );
or   ( new_n447_, new_n446_, new_n388_ );
or   ( new_n448_, new_n447_, new_n444_ );
and  ( new_n449_, new_n448_, new_n402_ );
and  ( new_n450_, new_n441_, new_n384_ );
or   ( new_n451_, new_n450_, new_n449_ );
or   ( new_n452_, new_n451_, new_n442_ );
or   ( new_n453_, new_n452_, new_n434_ );
or   ( new_n454_, new_n453_, new_n99_ );
and  ( new_n455_, new_n454_, new_n428_ );
or   ( new_n456_, new_n448_, new_n441_ );
and  ( new_n457_, new_n456_, new_n433_ );
and  ( new_n458_, new_n448_, new_n441_ );
or   ( new_n459_, new_n458_, new_n403_ );
and  ( new_n460_, new_n441_, new_n433_ );
and  ( new_n461_, new_n427_, new_n402_ );
or   ( new_n462_, new_n461_, new_n460_ );
and  ( new_n463_, new_n462_, new_n459_ );
and  ( new_n464_, new_n463_, RI2b1c4342d4e0_65 );
and  ( new_n465_, new_n464_, new_n457_ );
or   ( new_n466_, new_n465_, new_n455_ );
not  ( new_n467_, RI2b1c4342ca18_42 );
not  ( new_n468_, RI2b1c4342bb18_10 );
and  ( new_n469_, new_n138_, new_n468_ );
or   ( new_n470_, new_n469_, new_n467_ );
not  ( new_n471_, new_n413_ );
and  ( new_n472_, new_n471_, new_n412_ );
and  ( new_n473_, new_n138_, new_n416_ );
or   ( new_n474_, new_n473_, new_n412_ );
and  ( new_n475_, new_n474_, new_n411_ );
or   ( new_n476_, new_n475_, new_n472_ );
and  ( new_n477_, new_n138_, RI2b1c4342bb18_10 );
not  ( new_n478_, new_n477_ );
and  ( new_n479_, new_n478_, new_n467_ );
or   ( new_n480_, new_n479_, new_n476_ );
and  ( new_n481_, new_n480_, new_n470_ );
not  ( new_n482_, RI2b1c4342c9a0_41 );
and  ( new_n483_, new_n138_, RI2b1c4342baa0_9 );
xor  ( new_n484_, new_n483_, new_n482_ );
and  ( new_n485_, new_n484_, new_n481_ );
not  ( new_n486_, RI2b1c4342baa0_9 );
and  ( new_n487_, RI2b1c4342bb18_10, RI2b1c4342ca18_42 );
nor  ( new_n488_, new_n423_, new_n422_ );
and  ( new_n489_, new_n468_, new_n467_ );
nor  ( new_n490_, new_n489_, new_n488_ );
nor  ( new_n491_, new_n490_, new_n487_ );
and  ( new_n492_, new_n486_, new_n482_ );
nor  ( new_n493_, new_n492_, new_n491_ );
and  ( new_n494_, RI2b1c4342baa0_9, RI2b1c4342c9a0_41 );
nor  ( new_n495_, new_n494_, new_n137_ );
and  ( new_n496_, new_n495_, new_n493_ );
or   ( new_n497_, new_n496_, new_n486_ );
or   ( new_n498_, new_n497_, new_n485_ );
xor  ( new_n499_, RI2b1c4342bb18_10, RI2b1c4342ca18_42 );
nor  ( new_n500_, new_n499_, new_n488_ );
and  ( new_n501_, new_n499_, new_n476_ );
or   ( new_n502_, new_n501_, new_n500_ );
and  ( new_n503_, new_n502_, new_n477_ );
and  ( new_n504_, new_n503_, new_n433_ );
or   ( new_n505_, new_n504_, new_n498_ );
xor  ( new_n506_, RI2b1c4342baa0_9, RI2b1c4342c9a0_41 );
nor  ( new_n507_, new_n506_, new_n491_ );
and  ( new_n508_, new_n506_, new_n481_ );
or   ( new_n509_, new_n508_, new_n507_ );
and  ( new_n510_, new_n509_, new_n483_ );
and  ( new_n511_, new_n510_, new_n503_ );
and  ( new_n512_, new_n487_, new_n138_ );
or   ( new_n513_, new_n512_, new_n479_ );
and  ( new_n514_, new_n513_, new_n476_ );
nand ( new_n515_, new_n499_, new_n138_ );
nor  ( new_n516_, new_n515_, new_n488_ );
or   ( new_n517_, new_n516_, new_n468_ );
or   ( new_n518_, new_n517_, new_n514_ );
and  ( new_n519_, new_n518_, new_n498_ );
and  ( new_n520_, new_n503_, new_n427_ );
and  ( new_n521_, new_n518_, new_n433_ );
or   ( new_n522_, new_n521_, new_n520_ );
or   ( new_n523_, new_n522_, new_n519_ );
or   ( new_n524_, new_n523_, new_n511_ );
or   ( new_n525_, new_n524_, new_n112_ );
not  ( new_n526_, RI2b1c4342d558_66 );
and  ( new_n527_, new_n518_, new_n427_ );
or   ( new_n528_, new_n527_, new_n504_ );
or   ( new_n529_, new_n528_, new_n526_ );
and  ( new_n530_, new_n529_, new_n525_ );
and  ( new_n531_, new_n530_, new_n505_ );
or   ( new_n532_, new_n518_, new_n427_ );
and  ( new_n533_, new_n532_, new_n510_ );
and  ( new_n534_, new_n518_, new_n510_ );
and  ( new_n535_, new_n503_, new_n498_ );
or   ( new_n536_, new_n535_, new_n534_ );
and  ( new_n537_, new_n536_, new_n528_ );
and  ( new_n538_, new_n537_, RI2b1c4342d5d0_67 );
and  ( new_n539_, new_n522_, RI2b1c4342d558_66 );
or   ( new_n540_, new_n539_, new_n538_ );
and  ( new_n541_, new_n540_, new_n533_ );
or   ( new_n542_, new_n541_, new_n531_ );
and  ( new_n543_, new_n542_, new_n466_ );
and  ( new_n544_, new_n464_, new_n428_ );
and  ( new_n545_, new_n457_, new_n454_ );
or   ( new_n546_, new_n545_, new_n544_ );
and  ( new_n547_, new_n540_, new_n505_ );
and  ( new_n548_, new_n533_, new_n530_ );
or   ( new_n549_, new_n548_, new_n547_ );
and  ( new_n550_, new_n549_, new_n546_ );
or   ( new_n551_, new_n550_, new_n543_ );
not  ( new_n552_, RI2b1c4342c928_40 );
not  ( new_n553_, RI2b1c4342ba28_8 );
and  ( new_n554_, new_n138_, new_n553_ );
or   ( new_n555_, new_n554_, new_n552_ );
not  ( new_n556_, new_n483_ );
and  ( new_n557_, new_n556_, new_n482_ );
and  ( new_n558_, new_n138_, new_n486_ );
or   ( new_n559_, new_n558_, new_n482_ );
and  ( new_n560_, new_n559_, new_n481_ );
or   ( new_n561_, new_n560_, new_n557_ );
and  ( new_n562_, new_n138_, RI2b1c4342ba28_8 );
not  ( new_n563_, new_n562_ );
and  ( new_n564_, new_n563_, new_n552_ );
or   ( new_n565_, new_n564_, new_n561_ );
and  ( new_n566_, new_n565_, new_n555_ );
not  ( new_n567_, RI2b1c4342c8b0_39 );
and  ( new_n568_, new_n138_, RI2b1c4342b9b0_7 );
xor  ( new_n569_, new_n568_, new_n567_ );
and  ( new_n570_, new_n569_, new_n566_ );
not  ( new_n571_, RI2b1c4342b9b0_7 );
and  ( new_n572_, RI2b1c4342ba28_8, RI2b1c4342c928_40 );
nor  ( new_n573_, new_n494_, new_n493_ );
and  ( new_n574_, new_n553_, new_n552_ );
nor  ( new_n575_, new_n574_, new_n573_ );
nor  ( new_n576_, new_n575_, new_n572_ );
and  ( new_n577_, new_n571_, new_n567_ );
nor  ( new_n578_, new_n577_, new_n576_ );
and  ( new_n579_, RI2b1c4342b9b0_7, RI2b1c4342c8b0_39 );
nor  ( new_n580_, new_n579_, new_n137_ );
and  ( new_n581_, new_n580_, new_n578_ );
or   ( new_n582_, new_n581_, new_n571_ );
or   ( new_n583_, new_n582_, new_n570_ );
xor  ( new_n584_, RI2b1c4342ba28_8, RI2b1c4342c928_40 );
nor  ( new_n585_, new_n584_, new_n573_ );
and  ( new_n586_, new_n584_, new_n561_ );
or   ( new_n587_, new_n586_, new_n585_ );
and  ( new_n588_, new_n587_, new_n562_ );
and  ( new_n589_, new_n588_, new_n510_ );
or   ( new_n590_, new_n589_, new_n583_ );
not  ( new_n591_, RI2b1c4342d6c0_69 );
xor  ( new_n592_, RI2b1c4342b9b0_7, RI2b1c4342c8b0_39 );
nor  ( new_n593_, new_n592_, new_n576_ );
and  ( new_n594_, new_n592_, new_n566_ );
or   ( new_n595_, new_n594_, new_n593_ );
and  ( new_n596_, new_n595_, new_n568_ );
and  ( new_n597_, new_n596_, new_n588_ );
and  ( new_n598_, new_n572_, new_n138_ );
or   ( new_n599_, new_n598_, new_n564_ );
and  ( new_n600_, new_n599_, new_n561_ );
nand ( new_n601_, new_n584_, new_n138_ );
nor  ( new_n602_, new_n601_, new_n573_ );
or   ( new_n603_, new_n602_, new_n553_ );
or   ( new_n604_, new_n603_, new_n600_ );
and  ( new_n605_, new_n604_, new_n583_ );
and  ( new_n606_, new_n588_, new_n498_ );
and  ( new_n607_, new_n604_, new_n510_ );
or   ( new_n608_, new_n607_, new_n606_ );
or   ( new_n609_, new_n608_, new_n605_ );
or   ( new_n610_, new_n609_, new_n597_ );
or   ( new_n611_, new_n610_, new_n591_ );
not  ( new_n612_, RI2b1c4342d648_68 );
and  ( new_n613_, new_n604_, new_n498_ );
or   ( new_n614_, new_n613_, new_n589_ );
or   ( new_n615_, new_n614_, new_n612_ );
and  ( new_n616_, new_n615_, new_n611_ );
and  ( new_n617_, new_n616_, new_n590_ );
or   ( new_n618_, new_n604_, new_n498_ );
and  ( new_n619_, new_n618_, new_n596_ );
and  ( new_n620_, new_n604_, new_n596_ );
and  ( new_n621_, new_n588_, new_n583_ );
or   ( new_n622_, new_n621_, new_n620_ );
and  ( new_n623_, new_n622_, new_n614_ );
and  ( new_n624_, new_n623_, RI2b1c4342d6c0_69 );
and  ( new_n625_, new_n608_, RI2b1c4342d648_68 );
or   ( new_n626_, new_n625_, new_n624_ );
and  ( new_n627_, new_n626_, new_n619_ );
or   ( new_n628_, new_n627_, new_n617_ );
and  ( new_n629_, new_n628_, new_n551_ );
and  ( new_n630_, new_n546_, new_n542_ );
and  ( new_n631_, new_n549_, new_n466_ );
or   ( new_n632_, new_n631_, new_n630_ );
and  ( new_n633_, new_n626_, new_n590_ );
and  ( new_n634_, new_n619_, new_n616_ );
or   ( new_n635_, new_n634_, new_n633_ );
and  ( new_n636_, new_n635_, new_n632_ );
or   ( new_n637_, new_n636_, new_n629_ );
and  ( new_n638_, RI2b1c4342b758_2, RI2b1c4342c658_34 );
and  ( new_n639_, RI2b1c4342b7d0_3, RI2b1c4342c6d0_35 );
and  ( new_n640_, RI2b1c4342b848_4, RI2b1c4342c748_36 );
not  ( new_n641_, RI2b1c4342c748_36 );
not  ( new_n642_, RI2b1c4342b848_4 );
and  ( new_n643_, new_n642_, new_n641_ );
and  ( new_n644_, RI2b1c4342b8c0_5, RI2b1c4342c7c0_37 );
and  ( new_n645_, RI2b1c4342b938_6, RI2b1c4342c838_38 );
nor  ( new_n646_, new_n579_, new_n578_ );
not  ( new_n647_, RI2b1c4342c838_38 );
not  ( new_n648_, RI2b1c4342b938_6 );
and  ( new_n649_, new_n648_, new_n647_ );
nor  ( new_n650_, new_n649_, new_n646_ );
nor  ( new_n651_, new_n650_, new_n645_ );
not  ( new_n652_, RI2b1c4342c7c0_37 );
not  ( new_n653_, RI2b1c4342b8c0_5 );
and  ( new_n654_, new_n653_, new_n652_ );
nor  ( new_n655_, new_n654_, new_n651_ );
nor  ( new_n656_, new_n655_, new_n644_ );
nor  ( new_n657_, new_n656_, new_n643_ );
nor  ( new_n658_, new_n657_, new_n640_ );
not  ( new_n659_, RI2b1c4342c6d0_35 );
not  ( new_n660_, RI2b1c4342b7d0_3 );
and  ( new_n661_, new_n660_, new_n659_ );
nor  ( new_n662_, new_n661_, new_n658_ );
nor  ( new_n663_, new_n662_, new_n639_ );
not  ( new_n664_, RI2b1c4342c658_34 );
not  ( new_n665_, RI2b1c4342b758_2 );
and  ( new_n666_, new_n665_, new_n664_ );
nor  ( new_n667_, new_n666_, new_n663_ );
nor  ( new_n668_, new_n667_, new_n638_ );
nor  ( new_n669_, new_n668_, new_n137_ );
not  ( new_n670_, RI2b1c4342c5e0_33 );
and  ( new_n671_, new_n138_, RI2b1c4342b6e0_1 );
xor  ( new_n672_, new_n671_, new_n670_ );
and  ( new_n673_, new_n672_, new_n669_ );
and  ( new_n674_, new_n138_, new_n665_ );
or   ( new_n675_, new_n674_, new_n664_ );
and  ( new_n676_, new_n138_, RI2b1c4342b7d0_3 );
not  ( new_n677_, new_n676_ );
and  ( new_n678_, new_n677_, new_n659_ );
and  ( new_n679_, new_n138_, new_n642_ );
or   ( new_n680_, new_n679_, new_n641_ );
and  ( new_n681_, new_n138_, RI2b1c4342b848_4 );
not  ( new_n682_, new_n681_ );
and  ( new_n683_, new_n682_, new_n641_ );
and  ( new_n684_, new_n138_, RI2b1c4342b8c0_5 );
not  ( new_n685_, new_n684_ );
and  ( new_n686_, new_n685_, new_n652_ );
and  ( new_n687_, new_n138_, new_n648_ );
or   ( new_n688_, new_n687_, new_n647_ );
not  ( new_n689_, new_n568_ );
and  ( new_n690_, new_n689_, new_n567_ );
and  ( new_n691_, new_n138_, new_n571_ );
or   ( new_n692_, new_n691_, new_n567_ );
and  ( new_n693_, new_n692_, new_n566_ );
or   ( new_n694_, new_n693_, new_n690_ );
and  ( new_n695_, new_n138_, RI2b1c4342b938_6 );
not  ( new_n696_, new_n695_ );
and  ( new_n697_, new_n696_, new_n647_ );
or   ( new_n698_, new_n697_, new_n694_ );
and  ( new_n699_, new_n698_, new_n688_ );
and  ( new_n700_, new_n138_, new_n653_ );
or   ( new_n701_, new_n700_, new_n652_ );
and  ( new_n702_, new_n701_, new_n699_ );
or   ( new_n703_, new_n702_, new_n686_ );
or   ( new_n704_, new_n703_, new_n683_ );
and  ( new_n705_, new_n704_, new_n680_ );
and  ( new_n706_, new_n138_, new_n660_ );
or   ( new_n707_, new_n706_, new_n659_ );
and  ( new_n708_, new_n707_, new_n705_ );
or   ( new_n709_, new_n708_, new_n678_ );
and  ( new_n710_, new_n138_, RI2b1c4342b758_2 );
not  ( new_n711_, new_n710_ );
and  ( new_n712_, new_n711_, new_n664_ );
or   ( new_n713_, new_n712_, new_n709_ );
and  ( new_n714_, new_n713_, new_n675_ );
xor  ( new_n715_, RI2b1c4342b6e0_1, new_n670_ );
not  ( new_n716_, new_n715_ );
and  ( new_n717_, new_n716_, new_n138_ );
and  ( new_n718_, new_n717_, new_n714_ );
or   ( new_n719_, new_n718_, new_n673_ );
and  ( new_n720_, new_n719_, RI2b1c4342b6e0_1 );
and  ( new_n721_, new_n720_, RI2b1c4342da08_76 );
xor  ( new_n722_, new_n684_, new_n652_ );
and  ( new_n723_, new_n722_, new_n699_ );
nor  ( new_n724_, new_n644_, new_n137_ );
and  ( new_n725_, new_n724_, new_n655_ );
or   ( new_n726_, new_n725_, new_n653_ );
or   ( new_n727_, new_n726_, new_n723_ );
xor  ( new_n728_, RI2b1c4342b938_6, RI2b1c4342c838_38 );
nor  ( new_n729_, new_n728_, new_n646_ );
and  ( new_n730_, new_n728_, new_n694_ );
or   ( new_n731_, new_n730_, new_n729_ );
and  ( new_n732_, new_n731_, new_n695_ );
and  ( new_n733_, new_n732_, new_n596_ );
or   ( new_n734_, new_n733_, new_n727_ );
xor  ( new_n735_, RI2b1c4342b8c0_5, RI2b1c4342c7c0_37 );
nor  ( new_n736_, new_n735_, new_n651_ );
and  ( new_n737_, new_n735_, new_n699_ );
or   ( new_n738_, new_n737_, new_n736_ );
and  ( new_n739_, new_n738_, new_n684_ );
and  ( new_n740_, new_n739_, new_n732_ );
and  ( new_n741_, new_n645_, new_n138_ );
or   ( new_n742_, new_n741_, new_n697_ );
and  ( new_n743_, new_n742_, new_n694_ );
nand ( new_n744_, new_n728_, new_n138_ );
nor  ( new_n745_, new_n744_, new_n646_ );
or   ( new_n746_, new_n745_, new_n648_ );
or   ( new_n747_, new_n746_, new_n743_ );
and  ( new_n748_, new_n747_, new_n727_ );
and  ( new_n749_, new_n732_, new_n583_ );
and  ( new_n750_, new_n747_, new_n596_ );
or   ( new_n751_, new_n750_, new_n749_ );
or   ( new_n752_, new_n751_, new_n748_ );
or   ( new_n753_, new_n752_, new_n740_ );
or   ( new_n754_, new_n753_, new_n110_ );
not  ( new_n755_, RI2b1c4342d738_70 );
and  ( new_n756_, new_n747_, new_n583_ );
or   ( new_n757_, new_n756_, new_n733_ );
or   ( new_n758_, new_n757_, new_n755_ );
and  ( new_n759_, new_n758_, new_n754_ );
and  ( new_n760_, new_n759_, new_n734_ );
or   ( new_n761_, new_n747_, new_n583_ );
and  ( new_n762_, new_n761_, new_n739_ );
and  ( new_n763_, new_n747_, new_n739_ );
and  ( new_n764_, new_n732_, new_n727_ );
or   ( new_n765_, new_n764_, new_n763_ );
and  ( new_n766_, new_n765_, new_n757_ );
and  ( new_n767_, new_n766_, RI2b1c4342d7b0_71 );
and  ( new_n768_, new_n751_, RI2b1c4342d738_70 );
or   ( new_n769_, new_n768_, new_n767_ );
and  ( new_n770_, new_n769_, new_n762_ );
or   ( new_n771_, new_n770_, new_n760_ );
and  ( new_n772_, new_n639_, new_n138_ );
or   ( new_n773_, new_n772_, new_n678_ );
and  ( new_n774_, new_n773_, new_n705_ );
nor  ( new_n775_, new_n639_, new_n137_ );
and  ( new_n776_, new_n775_, new_n662_ );
or   ( new_n777_, new_n776_, new_n660_ );
or   ( new_n778_, new_n777_, new_n774_ );
xor  ( new_n779_, RI2b1c4342b848_4, RI2b1c4342c748_36 );
nor  ( new_n780_, new_n779_, new_n656_ );
and  ( new_n781_, new_n779_, new_n703_ );
or   ( new_n782_, new_n781_, new_n780_ );
and  ( new_n783_, new_n782_, new_n681_ );
and  ( new_n784_, new_n783_, new_n739_ );
or   ( new_n785_, new_n784_, new_n778_ );
xor  ( new_n786_, RI2b1c4342b7d0_3, RI2b1c4342c6d0_35 );
nor  ( new_n787_, new_n786_, new_n658_ );
and  ( new_n788_, new_n786_, new_n705_ );
or   ( new_n789_, new_n788_, new_n787_ );
and  ( new_n790_, new_n789_, new_n676_ );
and  ( new_n791_, new_n790_, new_n783_ );
and  ( new_n792_, new_n640_, new_n138_ );
or   ( new_n793_, new_n792_, new_n683_ );
and  ( new_n794_, new_n793_, new_n703_ );
nand ( new_n795_, new_n779_, new_n138_ );
nor  ( new_n796_, new_n795_, new_n656_ );
or   ( new_n797_, new_n796_, new_n642_ );
or   ( new_n798_, new_n797_, new_n794_ );
and  ( new_n799_, new_n798_, new_n778_ );
and  ( new_n800_, new_n783_, new_n727_ );
and  ( new_n801_, new_n798_, new_n739_ );
or   ( new_n802_, new_n801_, new_n800_ );
or   ( new_n803_, new_n802_, new_n799_ );
or   ( new_n804_, new_n803_, new_n791_ );
or   ( new_n805_, new_n804_, new_n105_ );
not  ( new_n806_, RI2b1c4342d828_72 );
and  ( new_n807_, new_n798_, new_n727_ );
or   ( new_n808_, new_n807_, new_n784_ );
or   ( new_n809_, new_n808_, new_n806_ );
and  ( new_n810_, new_n809_, new_n805_ );
and  ( new_n811_, new_n810_, new_n785_ );
or   ( new_n812_, new_n798_, new_n727_ );
and  ( new_n813_, new_n812_, new_n790_ );
and  ( new_n814_, new_n798_, new_n790_ );
and  ( new_n815_, new_n783_, new_n778_ );
or   ( new_n816_, new_n815_, new_n814_ );
and  ( new_n817_, new_n816_, new_n808_ );
and  ( new_n818_, new_n817_, RI2b1c4342d8a0_73 );
and  ( new_n819_, new_n802_, RI2b1c4342d828_72 );
or   ( new_n820_, new_n819_, new_n818_ );
and  ( new_n821_, new_n820_, new_n813_ );
or   ( new_n822_, new_n821_, new_n811_ );
and  ( new_n823_, new_n822_, new_n771_ );
and  ( new_n824_, new_n769_, new_n734_ );
and  ( new_n825_, new_n762_, new_n759_ );
or   ( new_n826_, new_n825_, new_n824_ );
and  ( new_n827_, new_n820_, new_n785_ );
and  ( new_n828_, new_n813_, new_n810_ );
or   ( new_n829_, new_n828_, new_n827_ );
and  ( new_n830_, new_n829_, new_n826_ );
or   ( new_n831_, new_n830_, new_n823_ );
xor  ( new_n832_, RI2b1c4342b758_2, RI2b1c4342c658_34 );
nor  ( new_n833_, new_n832_, new_n663_ );
and  ( new_n834_, new_n832_, new_n709_ );
or   ( new_n835_, new_n834_, new_n833_ );
and  ( new_n836_, new_n835_, new_n710_ );
and  ( new_n837_, new_n836_, new_n790_ );
and  ( new_n838_, new_n714_, new_n672_ );
nand ( new_n839_, new_n716_, new_n669_ );
nand ( new_n840_, new_n839_, RI2b1c4342b6e0_1 );
or   ( new_n841_, new_n840_, new_n838_ );
or   ( new_n842_, new_n841_, new_n837_ );
not  ( new_n843_, RI2b1c4342d990_75 );
and  ( new_n844_, new_n836_, new_n720_ );
and  ( new_n845_, new_n638_, new_n138_ );
or   ( new_n846_, new_n845_, new_n712_ );
and  ( new_n847_, new_n846_, new_n709_ );
nand ( new_n848_, new_n832_, new_n138_ );
nor  ( new_n849_, new_n848_, new_n663_ );
or   ( new_n850_, new_n849_, new_n665_ );
or   ( new_n851_, new_n850_, new_n847_ );
and  ( new_n852_, new_n851_, new_n841_ );
and  ( new_n853_, new_n836_, new_n778_ );
and  ( new_n854_, new_n851_, new_n790_ );
or   ( new_n855_, new_n854_, new_n853_ );
or   ( new_n856_, new_n855_, new_n852_ );
or   ( new_n857_, new_n856_, new_n844_ );
or   ( new_n858_, new_n857_, new_n843_ );
not  ( new_n859_, RI2b1c4342d918_74 );
and  ( new_n860_, new_n851_, new_n778_ );
or   ( new_n861_, new_n860_, new_n837_ );
or   ( new_n862_, new_n861_, new_n859_ );
and  ( new_n863_, new_n862_, new_n858_ );
and  ( new_n864_, new_n863_, new_n842_ );
or   ( new_n865_, new_n851_, new_n778_ );
and  ( new_n866_, new_n865_, new_n720_ );
and  ( new_n867_, new_n851_, new_n720_ );
and  ( new_n868_, new_n841_, new_n836_ );
or   ( new_n869_, new_n868_, new_n867_ );
and  ( new_n870_, new_n869_, new_n861_ );
and  ( new_n871_, new_n870_, RI2b1c4342d990_75 );
and  ( new_n872_, new_n855_, RI2b1c4342d918_74 );
or   ( new_n873_, new_n872_, new_n871_ );
and  ( new_n874_, new_n873_, new_n866_ );
or   ( new_n875_, new_n874_, new_n864_ );
and  ( new_n876_, new_n875_, new_n831_ );
and  ( new_n877_, new_n826_, new_n822_ );
and  ( new_n878_, new_n829_, new_n771_ );
or   ( new_n879_, new_n878_, new_n877_ );
and  ( new_n880_, new_n873_, new_n842_ );
and  ( new_n881_, new_n866_, new_n863_ );
or   ( new_n882_, new_n881_, new_n880_ );
and  ( new_n883_, new_n882_, new_n879_ );
or   ( new_n884_, new_n883_, new_n876_ );
and  ( new_n885_, new_n884_, new_n721_ );
not  ( new_n886_, RI2b1c4342da08_76 );
or   ( new_n887_, new_n841_, new_n886_ );
and  ( new_n888_, new_n879_, new_n875_ );
and  ( new_n889_, new_n882_, new_n831_ );
or   ( new_n890_, new_n889_, new_n888_ );
and  ( new_n891_, new_n890_, new_n887_ );
or   ( new_n892_, new_n891_, new_n885_ );
and  ( new_n893_, new_n892_, new_n637_ );
and  ( new_n894_, new_n632_, new_n628_ );
and  ( new_n895_, new_n635_, new_n551_ );
or   ( new_n896_, new_n895_, new_n894_ );
and  ( new_n897_, new_n887_, new_n884_ );
and  ( new_n898_, new_n890_, new_n721_ );
or   ( new_n899_, new_n898_, new_n897_ );
and  ( new_n900_, new_n899_, new_n896_ );
or   ( new_n901_, new_n900_, new_n893_ );
xor  ( new_n902_, RI2b1c4342bd70_15, RI2b1c4342cc70_47 );
nor  ( new_n903_, new_n902_, new_n250_ );
and  ( new_n904_, new_n902_, new_n375_ );
or   ( new_n905_, new_n904_, new_n903_ );
and  ( new_n906_, new_n905_, new_n265_ );
xor  ( new_n907_, RI2b1c4342bcf8_14, RI2b1c4342cbf8_46 );
nor  ( new_n908_, new_n907_, new_n255_ );
and  ( new_n909_, new_n907_, new_n379_ );
or   ( new_n910_, new_n909_, new_n908_ );
and  ( new_n911_, new_n910_, new_n262_ );
and  ( new_n912_, new_n911_, new_n906_ );
or   ( new_n913_, new_n912_, new_n448_ );
and  ( new_n914_, new_n911_, new_n384_ );
and  ( new_n915_, new_n140_, new_n138_ );
or   ( new_n916_, new_n915_, new_n264_ );
and  ( new_n917_, new_n916_, new_n379_ );
nand ( new_n918_, new_n907_, new_n138_ );
nor  ( new_n919_, new_n918_, new_n255_ );
or   ( new_n920_, new_n919_, new_n142_ );
or   ( new_n921_, new_n920_, new_n917_ );
and  ( new_n922_, new_n921_, new_n448_ );
and  ( new_n923_, new_n144_, new_n138_ );
or   ( new_n924_, new_n923_, new_n267_ );
and  ( new_n925_, new_n924_, new_n375_ );
nor  ( new_n926_, new_n144_, new_n137_ );
and  ( new_n927_, new_n926_, new_n254_ );
or   ( new_n928_, new_n927_, new_n252_ );
or   ( new_n929_, new_n928_, new_n925_ );
and  ( new_n930_, new_n929_, new_n911_ );
and  ( new_n931_, new_n921_, new_n906_ );
or   ( new_n932_, new_n931_, new_n930_ );
or   ( new_n933_, new_n932_, new_n922_ );
or   ( new_n934_, new_n933_, new_n914_ );
or   ( new_n935_, new_n934_, new_n99_ );
and  ( new_n936_, new_n935_, new_n913_ );
or   ( new_n937_, new_n929_, new_n921_ );
and  ( new_n938_, new_n937_, new_n384_ );
and  ( new_n939_, new_n929_, new_n921_ );
or   ( new_n940_, new_n939_, new_n912_ );
and  ( new_n941_, new_n921_, new_n384_ );
and  ( new_n942_, new_n911_, new_n448_ );
or   ( new_n943_, new_n942_, new_n941_ );
and  ( new_n944_, new_n943_, new_n940_ );
and  ( new_n945_, new_n944_, RI2b1c4342d4e0_65 );
and  ( new_n946_, new_n945_, new_n938_ );
or   ( new_n947_, new_n946_, new_n936_ );
or   ( new_n948_, new_n453_, new_n112_ );
or   ( new_n949_, new_n459_, new_n526_ );
and  ( new_n950_, new_n949_, new_n948_ );
and  ( new_n951_, new_n950_, new_n428_ );
and  ( new_n952_, new_n463_, RI2b1c4342d5d0_67 );
and  ( new_n953_, new_n451_, RI2b1c4342d558_66 );
or   ( new_n954_, new_n953_, new_n952_ );
and  ( new_n955_, new_n954_, new_n457_ );
or   ( new_n956_, new_n955_, new_n951_ );
and  ( new_n957_, new_n956_, new_n947_ );
or   ( new_n958_, new_n524_, new_n591_ );
or   ( new_n959_, new_n528_, new_n612_ );
and  ( new_n960_, new_n959_, new_n958_ );
and  ( new_n961_, new_n960_, new_n505_ );
and  ( new_n962_, new_n537_, RI2b1c4342d6c0_69 );
and  ( new_n963_, new_n522_, RI2b1c4342d648_68 );
or   ( new_n964_, new_n963_, new_n962_ );
and  ( new_n965_, new_n964_, new_n533_ );
or   ( new_n966_, new_n965_, new_n961_ );
or   ( new_n967_, new_n956_, new_n947_ );
and  ( new_n968_, new_n967_, new_n966_ );
or   ( new_n969_, new_n968_, new_n957_ );
or   ( new_n970_, new_n610_, new_n110_ );
or   ( new_n971_, new_n614_, new_n755_ );
and  ( new_n972_, new_n971_, new_n970_ );
and  ( new_n973_, new_n972_, new_n590_ );
and  ( new_n974_, new_n623_, RI2b1c4342d7b0_71 );
and  ( new_n975_, new_n608_, RI2b1c4342d738_70 );
or   ( new_n976_, new_n975_, new_n974_ );
and  ( new_n977_, new_n976_, new_n619_ );
or   ( new_n978_, new_n977_, new_n973_ );
or   ( new_n979_, new_n753_, new_n105_ );
or   ( new_n980_, new_n757_, new_n806_ );
and  ( new_n981_, new_n980_, new_n979_ );
and  ( new_n982_, new_n981_, new_n734_ );
and  ( new_n983_, new_n766_, RI2b1c4342d8a0_73 );
and  ( new_n984_, new_n751_, RI2b1c4342d828_72 );
or   ( new_n985_, new_n984_, new_n983_ );
and  ( new_n986_, new_n985_, new_n762_ );
or   ( new_n987_, new_n986_, new_n982_ );
and  ( new_n988_, new_n987_, new_n978_ );
or   ( new_n989_, new_n804_, new_n843_ );
or   ( new_n990_, new_n808_, new_n859_ );
and  ( new_n991_, new_n990_, new_n989_ );
and  ( new_n992_, new_n991_, new_n785_ );
and  ( new_n993_, new_n817_, RI2b1c4342d990_75 );
and  ( new_n994_, new_n802_, RI2b1c4342d918_74 );
or   ( new_n995_, new_n994_, new_n993_ );
and  ( new_n996_, new_n995_, new_n813_ );
or   ( new_n997_, new_n996_, new_n992_ );
or   ( new_n998_, new_n987_, new_n978_ );
and  ( new_n999_, new_n998_, new_n997_ );
or   ( new_n1000_, new_n999_, new_n988_ );
and  ( new_n1001_, new_n1000_, new_n969_ );
not  ( new_n1002_, RI2b1c4342daf8_78 );
or   ( new_n1003_, new_n841_, new_n1002_ );
not  ( new_n1004_, RI2b1c4342da80_77 );
or   ( new_n1005_, new_n857_, new_n1004_ );
or   ( new_n1006_, new_n861_, new_n886_ );
and  ( new_n1007_, new_n1006_, new_n1005_ );
and  ( new_n1008_, new_n1007_, new_n842_ );
and  ( new_n1009_, new_n870_, RI2b1c4342da80_77 );
and  ( new_n1010_, new_n855_, RI2b1c4342da08_76 );
or   ( new_n1011_, new_n1010_, new_n1009_ );
and  ( new_n1012_, new_n1011_, new_n866_ );
or   ( new_n1013_, new_n1012_, new_n1008_ );
and  ( new_n1014_, new_n1013_, new_n1003_ );
or   ( new_n1015_, new_n1000_, new_n969_ );
and  ( new_n1016_, new_n1015_, new_n1014_ );
or   ( new_n1017_, new_n1016_, new_n1001_ );
and  ( new_n1018_, new_n870_, RI2b1c4342da08_76 );
and  ( new_n1019_, new_n855_, RI2b1c4342d990_75 );
or   ( new_n1020_, new_n1019_, new_n1018_ );
and  ( new_n1021_, new_n1020_, new_n842_ );
or   ( new_n1022_, new_n857_, new_n886_ );
or   ( new_n1023_, new_n861_, new_n843_ );
and  ( new_n1024_, new_n1023_, new_n1022_ );
and  ( new_n1025_, new_n1024_, new_n866_ );
or   ( new_n1026_, new_n1025_, new_n1021_ );
and  ( new_n1027_, new_n720_, RI2b1c4342da80_77 );
and  ( new_n1028_, new_n1027_, new_n1026_ );
and  ( new_n1029_, new_n1024_, new_n842_ );
and  ( new_n1030_, new_n1020_, new_n866_ );
or   ( new_n1031_, new_n1030_, new_n1029_ );
or   ( new_n1032_, new_n841_, new_n1004_ );
and  ( new_n1033_, new_n1032_, new_n1031_ );
or   ( new_n1034_, new_n1033_, new_n1028_ );
or   ( new_n1035_, new_n804_, new_n859_ );
or   ( new_n1036_, new_n808_, new_n105_ );
and  ( new_n1037_, new_n1036_, new_n1035_ );
and  ( new_n1038_, new_n1037_, new_n785_ );
and  ( new_n1039_, new_n817_, RI2b1c4342d918_74 );
and  ( new_n1040_, new_n802_, RI2b1c4342d8a0_73 );
or   ( new_n1041_, new_n1040_, new_n1039_ );
and  ( new_n1042_, new_n1041_, new_n813_ );
or   ( new_n1043_, new_n1042_, new_n1038_ );
or   ( new_n1044_, new_n610_, new_n755_ );
or   ( new_n1045_, new_n614_, new_n591_ );
and  ( new_n1046_, new_n1045_, new_n1044_ );
and  ( new_n1047_, new_n1046_, new_n590_ );
and  ( new_n1048_, new_n623_, RI2b1c4342d738_70 );
and  ( new_n1049_, new_n608_, RI2b1c4342d6c0_69 );
or   ( new_n1050_, new_n1049_, new_n1048_ );
and  ( new_n1051_, new_n1050_, new_n619_ );
or   ( new_n1052_, new_n1051_, new_n1047_ );
or   ( new_n1053_, new_n753_, new_n806_ );
or   ( new_n1054_, new_n757_, new_n110_ );
and  ( new_n1055_, new_n1054_, new_n1053_ );
and  ( new_n1056_, new_n1055_, new_n734_ );
and  ( new_n1057_, new_n766_, RI2b1c4342d828_72 );
and  ( new_n1058_, new_n751_, RI2b1c4342d7b0_71 );
or   ( new_n1059_, new_n1058_, new_n1057_ );
and  ( new_n1060_, new_n1059_, new_n762_ );
or   ( new_n1061_, new_n1060_, new_n1056_ );
and  ( new_n1062_, new_n1061_, new_n1052_ );
and  ( new_n1063_, new_n1050_, new_n590_ );
and  ( new_n1064_, new_n1046_, new_n619_ );
or   ( new_n1065_, new_n1064_, new_n1063_ );
and  ( new_n1066_, new_n1059_, new_n734_ );
and  ( new_n1067_, new_n1055_, new_n762_ );
or   ( new_n1068_, new_n1067_, new_n1066_ );
and  ( new_n1069_, new_n1068_, new_n1065_ );
or   ( new_n1070_, new_n1069_, new_n1062_ );
and  ( new_n1071_, new_n1070_, new_n1043_ );
and  ( new_n1072_, new_n1041_, new_n785_ );
and  ( new_n1073_, new_n1037_, new_n813_ );
or   ( new_n1074_, new_n1073_, new_n1072_ );
and  ( new_n1075_, new_n1065_, new_n1061_ );
and  ( new_n1076_, new_n1068_, new_n1052_ );
or   ( new_n1077_, new_n1076_, new_n1075_ );
and  ( new_n1078_, new_n1077_, new_n1074_ );
or   ( new_n1079_, new_n1078_, new_n1071_ );
and  ( new_n1080_, new_n1079_, new_n1034_ );
or   ( new_n1081_, new_n1079_, new_n1034_ );
or   ( new_n1082_, new_n524_, new_n612_ );
or   ( new_n1083_, new_n528_, new_n112_ );
and  ( new_n1084_, new_n1083_, new_n1082_ );
and  ( new_n1085_, new_n1084_, new_n505_ );
and  ( new_n1086_, new_n537_, RI2b1c4342d648_68 );
and  ( new_n1087_, new_n522_, RI2b1c4342d5d0_67 );
or   ( new_n1088_, new_n1087_, new_n1086_ );
and  ( new_n1089_, new_n1088_, new_n533_ );
or   ( new_n1090_, new_n1089_, new_n1085_ );
or   ( new_n1091_, new_n453_, new_n526_ );
or   ( new_n1092_, new_n459_, new_n99_ );
and  ( new_n1093_, new_n1092_, new_n1091_ );
and  ( new_n1094_, new_n1093_, new_n428_ );
and  ( new_n1095_, new_n463_, RI2b1c4342d558_66 );
and  ( new_n1096_, new_n451_, RI2b1c4342d4e0_65 );
or   ( new_n1097_, new_n1096_, new_n1095_ );
and  ( new_n1098_, new_n1097_, new_n457_ );
or   ( new_n1099_, new_n1098_, new_n1094_ );
and  ( new_n1100_, new_n1099_, new_n938_ );
and  ( new_n1101_, new_n1097_, new_n428_ );
and  ( new_n1102_, new_n1093_, new_n457_ );
or   ( new_n1103_, new_n1102_, new_n1101_ );
and  ( new_n1104_, new_n1103_, new_n913_ );
or   ( new_n1105_, new_n1104_, new_n1100_ );
and  ( new_n1106_, new_n1105_, new_n1090_ );
and  ( new_n1107_, new_n1088_, new_n505_ );
and  ( new_n1108_, new_n1084_, new_n533_ );
or   ( new_n1109_, new_n1108_, new_n1107_ );
and  ( new_n1110_, new_n1099_, new_n913_ );
and  ( new_n1111_, new_n1103_, new_n938_ );
or   ( new_n1112_, new_n1111_, new_n1110_ );
and  ( new_n1113_, new_n1112_, new_n1109_ );
or   ( new_n1114_, new_n1113_, new_n1106_ );
and  ( new_n1115_, new_n1114_, new_n1081_ );
or   ( new_n1116_, new_n1115_, new_n1080_ );
and  ( new_n1117_, new_n1116_, new_n1017_ );
and  ( new_n1118_, new_n945_, new_n913_ );
and  ( new_n1119_, new_n938_, new_n935_ );
or   ( new_n1120_, new_n1119_, new_n1118_ );
and  ( new_n1121_, new_n954_, new_n428_ );
and  ( new_n1122_, new_n950_, new_n457_ );
or   ( new_n1123_, new_n1122_, new_n1121_ );
and  ( new_n1124_, new_n1123_, new_n1120_ );
and  ( new_n1125_, new_n964_, new_n505_ );
and  ( new_n1126_, new_n960_, new_n533_ );
or   ( new_n1127_, new_n1126_, new_n1125_ );
or   ( new_n1128_, new_n1123_, new_n1120_ );
and  ( new_n1129_, new_n1128_, new_n1127_ );
or   ( new_n1130_, new_n1129_, new_n1124_ );
and  ( new_n1131_, new_n976_, new_n590_ );
and  ( new_n1132_, new_n972_, new_n619_ );
or   ( new_n1133_, new_n1132_, new_n1131_ );
and  ( new_n1134_, new_n985_, new_n734_ );
and  ( new_n1135_, new_n981_, new_n762_ );
or   ( new_n1136_, new_n1135_, new_n1134_ );
and  ( new_n1137_, new_n1136_, new_n1133_ );
and  ( new_n1138_, new_n995_, new_n785_ );
and  ( new_n1139_, new_n991_, new_n813_ );
or   ( new_n1140_, new_n1139_, new_n1138_ );
or   ( new_n1141_, new_n1136_, new_n1133_ );
and  ( new_n1142_, new_n1141_, new_n1140_ );
or   ( new_n1143_, new_n1142_, new_n1137_ );
and  ( new_n1144_, new_n1143_, new_n1130_ );
or   ( new_n1145_, new_n1143_, new_n1130_ );
and  ( new_n1146_, new_n1011_, new_n842_ );
and  ( new_n1147_, new_n1007_, new_n866_ );
or   ( new_n1148_, new_n1147_, new_n1146_ );
and  ( new_n1149_, new_n720_, RI2b1c4342daf8_78 );
or   ( new_n1150_, new_n1149_, new_n1148_ );
and  ( new_n1151_, new_n1150_, new_n1145_ );
or   ( new_n1152_, new_n1151_, new_n1144_ );
and  ( new_n1153_, new_n1032_, new_n1026_ );
and  ( new_n1154_, new_n1031_, new_n1027_ );
or   ( new_n1155_, new_n1154_, new_n1153_ );
and  ( new_n1156_, new_n1077_, new_n1043_ );
and  ( new_n1157_, new_n1074_, new_n1070_ );
or   ( new_n1158_, new_n1157_, new_n1156_ );
and  ( new_n1159_, new_n1158_, new_n1155_ );
or   ( new_n1160_, new_n1158_, new_n1155_ );
and  ( new_n1161_, new_n1112_, new_n1090_ );
and  ( new_n1162_, new_n1109_, new_n1105_ );
or   ( new_n1163_, new_n1162_, new_n1161_ );
and  ( new_n1164_, new_n1163_, new_n1160_ );
or   ( new_n1165_, new_n1164_, new_n1159_ );
and  ( new_n1166_, new_n1165_, new_n1152_ );
or   ( new_n1167_, new_n1166_, new_n1117_ );
and  ( new_n1168_, new_n1167_, new_n901_ );
and  ( new_n1169_, new_n899_, new_n637_ );
and  ( new_n1170_, new_n896_, new_n892_ );
or   ( new_n1171_, new_n1170_, new_n1169_ );
and  ( new_n1172_, new_n1152_, new_n1116_ );
and  ( new_n1173_, new_n1165_, new_n1017_ );
or   ( new_n1174_, new_n1173_, new_n1172_ );
and  ( new_n1175_, new_n1174_, new_n1171_ );
or   ( new_n1176_, new_n1175_, new_n1168_ );
or   ( new_n1177_, new_n1032_, new_n1031_ );
or   ( new_n1178_, new_n1061_, new_n1052_ );
and  ( new_n1179_, new_n1178_, new_n1043_ );
or   ( new_n1180_, new_n1179_, new_n1062_ );
or   ( new_n1181_, new_n1099_, new_n938_ );
and  ( new_n1182_, new_n1181_, new_n1090_ );
or   ( new_n1183_, new_n1182_, new_n1100_ );
and  ( new_n1184_, new_n1183_, new_n1180_ );
or   ( new_n1185_, new_n1103_, new_n913_ );
and  ( new_n1186_, new_n1185_, new_n1109_ );
or   ( new_n1187_, new_n1186_, new_n1104_ );
or   ( new_n1188_, new_n1068_, new_n1065_ );
and  ( new_n1189_, new_n1188_, new_n1074_ );
or   ( new_n1190_, new_n1189_, new_n1069_ );
and  ( new_n1191_, new_n1190_, new_n1187_ );
or   ( new_n1192_, new_n1191_, new_n1184_ );
and  ( new_n1193_, new_n1192_, new_n1177_ );
and  ( new_n1194_, new_n1187_, new_n1180_ );
and  ( new_n1195_, new_n1190_, new_n1183_ );
or   ( new_n1196_, new_n1195_, new_n1194_ );
and  ( new_n1197_, new_n1196_, new_n1028_ );
or   ( new_n1198_, new_n1197_, new_n1193_ );
and  ( new_n1199_, new_n1148_, new_n1003_ );
and  ( new_n1200_, new_n1149_, new_n1013_ );
or   ( new_n1201_, new_n1200_, new_n1199_ );
or   ( new_n1202_, new_n1137_, new_n988_ );
and  ( new_n1203_, new_n1202_, new_n997_ );
and  ( new_n1204_, new_n1133_, new_n987_ );
and  ( new_n1205_, new_n1136_, new_n978_ );
or   ( new_n1206_, new_n1205_, new_n1204_ );
and  ( new_n1207_, new_n1206_, new_n1140_ );
or   ( new_n1208_, new_n1207_, new_n1203_ );
and  ( new_n1209_, new_n1208_, new_n1201_ );
or   ( new_n1210_, new_n1124_, new_n957_ );
and  ( new_n1211_, new_n1210_, new_n966_ );
and  ( new_n1212_, new_n1120_, new_n956_ );
and  ( new_n1213_, new_n1123_, new_n947_ );
or   ( new_n1214_, new_n1213_, new_n1212_ );
and  ( new_n1215_, new_n1214_, new_n1127_ );
or   ( new_n1216_, new_n1215_, new_n1211_ );
or   ( new_n1217_, new_n1208_, new_n1201_ );
and  ( new_n1218_, new_n1217_, new_n1216_ );
or   ( new_n1219_, new_n1218_, new_n1209_ );
or   ( new_n1220_, new_n524_, new_n755_ );
or   ( new_n1221_, new_n528_, new_n591_ );
and  ( new_n1222_, new_n1221_, new_n1220_ );
and  ( new_n1223_, new_n1222_, new_n505_ );
and  ( new_n1224_, new_n537_, RI2b1c4342d738_70 );
and  ( new_n1225_, new_n522_, RI2b1c4342d6c0_69 );
or   ( new_n1226_, new_n1225_, new_n1224_ );
and  ( new_n1227_, new_n1226_, new_n533_ );
or   ( new_n1228_, new_n1227_, new_n1223_ );
or   ( new_n1229_, new_n610_, new_n806_ );
or   ( new_n1230_, new_n614_, new_n110_ );
and  ( new_n1231_, new_n1230_, new_n1229_ );
and  ( new_n1232_, new_n1231_, new_n590_ );
and  ( new_n1233_, new_n623_, RI2b1c4342d828_72 );
and  ( new_n1234_, new_n608_, RI2b1c4342d7b0_71 );
or   ( new_n1235_, new_n1234_, new_n1233_ );
and  ( new_n1236_, new_n1235_, new_n619_ );
or   ( new_n1237_, new_n1236_, new_n1232_ );
and  ( new_n1238_, new_n1237_, new_n1228_ );
or   ( new_n1239_, new_n753_, new_n859_ );
or   ( new_n1240_, new_n757_, new_n105_ );
and  ( new_n1241_, new_n1240_, new_n1239_ );
and  ( new_n1242_, new_n1241_, new_n734_ );
and  ( new_n1243_, new_n766_, RI2b1c4342d918_74 );
and  ( new_n1244_, new_n751_, RI2b1c4342d8a0_73 );
or   ( new_n1245_, new_n1244_, new_n1243_ );
and  ( new_n1246_, new_n1245_, new_n762_ );
or   ( new_n1247_, new_n1246_, new_n1242_ );
or   ( new_n1248_, new_n1237_, new_n1228_ );
and  ( new_n1249_, new_n1248_, new_n1247_ );
or   ( new_n1250_, new_n1249_, new_n1238_ );
and  ( new_n1251_, new_n149_, new_n138_ );
or   ( new_n1252_, new_n1251_, new_n275_ );
and  ( new_n1253_, new_n1252_, new_n369_ );
nor  ( new_n1254_, new_n149_, new_n137_ );
and  ( new_n1255_, new_n1254_, new_n247_ );
or   ( new_n1256_, new_n1255_, new_n151_ );
or   ( new_n1257_, new_n1256_, new_n1253_ );
and  ( new_n1258_, new_n145_, new_n138_ );
or   ( new_n1259_, new_n1258_, new_n272_ );
and  ( new_n1260_, new_n1259_, new_n373_ );
xor  ( new_n1261_, RI2b1c4342bde8_16, RI2b1c4342cce8_48 );
nand ( new_n1262_, new_n1261_, new_n138_ );
nor  ( new_n1263_, new_n1262_, new_n248_ );
or   ( new_n1264_, new_n1263_, new_n147_ );
or   ( new_n1265_, new_n1264_, new_n1260_ );
or   ( new_n1266_, new_n1265_, new_n1257_ );
and  ( new_n1267_, new_n1266_, new_n906_ );
or   ( new_n1268_, new_n934_, new_n526_ );
or   ( new_n1269_, new_n940_, new_n99_ );
and  ( new_n1270_, new_n1269_, new_n1268_ );
and  ( new_n1271_, new_n1270_, new_n913_ );
and  ( new_n1272_, new_n944_, RI2b1c4342d558_66 );
and  ( new_n1273_, new_n932_, RI2b1c4342d4e0_65 );
or   ( new_n1274_, new_n1273_, new_n1272_ );
and  ( new_n1275_, new_n1274_, new_n938_ );
or   ( new_n1276_, new_n1275_, new_n1271_ );
and  ( new_n1277_, new_n1276_, new_n1267_ );
or   ( new_n1278_, new_n453_, new_n612_ );
or   ( new_n1279_, new_n459_, new_n112_ );
and  ( new_n1280_, new_n1279_, new_n1278_ );
and  ( new_n1281_, new_n1280_, new_n428_ );
and  ( new_n1282_, new_n463_, RI2b1c4342d648_68 );
and  ( new_n1283_, new_n451_, RI2b1c4342d5d0_67 );
or   ( new_n1284_, new_n1283_, new_n1282_ );
and  ( new_n1285_, new_n1284_, new_n457_ );
or   ( new_n1286_, new_n1285_, new_n1281_ );
or   ( new_n1287_, new_n1276_, new_n1267_ );
and  ( new_n1288_, new_n1287_, new_n1286_ );
or   ( new_n1289_, new_n1288_, new_n1277_ );
and  ( new_n1290_, new_n1289_, new_n1250_ );
or   ( new_n1291_, new_n804_, new_n886_ );
or   ( new_n1292_, new_n808_, new_n843_ );
and  ( new_n1293_, new_n1292_, new_n1291_ );
and  ( new_n1294_, new_n1293_, new_n785_ );
and  ( new_n1295_, new_n817_, RI2b1c4342da08_76 );
and  ( new_n1296_, new_n802_, RI2b1c4342d990_75 );
or   ( new_n1297_, new_n1296_, new_n1295_ );
and  ( new_n1298_, new_n1297_, new_n813_ );
or   ( new_n1299_, new_n1298_, new_n1294_ );
or   ( new_n1300_, new_n857_, new_n1002_ );
or   ( new_n1301_, new_n861_, new_n1004_ );
and  ( new_n1302_, new_n1301_, new_n1300_ );
and  ( new_n1303_, new_n1302_, new_n842_ );
and  ( new_n1304_, new_n870_, RI2b1c4342daf8_78 );
and  ( new_n1305_, new_n855_, RI2b1c4342da80_77 );
or   ( new_n1306_, new_n1305_, new_n1304_ );
and  ( new_n1307_, new_n1306_, new_n866_ );
or   ( new_n1308_, new_n1307_, new_n1303_ );
and  ( new_n1309_, new_n1308_, new_n1299_ );
not  ( new_n1310_, RI2b1c4342db70_79 );
or   ( new_n1311_, new_n841_, new_n1310_ );
or   ( new_n1312_, new_n1308_, new_n1299_ );
and  ( new_n1313_, new_n1312_, new_n1311_ );
or   ( new_n1314_, new_n1313_, new_n1309_ );
or   ( new_n1315_, new_n1289_, new_n1250_ );
and  ( new_n1316_, new_n1315_, new_n1314_ );
or   ( new_n1317_, new_n1316_, new_n1290_ );
and  ( new_n1318_, new_n1317_, new_n1219_ );
or   ( new_n1319_, new_n1317_, new_n1219_ );
or   ( new_n1320_, new_n1159_, new_n1080_ );
and  ( new_n1321_, new_n1320_, new_n1114_ );
and  ( new_n1322_, new_n1155_, new_n1079_ );
and  ( new_n1323_, new_n1158_, new_n1034_ );
or   ( new_n1324_, new_n1323_, new_n1322_ );
and  ( new_n1325_, new_n1324_, new_n1163_ );
or   ( new_n1326_, new_n1325_, new_n1321_ );
and  ( new_n1327_, new_n1326_, new_n1319_ );
or   ( new_n1328_, new_n1327_, new_n1318_ );
and  ( new_n1329_, new_n1328_, new_n1198_ );
and  ( new_n1330_, new_n1196_, new_n1177_ );
and  ( new_n1331_, new_n1192_, new_n1028_ );
or   ( new_n1332_, new_n1331_, new_n1330_ );
and  ( new_n1333_, new_n1149_, new_n1148_ );
or   ( new_n1334_, new_n1333_, new_n1014_ );
and  ( new_n1335_, new_n1206_, new_n997_ );
and  ( new_n1336_, new_n1202_, new_n1140_ );
or   ( new_n1337_, new_n1336_, new_n1335_ );
and  ( new_n1338_, new_n1337_, new_n1334_ );
and  ( new_n1339_, new_n1214_, new_n966_ );
and  ( new_n1340_, new_n1210_, new_n1127_ );
or   ( new_n1341_, new_n1340_, new_n1339_ );
or   ( new_n1342_, new_n1337_, new_n1334_ );
and  ( new_n1343_, new_n1342_, new_n1341_ );
or   ( new_n1344_, new_n1343_, new_n1338_ );
xor  ( new_n1345_, RI2b1c4342be60_17, RI2b1c4342cd60_49 );
nor  ( new_n1346_, new_n1345_, new_n246_ );
and  ( new_n1347_, new_n1345_, new_n369_ );
or   ( new_n1348_, new_n1347_, new_n1346_ );
and  ( new_n1349_, new_n1348_, new_n273_ );
nor  ( new_n1350_, new_n1261_, new_n248_ );
and  ( new_n1351_, new_n1261_, new_n373_ );
or   ( new_n1352_, new_n1351_, new_n1350_ );
and  ( new_n1353_, new_n1352_, new_n270_ );
and  ( new_n1354_, new_n1353_, new_n1349_ );
or   ( new_n1355_, new_n1354_, new_n929_ );
and  ( new_n1356_, new_n1274_, new_n913_ );
and  ( new_n1357_, new_n1270_, new_n938_ );
or   ( new_n1358_, new_n1357_, new_n1356_ );
and  ( new_n1359_, new_n1358_, new_n1355_ );
and  ( new_n1360_, new_n1284_, new_n428_ );
and  ( new_n1361_, new_n1280_, new_n457_ );
or   ( new_n1362_, new_n1361_, new_n1360_ );
or   ( new_n1363_, new_n1358_, new_n1355_ );
and  ( new_n1364_, new_n1363_, new_n1362_ );
or   ( new_n1365_, new_n1364_, new_n1359_ );
and  ( new_n1366_, new_n1226_, new_n505_ );
and  ( new_n1367_, new_n1222_, new_n533_ );
or   ( new_n1368_, new_n1367_, new_n1366_ );
and  ( new_n1369_, new_n1235_, new_n590_ );
and  ( new_n1370_, new_n1231_, new_n619_ );
or   ( new_n1371_, new_n1370_, new_n1369_ );
and  ( new_n1372_, new_n1371_, new_n1368_ );
and  ( new_n1373_, new_n1245_, new_n734_ );
and  ( new_n1374_, new_n1241_, new_n762_ );
or   ( new_n1375_, new_n1374_, new_n1373_ );
or   ( new_n1376_, new_n1371_, new_n1368_ );
and  ( new_n1377_, new_n1376_, new_n1375_ );
or   ( new_n1378_, new_n1377_, new_n1372_ );
or   ( new_n1379_, new_n1378_, new_n1365_ );
and  ( new_n1380_, new_n1378_, new_n1365_ );
and  ( new_n1381_, new_n1297_, new_n785_ );
and  ( new_n1382_, new_n1293_, new_n813_ );
or   ( new_n1383_, new_n1382_, new_n1381_ );
and  ( new_n1384_, new_n1306_, new_n842_ );
and  ( new_n1385_, new_n1302_, new_n866_ );
or   ( new_n1386_, new_n1385_, new_n1384_ );
or   ( new_n1387_, new_n1386_, new_n1383_ );
and  ( new_n1388_, new_n1386_, new_n1383_ );
and  ( new_n1389_, new_n720_, RI2b1c4342db70_79 );
or   ( new_n1390_, new_n1389_, new_n1388_ );
and  ( new_n1391_, new_n1390_, new_n1387_ );
or   ( new_n1392_, new_n1391_, new_n1380_ );
and  ( new_n1393_, new_n1392_, new_n1379_ );
or   ( new_n1394_, new_n1393_, new_n1344_ );
and  ( new_n1395_, new_n1393_, new_n1344_ );
and  ( new_n1396_, new_n1324_, new_n1114_ );
and  ( new_n1397_, new_n1320_, new_n1163_ );
or   ( new_n1398_, new_n1397_, new_n1396_ );
or   ( new_n1399_, new_n1398_, new_n1395_ );
and  ( new_n1400_, new_n1399_, new_n1394_ );
and  ( new_n1401_, new_n1400_, new_n1332_ );
or   ( new_n1402_, new_n1401_, new_n1329_ );
and  ( new_n1403_, new_n1402_, new_n1176_ );
and  ( new_n1404_, new_n1174_, new_n901_ );
and  ( new_n1405_, new_n1171_, new_n1167_ );
or   ( new_n1406_, new_n1405_, new_n1404_ );
and  ( new_n1407_, new_n1400_, new_n1198_ );
and  ( new_n1408_, new_n1332_, new_n1328_ );
or   ( new_n1409_, new_n1408_, new_n1407_ );
and  ( new_n1410_, new_n1409_, new_n1406_ );
or   ( new_n1411_, new_n1410_, new_n1403_ );
or   ( new_n1412_, new_n1144_, new_n1001_ );
and  ( new_n1413_, new_n1412_, new_n1014_ );
and  ( new_n1414_, new_n1130_, new_n1000_ );
and  ( new_n1415_, new_n1143_, new_n969_ );
or   ( new_n1416_, new_n1415_, new_n1414_ );
and  ( new_n1417_, new_n1416_, new_n1150_ );
or   ( new_n1418_, new_n1417_, new_n1413_ );
and  ( new_n1419_, new_n1353_, new_n906_ );
and  ( new_n1420_, new_n1265_, new_n929_ );
and  ( new_n1421_, new_n1353_, new_n1257_ );
and  ( new_n1422_, new_n1349_, new_n1265_ );
or   ( new_n1423_, new_n1422_, new_n1421_ );
or   ( new_n1424_, new_n1423_, new_n1420_ );
or   ( new_n1425_, new_n1424_, new_n1419_ );
or   ( new_n1426_, new_n1425_, new_n99_ );
and  ( new_n1427_, new_n1426_, new_n1355_ );
and  ( new_n1428_, new_n1265_, new_n1257_ );
or   ( new_n1429_, new_n1428_, new_n1354_ );
and  ( new_n1430_, new_n1265_, new_n906_ );
and  ( new_n1431_, new_n1353_, new_n929_ );
or   ( new_n1432_, new_n1431_, new_n1430_ );
and  ( new_n1433_, new_n1432_, new_n1429_ );
and  ( new_n1434_, new_n1433_, RI2b1c4342d4e0_65 );
and  ( new_n1435_, new_n1434_, new_n1267_ );
or   ( new_n1436_, new_n1435_, new_n1427_ );
or   ( new_n1437_, new_n934_, new_n112_ );
or   ( new_n1438_, new_n940_, new_n526_ );
and  ( new_n1439_, new_n1438_, new_n1437_ );
and  ( new_n1440_, new_n1439_, new_n913_ );
and  ( new_n1441_, new_n944_, RI2b1c4342d5d0_67 );
and  ( new_n1442_, new_n932_, RI2b1c4342d558_66 );
or   ( new_n1443_, new_n1442_, new_n1441_ );
and  ( new_n1444_, new_n1443_, new_n938_ );
or   ( new_n1445_, new_n1444_, new_n1440_ );
and  ( new_n1446_, new_n1445_, new_n1436_ );
or   ( new_n1447_, new_n1445_, new_n1436_ );
or   ( new_n1448_, new_n453_, new_n591_ );
or   ( new_n1449_, new_n459_, new_n612_ );
and  ( new_n1450_, new_n1449_, new_n1448_ );
and  ( new_n1451_, new_n1450_, new_n428_ );
and  ( new_n1452_, new_n463_, RI2b1c4342d6c0_69 );
and  ( new_n1453_, new_n451_, RI2b1c4342d648_68 );
or   ( new_n1454_, new_n1453_, new_n1452_ );
and  ( new_n1455_, new_n1454_, new_n457_ );
or   ( new_n1456_, new_n1455_, new_n1451_ );
and  ( new_n1457_, new_n1456_, new_n1447_ );
or   ( new_n1458_, new_n1457_, new_n1446_ );
or   ( new_n1459_, new_n524_, new_n110_ );
or   ( new_n1460_, new_n528_, new_n755_ );
and  ( new_n1461_, new_n1460_, new_n1459_ );
and  ( new_n1462_, new_n1461_, new_n505_ );
and  ( new_n1463_, new_n537_, RI2b1c4342d7b0_71 );
and  ( new_n1464_, new_n522_, RI2b1c4342d738_70 );
or   ( new_n1465_, new_n1464_, new_n1463_ );
and  ( new_n1466_, new_n1465_, new_n533_ );
or   ( new_n1467_, new_n1466_, new_n1462_ );
or   ( new_n1468_, new_n610_, new_n105_ );
or   ( new_n1469_, new_n614_, new_n806_ );
and  ( new_n1470_, new_n1469_, new_n1468_ );
and  ( new_n1471_, new_n1470_, new_n590_ );
and  ( new_n1472_, new_n623_, RI2b1c4342d8a0_73 );
and  ( new_n1473_, new_n608_, RI2b1c4342d828_72 );
or   ( new_n1474_, new_n1473_, new_n1472_ );
and  ( new_n1475_, new_n1474_, new_n619_ );
or   ( new_n1476_, new_n1475_, new_n1471_ );
and  ( new_n1477_, new_n1476_, new_n1467_ );
or   ( new_n1478_, new_n1476_, new_n1467_ );
or   ( new_n1479_, new_n753_, new_n843_ );
or   ( new_n1480_, new_n757_, new_n859_ );
and  ( new_n1481_, new_n1480_, new_n1479_ );
and  ( new_n1482_, new_n1481_, new_n734_ );
and  ( new_n1483_, new_n766_, RI2b1c4342d990_75 );
and  ( new_n1484_, new_n751_, RI2b1c4342d918_74 );
or   ( new_n1485_, new_n1484_, new_n1483_ );
and  ( new_n1486_, new_n1485_, new_n762_ );
or   ( new_n1487_, new_n1486_, new_n1482_ );
and  ( new_n1488_, new_n1487_, new_n1478_ );
or   ( new_n1489_, new_n1488_, new_n1477_ );
and  ( new_n1490_, new_n1489_, new_n1458_ );
or   ( new_n1491_, new_n857_, new_n1310_ );
or   ( new_n1492_, new_n861_, new_n1002_ );
and  ( new_n1493_, new_n1492_, new_n1491_ );
and  ( new_n1494_, new_n1493_, new_n842_ );
and  ( new_n1495_, new_n870_, RI2b1c4342db70_79 );
and  ( new_n1496_, new_n855_, RI2b1c4342daf8_78 );
or   ( new_n1497_, new_n1496_, new_n1495_ );
and  ( new_n1498_, new_n1497_, new_n866_ );
or   ( new_n1499_, new_n1498_, new_n1494_ );
or   ( new_n1500_, new_n804_, new_n1004_ );
or   ( new_n1501_, new_n808_, new_n886_ );
and  ( new_n1502_, new_n1501_, new_n1500_ );
and  ( new_n1503_, new_n1502_, new_n785_ );
and  ( new_n1504_, new_n817_, RI2b1c4342da80_77 );
and  ( new_n1505_, new_n802_, RI2b1c4342da08_76 );
or   ( new_n1506_, new_n1505_, new_n1504_ );
and  ( new_n1507_, new_n1506_, new_n813_ );
or   ( new_n1508_, new_n1507_, new_n1503_ );
and  ( new_n1509_, new_n1508_, new_n1499_ );
or   ( new_n1510_, new_n1508_, new_n1499_ );
not  ( new_n1511_, RI2b1c4342dbe8_80 );
or   ( new_n1512_, new_n841_, new_n1511_ );
and  ( new_n1513_, new_n1512_, new_n1510_ );
or   ( new_n1514_, new_n1513_, new_n1509_ );
or   ( new_n1515_, new_n1489_, new_n1458_ );
and  ( new_n1516_, new_n1515_, new_n1514_ );
or   ( new_n1517_, new_n1516_, new_n1490_ );
or   ( new_n1518_, new_n1388_, new_n1309_ );
and  ( new_n1519_, new_n1518_, new_n1311_ );
and  ( new_n1520_, new_n1383_, new_n1308_ );
and  ( new_n1521_, new_n1386_, new_n1299_ );
or   ( new_n1522_, new_n1521_, new_n1520_ );
and  ( new_n1523_, new_n1522_, new_n1389_ );
or   ( new_n1524_, new_n1523_, new_n1519_ );
or   ( new_n1525_, new_n1372_, new_n1238_ );
and  ( new_n1526_, new_n1525_, new_n1247_ );
and  ( new_n1527_, new_n1368_, new_n1237_ );
and  ( new_n1528_, new_n1371_, new_n1228_ );
or   ( new_n1529_, new_n1528_, new_n1527_ );
and  ( new_n1530_, new_n1529_, new_n1375_ );
or   ( new_n1531_, new_n1530_, new_n1526_ );
and  ( new_n1532_, new_n1531_, new_n1524_ );
or   ( new_n1533_, new_n1359_, new_n1277_ );
and  ( new_n1534_, new_n1533_, new_n1286_ );
and  ( new_n1535_, new_n1355_, new_n1276_ );
and  ( new_n1536_, new_n1358_, new_n1267_ );
or   ( new_n1537_, new_n1536_, new_n1535_ );
and  ( new_n1538_, new_n1537_, new_n1362_ );
or   ( new_n1539_, new_n1538_, new_n1534_ );
or   ( new_n1540_, new_n1531_, new_n1524_ );
and  ( new_n1541_, new_n1540_, new_n1539_ );
or   ( new_n1542_, new_n1541_, new_n1532_ );
and  ( new_n1543_, new_n1542_, new_n1517_ );
or   ( new_n1544_, new_n1338_, new_n1209_ );
and  ( new_n1545_, new_n1544_, new_n1216_ );
and  ( new_n1546_, new_n1334_, new_n1208_ );
and  ( new_n1547_, new_n1337_, new_n1201_ );
or   ( new_n1548_, new_n1547_, new_n1546_ );
and  ( new_n1549_, new_n1548_, new_n1341_ );
or   ( new_n1550_, new_n1549_, new_n1545_ );
or   ( new_n1551_, new_n1542_, new_n1517_ );
and  ( new_n1552_, new_n1551_, new_n1550_ );
or   ( new_n1553_, new_n1552_, new_n1543_ );
and  ( new_n1554_, new_n1553_, new_n1418_ );
or   ( new_n1555_, new_n1553_, new_n1418_ );
or   ( new_n1556_, new_n1395_, new_n1318_ );
and  ( new_n1557_, new_n1556_, new_n1326_ );
and  ( new_n1558_, new_n1393_, new_n1219_ );
and  ( new_n1559_, new_n1344_, new_n1317_ );
or   ( new_n1560_, new_n1559_, new_n1558_ );
and  ( new_n1561_, new_n1560_, new_n1398_ );
or   ( new_n1562_, new_n1561_, new_n1557_ );
and  ( new_n1563_, new_n1562_, new_n1555_ );
or   ( new_n1564_, new_n1563_, new_n1554_ );
and  ( new_n1565_, new_n1564_, new_n1411_ );
and  ( new_n1566_, new_n1409_, new_n1176_ );
and  ( new_n1567_, new_n1406_, new_n1402_ );
or   ( new_n1568_, new_n1567_, new_n1566_ );
and  ( new_n1569_, new_n1416_, new_n1014_ );
and  ( new_n1570_, new_n1412_, new_n1150_ );
or   ( new_n1571_, new_n1570_, new_n1569_ );
and  ( new_n1572_, new_n1522_, new_n1311_ );
and  ( new_n1573_, new_n1518_, new_n1389_ );
or   ( new_n1574_, new_n1573_, new_n1572_ );
and  ( new_n1575_, new_n1529_, new_n1247_ );
and  ( new_n1576_, new_n1525_, new_n1375_ );
or   ( new_n1577_, new_n1576_, new_n1575_ );
and  ( new_n1578_, new_n1577_, new_n1574_ );
and  ( new_n1579_, new_n1537_, new_n1286_ );
and  ( new_n1580_, new_n1533_, new_n1362_ );
or   ( new_n1581_, new_n1580_, new_n1579_ );
or   ( new_n1582_, new_n1577_, new_n1574_ );
and  ( new_n1583_, new_n1582_, new_n1581_ );
or   ( new_n1584_, new_n1583_, new_n1578_ );
and  ( new_n1585_, new_n1434_, new_n1355_ );
and  ( new_n1586_, new_n1426_, new_n1267_ );
or   ( new_n1587_, new_n1586_, new_n1585_ );
and  ( new_n1588_, new_n1443_, new_n913_ );
and  ( new_n1589_, new_n1439_, new_n938_ );
or   ( new_n1590_, new_n1589_, new_n1588_ );
and  ( new_n1591_, new_n1590_, new_n1587_ );
or   ( new_n1592_, new_n1590_, new_n1587_ );
and  ( new_n1593_, new_n1454_, new_n428_ );
and  ( new_n1594_, new_n1450_, new_n457_ );
or   ( new_n1595_, new_n1594_, new_n1593_ );
and  ( new_n1596_, new_n1595_, new_n1592_ );
or   ( new_n1597_, new_n1596_, new_n1591_ );
and  ( new_n1598_, new_n1465_, new_n505_ );
and  ( new_n1599_, new_n1461_, new_n533_ );
or   ( new_n1600_, new_n1599_, new_n1598_ );
and  ( new_n1601_, new_n1474_, new_n590_ );
and  ( new_n1602_, new_n1470_, new_n619_ );
or   ( new_n1603_, new_n1602_, new_n1601_ );
and  ( new_n1604_, new_n1603_, new_n1600_ );
or   ( new_n1605_, new_n1603_, new_n1600_ );
and  ( new_n1606_, new_n1485_, new_n734_ );
and  ( new_n1607_, new_n1481_, new_n762_ );
or   ( new_n1608_, new_n1607_, new_n1606_ );
and  ( new_n1609_, new_n1608_, new_n1605_ );
or   ( new_n1610_, new_n1609_, new_n1604_ );
or   ( new_n1611_, new_n1610_, new_n1597_ );
and  ( new_n1612_, new_n1610_, new_n1597_ );
and  ( new_n1613_, new_n1506_, new_n785_ );
and  ( new_n1614_, new_n1502_, new_n813_ );
or   ( new_n1615_, new_n1614_, new_n1613_ );
and  ( new_n1616_, new_n1497_, new_n842_ );
and  ( new_n1617_, new_n1493_, new_n866_ );
or   ( new_n1618_, new_n1617_, new_n1616_ );
or   ( new_n1619_, new_n1618_, new_n1615_ );
and  ( new_n1620_, new_n1618_, new_n1615_ );
and  ( new_n1621_, new_n720_, RI2b1c4342dbe8_80 );
or   ( new_n1622_, new_n1621_, new_n1620_ );
and  ( new_n1623_, new_n1622_, new_n1619_ );
or   ( new_n1624_, new_n1623_, new_n1612_ );
and  ( new_n1625_, new_n1624_, new_n1611_ );
or   ( new_n1626_, new_n1625_, new_n1584_ );
and  ( new_n1627_, new_n1625_, new_n1584_ );
and  ( new_n1628_, new_n1548_, new_n1216_ );
and  ( new_n1629_, new_n1544_, new_n1341_ );
or   ( new_n1630_, new_n1629_, new_n1628_ );
or   ( new_n1631_, new_n1630_, new_n1627_ );
and  ( new_n1632_, new_n1631_, new_n1626_ );
or   ( new_n1633_, new_n1632_, new_n1571_ );
and  ( new_n1634_, new_n1632_, new_n1571_ );
and  ( new_n1635_, new_n1560_, new_n1326_ );
and  ( new_n1636_, new_n1556_, new_n1398_ );
or   ( new_n1637_, new_n1636_, new_n1635_ );
or   ( new_n1638_, new_n1637_, new_n1634_ );
and  ( new_n1639_, new_n1638_, new_n1633_ );
and  ( new_n1640_, new_n1639_, new_n1568_ );
or   ( new_n1641_, new_n1640_, new_n1565_ );
or   ( new_n1642_, new_n1634_, new_n1554_ );
and  ( new_n1643_, new_n1642_, new_n1562_ );
and  ( new_n1644_, new_n1632_, new_n1418_ );
and  ( new_n1645_, new_n1571_, new_n1553_ );
or   ( new_n1646_, new_n1645_, new_n1644_ );
and  ( new_n1647_, new_n1646_, new_n1637_ );
or   ( new_n1648_, new_n1647_, new_n1643_ );
or   ( new_n1649_, new_n1380_, new_n1290_ );
and  ( new_n1650_, new_n1649_, new_n1314_ );
and  ( new_n1651_, new_n1365_, new_n1250_ );
and  ( new_n1652_, new_n1378_, new_n1289_ );
or   ( new_n1653_, new_n1652_, new_n1651_ );
and  ( new_n1654_, new_n1653_, new_n1391_ );
or   ( new_n1655_, new_n1654_, new_n1650_ );
or   ( new_n1656_, new_n1604_, new_n1477_ );
and  ( new_n1657_, new_n1656_, new_n1487_ );
and  ( new_n1658_, new_n1600_, new_n1476_ );
and  ( new_n1659_, new_n1603_, new_n1467_ );
or   ( new_n1660_, new_n1659_, new_n1658_ );
and  ( new_n1661_, new_n1660_, new_n1608_ );
or   ( new_n1662_, new_n1661_, new_n1657_ );
or   ( new_n1663_, new_n1620_, new_n1509_ );
and  ( new_n1664_, new_n1663_, new_n1512_ );
and  ( new_n1665_, new_n1615_, new_n1499_ );
and  ( new_n1666_, new_n1618_, new_n1508_ );
or   ( new_n1667_, new_n1666_, new_n1665_ );
and  ( new_n1668_, new_n1667_, new_n1621_ );
or   ( new_n1669_, new_n1668_, new_n1664_ );
and  ( new_n1670_, new_n1669_, new_n1662_ );
or   ( new_n1671_, new_n453_, new_n755_ );
or   ( new_n1672_, new_n459_, new_n591_ );
and  ( new_n1673_, new_n1672_, new_n1671_ );
and  ( new_n1674_, new_n1673_, new_n428_ );
and  ( new_n1675_, new_n463_, RI2b1c4342d738_70 );
and  ( new_n1676_, new_n451_, RI2b1c4342d6c0_69 );
or   ( new_n1677_, new_n1676_, new_n1675_ );
and  ( new_n1678_, new_n1677_, new_n457_ );
or   ( new_n1679_, new_n1678_, new_n1674_ );
or   ( new_n1680_, new_n524_, new_n806_ );
or   ( new_n1681_, new_n528_, new_n110_ );
and  ( new_n1682_, new_n1681_, new_n1680_ );
and  ( new_n1683_, new_n1682_, new_n505_ );
and  ( new_n1684_, new_n537_, RI2b1c4342d828_72 );
and  ( new_n1685_, new_n522_, RI2b1c4342d7b0_71 );
or   ( new_n1686_, new_n1685_, new_n1684_ );
and  ( new_n1687_, new_n1686_, new_n533_ );
or   ( new_n1688_, new_n1687_, new_n1683_ );
and  ( new_n1689_, new_n1688_, new_n1679_ );
or   ( new_n1690_, new_n610_, new_n859_ );
or   ( new_n1691_, new_n614_, new_n105_ );
and  ( new_n1692_, new_n1691_, new_n1690_ );
and  ( new_n1693_, new_n1692_, new_n590_ );
and  ( new_n1694_, new_n623_, RI2b1c4342d918_74 );
and  ( new_n1695_, new_n608_, RI2b1c4342d8a0_73 );
or   ( new_n1696_, new_n1695_, new_n1694_ );
and  ( new_n1697_, new_n1696_, new_n619_ );
or   ( new_n1698_, new_n1697_, new_n1693_ );
or   ( new_n1699_, new_n1688_, new_n1679_ );
and  ( new_n1700_, new_n1699_, new_n1698_ );
or   ( new_n1701_, new_n1700_, new_n1689_ );
xor  ( new_n1702_, new_n278_, new_n153_ );
and  ( new_n1703_, new_n1702_, new_n367_ );
xor  ( new_n1704_, RI2b1c4342bed8_18, RI2b1c4342cdd8_50 );
and  ( new_n1705_, new_n1704_, new_n138_ );
and  ( new_n1706_, new_n1705_, new_n243_ );
or   ( new_n1707_, new_n1706_, new_n154_ );
or   ( new_n1708_, new_n1707_, new_n1703_ );
xor  ( new_n1709_, new_n281_, new_n157_ );
and  ( new_n1710_, new_n1709_, new_n365_ );
xor  ( new_n1711_, RI2b1c4342bf50_19, RI2b1c4342ce50_51 );
and  ( new_n1712_, new_n1711_, new_n138_ );
and  ( new_n1713_, new_n1712_, new_n241_ );
or   ( new_n1714_, new_n1713_, new_n158_ );
or   ( new_n1715_, new_n1714_, new_n1710_ );
or   ( new_n1716_, new_n1715_, new_n1708_ );
and  ( new_n1717_, new_n1716_, new_n1349_ );
or   ( new_n1718_, new_n1425_, new_n526_ );
or   ( new_n1719_, new_n1429_, new_n99_ );
and  ( new_n1720_, new_n1719_, new_n1718_ );
and  ( new_n1721_, new_n1720_, new_n1355_ );
and  ( new_n1722_, new_n1433_, RI2b1c4342d558_66 );
and  ( new_n1723_, new_n1423_, RI2b1c4342d4e0_65 );
or   ( new_n1724_, new_n1723_, new_n1722_ );
and  ( new_n1725_, new_n1724_, new_n1267_ );
or   ( new_n1726_, new_n1725_, new_n1721_ );
and  ( new_n1727_, new_n1726_, new_n1717_ );
or   ( new_n1728_, new_n1726_, new_n1717_ );
or   ( new_n1729_, new_n934_, new_n612_ );
or   ( new_n1730_, new_n940_, new_n112_ );
and  ( new_n1731_, new_n1730_, new_n1729_ );
and  ( new_n1732_, new_n1731_, new_n913_ );
and  ( new_n1733_, new_n944_, RI2b1c4342d648_68 );
and  ( new_n1734_, new_n932_, RI2b1c4342d5d0_67 );
or   ( new_n1735_, new_n1734_, new_n1733_ );
and  ( new_n1736_, new_n1735_, new_n938_ );
or   ( new_n1737_, new_n1736_, new_n1732_ );
and  ( new_n1738_, new_n1737_, new_n1728_ );
or   ( new_n1739_, new_n1738_, new_n1727_ );
and  ( new_n1740_, new_n1739_, new_n1701_ );
or   ( new_n1741_, new_n1739_, new_n1701_ );
or   ( new_n1742_, new_n753_, new_n886_ );
or   ( new_n1743_, new_n757_, new_n843_ );
and  ( new_n1744_, new_n1743_, new_n1742_ );
and  ( new_n1745_, new_n1744_, new_n734_ );
and  ( new_n1746_, new_n766_, RI2b1c4342da08_76 );
and  ( new_n1747_, new_n751_, RI2b1c4342d990_75 );
or   ( new_n1748_, new_n1747_, new_n1746_ );
and  ( new_n1749_, new_n1748_, new_n762_ );
or   ( new_n1750_, new_n1749_, new_n1745_ );
or   ( new_n1751_, new_n804_, new_n1002_ );
or   ( new_n1752_, new_n808_, new_n1004_ );
and  ( new_n1753_, new_n1752_, new_n1751_ );
and  ( new_n1754_, new_n1753_, new_n785_ );
and  ( new_n1755_, new_n817_, RI2b1c4342daf8_78 );
and  ( new_n1756_, new_n802_, RI2b1c4342da80_77 );
or   ( new_n1757_, new_n1756_, new_n1755_ );
and  ( new_n1758_, new_n1757_, new_n813_ );
or   ( new_n1759_, new_n1758_, new_n1754_ );
and  ( new_n1760_, new_n1759_, new_n1750_ );
or   ( new_n1761_, new_n857_, new_n1511_ );
or   ( new_n1762_, new_n861_, new_n1310_ );
and  ( new_n1763_, new_n1762_, new_n1761_ );
and  ( new_n1764_, new_n1763_, new_n842_ );
and  ( new_n1765_, new_n870_, RI2b1c4342dbe8_80 );
and  ( new_n1766_, new_n855_, RI2b1c4342db70_79 );
or   ( new_n1767_, new_n1766_, new_n1765_ );
and  ( new_n1768_, new_n1767_, new_n866_ );
or   ( new_n1769_, new_n1768_, new_n1764_ );
or   ( new_n1770_, new_n1759_, new_n1750_ );
and  ( new_n1771_, new_n1770_, new_n1769_ );
or   ( new_n1772_, new_n1771_, new_n1760_ );
and  ( new_n1773_, new_n1772_, new_n1741_ );
or   ( new_n1774_, new_n1773_, new_n1740_ );
and  ( new_n1775_, new_n1774_, new_n1670_ );
or   ( new_n1776_, new_n1578_, new_n1532_ );
and  ( new_n1777_, new_n1776_, new_n1539_ );
and  ( new_n1778_, new_n1574_, new_n1531_ );
and  ( new_n1779_, new_n1577_, new_n1524_ );
or   ( new_n1780_, new_n1779_, new_n1778_ );
and  ( new_n1781_, new_n1780_, new_n1581_ );
or   ( new_n1782_, new_n1781_, new_n1777_ );
or   ( new_n1783_, new_n1774_, new_n1670_ );
and  ( new_n1784_, new_n1783_, new_n1782_ );
or   ( new_n1785_, new_n1784_, new_n1775_ );
and  ( new_n1786_, new_n1785_, new_n1655_ );
or   ( new_n1787_, new_n1627_, new_n1543_ );
and  ( new_n1788_, new_n1787_, new_n1550_ );
and  ( new_n1789_, new_n1625_, new_n1542_ );
and  ( new_n1790_, new_n1584_, new_n1517_ );
or   ( new_n1791_, new_n1790_, new_n1789_ );
and  ( new_n1792_, new_n1791_, new_n1630_ );
or   ( new_n1793_, new_n1792_, new_n1788_ );
or   ( new_n1794_, new_n1785_, new_n1655_ );
and  ( new_n1795_, new_n1794_, new_n1793_ );
or   ( new_n1796_, new_n1795_, new_n1786_ );
or   ( new_n1797_, new_n1796_, new_n1648_ );
and  ( new_n1798_, new_n1797_, new_n1641_ );
and  ( new_n1799_, new_n1796_, new_n1648_ );
and  ( new_n1800_, new_n1646_, new_n1562_ );
and  ( new_n1801_, new_n1642_, new_n1637_ );
or   ( new_n1802_, new_n1801_, new_n1800_ );
and  ( new_n1803_, new_n1653_, new_n1314_ );
and  ( new_n1804_, new_n1649_, new_n1391_ );
or   ( new_n1805_, new_n1804_, new_n1803_ );
and  ( new_n1806_, new_n1667_, new_n1512_ );
and  ( new_n1807_, new_n1663_, new_n1621_ );
or   ( new_n1808_, new_n1807_, new_n1806_ );
and  ( new_n1809_, new_n1660_, new_n1487_ );
and  ( new_n1810_, new_n1656_, new_n1608_ );
or   ( new_n1811_, new_n1810_, new_n1809_ );
or   ( new_n1812_, new_n1811_, new_n1808_ );
not  ( new_n1813_, new_n241_ );
nor  ( new_n1814_, new_n1711_, new_n1813_ );
and  ( new_n1815_, new_n1711_, new_n365_ );
or   ( new_n1816_, new_n1815_, new_n1814_ );
and  ( new_n1817_, new_n1816_, new_n281_ );
not  ( new_n1818_, new_n243_ );
nor  ( new_n1819_, new_n1704_, new_n1818_ );
and  ( new_n1820_, new_n1704_, new_n367_ );
or   ( new_n1821_, new_n1820_, new_n1819_ );
and  ( new_n1822_, new_n1821_, new_n278_ );
and  ( new_n1823_, new_n1822_, new_n1817_ );
or   ( new_n1824_, new_n1823_, new_n1257_ );
and  ( new_n1825_, new_n1724_, new_n1355_ );
and  ( new_n1826_, new_n1720_, new_n1267_ );
or   ( new_n1827_, new_n1826_, new_n1825_ );
and  ( new_n1828_, new_n1827_, new_n1824_ );
or   ( new_n1829_, new_n1827_, new_n1824_ );
and  ( new_n1830_, new_n1735_, new_n913_ );
and  ( new_n1831_, new_n1731_, new_n938_ );
or   ( new_n1832_, new_n1831_, new_n1830_ );
and  ( new_n1833_, new_n1832_, new_n1829_ );
or   ( new_n1834_, new_n1833_, new_n1828_ );
and  ( new_n1835_, new_n1677_, new_n428_ );
and  ( new_n1836_, new_n1673_, new_n457_ );
or   ( new_n1837_, new_n1836_, new_n1835_ );
and  ( new_n1838_, new_n1686_, new_n505_ );
and  ( new_n1839_, new_n1682_, new_n533_ );
or   ( new_n1840_, new_n1839_, new_n1838_ );
and  ( new_n1841_, new_n1840_, new_n1837_ );
and  ( new_n1842_, new_n1696_, new_n590_ );
and  ( new_n1843_, new_n1692_, new_n619_ );
or   ( new_n1844_, new_n1843_, new_n1842_ );
or   ( new_n1845_, new_n1840_, new_n1837_ );
and  ( new_n1846_, new_n1845_, new_n1844_ );
or   ( new_n1847_, new_n1846_, new_n1841_ );
and  ( new_n1848_, new_n1847_, new_n1834_ );
or   ( new_n1849_, new_n1847_, new_n1834_ );
and  ( new_n1850_, new_n1748_, new_n734_ );
and  ( new_n1851_, new_n1744_, new_n762_ );
or   ( new_n1852_, new_n1851_, new_n1850_ );
and  ( new_n1853_, new_n1757_, new_n785_ );
and  ( new_n1854_, new_n1753_, new_n813_ );
or   ( new_n1855_, new_n1854_, new_n1853_ );
and  ( new_n1856_, new_n1855_, new_n1852_ );
and  ( new_n1857_, new_n1767_, new_n842_ );
and  ( new_n1858_, new_n1763_, new_n866_ );
or   ( new_n1859_, new_n1858_, new_n1857_ );
or   ( new_n1860_, new_n1855_, new_n1852_ );
and  ( new_n1861_, new_n1860_, new_n1859_ );
or   ( new_n1862_, new_n1861_, new_n1856_ );
and  ( new_n1863_, new_n1862_, new_n1849_ );
or   ( new_n1864_, new_n1863_, new_n1848_ );
and  ( new_n1865_, new_n1864_, new_n1812_ );
and  ( new_n1866_, new_n1780_, new_n1539_ );
and  ( new_n1867_, new_n1776_, new_n1581_ );
or   ( new_n1868_, new_n1867_, new_n1866_ );
or   ( new_n1869_, new_n1864_, new_n1812_ );
and  ( new_n1870_, new_n1869_, new_n1868_ );
or   ( new_n1871_, new_n1870_, new_n1865_ );
and  ( new_n1872_, new_n1871_, new_n1805_ );
and  ( new_n1873_, new_n1791_, new_n1550_ );
and  ( new_n1874_, new_n1787_, new_n1630_ );
or   ( new_n1875_, new_n1874_, new_n1873_ );
or   ( new_n1876_, new_n1871_, new_n1805_ );
and  ( new_n1877_, new_n1876_, new_n1875_ );
or   ( new_n1878_, new_n1877_, new_n1872_ );
and  ( new_n1879_, new_n1878_, new_n1802_ );
or   ( new_n1880_, new_n1879_, new_n1799_ );
or   ( new_n1881_, new_n1848_, new_n1740_ );
and  ( new_n1882_, new_n1881_, new_n1772_ );
and  ( new_n1883_, new_n1834_, new_n1701_ );
and  ( new_n1884_, new_n1847_, new_n1739_ );
or   ( new_n1885_, new_n1884_, new_n1883_ );
and  ( new_n1886_, new_n1885_, new_n1862_ );
or   ( new_n1887_, new_n1886_, new_n1882_ );
or   ( new_n1888_, new_n1591_, new_n1446_ );
and  ( new_n1889_, new_n1888_, new_n1456_ );
and  ( new_n1890_, new_n1587_, new_n1445_ );
and  ( new_n1891_, new_n1590_, new_n1436_ );
or   ( new_n1892_, new_n1891_, new_n1890_ );
and  ( new_n1893_, new_n1892_, new_n1595_ );
or   ( new_n1894_, new_n1893_, new_n1889_ );
or   ( new_n1895_, new_n1425_, new_n112_ );
or   ( new_n1896_, new_n1429_, new_n526_ );
and  ( new_n1897_, new_n1896_, new_n1895_ );
and  ( new_n1898_, new_n1897_, new_n1355_ );
and  ( new_n1899_, new_n1433_, RI2b1c4342d5d0_67 );
and  ( new_n1900_, new_n1423_, RI2b1c4342d558_66 );
or   ( new_n1901_, new_n1900_, new_n1899_ );
and  ( new_n1902_, new_n1901_, new_n1267_ );
or   ( new_n1903_, new_n1902_, new_n1898_ );
and  ( new_n1904_, new_n1822_, new_n1349_ );
and  ( new_n1905_, new_n1708_, new_n1257_ );
and  ( new_n1906_, new_n1822_, new_n1715_ );
and  ( new_n1907_, new_n1817_, new_n1708_ );
or   ( new_n1908_, new_n1907_, new_n1906_ );
or   ( new_n1909_, new_n1908_, new_n1905_ );
or   ( new_n1910_, new_n1909_, new_n1904_ );
or   ( new_n1911_, new_n1910_, new_n99_ );
and  ( new_n1912_, new_n1911_, new_n1824_ );
and  ( new_n1913_, new_n1715_, new_n1708_ );
or   ( new_n1914_, new_n1913_, new_n1823_ );
and  ( new_n1915_, new_n1708_, new_n1349_ );
and  ( new_n1916_, new_n1822_, new_n1257_ );
or   ( new_n1917_, new_n1916_, new_n1915_ );
and  ( new_n1918_, new_n1917_, new_n1914_ );
and  ( new_n1919_, new_n1918_, RI2b1c4342d4e0_65 );
and  ( new_n1920_, new_n1919_, new_n1717_ );
or   ( new_n1921_, new_n1920_, new_n1912_ );
and  ( new_n1922_, new_n1921_, new_n1903_ );
or   ( new_n1923_, new_n934_, new_n591_ );
or   ( new_n1924_, new_n940_, new_n612_ );
and  ( new_n1925_, new_n1924_, new_n1923_ );
and  ( new_n1926_, new_n1925_, new_n913_ );
and  ( new_n1927_, new_n944_, RI2b1c4342d6c0_69 );
and  ( new_n1928_, new_n932_, RI2b1c4342d648_68 );
or   ( new_n1929_, new_n1928_, new_n1927_ );
and  ( new_n1930_, new_n1929_, new_n938_ );
or   ( new_n1931_, new_n1930_, new_n1926_ );
or   ( new_n1932_, new_n1921_, new_n1903_ );
and  ( new_n1933_, new_n1932_, new_n1931_ );
or   ( new_n1934_, new_n1933_, new_n1922_ );
or   ( new_n1935_, new_n524_, new_n105_ );
or   ( new_n1936_, new_n528_, new_n806_ );
and  ( new_n1937_, new_n1936_, new_n1935_ );
and  ( new_n1938_, new_n1937_, new_n505_ );
and  ( new_n1939_, new_n537_, RI2b1c4342d8a0_73 );
and  ( new_n1940_, new_n522_, RI2b1c4342d828_72 );
or   ( new_n1941_, new_n1940_, new_n1939_ );
and  ( new_n1942_, new_n1941_, new_n533_ );
or   ( new_n1943_, new_n1942_, new_n1938_ );
or   ( new_n1944_, new_n453_, new_n110_ );
or   ( new_n1945_, new_n459_, new_n755_ );
and  ( new_n1946_, new_n1945_, new_n1944_ );
and  ( new_n1947_, new_n1946_, new_n428_ );
and  ( new_n1948_, new_n463_, RI2b1c4342d7b0_71 );
and  ( new_n1949_, new_n451_, RI2b1c4342d738_70 );
or   ( new_n1950_, new_n1949_, new_n1948_ );
and  ( new_n1951_, new_n1950_, new_n457_ );
or   ( new_n1952_, new_n1951_, new_n1947_ );
and  ( new_n1953_, new_n1952_, new_n1943_ );
or   ( new_n1954_, new_n610_, new_n843_ );
or   ( new_n1955_, new_n614_, new_n859_ );
and  ( new_n1956_, new_n1955_, new_n1954_ );
and  ( new_n1957_, new_n1956_, new_n590_ );
and  ( new_n1958_, new_n623_, RI2b1c4342d990_75 );
and  ( new_n1959_, new_n608_, RI2b1c4342d918_74 );
or   ( new_n1960_, new_n1959_, new_n1958_ );
and  ( new_n1961_, new_n1960_, new_n619_ );
or   ( new_n1962_, new_n1961_, new_n1957_ );
or   ( new_n1963_, new_n1952_, new_n1943_ );
and  ( new_n1964_, new_n1963_, new_n1962_ );
or   ( new_n1965_, new_n1964_, new_n1953_ );
and  ( new_n1966_, new_n1965_, new_n1934_ );
or   ( new_n1967_, new_n1965_, new_n1934_ );
or   ( new_n1968_, new_n753_, new_n1004_ );
or   ( new_n1969_, new_n757_, new_n886_ );
and  ( new_n1970_, new_n1969_, new_n1968_ );
and  ( new_n1971_, new_n1970_, new_n734_ );
and  ( new_n1972_, new_n766_, RI2b1c4342da80_77 );
and  ( new_n1973_, new_n751_, RI2b1c4342da08_76 );
or   ( new_n1974_, new_n1973_, new_n1972_ );
and  ( new_n1975_, new_n1974_, new_n762_ );
or   ( new_n1976_, new_n1975_, new_n1971_ );
or   ( new_n1977_, new_n804_, new_n1310_ );
or   ( new_n1978_, new_n808_, new_n1002_ );
and  ( new_n1979_, new_n1978_, new_n1977_ );
and  ( new_n1980_, new_n1979_, new_n785_ );
and  ( new_n1981_, new_n817_, RI2b1c4342db70_79 );
and  ( new_n1982_, new_n802_, RI2b1c4342daf8_78 );
or   ( new_n1983_, new_n1982_, new_n1981_ );
and  ( new_n1984_, new_n1983_, new_n813_ );
or   ( new_n1985_, new_n1984_, new_n1980_ );
and  ( new_n1986_, new_n1985_, new_n1976_ );
or   ( new_n1987_, new_n857_, new_n126_ );
or   ( new_n1988_, new_n861_, new_n1511_ );
and  ( new_n1989_, new_n1988_, new_n1987_ );
and  ( new_n1990_, new_n1989_, new_n842_ );
and  ( new_n1991_, new_n870_, RI2b1c4342dc60_81 );
and  ( new_n1992_, new_n855_, RI2b1c4342dbe8_80 );
or   ( new_n1993_, new_n1992_, new_n1991_ );
and  ( new_n1994_, new_n1993_, new_n866_ );
or   ( new_n1995_, new_n1994_, new_n1990_ );
or   ( new_n1996_, new_n1985_, new_n1976_ );
and  ( new_n1997_, new_n1996_, new_n1995_ );
or   ( new_n1998_, new_n1997_, new_n1986_ );
and  ( new_n1999_, new_n1998_, new_n1967_ );
or   ( new_n2000_, new_n1999_, new_n1966_ );
or   ( new_n2001_, new_n841_, new_n126_ );
or   ( new_n2002_, new_n1856_, new_n1760_ );
and  ( new_n2003_, new_n2002_, new_n1769_ );
and  ( new_n2004_, new_n1852_, new_n1759_ );
and  ( new_n2005_, new_n1855_, new_n1750_ );
or   ( new_n2006_, new_n2005_, new_n2004_ );
and  ( new_n2007_, new_n2006_, new_n1859_ );
or   ( new_n2008_, new_n2007_, new_n2003_ );
and  ( new_n2009_, new_n2008_, new_n2001_ );
or   ( new_n2010_, new_n2008_, new_n2001_ );
or   ( new_n2011_, new_n1841_, new_n1689_ );
and  ( new_n2012_, new_n2011_, new_n1698_ );
and  ( new_n2013_, new_n1837_, new_n1688_ );
and  ( new_n2014_, new_n1840_, new_n1679_ );
or   ( new_n2015_, new_n2014_, new_n2013_ );
and  ( new_n2016_, new_n2015_, new_n1844_ );
or   ( new_n2017_, new_n2016_, new_n2012_ );
and  ( new_n2018_, new_n2017_, new_n2010_ );
or   ( new_n2019_, new_n2018_, new_n2009_ );
and  ( new_n2020_, new_n2019_, new_n2000_ );
and  ( new_n2021_, new_n1919_, new_n1824_ );
and  ( new_n2022_, new_n1911_, new_n1717_ );
or   ( new_n2023_, new_n2022_, new_n2021_ );
and  ( new_n2024_, new_n1901_, new_n1355_ );
and  ( new_n2025_, new_n1897_, new_n1267_ );
or   ( new_n2026_, new_n2025_, new_n2024_ );
and  ( new_n2027_, new_n2026_, new_n2023_ );
and  ( new_n2028_, new_n1929_, new_n913_ );
and  ( new_n2029_, new_n1925_, new_n938_ );
or   ( new_n2030_, new_n2029_, new_n2028_ );
or   ( new_n2031_, new_n2026_, new_n2023_ );
and  ( new_n2032_, new_n2031_, new_n2030_ );
or   ( new_n2033_, new_n2032_, new_n2027_ );
and  ( new_n2034_, new_n1950_, new_n428_ );
and  ( new_n2035_, new_n1946_, new_n457_ );
or   ( new_n2036_, new_n2035_, new_n2034_ );
and  ( new_n2037_, new_n1941_, new_n505_ );
and  ( new_n2038_, new_n1937_, new_n533_ );
or   ( new_n2039_, new_n2038_, new_n2037_ );
and  ( new_n2040_, new_n2039_, new_n2036_ );
and  ( new_n2041_, new_n1960_, new_n590_ );
and  ( new_n2042_, new_n1956_, new_n619_ );
or   ( new_n2043_, new_n2042_, new_n2041_ );
or   ( new_n2044_, new_n2039_, new_n2036_ );
and  ( new_n2045_, new_n2044_, new_n2043_ );
or   ( new_n2046_, new_n2045_, new_n2040_ );
and  ( new_n2047_, new_n2046_, new_n2033_ );
or   ( new_n2048_, new_n2046_, new_n2033_ );
and  ( new_n2049_, new_n1974_, new_n734_ );
and  ( new_n2050_, new_n1970_, new_n762_ );
or   ( new_n2051_, new_n2050_, new_n2049_ );
and  ( new_n2052_, new_n1983_, new_n785_ );
and  ( new_n2053_, new_n1979_, new_n813_ );
or   ( new_n2054_, new_n2053_, new_n2052_ );
and  ( new_n2055_, new_n2054_, new_n2051_ );
and  ( new_n2056_, new_n1993_, new_n842_ );
and  ( new_n2057_, new_n1989_, new_n866_ );
or   ( new_n2058_, new_n2057_, new_n2056_ );
or   ( new_n2059_, new_n2054_, new_n2051_ );
and  ( new_n2060_, new_n2059_, new_n2058_ );
or   ( new_n2061_, new_n2060_, new_n2055_ );
and  ( new_n2062_, new_n2061_, new_n2048_ );
or   ( new_n2063_, new_n2062_, new_n2047_ );
and  ( new_n2064_, new_n720_, RI2b1c4342dc60_81 );
and  ( new_n2065_, new_n2006_, new_n1769_ );
and  ( new_n2066_, new_n2002_, new_n1859_ );
or   ( new_n2067_, new_n2066_, new_n2065_ );
and  ( new_n2068_, new_n2067_, new_n2064_ );
or   ( new_n2069_, new_n2067_, new_n2064_ );
and  ( new_n2070_, new_n2015_, new_n1698_ );
and  ( new_n2071_, new_n2011_, new_n1844_ );
or   ( new_n2072_, new_n2071_, new_n2070_ );
and  ( new_n2073_, new_n2072_, new_n2069_ );
or   ( new_n2074_, new_n2073_, new_n2068_ );
and  ( new_n2075_, new_n2074_, new_n2063_ );
or   ( new_n2076_, new_n2075_, new_n2020_ );
and  ( new_n2077_, new_n2076_, new_n1894_ );
and  ( new_n2078_, new_n1892_, new_n1456_ );
and  ( new_n2079_, new_n1888_, new_n1595_ );
or   ( new_n2080_, new_n2079_, new_n2078_ );
and  ( new_n2081_, new_n2063_, new_n2019_ );
and  ( new_n2082_, new_n2074_, new_n2000_ );
or   ( new_n2083_, new_n2082_, new_n2081_ );
and  ( new_n2084_, new_n2083_, new_n2080_ );
or   ( new_n2085_, new_n2084_, new_n2077_ );
or   ( new_n2086_, new_n2085_, new_n1887_ );
or   ( new_n2087_, new_n1828_, new_n1727_ );
and  ( new_n2088_, new_n2087_, new_n1737_ );
and  ( new_n2089_, new_n1824_, new_n1726_ );
and  ( new_n2090_, new_n1827_, new_n1717_ );
or   ( new_n2091_, new_n2090_, new_n2089_ );
and  ( new_n2092_, new_n2091_, new_n1832_ );
or   ( new_n2093_, new_n2092_, new_n2088_ );
or   ( new_n2094_, new_n2068_, new_n2009_ );
and  ( new_n2095_, new_n2094_, new_n2017_ );
and  ( new_n2096_, new_n2064_, new_n2008_ );
and  ( new_n2097_, new_n2067_, new_n2001_ );
or   ( new_n2098_, new_n2097_, new_n2096_ );
and  ( new_n2099_, new_n2098_, new_n2072_ );
or   ( new_n2100_, new_n2099_, new_n2095_ );
and  ( new_n2101_, new_n2100_, new_n2093_ );
or   ( new_n2102_, new_n2100_, new_n2093_ );
or   ( new_n2103_, new_n2047_, new_n1966_ );
and  ( new_n2104_, new_n2103_, new_n1998_ );
and  ( new_n2105_, new_n2033_, new_n1965_ );
and  ( new_n2106_, new_n2046_, new_n1934_ );
or   ( new_n2107_, new_n2106_, new_n2105_ );
and  ( new_n2108_, new_n2107_, new_n2061_ );
or   ( new_n2109_, new_n2108_, new_n2104_ );
and  ( new_n2110_, new_n2109_, new_n2102_ );
or   ( new_n2111_, new_n2110_, new_n2101_ );
or   ( new_n2112_, new_n2055_, new_n1986_ );
and  ( new_n2113_, new_n2112_, new_n1995_ );
and  ( new_n2114_, new_n2051_, new_n1985_ );
and  ( new_n2115_, new_n2054_, new_n1976_ );
or   ( new_n2116_, new_n2115_, new_n2114_ );
and  ( new_n2117_, new_n2116_, new_n2058_ );
or   ( new_n2118_, new_n2117_, new_n2113_ );
not  ( new_n2119_, RI2b1c4342dcd8_82 );
or   ( new_n2120_, new_n841_, new_n2119_ );
and  ( new_n2121_, new_n2120_, new_n2118_ );
or   ( new_n2122_, new_n934_, new_n755_ );
or   ( new_n2123_, new_n940_, new_n591_ );
and  ( new_n2124_, new_n2123_, new_n2122_ );
and  ( new_n2125_, new_n2124_, new_n913_ );
and  ( new_n2126_, new_n944_, RI2b1c4342d738_70 );
and  ( new_n2127_, new_n932_, RI2b1c4342d6c0_69 );
or   ( new_n2128_, new_n2127_, new_n2126_ );
and  ( new_n2129_, new_n2128_, new_n938_ );
or   ( new_n2130_, new_n2129_, new_n2125_ );
or   ( new_n2131_, new_n453_, new_n806_ );
or   ( new_n2132_, new_n459_, new_n110_ );
and  ( new_n2133_, new_n2132_, new_n2131_ );
and  ( new_n2134_, new_n2133_, new_n428_ );
and  ( new_n2135_, new_n463_, RI2b1c4342d828_72 );
and  ( new_n2136_, new_n451_, RI2b1c4342d7b0_71 );
or   ( new_n2137_, new_n2136_, new_n2135_ );
and  ( new_n2138_, new_n2137_, new_n457_ );
or   ( new_n2139_, new_n2138_, new_n2134_ );
and  ( new_n2140_, new_n2139_, new_n2130_ );
or   ( new_n2141_, new_n524_, new_n859_ );
or   ( new_n2142_, new_n528_, new_n105_ );
and  ( new_n2143_, new_n2142_, new_n2141_ );
and  ( new_n2144_, new_n2143_, new_n505_ );
and  ( new_n2145_, new_n537_, RI2b1c4342d918_74 );
and  ( new_n2146_, new_n522_, RI2b1c4342d8a0_73 );
or   ( new_n2147_, new_n2146_, new_n2145_ );
and  ( new_n2148_, new_n2147_, new_n533_ );
or   ( new_n2149_, new_n2148_, new_n2144_ );
or   ( new_n2150_, new_n2139_, new_n2130_ );
and  ( new_n2151_, new_n2150_, new_n2149_ );
or   ( new_n2152_, new_n2151_, new_n2140_ );
xor  ( new_n2153_, new_n288_, new_n161_ );
and  ( new_n2154_, new_n2153_, new_n363_ );
xor  ( new_n2155_, RI2b1c4342bfc8_20, RI2b1c4342cec8_52 );
and  ( new_n2156_, new_n2155_, new_n138_ );
and  ( new_n2157_, new_n2156_, new_n239_ );
or   ( new_n2158_, new_n2157_, new_n162_ );
or   ( new_n2159_, new_n2158_, new_n2154_ );
xor  ( new_n2160_, new_n291_, new_n165_ );
and  ( new_n2161_, new_n2160_, new_n361_ );
xor  ( new_n2162_, RI2b1c4342c040_21, RI2b1c4342cf40_53 );
and  ( new_n2163_, new_n2162_, new_n138_ );
and  ( new_n2164_, new_n2163_, new_n237_ );
or   ( new_n2165_, new_n2164_, new_n166_ );
or   ( new_n2166_, new_n2165_, new_n2161_ );
or   ( new_n2167_, new_n2166_, new_n2159_ );
and  ( new_n2168_, new_n2167_, new_n1817_ );
or   ( new_n2169_, new_n1910_, new_n526_ );
or   ( new_n2170_, new_n1914_, new_n99_ );
and  ( new_n2171_, new_n2170_, new_n2169_ );
and  ( new_n2172_, new_n2171_, new_n1824_ );
and  ( new_n2173_, new_n1918_, RI2b1c4342d558_66 );
and  ( new_n2174_, new_n1908_, RI2b1c4342d4e0_65 );
or   ( new_n2175_, new_n2174_, new_n2173_ );
and  ( new_n2176_, new_n2175_, new_n1717_ );
or   ( new_n2177_, new_n2176_, new_n2172_ );
and  ( new_n2178_, new_n2177_, new_n2168_ );
or   ( new_n2179_, new_n1425_, new_n612_ );
or   ( new_n2180_, new_n1429_, new_n112_ );
and  ( new_n2181_, new_n2180_, new_n2179_ );
and  ( new_n2182_, new_n2181_, new_n1355_ );
and  ( new_n2183_, new_n1433_, RI2b1c4342d648_68 );
and  ( new_n2184_, new_n1423_, RI2b1c4342d5d0_67 );
or   ( new_n2185_, new_n2184_, new_n2183_ );
and  ( new_n2186_, new_n2185_, new_n1267_ );
or   ( new_n2187_, new_n2186_, new_n2182_ );
or   ( new_n2188_, new_n2177_, new_n2168_ );
and  ( new_n2189_, new_n2188_, new_n2187_ );
or   ( new_n2190_, new_n2189_, new_n2178_ );
and  ( new_n2191_, new_n2190_, new_n2152_ );
or   ( new_n2192_, new_n610_, new_n886_ );
or   ( new_n2193_, new_n614_, new_n843_ );
and  ( new_n2194_, new_n2193_, new_n2192_ );
and  ( new_n2195_, new_n2194_, new_n590_ );
and  ( new_n2196_, new_n623_, RI2b1c4342da08_76 );
and  ( new_n2197_, new_n608_, RI2b1c4342d990_75 );
or   ( new_n2198_, new_n2197_, new_n2196_ );
and  ( new_n2199_, new_n2198_, new_n619_ );
or   ( new_n2200_, new_n2199_, new_n2195_ );
or   ( new_n2201_, new_n753_, new_n1002_ );
or   ( new_n2202_, new_n757_, new_n1004_ );
and  ( new_n2203_, new_n2202_, new_n2201_ );
and  ( new_n2204_, new_n2203_, new_n734_ );
and  ( new_n2205_, new_n766_, RI2b1c4342daf8_78 );
and  ( new_n2206_, new_n751_, RI2b1c4342da80_77 );
or   ( new_n2207_, new_n2206_, new_n2205_ );
and  ( new_n2208_, new_n2207_, new_n762_ );
or   ( new_n2209_, new_n2208_, new_n2204_ );
and  ( new_n2210_, new_n2209_, new_n2200_ );
or   ( new_n2211_, new_n804_, new_n1511_ );
or   ( new_n2212_, new_n808_, new_n1310_ );
and  ( new_n2213_, new_n2212_, new_n2211_ );
and  ( new_n2214_, new_n2213_, new_n785_ );
and  ( new_n2215_, new_n817_, RI2b1c4342dbe8_80 );
and  ( new_n2216_, new_n802_, RI2b1c4342db70_79 );
or   ( new_n2217_, new_n2216_, new_n2215_ );
and  ( new_n2218_, new_n2217_, new_n813_ );
or   ( new_n2219_, new_n2218_, new_n2214_ );
or   ( new_n2220_, new_n2209_, new_n2200_ );
and  ( new_n2221_, new_n2220_, new_n2219_ );
or   ( new_n2222_, new_n2221_, new_n2210_ );
or   ( new_n2223_, new_n2190_, new_n2152_ );
and  ( new_n2224_, new_n2223_, new_n2222_ );
or   ( new_n2225_, new_n2224_, new_n2191_ );
and  ( new_n2226_, new_n2225_, new_n2121_ );
or   ( new_n2227_, new_n2225_, new_n2121_ );
or   ( new_n2228_, new_n2040_, new_n1953_ );
and  ( new_n2229_, new_n2228_, new_n1962_ );
and  ( new_n2230_, new_n2036_, new_n1943_ );
and  ( new_n2231_, new_n2039_, new_n1952_ );
or   ( new_n2232_, new_n2231_, new_n2230_ );
and  ( new_n2233_, new_n2232_, new_n2043_ );
or   ( new_n2234_, new_n2233_, new_n2229_ );
or   ( new_n2235_, new_n2027_, new_n1922_ );
and  ( new_n2236_, new_n2235_, new_n1931_ );
and  ( new_n2237_, new_n2023_, new_n1903_ );
and  ( new_n2238_, new_n2026_, new_n1921_ );
or   ( new_n2239_, new_n2238_, new_n2237_ );
and  ( new_n2240_, new_n2239_, new_n2030_ );
or   ( new_n2241_, new_n2240_, new_n2236_ );
or   ( new_n2242_, new_n2241_, new_n2234_ );
and  ( new_n2243_, new_n2242_, new_n2227_ );
or   ( new_n2244_, new_n2243_, new_n2226_ );
and  ( new_n2245_, new_n2244_, new_n2111_ );
or   ( new_n2246_, new_n2244_, new_n2111_ );
and  ( new_n2247_, new_n1808_, new_n1662_ );
and  ( new_n2248_, new_n1811_, new_n1669_ );
or   ( new_n2249_, new_n2248_, new_n2247_ );
and  ( new_n2250_, new_n2249_, new_n2246_ );
or   ( new_n2251_, new_n2250_, new_n2245_ );
and  ( new_n2252_, new_n2251_, new_n2086_ );
or   ( new_n2253_, new_n1612_, new_n1490_ );
and  ( new_n2254_, new_n2253_, new_n1514_ );
and  ( new_n2255_, new_n1597_, new_n1489_ );
and  ( new_n2256_, new_n1610_, new_n1458_ );
or   ( new_n2257_, new_n2256_, new_n2255_ );
and  ( new_n2258_, new_n2257_, new_n1623_ );
or   ( new_n2259_, new_n2258_, new_n2254_ );
or   ( new_n2260_, new_n2019_, new_n2000_ );
and  ( new_n2261_, new_n2260_, new_n1894_ );
or   ( new_n2262_, new_n2261_, new_n2020_ );
and  ( new_n2263_, new_n2262_, new_n2259_ );
and  ( new_n2264_, new_n2257_, new_n1514_ );
and  ( new_n2265_, new_n2253_, new_n1623_ );
or   ( new_n2266_, new_n2265_, new_n2264_ );
or   ( new_n2267_, new_n2074_, new_n2063_ );
and  ( new_n2268_, new_n2267_, new_n2080_ );
or   ( new_n2269_, new_n2268_, new_n2075_ );
and  ( new_n2270_, new_n2269_, new_n2266_ );
or   ( new_n2271_, new_n2270_, new_n2263_ );
or   ( new_n2272_, new_n1865_, new_n1775_ );
and  ( new_n2273_, new_n2272_, new_n1782_ );
and  ( new_n2274_, new_n1864_, new_n1670_ );
and  ( new_n2275_, new_n1812_, new_n1774_ );
or   ( new_n2276_, new_n2275_, new_n2274_ );
and  ( new_n2277_, new_n2276_, new_n1868_ );
or   ( new_n2278_, new_n2277_, new_n2273_ );
and  ( new_n2279_, new_n2278_, new_n2271_ );
and  ( new_n2280_, new_n2269_, new_n2259_ );
and  ( new_n2281_, new_n2266_, new_n2262_ );
or   ( new_n2282_, new_n2281_, new_n2280_ );
and  ( new_n2283_, new_n2276_, new_n1782_ );
and  ( new_n2284_, new_n2272_, new_n1868_ );
or   ( new_n2285_, new_n2284_, new_n2283_ );
and  ( new_n2286_, new_n2285_, new_n2282_ );
or   ( new_n2287_, new_n2286_, new_n2279_ );
or   ( new_n2288_, new_n2251_, new_n2086_ );
and  ( new_n2289_, new_n2288_, new_n2287_ );
or   ( new_n2290_, new_n2289_, new_n2252_ );
or   ( new_n2291_, new_n2262_, new_n2259_ );
and  ( new_n2292_, new_n2291_, new_n2278_ );
or   ( new_n2293_, new_n2292_, new_n2263_ );
and  ( new_n2294_, new_n2293_, new_n2290_ );
or   ( new_n2295_, new_n1872_, new_n1786_ );
and  ( new_n2296_, new_n2295_, new_n1793_ );
and  ( new_n2297_, new_n1871_, new_n1655_ );
and  ( new_n2298_, new_n1805_, new_n1785_ );
or   ( new_n2299_, new_n2298_, new_n2297_ );
and  ( new_n2300_, new_n2299_, new_n1875_ );
or   ( new_n2301_, new_n2300_, new_n2296_ );
or   ( new_n2302_, new_n2293_, new_n2290_ );
and  ( new_n2303_, new_n2302_, new_n2301_ );
or   ( new_n2304_, new_n2303_, new_n2294_ );
or   ( new_n2305_, new_n2304_, new_n1880_ );
or   ( new_n2306_, new_n1797_, new_n1641_ );
and  ( new_n2307_, new_n2306_, new_n2305_ );
or   ( new_n2308_, new_n2307_, new_n1798_ );
and  ( new_n2309_, new_n2304_, new_n1880_ );
or   ( new_n2310_, new_n2309_, new_n1798_ );
and  ( new_n2311_, new_n1885_, new_n1772_ );
and  ( new_n2312_, new_n1881_, new_n1862_ );
or   ( new_n2313_, new_n2312_, new_n2311_ );
and  ( new_n2314_, new_n2083_, new_n1894_ );
and  ( new_n2315_, new_n2080_, new_n2076_ );
or   ( new_n2316_, new_n2315_, new_n2314_ );
and  ( new_n2317_, new_n2316_, new_n2313_ );
and  ( new_n2318_, new_n720_, RI2b1c4342dcd8_82 );
and  ( new_n2319_, new_n2116_, new_n1995_ );
and  ( new_n2320_, new_n2112_, new_n2058_ );
or   ( new_n2321_, new_n2320_, new_n2319_ );
or   ( new_n2322_, new_n2321_, new_n2318_ );
not  ( new_n2323_, new_n237_ );
nor  ( new_n2324_, new_n2162_, new_n2323_ );
and  ( new_n2325_, new_n2162_, new_n361_ );
or   ( new_n2326_, new_n2325_, new_n2324_ );
and  ( new_n2327_, new_n2326_, new_n291_ );
not  ( new_n2328_, new_n239_ );
nor  ( new_n2329_, new_n2155_, new_n2328_ );
and  ( new_n2330_, new_n2155_, new_n363_ );
or   ( new_n2331_, new_n2330_, new_n2329_ );
and  ( new_n2332_, new_n2331_, new_n288_ );
and  ( new_n2333_, new_n2332_, new_n2327_ );
or   ( new_n2334_, new_n2333_, new_n1715_ );
and  ( new_n2335_, new_n2175_, new_n1824_ );
and  ( new_n2336_, new_n2171_, new_n1717_ );
or   ( new_n2337_, new_n2336_, new_n2335_ );
and  ( new_n2338_, new_n2337_, new_n2334_ );
and  ( new_n2339_, new_n2185_, new_n1355_ );
and  ( new_n2340_, new_n2181_, new_n1267_ );
or   ( new_n2341_, new_n2340_, new_n2339_ );
or   ( new_n2342_, new_n2337_, new_n2334_ );
and  ( new_n2343_, new_n2342_, new_n2341_ );
or   ( new_n2344_, new_n2343_, new_n2338_ );
and  ( new_n2345_, new_n2128_, new_n913_ );
and  ( new_n2346_, new_n2124_, new_n938_ );
or   ( new_n2347_, new_n2346_, new_n2345_ );
and  ( new_n2348_, new_n2137_, new_n428_ );
and  ( new_n2349_, new_n2133_, new_n457_ );
or   ( new_n2350_, new_n2349_, new_n2348_ );
and  ( new_n2351_, new_n2350_, new_n2347_ );
and  ( new_n2352_, new_n2147_, new_n505_ );
and  ( new_n2353_, new_n2143_, new_n533_ );
or   ( new_n2354_, new_n2353_, new_n2352_ );
or   ( new_n2355_, new_n2350_, new_n2347_ );
and  ( new_n2356_, new_n2355_, new_n2354_ );
or   ( new_n2357_, new_n2356_, new_n2351_ );
and  ( new_n2358_, new_n2357_, new_n2344_ );
and  ( new_n2359_, new_n2198_, new_n590_ );
and  ( new_n2360_, new_n2194_, new_n619_ );
or   ( new_n2361_, new_n2360_, new_n2359_ );
and  ( new_n2362_, new_n2207_, new_n734_ );
and  ( new_n2363_, new_n2203_, new_n762_ );
or   ( new_n2364_, new_n2363_, new_n2362_ );
and  ( new_n2365_, new_n2364_, new_n2361_ );
and  ( new_n2366_, new_n2217_, new_n785_ );
and  ( new_n2367_, new_n2213_, new_n813_ );
or   ( new_n2368_, new_n2367_, new_n2366_ );
or   ( new_n2369_, new_n2364_, new_n2361_ );
and  ( new_n2370_, new_n2369_, new_n2368_ );
or   ( new_n2371_, new_n2370_, new_n2365_ );
or   ( new_n2372_, new_n2357_, new_n2344_ );
and  ( new_n2373_, new_n2372_, new_n2371_ );
or   ( new_n2374_, new_n2373_, new_n2358_ );
and  ( new_n2375_, new_n2374_, new_n2322_ );
and  ( new_n2376_, new_n2232_, new_n1962_ );
and  ( new_n2377_, new_n2228_, new_n2043_ );
or   ( new_n2378_, new_n2377_, new_n2376_ );
and  ( new_n2379_, new_n2239_, new_n1931_ );
and  ( new_n2380_, new_n2235_, new_n2030_ );
or   ( new_n2381_, new_n2380_, new_n2379_ );
and  ( new_n2382_, new_n2381_, new_n2378_ );
or   ( new_n2383_, new_n2374_, new_n2322_ );
and  ( new_n2384_, new_n2383_, new_n2382_ );
or   ( new_n2385_, new_n2384_, new_n2375_ );
and  ( new_n2386_, new_n2091_, new_n1737_ );
and  ( new_n2387_, new_n2087_, new_n1832_ );
or   ( new_n2388_, new_n2387_, new_n2386_ );
and  ( new_n2389_, new_n2098_, new_n2017_ );
and  ( new_n2390_, new_n2094_, new_n2072_ );
or   ( new_n2391_, new_n2390_, new_n2389_ );
and  ( new_n2392_, new_n2391_, new_n2388_ );
or   ( new_n2393_, new_n2391_, new_n2388_ );
and  ( new_n2394_, new_n2107_, new_n1998_ );
and  ( new_n2395_, new_n2103_, new_n2061_ );
or   ( new_n2396_, new_n2395_, new_n2394_ );
and  ( new_n2397_, new_n2396_, new_n2393_ );
or   ( new_n2398_, new_n2397_, new_n2392_ );
and  ( new_n2399_, new_n2398_, new_n2385_ );
or   ( new_n2400_, new_n2398_, new_n2385_ );
and  ( new_n2401_, new_n1811_, new_n1808_ );
or   ( new_n2402_, new_n2401_, new_n1670_ );
and  ( new_n2403_, new_n2402_, new_n2400_ );
or   ( new_n2404_, new_n2403_, new_n2399_ );
and  ( new_n2405_, new_n2404_, new_n2317_ );
and  ( new_n2406_, new_n2282_, new_n2278_ );
and  ( new_n2407_, new_n2285_, new_n2271_ );
or   ( new_n2408_, new_n2407_, new_n2406_ );
or   ( new_n2409_, new_n2404_, new_n2317_ );
and  ( new_n2410_, new_n2409_, new_n2408_ );
or   ( new_n2411_, new_n2410_, new_n2405_ );
or   ( new_n2412_, new_n2269_, new_n2266_ );
and  ( new_n2413_, new_n2412_, new_n2285_ );
or   ( new_n2414_, new_n2413_, new_n2270_ );
and  ( new_n2415_, new_n2414_, new_n2411_ );
or   ( new_n2416_, new_n2415_, new_n2294_ );
and  ( new_n2417_, new_n2416_, new_n2301_ );
and  ( new_n2418_, new_n2299_, new_n1793_ );
and  ( new_n2419_, new_n2295_, new_n1875_ );
or   ( new_n2420_, new_n2419_, new_n2418_ );
and  ( new_n2421_, new_n2411_, new_n2293_ );
and  ( new_n2422_, new_n2414_, new_n2290_ );
or   ( new_n2423_, new_n2422_, new_n2421_ );
and  ( new_n2424_, new_n2423_, new_n2420_ );
or   ( new_n2425_, new_n2424_, new_n2417_ );
or   ( new_n2426_, new_n2405_, new_n2252_ );
and  ( new_n2427_, new_n2426_, new_n2287_ );
and  ( new_n2428_, new_n2404_, new_n2086_ );
and  ( new_n2429_, new_n2317_, new_n2251_ );
or   ( new_n2430_, new_n2429_, new_n2428_ );
and  ( new_n2431_, new_n2430_, new_n2408_ );
or   ( new_n2432_, new_n2431_, new_n2427_ );
and  ( new_n2433_, new_n2085_, new_n1887_ );
or   ( new_n2434_, new_n2433_, new_n2317_ );
or   ( new_n2435_, new_n1910_, new_n112_ );
or   ( new_n2436_, new_n1914_, new_n526_ );
and  ( new_n2437_, new_n2436_, new_n2435_ );
and  ( new_n2438_, new_n2437_, new_n1824_ );
and  ( new_n2439_, new_n1918_, RI2b1c4342d5d0_67 );
and  ( new_n2440_, new_n1908_, RI2b1c4342d558_66 );
or   ( new_n2441_, new_n2440_, new_n2439_ );
and  ( new_n2442_, new_n2441_, new_n1717_ );
or   ( new_n2443_, new_n2442_, new_n2438_ );
and  ( new_n2444_, new_n2332_, new_n1817_ );
and  ( new_n2445_, new_n2159_, new_n1715_ );
and  ( new_n2446_, new_n2332_, new_n2166_ );
and  ( new_n2447_, new_n2327_, new_n2159_ );
or   ( new_n2448_, new_n2447_, new_n2446_ );
or   ( new_n2449_, new_n2448_, new_n2445_ );
or   ( new_n2450_, new_n2449_, new_n2444_ );
or   ( new_n2451_, new_n2450_, new_n99_ );
and  ( new_n2452_, new_n2451_, new_n2334_ );
and  ( new_n2453_, new_n2166_, new_n2159_ );
or   ( new_n2454_, new_n2453_, new_n2333_ );
and  ( new_n2455_, new_n2159_, new_n1817_ );
and  ( new_n2456_, new_n2332_, new_n1715_ );
or   ( new_n2457_, new_n2456_, new_n2455_ );
and  ( new_n2458_, new_n2457_, new_n2454_ );
and  ( new_n2459_, new_n2458_, RI2b1c4342d4e0_65 );
and  ( new_n2460_, new_n2459_, new_n2168_ );
or   ( new_n2461_, new_n2460_, new_n2452_ );
and  ( new_n2462_, new_n2461_, new_n2443_ );
or   ( new_n2463_, new_n2461_, new_n2443_ );
or   ( new_n2464_, new_n1425_, new_n591_ );
or   ( new_n2465_, new_n1429_, new_n612_ );
and  ( new_n2466_, new_n2465_, new_n2464_ );
and  ( new_n2467_, new_n2466_, new_n1355_ );
and  ( new_n2468_, new_n1433_, RI2b1c4342d6c0_69 );
and  ( new_n2469_, new_n1423_, RI2b1c4342d648_68 );
or   ( new_n2470_, new_n2469_, new_n2468_ );
and  ( new_n2471_, new_n2470_, new_n1267_ );
or   ( new_n2472_, new_n2471_, new_n2467_ );
and  ( new_n2473_, new_n2472_, new_n2463_ );
or   ( new_n2474_, new_n2473_, new_n2462_ );
or   ( new_n2475_, new_n453_, new_n105_ );
or   ( new_n2476_, new_n459_, new_n806_ );
and  ( new_n2477_, new_n2476_, new_n2475_ );
and  ( new_n2478_, new_n2477_, new_n428_ );
and  ( new_n2479_, new_n463_, RI2b1c4342d8a0_73 );
and  ( new_n2480_, new_n451_, RI2b1c4342d828_72 );
or   ( new_n2481_, new_n2480_, new_n2479_ );
and  ( new_n2482_, new_n2481_, new_n457_ );
or   ( new_n2483_, new_n2482_, new_n2478_ );
or   ( new_n2484_, new_n934_, new_n110_ );
or   ( new_n2485_, new_n940_, new_n755_ );
and  ( new_n2486_, new_n2485_, new_n2484_ );
and  ( new_n2487_, new_n2486_, new_n913_ );
and  ( new_n2488_, new_n944_, RI2b1c4342d7b0_71 );
and  ( new_n2489_, new_n932_, RI2b1c4342d738_70 );
or   ( new_n2490_, new_n2489_, new_n2488_ );
and  ( new_n2491_, new_n2490_, new_n938_ );
or   ( new_n2492_, new_n2491_, new_n2487_ );
and  ( new_n2493_, new_n2492_, new_n2483_ );
or   ( new_n2494_, new_n2492_, new_n2483_ );
or   ( new_n2495_, new_n524_, new_n843_ );
or   ( new_n2496_, new_n528_, new_n859_ );
and  ( new_n2497_, new_n2496_, new_n2495_ );
and  ( new_n2498_, new_n2497_, new_n505_ );
and  ( new_n2499_, new_n537_, RI2b1c4342d990_75 );
and  ( new_n2500_, new_n522_, RI2b1c4342d918_74 );
or   ( new_n2501_, new_n2500_, new_n2499_ );
and  ( new_n2502_, new_n2501_, new_n533_ );
or   ( new_n2503_, new_n2502_, new_n2498_ );
and  ( new_n2504_, new_n2503_, new_n2494_ );
or   ( new_n2505_, new_n2504_, new_n2493_ );
and  ( new_n2506_, new_n2505_, new_n2474_ );
or   ( new_n2507_, new_n610_, new_n1004_ );
or   ( new_n2508_, new_n614_, new_n886_ );
and  ( new_n2509_, new_n2508_, new_n2507_ );
and  ( new_n2510_, new_n2509_, new_n590_ );
and  ( new_n2511_, new_n623_, RI2b1c4342da80_77 );
and  ( new_n2512_, new_n608_, RI2b1c4342da08_76 );
or   ( new_n2513_, new_n2512_, new_n2511_ );
and  ( new_n2514_, new_n2513_, new_n619_ );
or   ( new_n2515_, new_n2514_, new_n2510_ );
or   ( new_n2516_, new_n753_, new_n1310_ );
or   ( new_n2517_, new_n757_, new_n1002_ );
and  ( new_n2518_, new_n2517_, new_n2516_ );
and  ( new_n2519_, new_n2518_, new_n734_ );
and  ( new_n2520_, new_n766_, RI2b1c4342db70_79 );
and  ( new_n2521_, new_n751_, RI2b1c4342daf8_78 );
or   ( new_n2522_, new_n2521_, new_n2520_ );
and  ( new_n2523_, new_n2522_, new_n762_ );
or   ( new_n2524_, new_n2523_, new_n2519_ );
and  ( new_n2525_, new_n2524_, new_n2515_ );
or   ( new_n2526_, new_n2524_, new_n2515_ );
or   ( new_n2527_, new_n804_, new_n126_ );
or   ( new_n2528_, new_n808_, new_n1511_ );
and  ( new_n2529_, new_n2528_, new_n2527_ );
and  ( new_n2530_, new_n2529_, new_n785_ );
and  ( new_n2531_, new_n817_, RI2b1c4342dc60_81 );
and  ( new_n2532_, new_n802_, RI2b1c4342dbe8_80 );
or   ( new_n2533_, new_n2532_, new_n2531_ );
and  ( new_n2534_, new_n2533_, new_n813_ );
or   ( new_n2535_, new_n2534_, new_n2530_ );
and  ( new_n2536_, new_n2535_, new_n2526_ );
or   ( new_n2537_, new_n2536_, new_n2525_ );
or   ( new_n2538_, new_n2505_, new_n2474_ );
and  ( new_n2539_, new_n2538_, new_n2537_ );
or   ( new_n2540_, new_n2539_, new_n2506_ );
not  ( new_n2541_, RI2b1c4342ddc8_84 );
or   ( new_n2542_, new_n841_, new_n2541_ );
or   ( new_n2543_, new_n857_, new_n121_ );
or   ( new_n2544_, new_n861_, new_n2119_ );
and  ( new_n2545_, new_n2544_, new_n2543_ );
and  ( new_n2546_, new_n2545_, new_n842_ );
and  ( new_n2547_, new_n870_, RI2b1c4342dd50_83 );
and  ( new_n2548_, new_n855_, RI2b1c4342dcd8_82 );
or   ( new_n2549_, new_n2548_, new_n2547_ );
and  ( new_n2550_, new_n2549_, new_n866_ );
or   ( new_n2551_, new_n2550_, new_n2546_ );
and  ( new_n2552_, new_n2551_, new_n2542_ );
or   ( new_n2553_, new_n857_, new_n2119_ );
or   ( new_n2554_, new_n861_, new_n126_ );
and  ( new_n2555_, new_n2554_, new_n2553_ );
and  ( new_n2556_, new_n2555_, new_n842_ );
and  ( new_n2557_, new_n870_, RI2b1c4342dcd8_82 );
and  ( new_n2558_, new_n855_, RI2b1c4342dc60_81 );
or   ( new_n2559_, new_n2558_, new_n2557_ );
and  ( new_n2560_, new_n2559_, new_n866_ );
or   ( new_n2561_, new_n2560_, new_n2556_ );
and  ( new_n2562_, new_n2561_, new_n2552_ );
or   ( new_n2563_, new_n841_, new_n121_ );
or   ( new_n2564_, new_n2561_, new_n2552_ );
and  ( new_n2565_, new_n2564_, new_n2563_ );
or   ( new_n2566_, new_n2565_, new_n2562_ );
and  ( new_n2567_, new_n2566_, new_n2540_ );
or   ( new_n2568_, new_n2365_, new_n2210_ );
and  ( new_n2569_, new_n2568_, new_n2219_ );
and  ( new_n2570_, new_n2361_, new_n2209_ );
and  ( new_n2571_, new_n2364_, new_n2200_ );
or   ( new_n2572_, new_n2571_, new_n2570_ );
and  ( new_n2573_, new_n2572_, new_n2368_ );
or   ( new_n2574_, new_n2573_, new_n2569_ );
or   ( new_n2575_, new_n2351_, new_n2140_ );
and  ( new_n2576_, new_n2575_, new_n2149_ );
and  ( new_n2577_, new_n2347_, new_n2139_ );
and  ( new_n2578_, new_n2350_, new_n2130_ );
or   ( new_n2579_, new_n2578_, new_n2577_ );
and  ( new_n2580_, new_n2579_, new_n2354_ );
or   ( new_n2581_, new_n2580_, new_n2576_ );
and  ( new_n2582_, new_n2581_, new_n2574_ );
or   ( new_n2583_, new_n2338_, new_n2178_ );
and  ( new_n2584_, new_n2583_, new_n2187_ );
and  ( new_n2585_, new_n2334_, new_n2177_ );
and  ( new_n2586_, new_n2337_, new_n2168_ );
or   ( new_n2587_, new_n2586_, new_n2585_ );
and  ( new_n2588_, new_n2587_, new_n2341_ );
or   ( new_n2589_, new_n2588_, new_n2584_ );
or   ( new_n2590_, new_n2581_, new_n2574_ );
and  ( new_n2591_, new_n2590_, new_n2589_ );
or   ( new_n2592_, new_n2591_, new_n2582_ );
or   ( new_n2593_, new_n2566_, new_n2540_ );
and  ( new_n2594_, new_n2593_, new_n2592_ );
or   ( new_n2595_, new_n2594_, new_n2567_ );
and  ( new_n2596_, new_n2241_, new_n2234_ );
or   ( new_n2597_, new_n2596_, new_n2382_ );
and  ( new_n2598_, new_n2318_, new_n2118_ );
and  ( new_n2599_, new_n2321_, new_n2120_ );
or   ( new_n2600_, new_n2599_, new_n2598_ );
and  ( new_n2601_, new_n2600_, new_n2597_ );
or   ( new_n2602_, new_n2358_, new_n2191_ );
and  ( new_n2603_, new_n2602_, new_n2222_ );
and  ( new_n2604_, new_n2344_, new_n2152_ );
and  ( new_n2605_, new_n2357_, new_n2190_ );
or   ( new_n2606_, new_n2605_, new_n2604_ );
and  ( new_n2607_, new_n2606_, new_n2371_ );
or   ( new_n2608_, new_n2607_, new_n2603_ );
or   ( new_n2609_, new_n2600_, new_n2597_ );
and  ( new_n2610_, new_n2609_, new_n2608_ );
or   ( new_n2611_, new_n2610_, new_n2601_ );
and  ( new_n2612_, new_n2611_, new_n2595_ );
or   ( new_n2613_, new_n2611_, new_n2595_ );
or   ( new_n2614_, new_n2392_, new_n2101_ );
and  ( new_n2615_, new_n2614_, new_n2109_ );
and  ( new_n2616_, new_n2388_, new_n2100_ );
and  ( new_n2617_, new_n2391_, new_n2093_ );
or   ( new_n2618_, new_n2617_, new_n2616_ );
and  ( new_n2619_, new_n2618_, new_n2396_ );
or   ( new_n2620_, new_n2619_, new_n2615_ );
and  ( new_n2621_, new_n2620_, new_n2613_ );
or   ( new_n2622_, new_n2621_, new_n2612_ );
and  ( new_n2623_, new_n2622_, new_n2434_ );
or   ( new_n2624_, new_n2622_, new_n2434_ );
or   ( new_n2625_, new_n2399_, new_n2245_ );
and  ( new_n2626_, new_n2625_, new_n2249_ );
and  ( new_n2627_, new_n2385_, new_n2111_ );
and  ( new_n2628_, new_n2398_, new_n2244_ );
or   ( new_n2629_, new_n2628_, new_n2627_ );
and  ( new_n2630_, new_n2629_, new_n2402_ );
or   ( new_n2631_, new_n2630_, new_n2626_ );
and  ( new_n2632_, new_n2631_, new_n2624_ );
or   ( new_n2633_, new_n2632_, new_n2623_ );
or   ( new_n2634_, new_n2633_, new_n2432_ );
and  ( new_n2635_, new_n2634_, new_n2425_ );
or   ( new_n2636_, new_n2634_, new_n2425_ );
and  ( new_n2637_, new_n2633_, new_n2432_ );
and  ( new_n2638_, new_n2430_, new_n2287_ );
and  ( new_n2639_, new_n2426_, new_n2408_ );
or   ( new_n2640_, new_n2639_, new_n2638_ );
and  ( new_n2641_, new_n2313_, new_n2085_ );
and  ( new_n2642_, new_n2316_, new_n1887_ );
or   ( new_n2643_, new_n2642_, new_n2641_ );
and  ( new_n2644_, new_n2378_, new_n2241_ );
and  ( new_n2645_, new_n2381_, new_n2234_ );
or   ( new_n2646_, new_n2645_, new_n2644_ );
and  ( new_n2647_, new_n2321_, new_n2318_ );
or   ( new_n2648_, new_n2647_, new_n2121_ );
and  ( new_n2649_, new_n2648_, new_n2646_ );
and  ( new_n2650_, new_n2606_, new_n2222_ );
and  ( new_n2651_, new_n2602_, new_n2371_ );
or   ( new_n2652_, new_n2651_, new_n2650_ );
or   ( new_n2653_, new_n2648_, new_n2646_ );
and  ( new_n2654_, new_n2653_, new_n2652_ );
or   ( new_n2655_, new_n2654_, new_n2649_ );
and  ( new_n2656_, new_n2459_, new_n2334_ );
and  ( new_n2657_, new_n2451_, new_n2168_ );
or   ( new_n2658_, new_n2657_, new_n2656_ );
and  ( new_n2659_, new_n2441_, new_n1824_ );
and  ( new_n2660_, new_n2437_, new_n1717_ );
or   ( new_n2661_, new_n2660_, new_n2659_ );
and  ( new_n2662_, new_n2661_, new_n2658_ );
or   ( new_n2663_, new_n2661_, new_n2658_ );
and  ( new_n2664_, new_n2470_, new_n1355_ );
and  ( new_n2665_, new_n2466_, new_n1267_ );
or   ( new_n2666_, new_n2665_, new_n2664_ );
and  ( new_n2667_, new_n2666_, new_n2663_ );
or   ( new_n2668_, new_n2667_, new_n2662_ );
and  ( new_n2669_, new_n2490_, new_n913_ );
and  ( new_n2670_, new_n2486_, new_n938_ );
or   ( new_n2671_, new_n2670_, new_n2669_ );
and  ( new_n2672_, new_n2481_, new_n428_ );
and  ( new_n2673_, new_n2477_, new_n457_ );
or   ( new_n2674_, new_n2673_, new_n2672_ );
and  ( new_n2675_, new_n2674_, new_n2671_ );
or   ( new_n2676_, new_n2674_, new_n2671_ );
and  ( new_n2677_, new_n2501_, new_n505_ );
and  ( new_n2678_, new_n2497_, new_n533_ );
or   ( new_n2679_, new_n2678_, new_n2677_ );
and  ( new_n2680_, new_n2679_, new_n2676_ );
or   ( new_n2681_, new_n2680_, new_n2675_ );
and  ( new_n2682_, new_n2681_, new_n2668_ );
and  ( new_n2683_, new_n2513_, new_n590_ );
and  ( new_n2684_, new_n2509_, new_n619_ );
or   ( new_n2685_, new_n2684_, new_n2683_ );
and  ( new_n2686_, new_n2522_, new_n734_ );
and  ( new_n2687_, new_n2518_, new_n762_ );
or   ( new_n2688_, new_n2687_, new_n2686_ );
and  ( new_n2689_, new_n2688_, new_n2685_ );
or   ( new_n2690_, new_n2688_, new_n2685_ );
and  ( new_n2691_, new_n2533_, new_n785_ );
and  ( new_n2692_, new_n2529_, new_n813_ );
or   ( new_n2693_, new_n2692_, new_n2691_ );
and  ( new_n2694_, new_n2693_, new_n2690_ );
or   ( new_n2695_, new_n2694_, new_n2689_ );
or   ( new_n2696_, new_n2681_, new_n2668_ );
and  ( new_n2697_, new_n2696_, new_n2695_ );
or   ( new_n2698_, new_n2697_, new_n2682_ );
and  ( new_n2699_, new_n2549_, new_n842_ );
and  ( new_n2700_, new_n2545_, new_n866_ );
or   ( new_n2701_, new_n2700_, new_n2699_ );
and  ( new_n2702_, new_n720_, RI2b1c4342ddc8_84 );
or   ( new_n2703_, new_n2702_, new_n2701_ );
and  ( new_n2704_, new_n2559_, new_n842_ );
and  ( new_n2705_, new_n2555_, new_n866_ );
or   ( new_n2706_, new_n2705_, new_n2704_ );
or   ( new_n2707_, new_n2706_, new_n2703_ );
and  ( new_n2708_, new_n2706_, new_n2703_ );
and  ( new_n2709_, new_n720_, RI2b1c4342dd50_83 );
or   ( new_n2710_, new_n2709_, new_n2708_ );
and  ( new_n2711_, new_n2710_, new_n2707_ );
or   ( new_n2712_, new_n2711_, new_n2698_ );
and  ( new_n2713_, new_n2711_, new_n2698_ );
and  ( new_n2714_, new_n2572_, new_n2219_ );
and  ( new_n2715_, new_n2568_, new_n2368_ );
or   ( new_n2716_, new_n2715_, new_n2714_ );
and  ( new_n2717_, new_n2579_, new_n2149_ );
and  ( new_n2718_, new_n2575_, new_n2354_ );
or   ( new_n2719_, new_n2718_, new_n2717_ );
and  ( new_n2720_, new_n2719_, new_n2716_ );
and  ( new_n2721_, new_n2587_, new_n2187_ );
and  ( new_n2722_, new_n2583_, new_n2341_ );
or   ( new_n2723_, new_n2722_, new_n2721_ );
or   ( new_n2724_, new_n2719_, new_n2716_ );
and  ( new_n2725_, new_n2724_, new_n2723_ );
or   ( new_n2726_, new_n2725_, new_n2720_ );
or   ( new_n2727_, new_n2726_, new_n2713_ );
and  ( new_n2728_, new_n2727_, new_n2712_ );
or   ( new_n2729_, new_n2728_, new_n2655_ );
and  ( new_n2730_, new_n2728_, new_n2655_ );
and  ( new_n2731_, new_n2618_, new_n2109_ );
and  ( new_n2732_, new_n2614_, new_n2396_ );
or   ( new_n2733_, new_n2732_, new_n2731_ );
or   ( new_n2734_, new_n2733_, new_n2730_ );
and  ( new_n2735_, new_n2734_, new_n2729_ );
or   ( new_n2736_, new_n2735_, new_n2643_ );
and  ( new_n2737_, new_n2735_, new_n2643_ );
and  ( new_n2738_, new_n2629_, new_n2249_ );
and  ( new_n2739_, new_n2625_, new_n2402_ );
or   ( new_n2740_, new_n2739_, new_n2738_ );
or   ( new_n2741_, new_n2740_, new_n2737_ );
and  ( new_n2742_, new_n2741_, new_n2736_ );
and  ( new_n2743_, new_n2742_, new_n2640_ );
or   ( new_n2744_, new_n2743_, new_n2637_ );
or   ( new_n2745_, new_n2737_, new_n2623_ );
and  ( new_n2746_, new_n2745_, new_n2631_ );
and  ( new_n2747_, new_n2735_, new_n2434_ );
and  ( new_n2748_, new_n2643_, new_n2622_ );
or   ( new_n2749_, new_n2748_, new_n2747_ );
and  ( new_n2750_, new_n2749_, new_n2740_ );
or   ( new_n2751_, new_n2750_, new_n2746_ );
or   ( new_n2752_, new_n2375_, new_n2226_ );
and  ( new_n2753_, new_n2752_, new_n2242_ );
and  ( new_n2754_, new_n2374_, new_n2121_ );
and  ( new_n2755_, new_n2322_, new_n2225_ );
or   ( new_n2756_, new_n2755_, new_n2754_ );
and  ( new_n2757_, new_n2756_, new_n2382_ );
or   ( new_n2758_, new_n2757_, new_n2753_ );
or   ( new_n2759_, new_n2720_, new_n2582_ );
and  ( new_n2760_, new_n2759_, new_n2589_ );
and  ( new_n2761_, new_n2716_, new_n2581_ );
and  ( new_n2762_, new_n2719_, new_n2574_ );
or   ( new_n2763_, new_n2762_, new_n2761_ );
and  ( new_n2764_, new_n2763_, new_n2723_ );
or   ( new_n2765_, new_n2764_, new_n2760_ );
or   ( new_n2766_, new_n2708_, new_n2562_ );
and  ( new_n2767_, new_n2766_, new_n2563_ );
and  ( new_n2768_, new_n2703_, new_n2561_ );
and  ( new_n2769_, new_n2706_, new_n2552_ );
or   ( new_n2770_, new_n2769_, new_n2768_ );
and  ( new_n2771_, new_n2770_, new_n2709_ );
or   ( new_n2772_, new_n2771_, new_n2767_ );
and  ( new_n2773_, new_n2772_, new_n2765_ );
or   ( new_n2774_, new_n2682_, new_n2506_ );
and  ( new_n2775_, new_n2774_, new_n2537_ );
and  ( new_n2776_, new_n2668_, new_n2505_ );
and  ( new_n2777_, new_n2681_, new_n2474_ );
or   ( new_n2778_, new_n2777_, new_n2776_ );
and  ( new_n2779_, new_n2778_, new_n2695_ );
or   ( new_n2780_, new_n2779_, new_n2775_ );
or   ( new_n2781_, new_n2772_, new_n2765_ );
and  ( new_n2782_, new_n2781_, new_n2780_ );
or   ( new_n2783_, new_n2782_, new_n2773_ );
and  ( new_n2784_, new_n2701_, new_n2542_ );
and  ( new_n2785_, new_n2702_, new_n2551_ );
or   ( new_n2786_, new_n2785_, new_n2784_ );
or   ( new_n2787_, new_n804_, new_n2119_ );
or   ( new_n2788_, new_n808_, new_n126_ );
and  ( new_n2789_, new_n2788_, new_n2787_ );
and  ( new_n2790_, new_n2789_, new_n785_ );
and  ( new_n2791_, new_n817_, RI2b1c4342dcd8_82 );
and  ( new_n2792_, new_n802_, RI2b1c4342dc60_81 );
or   ( new_n2793_, new_n2792_, new_n2791_ );
and  ( new_n2794_, new_n2793_, new_n813_ );
or   ( new_n2795_, new_n2794_, new_n2790_ );
or   ( new_n2796_, new_n857_, new_n2541_ );
or   ( new_n2797_, new_n861_, new_n121_ );
and  ( new_n2798_, new_n2797_, new_n2796_ );
and  ( new_n2799_, new_n2798_, new_n842_ );
and  ( new_n2800_, new_n870_, RI2b1c4342ddc8_84 );
and  ( new_n2801_, new_n855_, RI2b1c4342dd50_83 );
or   ( new_n2802_, new_n2801_, new_n2800_ );
and  ( new_n2803_, new_n2802_, new_n866_ );
or   ( new_n2804_, new_n2803_, new_n2799_ );
and  ( new_n2805_, new_n2804_, new_n2795_ );
not  ( new_n2806_, RI2b1c4342de40_85 );
or   ( new_n2807_, new_n841_, new_n2806_ );
or   ( new_n2808_, new_n2804_, new_n2795_ );
and  ( new_n2809_, new_n2808_, new_n2807_ );
or   ( new_n2810_, new_n2809_, new_n2805_ );
and  ( new_n2811_, new_n2810_, new_n2786_ );
or   ( new_n2812_, new_n2689_, new_n2525_ );
and  ( new_n2813_, new_n2812_, new_n2535_ );
and  ( new_n2814_, new_n2685_, new_n2524_ );
and  ( new_n2815_, new_n2688_, new_n2515_ );
or   ( new_n2816_, new_n2815_, new_n2814_ );
and  ( new_n2817_, new_n2816_, new_n2693_ );
or   ( new_n2818_, new_n2817_, new_n2813_ );
or   ( new_n2819_, new_n2810_, new_n2786_ );
and  ( new_n2820_, new_n2819_, new_n2818_ );
or   ( new_n2821_, new_n2820_, new_n2811_ );
or   ( new_n2822_, new_n934_, new_n806_ );
or   ( new_n2823_, new_n940_, new_n110_ );
and  ( new_n2824_, new_n2823_, new_n2822_ );
and  ( new_n2825_, new_n2824_, new_n913_ );
and  ( new_n2826_, new_n944_, RI2b1c4342d828_72 );
and  ( new_n2827_, new_n932_, RI2b1c4342d7b0_71 );
or   ( new_n2828_, new_n2827_, new_n2826_ );
and  ( new_n2829_, new_n2828_, new_n938_ );
or   ( new_n2830_, new_n2829_, new_n2825_ );
or   ( new_n2831_, new_n1425_, new_n755_ );
or   ( new_n2832_, new_n1429_, new_n591_ );
and  ( new_n2833_, new_n2832_, new_n2831_ );
and  ( new_n2834_, new_n2833_, new_n1355_ );
and  ( new_n2835_, new_n1433_, RI2b1c4342d738_70 );
and  ( new_n2836_, new_n1423_, RI2b1c4342d6c0_69 );
or   ( new_n2837_, new_n2836_, new_n2835_ );
and  ( new_n2838_, new_n2837_, new_n1267_ );
or   ( new_n2839_, new_n2838_, new_n2834_ );
and  ( new_n2840_, new_n2839_, new_n2830_ );
or   ( new_n2841_, new_n453_, new_n859_ );
or   ( new_n2842_, new_n459_, new_n105_ );
and  ( new_n2843_, new_n2842_, new_n2841_ );
and  ( new_n2844_, new_n2843_, new_n428_ );
and  ( new_n2845_, new_n463_, RI2b1c4342d918_74 );
and  ( new_n2846_, new_n451_, RI2b1c4342d8a0_73 );
or   ( new_n2847_, new_n2846_, new_n2845_ );
and  ( new_n2848_, new_n2847_, new_n457_ );
or   ( new_n2849_, new_n2848_, new_n2844_ );
or   ( new_n2850_, new_n2839_, new_n2830_ );
and  ( new_n2851_, new_n2850_, new_n2849_ );
or   ( new_n2852_, new_n2851_, new_n2840_ );
xor  ( new_n2853_, new_n298_, new_n169_ );
and  ( new_n2854_, new_n2853_, new_n359_ );
xor  ( new_n2855_, RI2b1c4342c0b8_22, RI2b1c4342cfb8_54 );
and  ( new_n2856_, new_n2855_, new_n138_ );
and  ( new_n2857_, new_n2856_, new_n235_ );
or   ( new_n2858_, new_n2857_, new_n170_ );
or   ( new_n2859_, new_n2858_, new_n2854_ );
xor  ( new_n2860_, new_n301_, new_n173_ );
and  ( new_n2861_, new_n2860_, new_n357_ );
xor  ( new_n2862_, RI2b1c4342c130_23, RI2b1c4342d030_55 );
and  ( new_n2863_, new_n2862_, new_n138_ );
and  ( new_n2864_, new_n2863_, new_n233_ );
or   ( new_n2865_, new_n2864_, new_n174_ );
or   ( new_n2866_, new_n2865_, new_n2861_ );
or   ( new_n2867_, new_n2866_, new_n2859_ );
and  ( new_n2868_, new_n2867_, new_n2327_ );
or   ( new_n2869_, new_n2450_, new_n526_ );
or   ( new_n2870_, new_n2454_, new_n99_ );
and  ( new_n2871_, new_n2870_, new_n2869_ );
and  ( new_n2872_, new_n2871_, new_n2334_ );
and  ( new_n2873_, new_n2458_, RI2b1c4342d558_66 );
and  ( new_n2874_, new_n2448_, RI2b1c4342d4e0_65 );
or   ( new_n2875_, new_n2874_, new_n2873_ );
and  ( new_n2876_, new_n2875_, new_n2168_ );
or   ( new_n2877_, new_n2876_, new_n2872_ );
and  ( new_n2878_, new_n2877_, new_n2868_ );
or   ( new_n2879_, new_n1910_, new_n612_ );
or   ( new_n2880_, new_n1914_, new_n112_ );
and  ( new_n2881_, new_n2880_, new_n2879_ );
and  ( new_n2882_, new_n2881_, new_n1824_ );
and  ( new_n2883_, new_n1918_, RI2b1c4342d648_68 );
and  ( new_n2884_, new_n1908_, RI2b1c4342d5d0_67 );
or   ( new_n2885_, new_n2884_, new_n2883_ );
and  ( new_n2886_, new_n2885_, new_n1717_ );
or   ( new_n2887_, new_n2886_, new_n2882_ );
or   ( new_n2888_, new_n2877_, new_n2868_ );
and  ( new_n2889_, new_n2888_, new_n2887_ );
or   ( new_n2890_, new_n2889_, new_n2878_ );
and  ( new_n2891_, new_n2890_, new_n2852_ );
or   ( new_n2892_, new_n524_, new_n886_ );
or   ( new_n2893_, new_n528_, new_n843_ );
and  ( new_n2894_, new_n2893_, new_n2892_ );
and  ( new_n2895_, new_n2894_, new_n505_ );
and  ( new_n2896_, new_n537_, RI2b1c4342da08_76 );
and  ( new_n2897_, new_n522_, RI2b1c4342d990_75 );
or   ( new_n2898_, new_n2897_, new_n2896_ );
and  ( new_n2899_, new_n2898_, new_n533_ );
or   ( new_n2900_, new_n2899_, new_n2895_ );
or   ( new_n2901_, new_n610_, new_n1002_ );
or   ( new_n2902_, new_n614_, new_n1004_ );
and  ( new_n2903_, new_n2902_, new_n2901_ );
and  ( new_n2904_, new_n2903_, new_n590_ );
and  ( new_n2905_, new_n623_, RI2b1c4342daf8_78 );
and  ( new_n2906_, new_n608_, RI2b1c4342da80_77 );
or   ( new_n2907_, new_n2906_, new_n2905_ );
and  ( new_n2908_, new_n2907_, new_n619_ );
or   ( new_n2909_, new_n2908_, new_n2904_ );
and  ( new_n2910_, new_n2909_, new_n2900_ );
or   ( new_n2911_, new_n753_, new_n1511_ );
or   ( new_n2912_, new_n757_, new_n1310_ );
and  ( new_n2913_, new_n2912_, new_n2911_ );
and  ( new_n2914_, new_n2913_, new_n734_ );
and  ( new_n2915_, new_n766_, RI2b1c4342dbe8_80 );
and  ( new_n2916_, new_n751_, RI2b1c4342db70_79 );
or   ( new_n2917_, new_n2916_, new_n2915_ );
and  ( new_n2918_, new_n2917_, new_n762_ );
or   ( new_n2919_, new_n2918_, new_n2914_ );
or   ( new_n2920_, new_n2909_, new_n2900_ );
and  ( new_n2921_, new_n2920_, new_n2919_ );
or   ( new_n2922_, new_n2921_, new_n2910_ );
or   ( new_n2923_, new_n2890_, new_n2852_ );
and  ( new_n2924_, new_n2923_, new_n2922_ );
or   ( new_n2925_, new_n2924_, new_n2891_ );
and  ( new_n2926_, new_n2925_, new_n2821_ );
or   ( new_n2927_, new_n2675_, new_n2493_ );
and  ( new_n2928_, new_n2927_, new_n2503_ );
and  ( new_n2929_, new_n2671_, new_n2483_ );
and  ( new_n2930_, new_n2674_, new_n2492_ );
or   ( new_n2931_, new_n2930_, new_n2929_ );
and  ( new_n2932_, new_n2931_, new_n2679_ );
or   ( new_n2933_, new_n2932_, new_n2928_ );
or   ( new_n2934_, new_n2662_, new_n2462_ );
and  ( new_n2935_, new_n2934_, new_n2472_ );
and  ( new_n2936_, new_n2658_, new_n2443_ );
and  ( new_n2937_, new_n2661_, new_n2461_ );
or   ( new_n2938_, new_n2937_, new_n2936_ );
and  ( new_n2939_, new_n2938_, new_n2666_ );
or   ( new_n2940_, new_n2939_, new_n2935_ );
or   ( new_n2941_, new_n2940_, new_n2933_ );
or   ( new_n2942_, new_n2925_, new_n2821_ );
and  ( new_n2943_, new_n2942_, new_n2941_ );
or   ( new_n2944_, new_n2943_, new_n2926_ );
and  ( new_n2945_, new_n2944_, new_n2783_ );
or   ( new_n2946_, new_n2649_, new_n2601_ );
and  ( new_n2947_, new_n2946_, new_n2608_ );
and  ( new_n2948_, new_n2646_, new_n2600_ );
and  ( new_n2949_, new_n2648_, new_n2597_ );
or   ( new_n2950_, new_n2949_, new_n2948_ );
and  ( new_n2951_, new_n2950_, new_n2652_ );
or   ( new_n2952_, new_n2951_, new_n2947_ );
or   ( new_n2953_, new_n2944_, new_n2783_ );
and  ( new_n2954_, new_n2953_, new_n2952_ );
or   ( new_n2955_, new_n2954_, new_n2945_ );
and  ( new_n2956_, new_n2955_, new_n2758_ );
or   ( new_n2957_, new_n2955_, new_n2758_ );
or   ( new_n2958_, new_n2730_, new_n2612_ );
and  ( new_n2959_, new_n2958_, new_n2620_ );
and  ( new_n2960_, new_n2728_, new_n2611_ );
and  ( new_n2961_, new_n2655_, new_n2595_ );
or   ( new_n2962_, new_n2961_, new_n2960_ );
and  ( new_n2963_, new_n2962_, new_n2733_ );
or   ( new_n2964_, new_n2963_, new_n2959_ );
and  ( new_n2965_, new_n2964_, new_n2957_ );
or   ( new_n2966_, new_n2965_, new_n2956_ );
or   ( new_n2967_, new_n2966_, new_n2751_ );
or   ( new_n2968_, new_n2967_, new_n2744_ );
and  ( new_n2969_, new_n2968_, new_n2636_ );
or   ( new_n2970_, new_n2969_, new_n2635_ );
or   ( new_n2971_, new_n2970_, new_n2310_ );
and  ( new_n2972_, new_n2971_, new_n2308_ );
and  ( new_n2973_, new_n2966_, new_n2751_ );
and  ( new_n2974_, new_n2749_, new_n2631_ );
and  ( new_n2975_, new_n2745_, new_n2740_ );
or   ( new_n2976_, new_n2975_, new_n2974_ );
and  ( new_n2977_, new_n2756_, new_n2242_ );
and  ( new_n2978_, new_n2752_, new_n2382_ );
or   ( new_n2979_, new_n2978_, new_n2977_ );
and  ( new_n2980_, new_n2763_, new_n2589_ );
and  ( new_n2981_, new_n2759_, new_n2723_ );
or   ( new_n2982_, new_n2981_, new_n2980_ );
and  ( new_n2983_, new_n2770_, new_n2563_ );
and  ( new_n2984_, new_n2766_, new_n2709_ );
or   ( new_n2985_, new_n2984_, new_n2983_ );
and  ( new_n2986_, new_n2985_, new_n2982_ );
and  ( new_n2987_, new_n2778_, new_n2537_ );
and  ( new_n2988_, new_n2774_, new_n2695_ );
or   ( new_n2989_, new_n2988_, new_n2987_ );
or   ( new_n2990_, new_n2985_, new_n2982_ );
and  ( new_n2991_, new_n2990_, new_n2989_ );
or   ( new_n2992_, new_n2991_, new_n2986_ );
not  ( new_n2993_, new_n233_ );
nor  ( new_n2994_, new_n2862_, new_n2993_ );
and  ( new_n2995_, new_n2862_, new_n357_ );
or   ( new_n2996_, new_n2995_, new_n2994_ );
and  ( new_n2997_, new_n2996_, new_n301_ );
not  ( new_n2998_, new_n235_ );
nor  ( new_n2999_, new_n2855_, new_n2998_ );
and  ( new_n3000_, new_n2855_, new_n359_ );
or   ( new_n3001_, new_n3000_, new_n2999_ );
and  ( new_n3002_, new_n3001_, new_n298_ );
and  ( new_n3003_, new_n3002_, new_n2997_ );
or   ( new_n3004_, new_n3003_, new_n2166_ );
and  ( new_n3005_, new_n2875_, new_n2334_ );
and  ( new_n3006_, new_n2871_, new_n2168_ );
or   ( new_n3007_, new_n3006_, new_n3005_ );
and  ( new_n3008_, new_n3007_, new_n3004_ );
and  ( new_n3009_, new_n2885_, new_n1824_ );
and  ( new_n3010_, new_n2881_, new_n1717_ );
or   ( new_n3011_, new_n3010_, new_n3009_ );
or   ( new_n3012_, new_n3007_, new_n3004_ );
and  ( new_n3013_, new_n3012_, new_n3011_ );
or   ( new_n3014_, new_n3013_, new_n3008_ );
and  ( new_n3015_, new_n2837_, new_n1355_ );
and  ( new_n3016_, new_n2833_, new_n1267_ );
or   ( new_n3017_, new_n3016_, new_n3015_ );
and  ( new_n3018_, new_n2828_, new_n913_ );
and  ( new_n3019_, new_n2824_, new_n938_ );
or   ( new_n3020_, new_n3019_, new_n3018_ );
and  ( new_n3021_, new_n3020_, new_n3017_ );
and  ( new_n3022_, new_n2847_, new_n428_ );
and  ( new_n3023_, new_n2843_, new_n457_ );
or   ( new_n3024_, new_n3023_, new_n3022_ );
or   ( new_n3025_, new_n3020_, new_n3017_ );
and  ( new_n3026_, new_n3025_, new_n3024_ );
or   ( new_n3027_, new_n3026_, new_n3021_ );
and  ( new_n3028_, new_n3027_, new_n3014_ );
and  ( new_n3029_, new_n2898_, new_n505_ );
and  ( new_n3030_, new_n2894_, new_n533_ );
or   ( new_n3031_, new_n3030_, new_n3029_ );
and  ( new_n3032_, new_n2907_, new_n590_ );
and  ( new_n3033_, new_n2903_, new_n619_ );
or   ( new_n3034_, new_n3033_, new_n3032_ );
and  ( new_n3035_, new_n3034_, new_n3031_ );
and  ( new_n3036_, new_n2917_, new_n734_ );
and  ( new_n3037_, new_n2913_, new_n762_ );
or   ( new_n3038_, new_n3037_, new_n3036_ );
or   ( new_n3039_, new_n3034_, new_n3031_ );
and  ( new_n3040_, new_n3039_, new_n3038_ );
or   ( new_n3041_, new_n3040_, new_n3035_ );
or   ( new_n3042_, new_n3027_, new_n3014_ );
and  ( new_n3043_, new_n3042_, new_n3041_ );
or   ( new_n3044_, new_n3043_, new_n3028_ );
and  ( new_n3045_, new_n2702_, new_n2701_ );
or   ( new_n3046_, new_n3045_, new_n2552_ );
and  ( new_n3047_, new_n2793_, new_n785_ );
and  ( new_n3048_, new_n2789_, new_n813_ );
or   ( new_n3049_, new_n3048_, new_n3047_ );
and  ( new_n3050_, new_n2802_, new_n842_ );
and  ( new_n3051_, new_n2798_, new_n866_ );
or   ( new_n3052_, new_n3051_, new_n3050_ );
or   ( new_n3053_, new_n3052_, new_n3049_ );
and  ( new_n3054_, new_n3052_, new_n3049_ );
and  ( new_n3055_, new_n720_, RI2b1c4342de40_85 );
or   ( new_n3056_, new_n3055_, new_n3054_ );
and  ( new_n3057_, new_n3056_, new_n3053_ );
or   ( new_n3058_, new_n3057_, new_n3046_ );
and  ( new_n3059_, new_n3057_, new_n3046_ );
and  ( new_n3060_, new_n2816_, new_n2535_ );
and  ( new_n3061_, new_n2812_, new_n2693_ );
or   ( new_n3062_, new_n3061_, new_n3060_ );
or   ( new_n3063_, new_n3062_, new_n3059_ );
and  ( new_n3064_, new_n3063_, new_n3058_ );
or   ( new_n3065_, new_n3064_, new_n3044_ );
and  ( new_n3066_, new_n2931_, new_n2503_ );
and  ( new_n3067_, new_n2927_, new_n2679_ );
or   ( new_n3068_, new_n3067_, new_n3066_ );
and  ( new_n3069_, new_n2938_, new_n2472_ );
and  ( new_n3070_, new_n2934_, new_n2666_ );
or   ( new_n3071_, new_n3070_, new_n3069_ );
and  ( new_n3072_, new_n3071_, new_n3068_ );
and  ( new_n3073_, new_n3064_, new_n3044_ );
or   ( new_n3074_, new_n3073_, new_n3072_ );
and  ( new_n3075_, new_n3074_, new_n3065_ );
or   ( new_n3076_, new_n3075_, new_n2992_ );
and  ( new_n3077_, new_n3075_, new_n2992_ );
and  ( new_n3078_, new_n2950_, new_n2608_ );
and  ( new_n3079_, new_n2946_, new_n2652_ );
or   ( new_n3080_, new_n3079_, new_n3078_ );
or   ( new_n3081_, new_n3080_, new_n3077_ );
and  ( new_n3082_, new_n3081_, new_n3076_ );
or   ( new_n3083_, new_n3082_, new_n2979_ );
and  ( new_n3084_, new_n3082_, new_n2979_ );
and  ( new_n3085_, new_n2962_, new_n2620_ );
and  ( new_n3086_, new_n2958_, new_n2733_ );
or   ( new_n3087_, new_n3086_, new_n3085_ );
or   ( new_n3088_, new_n3087_, new_n3084_ );
and  ( new_n3089_, new_n3088_, new_n3083_ );
and  ( new_n3090_, new_n3089_, new_n2976_ );
or   ( new_n3091_, new_n3090_, new_n2973_ );
or   ( new_n3092_, new_n3084_, new_n2956_ );
and  ( new_n3093_, new_n3092_, new_n2964_ );
and  ( new_n3094_, new_n3082_, new_n2758_ );
and  ( new_n3095_, new_n2979_, new_n2955_ );
or   ( new_n3096_, new_n3095_, new_n3094_ );
and  ( new_n3097_, new_n3096_, new_n3087_ );
or   ( new_n3098_, new_n3097_, new_n3093_ );
or   ( new_n3099_, new_n2713_, new_n2567_ );
and  ( new_n3100_, new_n3099_, new_n2592_ );
and  ( new_n3101_, new_n2698_, new_n2566_ );
and  ( new_n3102_, new_n2711_, new_n2540_ );
or   ( new_n3103_, new_n3102_, new_n3101_ );
and  ( new_n3104_, new_n3103_, new_n2726_ );
or   ( new_n3105_, new_n3104_, new_n3100_ );
and  ( new_n3106_, new_n3002_, new_n2327_ );
and  ( new_n3107_, new_n2859_, new_n2166_ );
and  ( new_n3108_, new_n3002_, new_n2866_ );
and  ( new_n3109_, new_n2997_, new_n2859_ );
or   ( new_n3110_, new_n3109_, new_n3108_ );
or   ( new_n3111_, new_n3110_, new_n3107_ );
or   ( new_n3112_, new_n3111_, new_n3106_ );
or   ( new_n3113_, new_n3112_, new_n99_ );
and  ( new_n3114_, new_n3113_, new_n3004_ );
and  ( new_n3115_, new_n2866_, new_n2859_ );
or   ( new_n3116_, new_n3115_, new_n3003_ );
and  ( new_n3117_, new_n2859_, new_n2327_ );
and  ( new_n3118_, new_n3002_, new_n2166_ );
or   ( new_n3119_, new_n3118_, new_n3117_ );
and  ( new_n3120_, new_n3119_, new_n3116_ );
and  ( new_n3121_, new_n3120_, RI2b1c4342d4e0_65 );
and  ( new_n3122_, new_n3121_, new_n2868_ );
or   ( new_n3123_, new_n3122_, new_n3114_ );
or   ( new_n3124_, new_n2450_, new_n112_ );
or   ( new_n3125_, new_n2454_, new_n526_ );
and  ( new_n3126_, new_n3125_, new_n3124_ );
and  ( new_n3127_, new_n3126_, new_n2334_ );
and  ( new_n3128_, new_n2458_, RI2b1c4342d5d0_67 );
and  ( new_n3129_, new_n2448_, RI2b1c4342d558_66 );
or   ( new_n3130_, new_n3129_, new_n3128_ );
and  ( new_n3131_, new_n3130_, new_n2168_ );
or   ( new_n3132_, new_n3131_, new_n3127_ );
and  ( new_n3133_, new_n3132_, new_n3123_ );
or   ( new_n3134_, new_n3132_, new_n3123_ );
or   ( new_n3135_, new_n1910_, new_n591_ );
or   ( new_n3136_, new_n1914_, new_n612_ );
and  ( new_n3137_, new_n3136_, new_n3135_ );
and  ( new_n3138_, new_n3137_, new_n1824_ );
and  ( new_n3139_, new_n1918_, RI2b1c4342d6c0_69 );
and  ( new_n3140_, new_n1908_, RI2b1c4342d648_68 );
or   ( new_n3141_, new_n3140_, new_n3139_ );
and  ( new_n3142_, new_n3141_, new_n1717_ );
or   ( new_n3143_, new_n3142_, new_n3138_ );
and  ( new_n3144_, new_n3143_, new_n3134_ );
or   ( new_n3145_, new_n3144_, new_n3133_ );
or   ( new_n3146_, new_n1425_, new_n110_ );
or   ( new_n3147_, new_n1429_, new_n755_ );
and  ( new_n3148_, new_n3147_, new_n3146_ );
and  ( new_n3149_, new_n3148_, new_n1355_ );
and  ( new_n3150_, new_n1433_, RI2b1c4342d7b0_71 );
and  ( new_n3151_, new_n1423_, RI2b1c4342d738_70 );
or   ( new_n3152_, new_n3151_, new_n3150_ );
and  ( new_n3153_, new_n3152_, new_n1267_ );
or   ( new_n3154_, new_n3153_, new_n3149_ );
or   ( new_n3155_, new_n934_, new_n105_ );
or   ( new_n3156_, new_n940_, new_n806_ );
and  ( new_n3157_, new_n3156_, new_n3155_ );
and  ( new_n3158_, new_n3157_, new_n913_ );
and  ( new_n3159_, new_n944_, RI2b1c4342d8a0_73 );
and  ( new_n3160_, new_n932_, RI2b1c4342d828_72 );
or   ( new_n3161_, new_n3160_, new_n3159_ );
and  ( new_n3162_, new_n3161_, new_n938_ );
or   ( new_n3163_, new_n3162_, new_n3158_ );
and  ( new_n3164_, new_n3163_, new_n3154_ );
or   ( new_n3165_, new_n3163_, new_n3154_ );
or   ( new_n3166_, new_n453_, new_n843_ );
or   ( new_n3167_, new_n459_, new_n859_ );
and  ( new_n3168_, new_n3167_, new_n3166_ );
and  ( new_n3169_, new_n3168_, new_n428_ );
and  ( new_n3170_, new_n463_, RI2b1c4342d990_75 );
and  ( new_n3171_, new_n451_, RI2b1c4342d918_74 );
or   ( new_n3172_, new_n3171_, new_n3170_ );
and  ( new_n3173_, new_n3172_, new_n457_ );
or   ( new_n3174_, new_n3173_, new_n3169_ );
and  ( new_n3175_, new_n3174_, new_n3165_ );
or   ( new_n3176_, new_n3175_, new_n3164_ );
and  ( new_n3177_, new_n3176_, new_n3145_ );
or   ( new_n3178_, new_n3176_, new_n3145_ );
or   ( new_n3179_, new_n524_, new_n1004_ );
or   ( new_n3180_, new_n528_, new_n886_ );
and  ( new_n3181_, new_n3180_, new_n3179_ );
and  ( new_n3182_, new_n3181_, new_n505_ );
and  ( new_n3183_, new_n537_, RI2b1c4342da80_77 );
and  ( new_n3184_, new_n522_, RI2b1c4342da08_76 );
or   ( new_n3185_, new_n3184_, new_n3183_ );
and  ( new_n3186_, new_n3185_, new_n533_ );
or   ( new_n3187_, new_n3186_, new_n3182_ );
or   ( new_n3188_, new_n610_, new_n1310_ );
or   ( new_n3189_, new_n614_, new_n1002_ );
and  ( new_n3190_, new_n3189_, new_n3188_ );
and  ( new_n3191_, new_n3190_, new_n590_ );
and  ( new_n3192_, new_n623_, RI2b1c4342db70_79 );
and  ( new_n3193_, new_n608_, RI2b1c4342daf8_78 );
or   ( new_n3194_, new_n3193_, new_n3192_ );
and  ( new_n3195_, new_n3194_, new_n619_ );
or   ( new_n3196_, new_n3195_, new_n3191_ );
and  ( new_n3197_, new_n3196_, new_n3187_ );
or   ( new_n3198_, new_n3196_, new_n3187_ );
or   ( new_n3199_, new_n753_, new_n126_ );
or   ( new_n3200_, new_n757_, new_n1511_ );
and  ( new_n3201_, new_n3200_, new_n3199_ );
and  ( new_n3202_, new_n3201_, new_n734_ );
and  ( new_n3203_, new_n766_, RI2b1c4342dc60_81 );
and  ( new_n3204_, new_n751_, RI2b1c4342dbe8_80 );
or   ( new_n3205_, new_n3204_, new_n3203_ );
and  ( new_n3206_, new_n3205_, new_n762_ );
or   ( new_n3207_, new_n3206_, new_n3202_ );
and  ( new_n3208_, new_n3207_, new_n3198_ );
or   ( new_n3209_, new_n3208_, new_n3197_ );
and  ( new_n3210_, new_n3209_, new_n3178_ );
or   ( new_n3211_, new_n3210_, new_n3177_ );
or   ( new_n3212_, new_n3054_, new_n2805_ );
and  ( new_n3213_, new_n3212_, new_n2807_ );
and  ( new_n3214_, new_n3049_, new_n2804_ );
and  ( new_n3215_, new_n3052_, new_n2795_ );
or   ( new_n3216_, new_n3215_, new_n3214_ );
and  ( new_n3217_, new_n3216_, new_n3055_ );
or   ( new_n3218_, new_n3217_, new_n3213_ );
or   ( new_n3219_, new_n804_, new_n121_ );
or   ( new_n3220_, new_n808_, new_n2119_ );
and  ( new_n3221_, new_n3220_, new_n3219_ );
and  ( new_n3222_, new_n3221_, new_n785_ );
and  ( new_n3223_, new_n817_, RI2b1c4342dd50_83 );
and  ( new_n3224_, new_n802_, RI2b1c4342dcd8_82 );
or   ( new_n3225_, new_n3224_, new_n3223_ );
and  ( new_n3226_, new_n3225_, new_n813_ );
or   ( new_n3227_, new_n3226_, new_n3222_ );
or   ( new_n3228_, new_n857_, new_n2806_ );
or   ( new_n3229_, new_n861_, new_n2541_ );
and  ( new_n3230_, new_n3229_, new_n3228_ );
and  ( new_n3231_, new_n3230_, new_n842_ );
and  ( new_n3232_, new_n870_, RI2b1c4342de40_85 );
and  ( new_n3233_, new_n855_, RI2b1c4342ddc8_84 );
or   ( new_n3234_, new_n3233_, new_n3232_ );
and  ( new_n3235_, new_n3234_, new_n866_ );
or   ( new_n3236_, new_n3235_, new_n3231_ );
and  ( new_n3237_, new_n3236_, new_n3227_ );
or   ( new_n3238_, new_n3236_, new_n3227_ );
not  ( new_n3239_, RI2b1c4342deb8_86 );
or   ( new_n3240_, new_n841_, new_n3239_ );
and  ( new_n3241_, new_n3240_, new_n3238_ );
or   ( new_n3242_, new_n3241_, new_n3237_ );
and  ( new_n3243_, new_n3242_, new_n3218_ );
or   ( new_n3244_, new_n3242_, new_n3218_ );
or   ( new_n3245_, new_n3035_, new_n2910_ );
and  ( new_n3246_, new_n3245_, new_n2919_ );
and  ( new_n3247_, new_n3031_, new_n2909_ );
and  ( new_n3248_, new_n3034_, new_n2900_ );
or   ( new_n3249_, new_n3248_, new_n3247_ );
and  ( new_n3250_, new_n3249_, new_n3038_ );
or   ( new_n3251_, new_n3250_, new_n3246_ );
and  ( new_n3252_, new_n3251_, new_n3244_ );
or   ( new_n3253_, new_n3252_, new_n3243_ );
and  ( new_n3254_, new_n3253_, new_n3211_ );
or   ( new_n3255_, new_n3253_, new_n3211_ );
or   ( new_n3256_, new_n3021_, new_n2840_ );
and  ( new_n3257_, new_n3256_, new_n2849_ );
and  ( new_n3258_, new_n3017_, new_n2830_ );
and  ( new_n3259_, new_n3020_, new_n2839_ );
or   ( new_n3260_, new_n3259_, new_n3258_ );
and  ( new_n3261_, new_n3260_, new_n3024_ );
or   ( new_n3262_, new_n3261_, new_n3257_ );
or   ( new_n3263_, new_n3008_, new_n2878_ );
and  ( new_n3264_, new_n3263_, new_n2887_ );
and  ( new_n3265_, new_n3004_, new_n2877_ );
and  ( new_n3266_, new_n3007_, new_n2868_ );
or   ( new_n3267_, new_n3266_, new_n3265_ );
and  ( new_n3268_, new_n3267_, new_n3011_ );
or   ( new_n3269_, new_n3268_, new_n3264_ );
or   ( new_n3270_, new_n3269_, new_n3262_ );
and  ( new_n3271_, new_n3270_, new_n3255_ );
or   ( new_n3272_, new_n3271_, new_n3254_ );
and  ( new_n3273_, new_n2940_, new_n2933_ );
or   ( new_n3274_, new_n3273_, new_n3072_ );
or   ( new_n3275_, new_n3059_, new_n2811_ );
and  ( new_n3276_, new_n3275_, new_n2818_ );
and  ( new_n3277_, new_n3057_, new_n2786_ );
and  ( new_n3278_, new_n3046_, new_n2810_ );
or   ( new_n3279_, new_n3278_, new_n3277_ );
and  ( new_n3280_, new_n3279_, new_n3062_ );
or   ( new_n3281_, new_n3280_, new_n3276_ );
and  ( new_n3282_, new_n3281_, new_n3274_ );
or   ( new_n3283_, new_n3281_, new_n3274_ );
or   ( new_n3284_, new_n3028_, new_n2891_ );
and  ( new_n3285_, new_n3284_, new_n2922_ );
and  ( new_n3286_, new_n3014_, new_n2852_ );
and  ( new_n3287_, new_n3027_, new_n2890_ );
or   ( new_n3288_, new_n3287_, new_n3286_ );
and  ( new_n3289_, new_n3288_, new_n3041_ );
or   ( new_n3290_, new_n3289_, new_n3285_ );
and  ( new_n3291_, new_n3290_, new_n3283_ );
or   ( new_n3292_, new_n3291_, new_n3282_ );
and  ( new_n3293_, new_n3292_, new_n3272_ );
or   ( new_n3294_, new_n2986_, new_n2773_ );
and  ( new_n3295_, new_n3294_, new_n2780_ );
and  ( new_n3296_, new_n2982_, new_n2772_ );
and  ( new_n3297_, new_n2985_, new_n2765_ );
or   ( new_n3298_, new_n3297_, new_n3296_ );
and  ( new_n3299_, new_n3298_, new_n2989_ );
or   ( new_n3300_, new_n3299_, new_n3295_ );
or   ( new_n3301_, new_n3292_, new_n3272_ );
and  ( new_n3302_, new_n3301_, new_n3300_ );
or   ( new_n3303_, new_n3302_, new_n3293_ );
and  ( new_n3304_, new_n3303_, new_n3105_ );
or   ( new_n3305_, new_n3077_, new_n2945_ );
and  ( new_n3306_, new_n3305_, new_n2952_ );
and  ( new_n3307_, new_n3075_, new_n2783_ );
and  ( new_n3308_, new_n2992_, new_n2944_ );
or   ( new_n3309_, new_n3308_, new_n3307_ );
and  ( new_n3310_, new_n3309_, new_n3080_ );
or   ( new_n3311_, new_n3310_, new_n3306_ );
or   ( new_n3312_, new_n3303_, new_n3105_ );
and  ( new_n3313_, new_n3312_, new_n3311_ );
or   ( new_n3314_, new_n3313_, new_n3304_ );
or   ( new_n3315_, new_n3314_, new_n3098_ );
and  ( new_n3316_, new_n3315_, new_n3091_ );
or   ( new_n3317_, new_n3315_, new_n3091_ );
and  ( new_n3318_, new_n3314_, new_n3098_ );
and  ( new_n3319_, new_n3096_, new_n2964_ );
and  ( new_n3320_, new_n3092_, new_n3087_ );
or   ( new_n3321_, new_n3320_, new_n3319_ );
and  ( new_n3322_, new_n3103_, new_n2592_ );
and  ( new_n3323_, new_n3099_, new_n2726_ );
or   ( new_n3324_, new_n3323_, new_n3322_ );
and  ( new_n3325_, new_n3068_, new_n2940_ );
and  ( new_n3326_, new_n3071_, new_n2933_ );
or   ( new_n3327_, new_n3326_, new_n3325_ );
and  ( new_n3328_, new_n3279_, new_n2818_ );
and  ( new_n3329_, new_n3275_, new_n3062_ );
or   ( new_n3330_, new_n3329_, new_n3328_ );
and  ( new_n3331_, new_n3330_, new_n3327_ );
or   ( new_n3332_, new_n3330_, new_n3327_ );
and  ( new_n3333_, new_n3288_, new_n2922_ );
and  ( new_n3334_, new_n3284_, new_n3041_ );
or   ( new_n3335_, new_n3334_, new_n3333_ );
and  ( new_n3336_, new_n3335_, new_n3332_ );
or   ( new_n3337_, new_n3336_, new_n3331_ );
and  ( new_n3338_, new_n3121_, new_n3004_ );
and  ( new_n3339_, new_n3113_, new_n2868_ );
or   ( new_n3340_, new_n3339_, new_n3338_ );
and  ( new_n3341_, new_n3130_, new_n2334_ );
and  ( new_n3342_, new_n3126_, new_n2168_ );
or   ( new_n3343_, new_n3342_, new_n3341_ );
and  ( new_n3344_, new_n3343_, new_n3340_ );
or   ( new_n3345_, new_n3343_, new_n3340_ );
and  ( new_n3346_, new_n3141_, new_n1824_ );
and  ( new_n3347_, new_n3137_, new_n1717_ );
or   ( new_n3348_, new_n3347_, new_n3346_ );
and  ( new_n3349_, new_n3348_, new_n3345_ );
or   ( new_n3350_, new_n3349_, new_n3344_ );
and  ( new_n3351_, new_n3152_, new_n1355_ );
and  ( new_n3352_, new_n3148_, new_n1267_ );
or   ( new_n3353_, new_n3352_, new_n3351_ );
and  ( new_n3354_, new_n3161_, new_n913_ );
and  ( new_n3355_, new_n3157_, new_n938_ );
or   ( new_n3356_, new_n3355_, new_n3354_ );
and  ( new_n3357_, new_n3356_, new_n3353_ );
or   ( new_n3358_, new_n3356_, new_n3353_ );
and  ( new_n3359_, new_n3172_, new_n428_ );
and  ( new_n3360_, new_n3168_, new_n457_ );
or   ( new_n3361_, new_n3360_, new_n3359_ );
and  ( new_n3362_, new_n3361_, new_n3358_ );
or   ( new_n3363_, new_n3362_, new_n3357_ );
and  ( new_n3364_, new_n3363_, new_n3350_ );
or   ( new_n3365_, new_n3363_, new_n3350_ );
and  ( new_n3366_, new_n3185_, new_n505_ );
and  ( new_n3367_, new_n3181_, new_n533_ );
or   ( new_n3368_, new_n3367_, new_n3366_ );
and  ( new_n3369_, new_n3194_, new_n590_ );
and  ( new_n3370_, new_n3190_, new_n619_ );
or   ( new_n3371_, new_n3370_, new_n3369_ );
and  ( new_n3372_, new_n3371_, new_n3368_ );
or   ( new_n3373_, new_n3371_, new_n3368_ );
and  ( new_n3374_, new_n3205_, new_n734_ );
and  ( new_n3375_, new_n3201_, new_n762_ );
or   ( new_n3376_, new_n3375_, new_n3374_ );
and  ( new_n3377_, new_n3376_, new_n3373_ );
or   ( new_n3378_, new_n3377_, new_n3372_ );
and  ( new_n3379_, new_n3378_, new_n3365_ );
or   ( new_n3380_, new_n3379_, new_n3364_ );
and  ( new_n3381_, new_n3216_, new_n2807_ );
and  ( new_n3382_, new_n3212_, new_n3055_ );
or   ( new_n3383_, new_n3382_, new_n3381_ );
and  ( new_n3384_, new_n3225_, new_n785_ );
and  ( new_n3385_, new_n3221_, new_n813_ );
or   ( new_n3386_, new_n3385_, new_n3384_ );
and  ( new_n3387_, new_n3234_, new_n842_ );
and  ( new_n3388_, new_n3230_, new_n866_ );
or   ( new_n3389_, new_n3388_, new_n3387_ );
or   ( new_n3390_, new_n3389_, new_n3386_ );
and  ( new_n3391_, new_n3389_, new_n3386_ );
and  ( new_n3392_, new_n720_, RI2b1c4342deb8_86 );
or   ( new_n3393_, new_n3392_, new_n3391_ );
and  ( new_n3394_, new_n3393_, new_n3390_ );
or   ( new_n3395_, new_n3394_, new_n3383_ );
and  ( new_n3396_, new_n3394_, new_n3383_ );
and  ( new_n3397_, new_n3249_, new_n2919_ );
and  ( new_n3398_, new_n3245_, new_n3038_ );
or   ( new_n3399_, new_n3398_, new_n3397_ );
or   ( new_n3400_, new_n3399_, new_n3396_ );
and  ( new_n3401_, new_n3400_, new_n3395_ );
or   ( new_n3402_, new_n3401_, new_n3380_ );
and  ( new_n3403_, new_n3401_, new_n3380_ );
and  ( new_n3404_, new_n3260_, new_n2849_ );
and  ( new_n3405_, new_n3256_, new_n3024_ );
or   ( new_n3406_, new_n3405_, new_n3404_ );
and  ( new_n3407_, new_n3267_, new_n2887_ );
and  ( new_n3408_, new_n3263_, new_n3011_ );
or   ( new_n3409_, new_n3408_, new_n3407_ );
and  ( new_n3410_, new_n3409_, new_n3406_ );
or   ( new_n3411_, new_n3410_, new_n3403_ );
and  ( new_n3412_, new_n3411_, new_n3402_ );
or   ( new_n3413_, new_n3412_, new_n3337_ );
and  ( new_n3414_, new_n3412_, new_n3337_ );
and  ( new_n3415_, new_n3298_, new_n2780_ );
and  ( new_n3416_, new_n3294_, new_n2989_ );
or   ( new_n3417_, new_n3416_, new_n3415_ );
or   ( new_n3418_, new_n3417_, new_n3414_ );
and  ( new_n3419_, new_n3418_, new_n3413_ );
or   ( new_n3420_, new_n3419_, new_n3324_ );
and  ( new_n3421_, new_n3419_, new_n3324_ );
and  ( new_n3422_, new_n3309_, new_n2952_ );
and  ( new_n3423_, new_n3305_, new_n3080_ );
or   ( new_n3424_, new_n3423_, new_n3422_ );
or   ( new_n3425_, new_n3424_, new_n3421_ );
and  ( new_n3426_, new_n3425_, new_n3420_ );
and  ( new_n3427_, new_n3426_, new_n3321_ );
or   ( new_n3428_, new_n3427_, new_n3318_ );
or   ( new_n3429_, new_n3421_, new_n3304_ );
and  ( new_n3430_, new_n3429_, new_n3311_ );
and  ( new_n3431_, new_n3419_, new_n3105_ );
and  ( new_n3432_, new_n3324_, new_n3303_ );
or   ( new_n3433_, new_n3432_, new_n3431_ );
and  ( new_n3434_, new_n3433_, new_n3424_ );
or   ( new_n3435_, new_n3434_, new_n3430_ );
or   ( new_n3436_, new_n3073_, new_n2926_ );
and  ( new_n3437_, new_n3436_, new_n2941_ );
and  ( new_n3438_, new_n3044_, new_n2821_ );
and  ( new_n3439_, new_n3064_, new_n2925_ );
or   ( new_n3440_, new_n3439_, new_n3438_ );
and  ( new_n3441_, new_n3440_, new_n3072_ );
or   ( new_n3442_, new_n3441_, new_n3437_ );
and  ( new_n3443_, new_n3269_, new_n3262_ );
or   ( new_n3444_, new_n3443_, new_n3410_ );
or   ( new_n3445_, new_n3396_, new_n3243_ );
and  ( new_n3446_, new_n3445_, new_n3251_ );
and  ( new_n3447_, new_n3394_, new_n3218_ );
and  ( new_n3448_, new_n3383_, new_n3242_ );
or   ( new_n3449_, new_n3448_, new_n3447_ );
and  ( new_n3450_, new_n3449_, new_n3399_ );
or   ( new_n3451_, new_n3450_, new_n3446_ );
and  ( new_n3452_, new_n3451_, new_n3444_ );
or   ( new_n3453_, new_n3451_, new_n3444_ );
or   ( new_n3454_, new_n3364_, new_n3177_ );
and  ( new_n3455_, new_n3454_, new_n3209_ );
and  ( new_n3456_, new_n3350_, new_n3176_ );
and  ( new_n3457_, new_n3363_, new_n3145_ );
or   ( new_n3458_, new_n3457_, new_n3456_ );
and  ( new_n3459_, new_n3458_, new_n3378_ );
or   ( new_n3460_, new_n3459_, new_n3455_ );
and  ( new_n3461_, new_n3460_, new_n3453_ );
or   ( new_n3462_, new_n3461_, new_n3452_ );
or   ( new_n3463_, new_n3391_, new_n3237_ );
and  ( new_n3464_, new_n3463_, new_n3240_ );
and  ( new_n3465_, new_n3386_, new_n3236_ );
and  ( new_n3466_, new_n3389_, new_n3227_ );
or   ( new_n3467_, new_n3466_, new_n3465_ );
and  ( new_n3468_, new_n3467_, new_n3392_ );
or   ( new_n3469_, new_n3468_, new_n3464_ );
or   ( new_n3470_, new_n753_, new_n2119_ );
or   ( new_n3471_, new_n757_, new_n126_ );
and  ( new_n3472_, new_n3471_, new_n3470_ );
and  ( new_n3473_, new_n3472_, new_n734_ );
and  ( new_n3474_, new_n766_, RI2b1c4342dcd8_82 );
and  ( new_n3475_, new_n751_, RI2b1c4342dc60_81 );
or   ( new_n3476_, new_n3475_, new_n3474_ );
and  ( new_n3477_, new_n3476_, new_n762_ );
or   ( new_n3478_, new_n3477_, new_n3473_ );
or   ( new_n3479_, new_n804_, new_n2541_ );
or   ( new_n3480_, new_n808_, new_n121_ );
and  ( new_n3481_, new_n3480_, new_n3479_ );
and  ( new_n3482_, new_n3481_, new_n785_ );
and  ( new_n3483_, new_n817_, RI2b1c4342ddc8_84 );
and  ( new_n3484_, new_n802_, RI2b1c4342dd50_83 );
or   ( new_n3485_, new_n3484_, new_n3483_ );
and  ( new_n3486_, new_n3485_, new_n813_ );
or   ( new_n3487_, new_n3486_, new_n3482_ );
and  ( new_n3488_, new_n3487_, new_n3478_ );
or   ( new_n3489_, new_n3487_, new_n3478_ );
or   ( new_n3490_, new_n857_, new_n3239_ );
or   ( new_n3491_, new_n861_, new_n2806_ );
and  ( new_n3492_, new_n3491_, new_n3490_ );
and  ( new_n3493_, new_n3492_, new_n842_ );
and  ( new_n3494_, new_n870_, RI2b1c4342deb8_86 );
and  ( new_n3495_, new_n855_, RI2b1c4342de40_85 );
or   ( new_n3496_, new_n3495_, new_n3494_ );
and  ( new_n3497_, new_n3496_, new_n866_ );
or   ( new_n3498_, new_n3497_, new_n3493_ );
and  ( new_n3499_, new_n3498_, new_n3489_ );
or   ( new_n3500_, new_n3499_, new_n3488_ );
and  ( new_n3501_, new_n3500_, new_n3469_ );
or   ( new_n3502_, new_n1910_, new_n755_ );
or   ( new_n3503_, new_n1914_, new_n591_ );
and  ( new_n3504_, new_n3503_, new_n3502_ );
and  ( new_n3505_, new_n3504_, new_n1824_ );
and  ( new_n3506_, new_n1918_, RI2b1c4342d738_70 );
and  ( new_n3507_, new_n1908_, RI2b1c4342d6c0_69 );
or   ( new_n3508_, new_n3507_, new_n3506_ );
and  ( new_n3509_, new_n3508_, new_n1717_ );
or   ( new_n3510_, new_n3509_, new_n3505_ );
or   ( new_n3511_, new_n1425_, new_n806_ );
or   ( new_n3512_, new_n1429_, new_n110_ );
and  ( new_n3513_, new_n3512_, new_n3511_ );
and  ( new_n3514_, new_n3513_, new_n1355_ );
and  ( new_n3515_, new_n1433_, RI2b1c4342d828_72 );
and  ( new_n3516_, new_n1423_, RI2b1c4342d7b0_71 );
or   ( new_n3517_, new_n3516_, new_n3515_ );
and  ( new_n3518_, new_n3517_, new_n1267_ );
or   ( new_n3519_, new_n3518_, new_n3514_ );
and  ( new_n3520_, new_n3519_, new_n3510_ );
or   ( new_n3521_, new_n3519_, new_n3510_ );
or   ( new_n3522_, new_n934_, new_n859_ );
or   ( new_n3523_, new_n940_, new_n105_ );
and  ( new_n3524_, new_n3523_, new_n3522_ );
and  ( new_n3525_, new_n3524_, new_n913_ );
and  ( new_n3526_, new_n944_, RI2b1c4342d918_74 );
and  ( new_n3527_, new_n932_, RI2b1c4342d8a0_73 );
or   ( new_n3528_, new_n3527_, new_n3526_ );
and  ( new_n3529_, new_n3528_, new_n938_ );
or   ( new_n3530_, new_n3529_, new_n3525_ );
and  ( new_n3531_, new_n3530_, new_n3521_ );
or   ( new_n3532_, new_n3531_, new_n3520_ );
xor  ( new_n3533_, new_n309_, new_n182_ );
and  ( new_n3534_, new_n3533_, new_n352_ );
xor  ( new_n3535_, RI2b1c4342c220_25, RI2b1c4342d120_57 );
and  ( new_n3536_, new_n3535_, new_n228_ );
and  ( new_n3537_, new_n3536_, new_n138_ );
or   ( new_n3538_, new_n3537_, new_n183_ );
or   ( new_n3539_, new_n3538_, new_n3534_ );
xor  ( new_n3540_, new_n306_, new_n177_ );
and  ( new_n3541_, new_n3540_, new_n354_ );
xor  ( new_n3542_, RI2b1c4342c1a8_24, RI2b1c4342d0a8_56 );
and  ( new_n3543_, new_n3542_, new_n138_ );
and  ( new_n3544_, new_n3543_, new_n230_ );
or   ( new_n3545_, new_n3544_, new_n178_ );
or   ( new_n3546_, new_n3545_, new_n3541_ );
or   ( new_n3547_, new_n3546_, new_n3539_ );
and  ( new_n3548_, new_n3547_, new_n2997_ );
or   ( new_n3549_, new_n3112_, new_n526_ );
or   ( new_n3550_, new_n3116_, new_n99_ );
and  ( new_n3551_, new_n3550_, new_n3549_ );
and  ( new_n3552_, new_n3551_, new_n3004_ );
and  ( new_n3553_, new_n3120_, RI2b1c4342d558_66 );
and  ( new_n3554_, new_n3110_, RI2b1c4342d4e0_65 );
or   ( new_n3555_, new_n3554_, new_n3553_ );
and  ( new_n3556_, new_n3555_, new_n2868_ );
or   ( new_n3557_, new_n3556_, new_n3552_ );
and  ( new_n3558_, new_n3557_, new_n3548_ );
or   ( new_n3559_, new_n3557_, new_n3548_ );
or   ( new_n3560_, new_n2450_, new_n612_ );
or   ( new_n3561_, new_n2454_, new_n112_ );
and  ( new_n3562_, new_n3561_, new_n3560_ );
and  ( new_n3563_, new_n3562_, new_n2334_ );
and  ( new_n3564_, new_n2458_, RI2b1c4342d648_68 );
and  ( new_n3565_, new_n2448_, RI2b1c4342d5d0_67 );
or   ( new_n3566_, new_n3565_, new_n3564_ );
and  ( new_n3567_, new_n3566_, new_n2168_ );
or   ( new_n3568_, new_n3567_, new_n3563_ );
and  ( new_n3569_, new_n3568_, new_n3559_ );
or   ( new_n3570_, new_n3569_, new_n3558_ );
and  ( new_n3571_, new_n3570_, new_n3532_ );
or   ( new_n3572_, new_n3570_, new_n3532_ );
or   ( new_n3573_, new_n453_, new_n886_ );
or   ( new_n3574_, new_n459_, new_n843_ );
and  ( new_n3575_, new_n3574_, new_n3573_ );
and  ( new_n3576_, new_n3575_, new_n428_ );
and  ( new_n3577_, new_n463_, RI2b1c4342da08_76 );
and  ( new_n3578_, new_n451_, RI2b1c4342d990_75 );
or   ( new_n3579_, new_n3578_, new_n3577_ );
and  ( new_n3580_, new_n3579_, new_n457_ );
or   ( new_n3581_, new_n3580_, new_n3576_ );
or   ( new_n3582_, new_n524_, new_n1002_ );
or   ( new_n3583_, new_n528_, new_n1004_ );
and  ( new_n3584_, new_n3583_, new_n3582_ );
and  ( new_n3585_, new_n3584_, new_n505_ );
and  ( new_n3586_, new_n537_, RI2b1c4342daf8_78 );
and  ( new_n3587_, new_n522_, RI2b1c4342da80_77 );
or   ( new_n3588_, new_n3587_, new_n3586_ );
and  ( new_n3589_, new_n3588_, new_n533_ );
or   ( new_n3590_, new_n3589_, new_n3585_ );
and  ( new_n3591_, new_n3590_, new_n3581_ );
or   ( new_n3592_, new_n3590_, new_n3581_ );
or   ( new_n3593_, new_n610_, new_n1511_ );
or   ( new_n3594_, new_n614_, new_n1310_ );
and  ( new_n3595_, new_n3594_, new_n3593_ );
and  ( new_n3596_, new_n3595_, new_n590_ );
and  ( new_n3597_, new_n623_, RI2b1c4342dbe8_80 );
and  ( new_n3598_, new_n608_, RI2b1c4342db70_79 );
or   ( new_n3599_, new_n3598_, new_n3597_ );
and  ( new_n3600_, new_n3599_, new_n619_ );
or   ( new_n3601_, new_n3600_, new_n3596_ );
and  ( new_n3602_, new_n3601_, new_n3592_ );
or   ( new_n3603_, new_n3602_, new_n3591_ );
and  ( new_n3604_, new_n3603_, new_n3572_ );
or   ( new_n3605_, new_n3604_, new_n3571_ );
and  ( new_n3606_, new_n3605_, new_n3501_ );
or   ( new_n3607_, new_n3605_, new_n3501_ );
or   ( new_n3608_, new_n3372_, new_n3197_ );
and  ( new_n3609_, new_n3608_, new_n3207_ );
and  ( new_n3610_, new_n3368_, new_n3196_ );
and  ( new_n3611_, new_n3371_, new_n3187_ );
or   ( new_n3612_, new_n3611_, new_n3610_ );
and  ( new_n3613_, new_n3612_, new_n3376_ );
or   ( new_n3614_, new_n3613_, new_n3609_ );
or   ( new_n3615_, new_n3357_, new_n3164_ );
and  ( new_n3616_, new_n3615_, new_n3174_ );
and  ( new_n3617_, new_n3353_, new_n3163_ );
and  ( new_n3618_, new_n3356_, new_n3154_ );
or   ( new_n3619_, new_n3618_, new_n3617_ );
and  ( new_n3620_, new_n3619_, new_n3361_ );
or   ( new_n3621_, new_n3620_, new_n3616_ );
and  ( new_n3622_, new_n3621_, new_n3614_ );
or   ( new_n3623_, new_n3621_, new_n3614_ );
or   ( new_n3624_, new_n3344_, new_n3133_ );
and  ( new_n3625_, new_n3624_, new_n3143_ );
and  ( new_n3626_, new_n3340_, new_n3132_ );
and  ( new_n3627_, new_n3343_, new_n3123_ );
or   ( new_n3628_, new_n3627_, new_n3626_ );
and  ( new_n3629_, new_n3628_, new_n3348_ );
or   ( new_n3630_, new_n3629_, new_n3625_ );
and  ( new_n3631_, new_n3630_, new_n3623_ );
or   ( new_n3632_, new_n3631_, new_n3622_ );
and  ( new_n3633_, new_n3632_, new_n3607_ );
or   ( new_n3634_, new_n3633_, new_n3606_ );
and  ( new_n3635_, new_n3634_, new_n3462_ );
or   ( new_n3636_, new_n3634_, new_n3462_ );
or   ( new_n3637_, new_n3331_, new_n3282_ );
and  ( new_n3638_, new_n3637_, new_n3290_ );
and  ( new_n3639_, new_n3327_, new_n3281_ );
and  ( new_n3640_, new_n3330_, new_n3274_ );
or   ( new_n3641_, new_n3640_, new_n3639_ );
and  ( new_n3642_, new_n3641_, new_n3335_ );
or   ( new_n3643_, new_n3642_, new_n3638_ );
and  ( new_n3644_, new_n3643_, new_n3636_ );
or   ( new_n3645_, new_n3644_, new_n3635_ );
and  ( new_n3646_, new_n3645_, new_n3442_ );
or   ( new_n3647_, new_n3414_, new_n3293_ );
and  ( new_n3648_, new_n3647_, new_n3300_ );
and  ( new_n3649_, new_n3412_, new_n3292_ );
and  ( new_n3650_, new_n3337_, new_n3272_ );
or   ( new_n3651_, new_n3650_, new_n3649_ );
and  ( new_n3652_, new_n3651_, new_n3417_ );
or   ( new_n3653_, new_n3652_, new_n3648_ );
or   ( new_n3654_, new_n3645_, new_n3442_ );
and  ( new_n3655_, new_n3654_, new_n3653_ );
or   ( new_n3656_, new_n3655_, new_n3646_ );
or   ( new_n3657_, new_n3656_, new_n3435_ );
or   ( new_n3658_, new_n3657_, new_n3428_ );
and  ( new_n3659_, new_n3658_, new_n3317_ );
or   ( new_n3660_, new_n3659_, new_n3316_ );
and  ( new_n3661_, new_n3656_, new_n3435_ );
and  ( new_n3662_, new_n3433_, new_n3311_ );
and  ( new_n3663_, new_n3429_, new_n3424_ );
or   ( new_n3664_, new_n3663_, new_n3662_ );
and  ( new_n3665_, new_n3440_, new_n2941_ );
and  ( new_n3666_, new_n3436_, new_n3072_ );
or   ( new_n3667_, new_n3666_, new_n3665_ );
and  ( new_n3668_, new_n3467_, new_n3240_ );
and  ( new_n3669_, new_n3463_, new_n3392_ );
or   ( new_n3670_, new_n3669_, new_n3668_ );
and  ( new_n3671_, new_n3476_, new_n734_ );
and  ( new_n3672_, new_n3472_, new_n762_ );
or   ( new_n3673_, new_n3672_, new_n3671_ );
and  ( new_n3674_, new_n3485_, new_n785_ );
and  ( new_n3675_, new_n3481_, new_n813_ );
or   ( new_n3676_, new_n3675_, new_n3674_ );
and  ( new_n3677_, new_n3676_, new_n3673_ );
or   ( new_n3678_, new_n3676_, new_n3673_ );
and  ( new_n3679_, new_n3496_, new_n842_ );
and  ( new_n3680_, new_n3492_, new_n866_ );
or   ( new_n3681_, new_n3680_, new_n3679_ );
and  ( new_n3682_, new_n3681_, new_n3678_ );
or   ( new_n3683_, new_n3682_, new_n3677_ );
or   ( new_n3684_, new_n3683_, new_n3670_ );
not  ( new_n3685_, new_n228_ );
nor  ( new_n3686_, new_n3535_, new_n3685_ );
and  ( new_n3687_, new_n3535_, new_n352_ );
or   ( new_n3688_, new_n3687_, new_n3686_ );
and  ( new_n3689_, new_n3688_, new_n309_ );
nor  ( new_n3690_, new_n3542_, new_n231_ );
and  ( new_n3691_, new_n3542_, new_n354_ );
or   ( new_n3692_, new_n3691_, new_n3690_ );
and  ( new_n3693_, new_n3692_, new_n306_ );
and  ( new_n3694_, new_n3693_, new_n3689_ );
or   ( new_n3695_, new_n3694_, new_n2866_ );
and  ( new_n3696_, new_n3555_, new_n3004_ );
and  ( new_n3697_, new_n3551_, new_n2868_ );
or   ( new_n3698_, new_n3697_, new_n3696_ );
and  ( new_n3699_, new_n3698_, new_n3695_ );
or   ( new_n3700_, new_n3698_, new_n3695_ );
and  ( new_n3701_, new_n3566_, new_n2334_ );
and  ( new_n3702_, new_n3562_, new_n2168_ );
or   ( new_n3703_, new_n3702_, new_n3701_ );
and  ( new_n3704_, new_n3703_, new_n3700_ );
or   ( new_n3705_, new_n3704_, new_n3699_ );
and  ( new_n3706_, new_n3508_, new_n1824_ );
and  ( new_n3707_, new_n3504_, new_n1717_ );
or   ( new_n3708_, new_n3707_, new_n3706_ );
and  ( new_n3709_, new_n3517_, new_n1355_ );
and  ( new_n3710_, new_n3513_, new_n1267_ );
or   ( new_n3711_, new_n3710_, new_n3709_ );
and  ( new_n3712_, new_n3711_, new_n3708_ );
or   ( new_n3713_, new_n3711_, new_n3708_ );
and  ( new_n3714_, new_n3528_, new_n913_ );
and  ( new_n3715_, new_n3524_, new_n938_ );
or   ( new_n3716_, new_n3715_, new_n3714_ );
and  ( new_n3717_, new_n3716_, new_n3713_ );
or   ( new_n3718_, new_n3717_, new_n3712_ );
and  ( new_n3719_, new_n3718_, new_n3705_ );
or   ( new_n3720_, new_n3718_, new_n3705_ );
and  ( new_n3721_, new_n3579_, new_n428_ );
and  ( new_n3722_, new_n3575_, new_n457_ );
or   ( new_n3723_, new_n3722_, new_n3721_ );
and  ( new_n3724_, new_n3588_, new_n505_ );
and  ( new_n3725_, new_n3584_, new_n533_ );
or   ( new_n3726_, new_n3725_, new_n3724_ );
and  ( new_n3727_, new_n3726_, new_n3723_ );
or   ( new_n3728_, new_n3726_, new_n3723_ );
and  ( new_n3729_, new_n3599_, new_n590_ );
and  ( new_n3730_, new_n3595_, new_n619_ );
or   ( new_n3731_, new_n3730_, new_n3729_ );
and  ( new_n3732_, new_n3731_, new_n3728_ );
or   ( new_n3733_, new_n3732_, new_n3727_ );
and  ( new_n3734_, new_n3733_, new_n3720_ );
or   ( new_n3735_, new_n3734_, new_n3719_ );
and  ( new_n3736_, new_n3735_, new_n3684_ );
or   ( new_n3737_, new_n3735_, new_n3684_ );
and  ( new_n3738_, new_n3612_, new_n3207_ );
and  ( new_n3739_, new_n3608_, new_n3376_ );
or   ( new_n3740_, new_n3739_, new_n3738_ );
and  ( new_n3741_, new_n3619_, new_n3174_ );
and  ( new_n3742_, new_n3615_, new_n3361_ );
or   ( new_n3743_, new_n3742_, new_n3741_ );
and  ( new_n3744_, new_n3743_, new_n3740_ );
or   ( new_n3745_, new_n3743_, new_n3740_ );
and  ( new_n3746_, new_n3628_, new_n3143_ );
and  ( new_n3747_, new_n3624_, new_n3348_ );
or   ( new_n3748_, new_n3747_, new_n3746_ );
and  ( new_n3749_, new_n3748_, new_n3745_ );
or   ( new_n3750_, new_n3749_, new_n3744_ );
and  ( new_n3751_, new_n3750_, new_n3737_ );
or   ( new_n3752_, new_n3751_, new_n3736_ );
and  ( new_n3753_, new_n3406_, new_n3269_ );
and  ( new_n3754_, new_n3409_, new_n3262_ );
or   ( new_n3755_, new_n3754_, new_n3753_ );
and  ( new_n3756_, new_n3449_, new_n3251_ );
and  ( new_n3757_, new_n3445_, new_n3399_ );
or   ( new_n3758_, new_n3757_, new_n3756_ );
and  ( new_n3759_, new_n3758_, new_n3755_ );
or   ( new_n3760_, new_n3758_, new_n3755_ );
and  ( new_n3761_, new_n3458_, new_n3209_ );
and  ( new_n3762_, new_n3454_, new_n3378_ );
or   ( new_n3763_, new_n3762_, new_n3761_ );
and  ( new_n3764_, new_n3763_, new_n3760_ );
or   ( new_n3765_, new_n3764_, new_n3759_ );
and  ( new_n3766_, new_n3765_, new_n3752_ );
or   ( new_n3767_, new_n3765_, new_n3752_ );
and  ( new_n3768_, new_n3641_, new_n3290_ );
and  ( new_n3769_, new_n3637_, new_n3335_ );
or   ( new_n3770_, new_n3769_, new_n3768_ );
and  ( new_n3771_, new_n3770_, new_n3767_ );
or   ( new_n3772_, new_n3771_, new_n3766_ );
and  ( new_n3773_, new_n3772_, new_n3667_ );
and  ( new_n3774_, new_n3651_, new_n3300_ );
and  ( new_n3775_, new_n3647_, new_n3417_ );
or   ( new_n3776_, new_n3775_, new_n3774_ );
or   ( new_n3777_, new_n3772_, new_n3667_ );
and  ( new_n3778_, new_n3777_, new_n3776_ );
or   ( new_n3779_, new_n3778_, new_n3773_ );
and  ( new_n3780_, new_n3779_, new_n3664_ );
or   ( new_n3781_, new_n3780_, new_n3661_ );
or   ( new_n3782_, new_n3773_, new_n3646_ );
and  ( new_n3783_, new_n3782_, new_n3653_ );
and  ( new_n3784_, new_n3772_, new_n3442_ );
and  ( new_n3785_, new_n3667_, new_n3645_ );
or   ( new_n3786_, new_n3785_, new_n3784_ );
and  ( new_n3787_, new_n3786_, new_n3776_ );
or   ( new_n3788_, new_n3787_, new_n3783_ );
or   ( new_n3789_, new_n3403_, new_n3254_ );
and  ( new_n3790_, new_n3789_, new_n3270_ );
and  ( new_n3791_, new_n3380_, new_n3253_ );
and  ( new_n3792_, new_n3401_, new_n3211_ );
or   ( new_n3793_, new_n3792_, new_n3791_ );
and  ( new_n3794_, new_n3793_, new_n3410_ );
or   ( new_n3795_, new_n3794_, new_n3790_ );
and  ( new_n3796_, new_n3693_, new_n2997_ );
and  ( new_n3797_, new_n3546_, new_n2866_ );
and  ( new_n3798_, new_n3693_, new_n3539_ );
and  ( new_n3799_, new_n3689_, new_n3546_ );
or   ( new_n3800_, new_n3799_, new_n3798_ );
or   ( new_n3801_, new_n3800_, new_n3797_ );
or   ( new_n3802_, new_n3801_, new_n3796_ );
or   ( new_n3803_, new_n3802_, new_n99_ );
and  ( new_n3804_, new_n3803_, new_n3695_ );
and  ( new_n3805_, new_n3546_, new_n3539_ );
or   ( new_n3806_, new_n3805_, new_n3694_ );
and  ( new_n3807_, new_n3546_, new_n2997_ );
and  ( new_n3808_, new_n3693_, new_n2866_ );
or   ( new_n3809_, new_n3808_, new_n3807_ );
and  ( new_n3810_, new_n3809_, new_n3806_ );
and  ( new_n3811_, new_n3810_, RI2b1c4342d4e0_65 );
and  ( new_n3812_, new_n3811_, new_n3548_ );
or   ( new_n3813_, new_n3812_, new_n3804_ );
or   ( new_n3814_, new_n3112_, new_n112_ );
or   ( new_n3815_, new_n3116_, new_n526_ );
and  ( new_n3816_, new_n3815_, new_n3814_ );
and  ( new_n3817_, new_n3816_, new_n3004_ );
and  ( new_n3818_, new_n3120_, RI2b1c4342d5d0_67 );
and  ( new_n3819_, new_n3110_, RI2b1c4342d558_66 );
or   ( new_n3820_, new_n3819_, new_n3818_ );
and  ( new_n3821_, new_n3820_, new_n2868_ );
or   ( new_n3822_, new_n3821_, new_n3817_ );
and  ( new_n3823_, new_n3822_, new_n3813_ );
or   ( new_n3824_, new_n3822_, new_n3813_ );
or   ( new_n3825_, new_n2450_, new_n591_ );
or   ( new_n3826_, new_n2454_, new_n612_ );
and  ( new_n3827_, new_n3826_, new_n3825_ );
and  ( new_n3828_, new_n3827_, new_n2334_ );
and  ( new_n3829_, new_n2458_, RI2b1c4342d6c0_69 );
and  ( new_n3830_, new_n2448_, RI2b1c4342d648_68 );
or   ( new_n3831_, new_n3830_, new_n3829_ );
and  ( new_n3832_, new_n3831_, new_n2168_ );
or   ( new_n3833_, new_n3832_, new_n3828_ );
and  ( new_n3834_, new_n3833_, new_n3824_ );
or   ( new_n3835_, new_n3834_, new_n3823_ );
or   ( new_n3836_, new_n1910_, new_n110_ );
or   ( new_n3837_, new_n1914_, new_n755_ );
and  ( new_n3838_, new_n3837_, new_n3836_ );
and  ( new_n3839_, new_n3838_, new_n1824_ );
and  ( new_n3840_, new_n1918_, RI2b1c4342d7b0_71 );
and  ( new_n3841_, new_n1908_, RI2b1c4342d738_70 );
or   ( new_n3842_, new_n3841_, new_n3840_ );
and  ( new_n3843_, new_n3842_, new_n1717_ );
or   ( new_n3844_, new_n3843_, new_n3839_ );
or   ( new_n3845_, new_n1425_, new_n105_ );
or   ( new_n3846_, new_n1429_, new_n806_ );
and  ( new_n3847_, new_n3846_, new_n3845_ );
and  ( new_n3848_, new_n3847_, new_n1355_ );
and  ( new_n3849_, new_n1433_, RI2b1c4342d8a0_73 );
and  ( new_n3850_, new_n1423_, RI2b1c4342d828_72 );
or   ( new_n3851_, new_n3850_, new_n3849_ );
and  ( new_n3852_, new_n3851_, new_n1267_ );
or   ( new_n3853_, new_n3852_, new_n3848_ );
and  ( new_n3854_, new_n3853_, new_n3844_ );
or   ( new_n3855_, new_n3853_, new_n3844_ );
or   ( new_n3856_, new_n934_, new_n843_ );
or   ( new_n3857_, new_n940_, new_n859_ );
and  ( new_n3858_, new_n3857_, new_n3856_ );
and  ( new_n3859_, new_n3858_, new_n913_ );
and  ( new_n3860_, new_n944_, RI2b1c4342d990_75 );
and  ( new_n3861_, new_n932_, RI2b1c4342d918_74 );
or   ( new_n3862_, new_n3861_, new_n3860_ );
and  ( new_n3863_, new_n3862_, new_n938_ );
or   ( new_n3864_, new_n3863_, new_n3859_ );
and  ( new_n3865_, new_n3864_, new_n3855_ );
or   ( new_n3866_, new_n3865_, new_n3854_ );
and  ( new_n3867_, new_n3866_, new_n3835_ );
or   ( new_n3868_, new_n3866_, new_n3835_ );
or   ( new_n3869_, new_n453_, new_n1004_ );
or   ( new_n3870_, new_n459_, new_n886_ );
and  ( new_n3871_, new_n3870_, new_n3869_ );
and  ( new_n3872_, new_n3871_, new_n428_ );
and  ( new_n3873_, new_n463_, RI2b1c4342da80_77 );
and  ( new_n3874_, new_n451_, RI2b1c4342da08_76 );
or   ( new_n3875_, new_n3874_, new_n3873_ );
and  ( new_n3876_, new_n3875_, new_n457_ );
or   ( new_n3877_, new_n3876_, new_n3872_ );
or   ( new_n3878_, new_n524_, new_n1310_ );
or   ( new_n3879_, new_n528_, new_n1002_ );
and  ( new_n3880_, new_n3879_, new_n3878_ );
and  ( new_n3881_, new_n3880_, new_n505_ );
and  ( new_n3882_, new_n537_, RI2b1c4342db70_79 );
and  ( new_n3883_, new_n522_, RI2b1c4342daf8_78 );
or   ( new_n3884_, new_n3883_, new_n3882_ );
and  ( new_n3885_, new_n3884_, new_n533_ );
or   ( new_n3886_, new_n3885_, new_n3881_ );
and  ( new_n3887_, new_n3886_, new_n3877_ );
or   ( new_n3888_, new_n3886_, new_n3877_ );
or   ( new_n3889_, new_n610_, new_n126_ );
or   ( new_n3890_, new_n614_, new_n1511_ );
and  ( new_n3891_, new_n3890_, new_n3889_ );
and  ( new_n3892_, new_n3891_, new_n590_ );
and  ( new_n3893_, new_n623_, RI2b1c4342dc60_81 );
and  ( new_n3894_, new_n608_, RI2b1c4342dbe8_80 );
or   ( new_n3895_, new_n3894_, new_n3893_ );
and  ( new_n3896_, new_n3895_, new_n619_ );
or   ( new_n3897_, new_n3896_, new_n3892_ );
and  ( new_n3898_, new_n3897_, new_n3888_ );
or   ( new_n3899_, new_n3898_, new_n3887_ );
and  ( new_n3900_, new_n3899_, new_n3868_ );
or   ( new_n3901_, new_n3900_, new_n3867_ );
not  ( new_n3902_, RI2b1c4342dfa8_88 );
or   ( new_n3903_, new_n841_, new_n3902_ );
or   ( new_n3904_, new_n753_, new_n121_ );
or   ( new_n3905_, new_n757_, new_n2119_ );
and  ( new_n3906_, new_n3905_, new_n3904_ );
and  ( new_n3907_, new_n3906_, new_n734_ );
and  ( new_n3908_, new_n766_, RI2b1c4342dd50_83 );
and  ( new_n3909_, new_n751_, RI2b1c4342dcd8_82 );
or   ( new_n3910_, new_n3909_, new_n3908_ );
and  ( new_n3911_, new_n3910_, new_n762_ );
or   ( new_n3912_, new_n3911_, new_n3907_ );
or   ( new_n3913_, new_n804_, new_n2806_ );
or   ( new_n3914_, new_n808_, new_n2541_ );
and  ( new_n3915_, new_n3914_, new_n3913_ );
and  ( new_n3916_, new_n3915_, new_n785_ );
and  ( new_n3917_, new_n817_, RI2b1c4342de40_85 );
and  ( new_n3918_, new_n802_, RI2b1c4342ddc8_84 );
or   ( new_n3919_, new_n3918_, new_n3917_ );
and  ( new_n3920_, new_n3919_, new_n813_ );
or   ( new_n3921_, new_n3920_, new_n3916_ );
and  ( new_n3922_, new_n3921_, new_n3912_ );
or   ( new_n3923_, new_n3921_, new_n3912_ );
not  ( new_n3924_, RI2b1c4342df30_87 );
or   ( new_n3925_, new_n857_, new_n3924_ );
or   ( new_n3926_, new_n861_, new_n3239_ );
and  ( new_n3927_, new_n3926_, new_n3925_ );
and  ( new_n3928_, new_n3927_, new_n842_ );
and  ( new_n3929_, new_n870_, RI2b1c4342df30_87 );
and  ( new_n3930_, new_n855_, RI2b1c4342deb8_86 );
or   ( new_n3931_, new_n3930_, new_n3929_ );
and  ( new_n3932_, new_n3931_, new_n866_ );
or   ( new_n3933_, new_n3932_, new_n3928_ );
and  ( new_n3934_, new_n3933_, new_n3923_ );
or   ( new_n3935_, new_n3934_, new_n3922_ );
and  ( new_n3936_, new_n3935_, new_n3903_ );
or   ( new_n3937_, new_n3935_, new_n3903_ );
or   ( new_n3938_, new_n841_, new_n3924_ );
and  ( new_n3939_, new_n3938_, new_n3937_ );
or   ( new_n3940_, new_n3939_, new_n3936_ );
and  ( new_n3941_, new_n3940_, new_n3901_ );
or   ( new_n3942_, new_n3940_, new_n3901_ );
or   ( new_n3943_, new_n3677_, new_n3488_ );
and  ( new_n3944_, new_n3943_, new_n3498_ );
and  ( new_n3945_, new_n3673_, new_n3487_ );
and  ( new_n3946_, new_n3676_, new_n3478_ );
or   ( new_n3947_, new_n3946_, new_n3945_ );
and  ( new_n3948_, new_n3947_, new_n3681_ );
or   ( new_n3949_, new_n3948_, new_n3944_ );
or   ( new_n3950_, new_n3727_, new_n3591_ );
and  ( new_n3951_, new_n3950_, new_n3601_ );
and  ( new_n3952_, new_n3723_, new_n3590_ );
and  ( new_n3953_, new_n3726_, new_n3581_ );
or   ( new_n3954_, new_n3953_, new_n3952_ );
and  ( new_n3955_, new_n3954_, new_n3731_ );
or   ( new_n3956_, new_n3955_, new_n3951_ );
and  ( new_n3957_, new_n3956_, new_n3949_ );
or   ( new_n3958_, new_n3956_, new_n3949_ );
or   ( new_n3959_, new_n3712_, new_n3520_ );
and  ( new_n3960_, new_n3959_, new_n3530_ );
and  ( new_n3961_, new_n3708_, new_n3519_ );
and  ( new_n3962_, new_n3711_, new_n3510_ );
or   ( new_n3963_, new_n3962_, new_n3961_ );
and  ( new_n3964_, new_n3963_, new_n3716_ );
or   ( new_n3965_, new_n3964_, new_n3960_ );
and  ( new_n3966_, new_n3965_, new_n3958_ );
or   ( new_n3967_, new_n3966_, new_n3957_ );
and  ( new_n3968_, new_n3967_, new_n3942_ );
or   ( new_n3969_, new_n3968_, new_n3941_ );
or   ( new_n3970_, new_n3744_, new_n3622_ );
and  ( new_n3971_, new_n3970_, new_n3630_ );
and  ( new_n3972_, new_n3740_, new_n3621_ );
and  ( new_n3973_, new_n3743_, new_n3614_ );
or   ( new_n3974_, new_n3973_, new_n3972_ );
and  ( new_n3975_, new_n3974_, new_n3748_ );
or   ( new_n3976_, new_n3975_, new_n3971_ );
and  ( new_n3977_, new_n3683_, new_n3469_ );
and  ( new_n3978_, new_n3670_, new_n3500_ );
or   ( new_n3979_, new_n3978_, new_n3977_ );
and  ( new_n3980_, new_n3979_, new_n3976_ );
or   ( new_n3981_, new_n3979_, new_n3976_ );
or   ( new_n3982_, new_n3719_, new_n3571_ );
and  ( new_n3983_, new_n3982_, new_n3603_ );
and  ( new_n3984_, new_n3705_, new_n3532_ );
and  ( new_n3985_, new_n3718_, new_n3570_ );
or   ( new_n3986_, new_n3985_, new_n3984_ );
and  ( new_n3987_, new_n3986_, new_n3733_ );
or   ( new_n3988_, new_n3987_, new_n3983_ );
and  ( new_n3989_, new_n3988_, new_n3981_ );
or   ( new_n3990_, new_n3989_, new_n3980_ );
and  ( new_n3991_, new_n3990_, new_n3969_ );
or   ( new_n3992_, new_n3990_, new_n3969_ );
or   ( new_n3993_, new_n3759_, new_n3452_ );
and  ( new_n3994_, new_n3993_, new_n3460_ );
and  ( new_n3995_, new_n3755_, new_n3451_ );
and  ( new_n3996_, new_n3758_, new_n3444_ );
or   ( new_n3997_, new_n3996_, new_n3995_ );
and  ( new_n3998_, new_n3997_, new_n3763_ );
or   ( new_n3999_, new_n3998_, new_n3994_ );
and  ( new_n4000_, new_n3999_, new_n3992_ );
or   ( new_n4001_, new_n4000_, new_n3991_ );
and  ( new_n4002_, new_n4001_, new_n3795_ );
or   ( new_n4003_, new_n4001_, new_n3795_ );
or   ( new_n4004_, new_n3766_, new_n3635_ );
and  ( new_n4005_, new_n4004_, new_n3643_ );
and  ( new_n4006_, new_n3752_, new_n3462_ );
and  ( new_n4007_, new_n3765_, new_n3634_ );
or   ( new_n4008_, new_n4007_, new_n4006_ );
and  ( new_n4009_, new_n4008_, new_n3770_ );
or   ( new_n4010_, new_n4009_, new_n4005_ );
and  ( new_n4011_, new_n4010_, new_n4003_ );
or   ( new_n4012_, new_n4011_, new_n4002_ );
or   ( new_n4013_, new_n4012_, new_n3788_ );
and  ( new_n4014_, new_n4013_, new_n3781_ );
or   ( new_n4015_, new_n4013_, new_n3781_ );
and  ( new_n4016_, new_n4012_, new_n3788_ );
and  ( new_n4017_, new_n3786_, new_n3653_ );
and  ( new_n4018_, new_n3782_, new_n3776_ );
or   ( new_n4019_, new_n4018_, new_n4017_ );
and  ( new_n4020_, new_n3793_, new_n3270_ );
and  ( new_n4021_, new_n3789_, new_n3410_ );
or   ( new_n4022_, new_n4021_, new_n4020_ );
and  ( new_n4023_, new_n3811_, new_n3695_ );
and  ( new_n4024_, new_n3803_, new_n3548_ );
or   ( new_n4025_, new_n4024_, new_n4023_ );
and  ( new_n4026_, new_n3820_, new_n3004_ );
and  ( new_n4027_, new_n3816_, new_n2868_ );
or   ( new_n4028_, new_n4027_, new_n4026_ );
and  ( new_n4029_, new_n4028_, new_n4025_ );
or   ( new_n4030_, new_n4028_, new_n4025_ );
and  ( new_n4031_, new_n3831_, new_n2334_ );
and  ( new_n4032_, new_n3827_, new_n2168_ );
or   ( new_n4033_, new_n4032_, new_n4031_ );
and  ( new_n4034_, new_n4033_, new_n4030_ );
or   ( new_n4035_, new_n4034_, new_n4029_ );
and  ( new_n4036_, new_n3842_, new_n1824_ );
and  ( new_n4037_, new_n3838_, new_n1717_ );
or   ( new_n4038_, new_n4037_, new_n4036_ );
and  ( new_n4039_, new_n3851_, new_n1355_ );
and  ( new_n4040_, new_n3847_, new_n1267_ );
or   ( new_n4041_, new_n4040_, new_n4039_ );
and  ( new_n4042_, new_n4041_, new_n4038_ );
or   ( new_n4043_, new_n4041_, new_n4038_ );
and  ( new_n4044_, new_n3862_, new_n913_ );
and  ( new_n4045_, new_n3858_, new_n938_ );
or   ( new_n4046_, new_n4045_, new_n4044_ );
and  ( new_n4047_, new_n4046_, new_n4043_ );
or   ( new_n4048_, new_n4047_, new_n4042_ );
and  ( new_n4049_, new_n4048_, new_n4035_ );
or   ( new_n4050_, new_n4048_, new_n4035_ );
and  ( new_n4051_, new_n3875_, new_n428_ );
and  ( new_n4052_, new_n3871_, new_n457_ );
or   ( new_n4053_, new_n4052_, new_n4051_ );
and  ( new_n4054_, new_n3884_, new_n505_ );
and  ( new_n4055_, new_n3880_, new_n533_ );
or   ( new_n4056_, new_n4055_, new_n4054_ );
and  ( new_n4057_, new_n4056_, new_n4053_ );
or   ( new_n4058_, new_n4056_, new_n4053_ );
and  ( new_n4059_, new_n3895_, new_n590_ );
and  ( new_n4060_, new_n3891_, new_n619_ );
or   ( new_n4061_, new_n4060_, new_n4059_ );
and  ( new_n4062_, new_n4061_, new_n4058_ );
or   ( new_n4063_, new_n4062_, new_n4057_ );
and  ( new_n4064_, new_n4063_, new_n4050_ );
or   ( new_n4065_, new_n4064_, new_n4049_ );
and  ( new_n4066_, new_n720_, RI2b1c4342dfa8_88 );
and  ( new_n4067_, new_n3910_, new_n734_ );
and  ( new_n4068_, new_n3906_, new_n762_ );
or   ( new_n4069_, new_n4068_, new_n4067_ );
and  ( new_n4070_, new_n3919_, new_n785_ );
and  ( new_n4071_, new_n3915_, new_n813_ );
or   ( new_n4072_, new_n4071_, new_n4070_ );
and  ( new_n4073_, new_n4072_, new_n4069_ );
or   ( new_n4074_, new_n4072_, new_n4069_ );
and  ( new_n4075_, new_n3931_, new_n842_ );
and  ( new_n4076_, new_n3927_, new_n866_ );
or   ( new_n4077_, new_n4076_, new_n4075_ );
and  ( new_n4078_, new_n4077_, new_n4074_ );
or   ( new_n4079_, new_n4078_, new_n4073_ );
and  ( new_n4080_, new_n4079_, new_n4066_ );
or   ( new_n4081_, new_n4079_, new_n4066_ );
and  ( new_n4082_, new_n720_, RI2b1c4342df30_87 );
and  ( new_n4083_, new_n4082_, new_n4081_ );
or   ( new_n4084_, new_n4083_, new_n4080_ );
and  ( new_n4085_, new_n4084_, new_n4065_ );
or   ( new_n4086_, new_n4084_, new_n4065_ );
and  ( new_n4087_, new_n3947_, new_n3498_ );
and  ( new_n4088_, new_n3943_, new_n3681_ );
or   ( new_n4089_, new_n4088_, new_n4087_ );
and  ( new_n4090_, new_n3954_, new_n3601_ );
and  ( new_n4091_, new_n3950_, new_n3731_ );
or   ( new_n4092_, new_n4091_, new_n4090_ );
and  ( new_n4093_, new_n4092_, new_n4089_ );
or   ( new_n4094_, new_n4092_, new_n4089_ );
and  ( new_n4095_, new_n3963_, new_n3530_ );
and  ( new_n4096_, new_n3959_, new_n3716_ );
or   ( new_n4097_, new_n4096_, new_n4095_ );
and  ( new_n4098_, new_n4097_, new_n4094_ );
or   ( new_n4099_, new_n4098_, new_n4093_ );
and  ( new_n4100_, new_n4099_, new_n4086_ );
or   ( new_n4101_, new_n4100_, new_n4085_ );
and  ( new_n4102_, new_n3974_, new_n3630_ );
and  ( new_n4103_, new_n3970_, new_n3748_ );
or   ( new_n4104_, new_n4103_, new_n4102_ );
and  ( new_n4105_, new_n3683_, new_n3670_ );
or   ( new_n4106_, new_n4105_, new_n3501_ );
and  ( new_n4107_, new_n4106_, new_n4104_ );
or   ( new_n4108_, new_n4106_, new_n4104_ );
and  ( new_n4109_, new_n3986_, new_n3603_ );
and  ( new_n4110_, new_n3982_, new_n3733_ );
or   ( new_n4111_, new_n4110_, new_n4109_ );
and  ( new_n4112_, new_n4111_, new_n4108_ );
or   ( new_n4113_, new_n4112_, new_n4107_ );
and  ( new_n4114_, new_n4113_, new_n4101_ );
or   ( new_n4115_, new_n4113_, new_n4101_ );
and  ( new_n4116_, new_n3997_, new_n3460_ );
and  ( new_n4117_, new_n3993_, new_n3763_ );
or   ( new_n4118_, new_n4117_, new_n4116_ );
and  ( new_n4119_, new_n4118_, new_n4115_ );
or   ( new_n4120_, new_n4119_, new_n4114_ );
and  ( new_n4121_, new_n4120_, new_n4022_ );
or   ( new_n4122_, new_n4120_, new_n4022_ );
and  ( new_n4123_, new_n4008_, new_n3643_ );
and  ( new_n4124_, new_n4004_, new_n3770_ );
or   ( new_n4125_, new_n4124_, new_n4123_ );
and  ( new_n4126_, new_n4125_, new_n4122_ );
or   ( new_n4127_, new_n4126_, new_n4121_ );
and  ( new_n4128_, new_n4127_, new_n4019_ );
or   ( new_n4129_, new_n4128_, new_n4016_ );
or   ( new_n4130_, new_n4121_, new_n4002_ );
and  ( new_n4131_, new_n4130_, new_n4010_ );
and  ( new_n4132_, new_n4120_, new_n3795_ );
and  ( new_n4133_, new_n4022_, new_n4001_ );
or   ( new_n4134_, new_n4133_, new_n4132_ );
and  ( new_n4135_, new_n4134_, new_n4125_ );
or   ( new_n4136_, new_n4135_, new_n4131_ );
or   ( new_n4137_, new_n3736_, new_n3606_ );
and  ( new_n4138_, new_n4137_, new_n3632_ );
and  ( new_n4139_, new_n3735_, new_n3501_ );
and  ( new_n4140_, new_n3684_, new_n3605_ );
or   ( new_n4141_, new_n4140_, new_n4139_ );
and  ( new_n4142_, new_n4141_, new_n3750_ );
or   ( new_n4143_, new_n4142_, new_n4138_ );
or   ( new_n4144_, new_n3699_, new_n3558_ );
and  ( new_n4145_, new_n4144_, new_n3568_ );
and  ( new_n4146_, new_n3695_, new_n3557_ );
and  ( new_n4147_, new_n3698_, new_n3548_ );
or   ( new_n4148_, new_n4147_, new_n4146_ );
and  ( new_n4149_, new_n4148_, new_n3703_ );
or   ( new_n4150_, new_n4149_, new_n4145_ );
or   ( new_n4151_, new_n4093_, new_n3957_ );
and  ( new_n4152_, new_n4151_, new_n3965_ );
and  ( new_n4153_, new_n4089_, new_n3956_ );
and  ( new_n4154_, new_n4092_, new_n3949_ );
or   ( new_n4155_, new_n4154_, new_n4153_ );
and  ( new_n4156_, new_n4155_, new_n4097_ );
or   ( new_n4157_, new_n4156_, new_n4152_ );
and  ( new_n4158_, new_n4157_, new_n4150_ );
or   ( new_n4159_, new_n4157_, new_n4150_ );
or   ( new_n4160_, new_n4080_, new_n3936_ );
and  ( new_n4161_, new_n4160_, new_n3938_ );
and  ( new_n4162_, new_n4079_, new_n3903_ );
and  ( new_n4163_, new_n4066_, new_n3935_ );
or   ( new_n4164_, new_n4163_, new_n4162_ );
and  ( new_n4165_, new_n4164_, new_n4082_ );
or   ( new_n4166_, new_n4165_, new_n4161_ );
and  ( new_n4167_, new_n4166_, new_n4159_ );
or   ( new_n4168_, new_n4167_, new_n4158_ );
or   ( new_n4169_, new_n2450_, new_n755_ );
or   ( new_n4170_, new_n2454_, new_n591_ );
and  ( new_n4171_, new_n4170_, new_n4169_ );
and  ( new_n4172_, new_n4171_, new_n2334_ );
and  ( new_n4173_, new_n2458_, RI2b1c4342d738_70 );
and  ( new_n4174_, new_n2448_, RI2b1c4342d6c0_69 );
or   ( new_n4175_, new_n4174_, new_n4173_ );
and  ( new_n4176_, new_n4175_, new_n2168_ );
or   ( new_n4177_, new_n4176_, new_n4172_ );
or   ( new_n4178_, new_n1910_, new_n806_ );
or   ( new_n4179_, new_n1914_, new_n110_ );
and  ( new_n4180_, new_n4179_, new_n4178_ );
and  ( new_n4181_, new_n4180_, new_n1824_ );
and  ( new_n4182_, new_n1918_, RI2b1c4342d828_72 );
and  ( new_n4183_, new_n1908_, RI2b1c4342d7b0_71 );
or   ( new_n4184_, new_n4183_, new_n4182_ );
and  ( new_n4185_, new_n4184_, new_n1717_ );
or   ( new_n4186_, new_n4185_, new_n4181_ );
and  ( new_n4187_, new_n4186_, new_n4177_ );
or   ( new_n4188_, new_n4186_, new_n4177_ );
or   ( new_n4189_, new_n1425_, new_n859_ );
or   ( new_n4190_, new_n1429_, new_n105_ );
and  ( new_n4191_, new_n4190_, new_n4189_ );
and  ( new_n4192_, new_n4191_, new_n1355_ );
and  ( new_n4193_, new_n1433_, RI2b1c4342d918_74 );
and  ( new_n4194_, new_n1423_, RI2b1c4342d8a0_73 );
or   ( new_n4195_, new_n4194_, new_n4193_ );
and  ( new_n4196_, new_n4195_, new_n1267_ );
or   ( new_n4197_, new_n4196_, new_n4192_ );
and  ( new_n4198_, new_n4197_, new_n4188_ );
or   ( new_n4199_, new_n4198_, new_n4187_ );
xor  ( new_n4200_, new_n317_, new_n191_ );
and  ( new_n4201_, new_n4200_, new_n347_ );
xor  ( new_n4202_, RI2b1c4342c310_27, RI2b1c4342d210_59 );
and  ( new_n4203_, new_n4202_, new_n223_ );
and  ( new_n4204_, new_n4203_, new_n138_ );
or   ( new_n4205_, new_n4204_, new_n192_ );
or   ( new_n4206_, new_n4205_, new_n4201_ );
xor  ( new_n4207_, new_n314_, new_n186_ );
and  ( new_n4208_, new_n4207_, new_n349_ );
xor  ( new_n4209_, RI2b1c4342c298_26, RI2b1c4342d198_58 );
and  ( new_n4210_, new_n4209_, new_n225_ );
and  ( new_n4211_, new_n4210_, new_n138_ );
or   ( new_n4212_, new_n4211_, new_n187_ );
or   ( new_n4213_, new_n4212_, new_n4208_ );
or   ( new_n4214_, new_n4213_, new_n4206_ );
and  ( new_n4215_, new_n4214_, new_n3689_ );
or   ( new_n4216_, new_n3802_, new_n526_ );
or   ( new_n4217_, new_n3806_, new_n99_ );
and  ( new_n4218_, new_n4217_, new_n4216_ );
and  ( new_n4219_, new_n4218_, new_n3695_ );
and  ( new_n4220_, new_n3810_, RI2b1c4342d558_66 );
and  ( new_n4221_, new_n3800_, RI2b1c4342d4e0_65 );
or   ( new_n4222_, new_n4221_, new_n4220_ );
and  ( new_n4223_, new_n4222_, new_n3548_ );
or   ( new_n4224_, new_n4223_, new_n4219_ );
and  ( new_n4225_, new_n4224_, new_n4215_ );
or   ( new_n4226_, new_n4224_, new_n4215_ );
or   ( new_n4227_, new_n3112_, new_n612_ );
or   ( new_n4228_, new_n3116_, new_n112_ );
and  ( new_n4229_, new_n4228_, new_n4227_ );
and  ( new_n4230_, new_n4229_, new_n3004_ );
and  ( new_n4231_, new_n3120_, RI2b1c4342d648_68 );
and  ( new_n4232_, new_n3110_, RI2b1c4342d5d0_67 );
or   ( new_n4233_, new_n4232_, new_n4231_ );
and  ( new_n4234_, new_n4233_, new_n2868_ );
or   ( new_n4235_, new_n4234_, new_n4230_ );
and  ( new_n4236_, new_n4235_, new_n4226_ );
or   ( new_n4237_, new_n4236_, new_n4225_ );
and  ( new_n4238_, new_n4237_, new_n4199_ );
or   ( new_n4239_, new_n4237_, new_n4199_ );
or   ( new_n4240_, new_n934_, new_n886_ );
or   ( new_n4241_, new_n940_, new_n843_ );
and  ( new_n4242_, new_n4241_, new_n4240_ );
and  ( new_n4243_, new_n4242_, new_n913_ );
and  ( new_n4244_, new_n944_, RI2b1c4342da08_76 );
and  ( new_n4245_, new_n932_, RI2b1c4342d990_75 );
or   ( new_n4246_, new_n4245_, new_n4244_ );
and  ( new_n4247_, new_n4246_, new_n938_ );
or   ( new_n4248_, new_n4247_, new_n4243_ );
or   ( new_n4249_, new_n453_, new_n1002_ );
or   ( new_n4250_, new_n459_, new_n1004_ );
and  ( new_n4251_, new_n4250_, new_n4249_ );
and  ( new_n4252_, new_n4251_, new_n428_ );
and  ( new_n4253_, new_n463_, RI2b1c4342daf8_78 );
and  ( new_n4254_, new_n451_, RI2b1c4342da80_77 );
or   ( new_n4255_, new_n4254_, new_n4253_ );
and  ( new_n4256_, new_n4255_, new_n457_ );
or   ( new_n4257_, new_n4256_, new_n4252_ );
and  ( new_n4258_, new_n4257_, new_n4248_ );
or   ( new_n4259_, new_n4257_, new_n4248_ );
or   ( new_n4260_, new_n524_, new_n1511_ );
or   ( new_n4261_, new_n528_, new_n1310_ );
and  ( new_n4262_, new_n4261_, new_n4260_ );
and  ( new_n4263_, new_n4262_, new_n505_ );
and  ( new_n4264_, new_n537_, RI2b1c4342dbe8_80 );
and  ( new_n4265_, new_n522_, RI2b1c4342db70_79 );
or   ( new_n4266_, new_n4265_, new_n4264_ );
and  ( new_n4267_, new_n4266_, new_n533_ );
or   ( new_n4268_, new_n4267_, new_n4263_ );
and  ( new_n4269_, new_n4268_, new_n4259_ );
or   ( new_n4270_, new_n4269_, new_n4258_ );
and  ( new_n4271_, new_n4270_, new_n4239_ );
or   ( new_n4272_, new_n4271_, new_n4238_ );
or   ( new_n4273_, new_n610_, new_n2119_ );
or   ( new_n4274_, new_n614_, new_n126_ );
and  ( new_n4275_, new_n4274_, new_n4273_ );
and  ( new_n4276_, new_n4275_, new_n590_ );
and  ( new_n4277_, new_n623_, RI2b1c4342dcd8_82 );
and  ( new_n4278_, new_n608_, RI2b1c4342dc60_81 );
or   ( new_n4279_, new_n4278_, new_n4277_ );
and  ( new_n4280_, new_n4279_, new_n619_ );
or   ( new_n4281_, new_n4280_, new_n4276_ );
or   ( new_n4282_, new_n753_, new_n2541_ );
or   ( new_n4283_, new_n757_, new_n121_ );
and  ( new_n4284_, new_n4283_, new_n4282_ );
and  ( new_n4285_, new_n4284_, new_n734_ );
and  ( new_n4286_, new_n766_, RI2b1c4342ddc8_84 );
and  ( new_n4287_, new_n751_, RI2b1c4342dd50_83 );
or   ( new_n4288_, new_n4287_, new_n4286_ );
and  ( new_n4289_, new_n4288_, new_n762_ );
or   ( new_n4290_, new_n4289_, new_n4285_ );
and  ( new_n4291_, new_n4290_, new_n4281_ );
or   ( new_n4292_, new_n4290_, new_n4281_ );
or   ( new_n4293_, new_n804_, new_n3239_ );
or   ( new_n4294_, new_n808_, new_n2806_ );
and  ( new_n4295_, new_n4294_, new_n4293_ );
and  ( new_n4296_, new_n4295_, new_n785_ );
and  ( new_n4297_, new_n817_, RI2b1c4342deb8_86 );
and  ( new_n4298_, new_n802_, RI2b1c4342de40_85 );
or   ( new_n4299_, new_n4298_, new_n4297_ );
and  ( new_n4300_, new_n4299_, new_n813_ );
or   ( new_n4301_, new_n4300_, new_n4296_ );
and  ( new_n4302_, new_n4301_, new_n4292_ );
or   ( new_n4303_, new_n4302_, new_n4291_ );
or   ( new_n4304_, new_n4303_, new_n4066_ );
and  ( new_n4305_, new_n4303_, new_n4066_ );
or   ( new_n4306_, new_n4073_, new_n3922_ );
and  ( new_n4307_, new_n4306_, new_n3933_ );
and  ( new_n4308_, new_n4069_, new_n3921_ );
and  ( new_n4309_, new_n4072_, new_n3912_ );
or   ( new_n4310_, new_n4309_, new_n4308_ );
and  ( new_n4311_, new_n4310_, new_n4077_ );
or   ( new_n4312_, new_n4311_, new_n4307_ );
or   ( new_n4313_, new_n4312_, new_n4305_ );
and  ( new_n4314_, new_n4313_, new_n4304_ );
and  ( new_n4315_, new_n4314_, new_n4272_ );
or   ( new_n4316_, new_n4314_, new_n4272_ );
or   ( new_n4317_, new_n4057_, new_n3887_ );
and  ( new_n4318_, new_n4317_, new_n3897_ );
and  ( new_n4319_, new_n4053_, new_n3886_ );
and  ( new_n4320_, new_n4056_, new_n3877_ );
or   ( new_n4321_, new_n4320_, new_n4319_ );
and  ( new_n4322_, new_n4321_, new_n4061_ );
or   ( new_n4323_, new_n4322_, new_n4318_ );
or   ( new_n4324_, new_n4042_, new_n3854_ );
and  ( new_n4325_, new_n4324_, new_n3864_ );
and  ( new_n4326_, new_n4038_, new_n3853_ );
and  ( new_n4327_, new_n4041_, new_n3844_ );
or   ( new_n4328_, new_n4327_, new_n4326_ );
and  ( new_n4329_, new_n4328_, new_n4046_ );
or   ( new_n4330_, new_n4329_, new_n4325_ );
and  ( new_n4331_, new_n4330_, new_n4323_ );
or   ( new_n4332_, new_n4330_, new_n4323_ );
or   ( new_n4333_, new_n4029_, new_n3823_ );
and  ( new_n4334_, new_n4333_, new_n3833_ );
and  ( new_n4335_, new_n4025_, new_n3822_ );
and  ( new_n4336_, new_n4028_, new_n3813_ );
or   ( new_n4337_, new_n4336_, new_n4335_ );
and  ( new_n4338_, new_n4337_, new_n4033_ );
or   ( new_n4339_, new_n4338_, new_n4334_ );
and  ( new_n4340_, new_n4339_, new_n4332_ );
or   ( new_n4341_, new_n4340_, new_n4331_ );
and  ( new_n4342_, new_n4341_, new_n4316_ );
or   ( new_n4343_, new_n4342_, new_n4315_ );
and  ( new_n4344_, new_n4343_, new_n4168_ );
or   ( new_n4345_, new_n4343_, new_n4168_ );
or   ( new_n4346_, new_n4107_, new_n3980_ );
and  ( new_n4347_, new_n4346_, new_n3988_ );
and  ( new_n4348_, new_n4104_, new_n3979_ );
and  ( new_n4349_, new_n4106_, new_n3976_ );
or   ( new_n4350_, new_n4349_, new_n4348_ );
and  ( new_n4351_, new_n4350_, new_n4111_ );
or   ( new_n4352_, new_n4351_, new_n4347_ );
and  ( new_n4353_, new_n4352_, new_n4345_ );
or   ( new_n4354_, new_n4353_, new_n4344_ );
and  ( new_n4355_, new_n4354_, new_n4143_ );
or   ( new_n4356_, new_n4354_, new_n4143_ );
or   ( new_n4357_, new_n4114_, new_n3991_ );
and  ( new_n4358_, new_n4357_, new_n3999_ );
and  ( new_n4359_, new_n4101_, new_n3990_ );
and  ( new_n4360_, new_n4113_, new_n3969_ );
or   ( new_n4361_, new_n4360_, new_n4359_ );
and  ( new_n4362_, new_n4361_, new_n4118_ );
or   ( new_n4363_, new_n4362_, new_n4358_ );
and  ( new_n4364_, new_n4363_, new_n4356_ );
or   ( new_n4365_, new_n4364_, new_n4355_ );
or   ( new_n4366_, new_n4365_, new_n4136_ );
or   ( new_n4367_, new_n4366_, new_n4129_ );
and  ( new_n4368_, new_n4367_, new_n4015_ );
or   ( new_n4369_, new_n4368_, new_n4014_ );
and  ( new_n4370_, new_n3657_, new_n3428_ );
or   ( new_n4371_, new_n4370_, new_n3316_ );
or   ( new_n4372_, new_n4371_, new_n4369_ );
and  ( new_n4373_, new_n4372_, new_n3660_ );
and  ( new_n4374_, new_n2967_, new_n2744_ );
or   ( new_n4375_, new_n4374_, new_n2635_ );
or   ( new_n4376_, new_n4375_, new_n2310_ );
or   ( new_n4377_, new_n4376_, new_n4373_ );
and  ( new_n4378_, new_n4377_, new_n2972_ );
and  ( new_n4379_, new_n4366_, new_n4129_ );
or   ( new_n4380_, new_n4379_, new_n4014_ );
or   ( new_n4381_, new_n4380_, new_n4371_ );
or   ( new_n4382_, new_n4381_, new_n4376_ );
and  ( new_n4383_, new_n4365_, new_n4136_ );
and  ( new_n4384_, new_n4134_, new_n4010_ );
and  ( new_n4385_, new_n4130_, new_n4125_ );
or   ( new_n4386_, new_n4385_, new_n4384_ );
and  ( new_n4387_, new_n4141_, new_n3632_ );
and  ( new_n4388_, new_n4137_, new_n3750_ );
or   ( new_n4389_, new_n4388_, new_n4387_ );
not  ( new_n4390_, new_n223_ );
nor  ( new_n4391_, new_n4202_, new_n4390_ );
and  ( new_n4392_, new_n4202_, new_n347_ );
or   ( new_n4393_, new_n4392_, new_n4391_ );
and  ( new_n4394_, new_n4393_, new_n317_ );
nor  ( new_n4395_, new_n4209_, new_n226_ );
and  ( new_n4396_, new_n4209_, new_n349_ );
or   ( new_n4397_, new_n4396_, new_n4395_ );
and  ( new_n4398_, new_n4397_, new_n314_ );
and  ( new_n4399_, new_n4398_, new_n4394_ );
or   ( new_n4400_, new_n4399_, new_n3539_ );
and  ( new_n4401_, new_n4222_, new_n3695_ );
and  ( new_n4402_, new_n4218_, new_n3548_ );
or   ( new_n4403_, new_n4402_, new_n4401_ );
and  ( new_n4404_, new_n4403_, new_n4400_ );
or   ( new_n4405_, new_n4403_, new_n4400_ );
and  ( new_n4406_, new_n4233_, new_n3004_ );
and  ( new_n4407_, new_n4229_, new_n2868_ );
or   ( new_n4408_, new_n4407_, new_n4406_ );
and  ( new_n4409_, new_n4408_, new_n4405_ );
or   ( new_n4410_, new_n4409_, new_n4404_ );
and  ( new_n4411_, new_n4175_, new_n2334_ );
and  ( new_n4412_, new_n4171_, new_n2168_ );
or   ( new_n4413_, new_n4412_, new_n4411_ );
and  ( new_n4414_, new_n4184_, new_n1824_ );
and  ( new_n4415_, new_n4180_, new_n1717_ );
or   ( new_n4416_, new_n4415_, new_n4414_ );
and  ( new_n4417_, new_n4416_, new_n4413_ );
or   ( new_n4418_, new_n4416_, new_n4413_ );
and  ( new_n4419_, new_n4195_, new_n1355_ );
and  ( new_n4420_, new_n4191_, new_n1267_ );
or   ( new_n4421_, new_n4420_, new_n4419_ );
and  ( new_n4422_, new_n4421_, new_n4418_ );
or   ( new_n4423_, new_n4422_, new_n4417_ );
and  ( new_n4424_, new_n4423_, new_n4410_ );
or   ( new_n4425_, new_n4423_, new_n4410_ );
and  ( new_n4426_, new_n4246_, new_n913_ );
and  ( new_n4427_, new_n4242_, new_n938_ );
or   ( new_n4428_, new_n4427_, new_n4426_ );
and  ( new_n4429_, new_n4255_, new_n428_ );
and  ( new_n4430_, new_n4251_, new_n457_ );
or   ( new_n4431_, new_n4430_, new_n4429_ );
and  ( new_n4432_, new_n4431_, new_n4428_ );
or   ( new_n4433_, new_n4431_, new_n4428_ );
and  ( new_n4434_, new_n4266_, new_n505_ );
and  ( new_n4435_, new_n4262_, new_n533_ );
or   ( new_n4436_, new_n4435_, new_n4434_ );
and  ( new_n4437_, new_n4436_, new_n4433_ );
or   ( new_n4438_, new_n4437_, new_n4432_ );
and  ( new_n4439_, new_n4438_, new_n4425_ );
or   ( new_n4440_, new_n4439_, new_n4424_ );
and  ( new_n4441_, new_n4279_, new_n590_ );
and  ( new_n4442_, new_n4275_, new_n619_ );
or   ( new_n4443_, new_n4442_, new_n4441_ );
and  ( new_n4444_, new_n4288_, new_n734_ );
and  ( new_n4445_, new_n4284_, new_n762_ );
or   ( new_n4446_, new_n4445_, new_n4444_ );
and  ( new_n4447_, new_n4446_, new_n4443_ );
or   ( new_n4448_, new_n4446_, new_n4443_ );
and  ( new_n4449_, new_n4299_, new_n785_ );
and  ( new_n4450_, new_n4295_, new_n813_ );
or   ( new_n4451_, new_n4450_, new_n4449_ );
and  ( new_n4452_, new_n4451_, new_n4448_ );
or   ( new_n4453_, new_n4452_, new_n4447_ );
and  ( new_n4454_, new_n4453_, new_n3903_ );
or   ( new_n4455_, new_n4453_, new_n3903_ );
and  ( new_n4456_, new_n4310_, new_n3933_ );
and  ( new_n4457_, new_n4306_, new_n4077_ );
or   ( new_n4458_, new_n4457_, new_n4456_ );
and  ( new_n4459_, new_n4458_, new_n4455_ );
or   ( new_n4460_, new_n4459_, new_n4454_ );
and  ( new_n4461_, new_n4460_, new_n4440_ );
or   ( new_n4462_, new_n4460_, new_n4440_ );
and  ( new_n4463_, new_n4321_, new_n3897_ );
and  ( new_n4464_, new_n4317_, new_n4061_ );
or   ( new_n4465_, new_n4464_, new_n4463_ );
and  ( new_n4466_, new_n4328_, new_n3864_ );
and  ( new_n4467_, new_n4324_, new_n4046_ );
or   ( new_n4468_, new_n4467_, new_n4466_ );
and  ( new_n4469_, new_n4468_, new_n4465_ );
or   ( new_n4470_, new_n4468_, new_n4465_ );
and  ( new_n4471_, new_n4337_, new_n3833_ );
and  ( new_n4472_, new_n4333_, new_n4033_ );
or   ( new_n4473_, new_n4472_, new_n4471_ );
and  ( new_n4474_, new_n4473_, new_n4470_ );
or   ( new_n4475_, new_n4474_, new_n4469_ );
and  ( new_n4476_, new_n4475_, new_n4462_ );
or   ( new_n4477_, new_n4476_, new_n4461_ );
and  ( new_n4478_, new_n4148_, new_n3568_ );
and  ( new_n4479_, new_n4144_, new_n3703_ );
or   ( new_n4480_, new_n4479_, new_n4478_ );
and  ( new_n4481_, new_n4155_, new_n3965_ );
and  ( new_n4482_, new_n4151_, new_n4097_ );
or   ( new_n4483_, new_n4482_, new_n4481_ );
and  ( new_n4484_, new_n4483_, new_n4480_ );
or   ( new_n4485_, new_n4483_, new_n4480_ );
and  ( new_n4486_, new_n4164_, new_n3938_ );
and  ( new_n4487_, new_n4160_, new_n4082_ );
or   ( new_n4488_, new_n4487_, new_n4486_ );
and  ( new_n4489_, new_n4488_, new_n4485_ );
or   ( new_n4490_, new_n4489_, new_n4484_ );
and  ( new_n4491_, new_n4490_, new_n4477_ );
or   ( new_n4492_, new_n4490_, new_n4477_ );
and  ( new_n4493_, new_n4350_, new_n3988_ );
and  ( new_n4494_, new_n4346_, new_n4111_ );
or   ( new_n4495_, new_n4494_, new_n4493_ );
and  ( new_n4496_, new_n4495_, new_n4492_ );
or   ( new_n4497_, new_n4496_, new_n4491_ );
and  ( new_n4498_, new_n4497_, new_n4389_ );
or   ( new_n4499_, new_n4497_, new_n4389_ );
and  ( new_n4500_, new_n4361_, new_n3999_ );
and  ( new_n4501_, new_n4357_, new_n4118_ );
or   ( new_n4502_, new_n4501_, new_n4500_ );
and  ( new_n4503_, new_n4502_, new_n4499_ );
or   ( new_n4504_, new_n4503_, new_n4498_ );
and  ( new_n4505_, new_n4504_, new_n4386_ );
or   ( new_n4506_, new_n4505_, new_n4383_ );
or   ( new_n4507_, new_n4498_, new_n4355_ );
and  ( new_n4508_, new_n4507_, new_n4363_ );
and  ( new_n4509_, new_n4497_, new_n4143_ );
and  ( new_n4510_, new_n4389_, new_n4354_ );
or   ( new_n4511_, new_n4510_, new_n4509_ );
and  ( new_n4512_, new_n4511_, new_n4502_ );
or   ( new_n4513_, new_n4512_, new_n4508_ );
or   ( new_n4514_, new_n4484_, new_n4158_ );
and  ( new_n4515_, new_n4514_, new_n4166_ );
and  ( new_n4516_, new_n4480_, new_n4157_ );
and  ( new_n4517_, new_n4483_, new_n4150_ );
or   ( new_n4518_, new_n4517_, new_n4516_ );
and  ( new_n4519_, new_n4518_, new_n4488_ );
or   ( new_n4520_, new_n4519_, new_n4515_ );
or   ( new_n4521_, new_n4461_, new_n4315_ );
and  ( new_n4522_, new_n4521_, new_n4341_ );
and  ( new_n4523_, new_n4440_, new_n4314_ );
and  ( new_n4524_, new_n4460_, new_n4272_ );
or   ( new_n4525_, new_n4524_, new_n4523_ );
and  ( new_n4526_, new_n4525_, new_n4475_ );
or   ( new_n4527_, new_n4526_, new_n4522_ );
or   ( new_n4528_, new_n4527_, new_n4520_ );
and  ( new_n4529_, new_n4398_, new_n3689_ );
and  ( new_n4530_, new_n4213_, new_n3539_ );
and  ( new_n4531_, new_n4398_, new_n4206_ );
and  ( new_n4532_, new_n4394_, new_n4213_ );
or   ( new_n4533_, new_n4532_, new_n4531_ );
or   ( new_n4534_, new_n4533_, new_n4530_ );
or   ( new_n4535_, new_n4534_, new_n4529_ );
or   ( new_n4536_, new_n4535_, new_n99_ );
and  ( new_n4537_, new_n4536_, new_n4400_ );
and  ( new_n4538_, new_n4213_, new_n4206_ );
or   ( new_n4539_, new_n4538_, new_n4399_ );
and  ( new_n4540_, new_n4213_, new_n3689_ );
and  ( new_n4541_, new_n4398_, new_n3539_ );
or   ( new_n4542_, new_n4541_, new_n4540_ );
and  ( new_n4543_, new_n4542_, new_n4539_ );
and  ( new_n4544_, new_n4543_, RI2b1c4342d4e0_65 );
and  ( new_n4545_, new_n4544_, new_n4215_ );
or   ( new_n4546_, new_n4545_, new_n4537_ );
or   ( new_n4547_, new_n3802_, new_n112_ );
or   ( new_n4548_, new_n3806_, new_n526_ );
and  ( new_n4549_, new_n4548_, new_n4547_ );
and  ( new_n4550_, new_n4549_, new_n3695_ );
and  ( new_n4551_, new_n3810_, RI2b1c4342d5d0_67 );
and  ( new_n4552_, new_n3800_, RI2b1c4342d558_66 );
or   ( new_n4553_, new_n4552_, new_n4551_ );
and  ( new_n4554_, new_n4553_, new_n3548_ );
or   ( new_n4555_, new_n4554_, new_n4550_ );
and  ( new_n4556_, new_n4555_, new_n4546_ );
or   ( new_n4557_, new_n4555_, new_n4546_ );
or   ( new_n4558_, new_n3112_, new_n591_ );
or   ( new_n4559_, new_n3116_, new_n612_ );
and  ( new_n4560_, new_n4559_, new_n4558_ );
and  ( new_n4561_, new_n4560_, new_n3004_ );
and  ( new_n4562_, new_n3120_, RI2b1c4342d6c0_69 );
and  ( new_n4563_, new_n3110_, RI2b1c4342d648_68 );
or   ( new_n4564_, new_n4563_, new_n4562_ );
and  ( new_n4565_, new_n4564_, new_n2868_ );
or   ( new_n4566_, new_n4565_, new_n4561_ );
and  ( new_n4567_, new_n4566_, new_n4557_ );
or   ( new_n4568_, new_n4567_, new_n4556_ );
or   ( new_n4569_, new_n2450_, new_n110_ );
or   ( new_n4570_, new_n2454_, new_n755_ );
and  ( new_n4571_, new_n4570_, new_n4569_ );
and  ( new_n4572_, new_n4571_, new_n2334_ );
and  ( new_n4573_, new_n2458_, RI2b1c4342d7b0_71 );
and  ( new_n4574_, new_n2448_, RI2b1c4342d738_70 );
or   ( new_n4575_, new_n4574_, new_n4573_ );
and  ( new_n4576_, new_n4575_, new_n2168_ );
or   ( new_n4577_, new_n4576_, new_n4572_ );
or   ( new_n4578_, new_n1910_, new_n105_ );
or   ( new_n4579_, new_n1914_, new_n806_ );
and  ( new_n4580_, new_n4579_, new_n4578_ );
and  ( new_n4581_, new_n4580_, new_n1824_ );
and  ( new_n4582_, new_n1918_, RI2b1c4342d8a0_73 );
and  ( new_n4583_, new_n1908_, RI2b1c4342d828_72 );
or   ( new_n4584_, new_n4583_, new_n4582_ );
and  ( new_n4585_, new_n4584_, new_n1717_ );
or   ( new_n4586_, new_n4585_, new_n4581_ );
and  ( new_n4587_, new_n4586_, new_n4577_ );
or   ( new_n4588_, new_n4586_, new_n4577_ );
or   ( new_n4589_, new_n1425_, new_n843_ );
or   ( new_n4590_, new_n1429_, new_n859_ );
and  ( new_n4591_, new_n4590_, new_n4589_ );
and  ( new_n4592_, new_n4591_, new_n1355_ );
and  ( new_n4593_, new_n1433_, RI2b1c4342d990_75 );
and  ( new_n4594_, new_n1423_, RI2b1c4342d918_74 );
or   ( new_n4595_, new_n4594_, new_n4593_ );
and  ( new_n4596_, new_n4595_, new_n1267_ );
or   ( new_n4597_, new_n4596_, new_n4592_ );
and  ( new_n4598_, new_n4597_, new_n4588_ );
or   ( new_n4599_, new_n4598_, new_n4587_ );
and  ( new_n4600_, new_n4599_, new_n4568_ );
or   ( new_n4601_, new_n4599_, new_n4568_ );
or   ( new_n4602_, new_n934_, new_n1004_ );
or   ( new_n4603_, new_n940_, new_n886_ );
and  ( new_n4604_, new_n4603_, new_n4602_ );
and  ( new_n4605_, new_n4604_, new_n913_ );
and  ( new_n4606_, new_n944_, RI2b1c4342da80_77 );
and  ( new_n4607_, new_n932_, RI2b1c4342da08_76 );
or   ( new_n4608_, new_n4607_, new_n4606_ );
and  ( new_n4609_, new_n4608_, new_n938_ );
or   ( new_n4610_, new_n4609_, new_n4605_ );
or   ( new_n4611_, new_n453_, new_n1310_ );
or   ( new_n4612_, new_n459_, new_n1002_ );
and  ( new_n4613_, new_n4612_, new_n4611_ );
and  ( new_n4614_, new_n4613_, new_n428_ );
and  ( new_n4615_, new_n463_, RI2b1c4342db70_79 );
and  ( new_n4616_, new_n451_, RI2b1c4342daf8_78 );
or   ( new_n4617_, new_n4616_, new_n4615_ );
and  ( new_n4618_, new_n4617_, new_n457_ );
or   ( new_n4619_, new_n4618_, new_n4614_ );
and  ( new_n4620_, new_n4619_, new_n4610_ );
or   ( new_n4621_, new_n4619_, new_n4610_ );
or   ( new_n4622_, new_n524_, new_n126_ );
or   ( new_n4623_, new_n528_, new_n1511_ );
and  ( new_n4624_, new_n4623_, new_n4622_ );
and  ( new_n4625_, new_n4624_, new_n505_ );
and  ( new_n4626_, new_n537_, RI2b1c4342dc60_81 );
and  ( new_n4627_, new_n522_, RI2b1c4342dbe8_80 );
or   ( new_n4628_, new_n4627_, new_n4626_ );
and  ( new_n4629_, new_n4628_, new_n533_ );
or   ( new_n4630_, new_n4629_, new_n4625_ );
and  ( new_n4631_, new_n4630_, new_n4621_ );
or   ( new_n4632_, new_n4631_, new_n4620_ );
and  ( new_n4633_, new_n4632_, new_n4601_ );
or   ( new_n4634_, new_n4633_, new_n4600_ );
not  ( new_n4635_, RI2b1c4342e098_90 );
or   ( new_n4636_, new_n841_, new_n4635_ );
or   ( new_n4637_, new_n857_, new_n132_ );
or   ( new_n4638_, new_n861_, new_n3902_ );
and  ( new_n4639_, new_n4638_, new_n4637_ );
and  ( new_n4640_, new_n4639_, new_n842_ );
and  ( new_n4641_, new_n870_, RI2b1c4342e020_89 );
and  ( new_n4642_, new_n855_, RI2b1c4342dfa8_88 );
or   ( new_n4643_, new_n4642_, new_n4641_ );
and  ( new_n4644_, new_n4643_, new_n866_ );
or   ( new_n4645_, new_n4644_, new_n4640_ );
and  ( new_n4646_, new_n4645_, new_n4636_ );
or   ( new_n4647_, new_n610_, new_n121_ );
or   ( new_n4648_, new_n614_, new_n2119_ );
and  ( new_n4649_, new_n4648_, new_n4647_ );
and  ( new_n4650_, new_n4649_, new_n590_ );
and  ( new_n4651_, new_n623_, RI2b1c4342dd50_83 );
and  ( new_n4652_, new_n608_, RI2b1c4342dcd8_82 );
or   ( new_n4653_, new_n4652_, new_n4651_ );
and  ( new_n4654_, new_n4653_, new_n619_ );
or   ( new_n4655_, new_n4654_, new_n4650_ );
or   ( new_n4656_, new_n753_, new_n2806_ );
or   ( new_n4657_, new_n757_, new_n2541_ );
and  ( new_n4658_, new_n4657_, new_n4656_ );
and  ( new_n4659_, new_n4658_, new_n734_ );
and  ( new_n4660_, new_n766_, RI2b1c4342de40_85 );
and  ( new_n4661_, new_n751_, RI2b1c4342ddc8_84 );
or   ( new_n4662_, new_n4661_, new_n4660_ );
and  ( new_n4663_, new_n4662_, new_n762_ );
or   ( new_n4664_, new_n4663_, new_n4659_ );
and  ( new_n4665_, new_n4664_, new_n4655_ );
or   ( new_n4666_, new_n4664_, new_n4655_ );
or   ( new_n4667_, new_n804_, new_n3924_ );
or   ( new_n4668_, new_n808_, new_n3239_ );
and  ( new_n4669_, new_n4668_, new_n4667_ );
and  ( new_n4670_, new_n4669_, new_n785_ );
and  ( new_n4671_, new_n817_, RI2b1c4342df30_87 );
and  ( new_n4672_, new_n802_, RI2b1c4342deb8_86 );
or   ( new_n4673_, new_n4672_, new_n4671_ );
and  ( new_n4674_, new_n4673_, new_n813_ );
or   ( new_n4675_, new_n4674_, new_n4670_ );
and  ( new_n4676_, new_n4675_, new_n4666_ );
or   ( new_n4677_, new_n4676_, new_n4665_ );
and  ( new_n4678_, new_n4677_, new_n4646_ );
or   ( new_n4679_, new_n4677_, new_n4646_ );
or   ( new_n4680_, new_n857_, new_n3902_ );
or   ( new_n4681_, new_n861_, new_n3924_ );
and  ( new_n4682_, new_n4681_, new_n4680_ );
and  ( new_n4683_, new_n4682_, new_n842_ );
and  ( new_n4684_, new_n870_, RI2b1c4342dfa8_88 );
and  ( new_n4685_, new_n855_, RI2b1c4342df30_87 );
or   ( new_n4686_, new_n4685_, new_n4684_ );
and  ( new_n4687_, new_n4686_, new_n866_ );
or   ( new_n4688_, new_n4687_, new_n4683_ );
and  ( new_n4689_, new_n4688_, new_n4679_ );
or   ( new_n4690_, new_n4689_, new_n4678_ );
and  ( new_n4691_, new_n4690_, new_n4634_ );
or   ( new_n4692_, new_n4690_, new_n4634_ );
or   ( new_n4693_, new_n841_, new_n132_ );
or   ( new_n4694_, new_n4447_, new_n4291_ );
and  ( new_n4695_, new_n4694_, new_n4301_ );
and  ( new_n4696_, new_n4443_, new_n4290_ );
and  ( new_n4697_, new_n4446_, new_n4281_ );
or   ( new_n4698_, new_n4697_, new_n4696_ );
and  ( new_n4699_, new_n4698_, new_n4451_ );
or   ( new_n4700_, new_n4699_, new_n4695_ );
and  ( new_n4701_, new_n4700_, new_n4693_ );
or   ( new_n4702_, new_n4700_, new_n4693_ );
or   ( new_n4703_, new_n4432_, new_n4258_ );
and  ( new_n4704_, new_n4703_, new_n4268_ );
and  ( new_n4705_, new_n4428_, new_n4257_ );
and  ( new_n4706_, new_n4431_, new_n4248_ );
or   ( new_n4707_, new_n4706_, new_n4705_ );
and  ( new_n4708_, new_n4707_, new_n4436_ );
or   ( new_n4709_, new_n4708_, new_n4704_ );
and  ( new_n4710_, new_n4709_, new_n4702_ );
or   ( new_n4711_, new_n4710_, new_n4701_ );
and  ( new_n4712_, new_n4711_, new_n4692_ );
or   ( new_n4713_, new_n4712_, new_n4691_ );
or   ( new_n4714_, new_n4469_, new_n4331_ );
and  ( new_n4715_, new_n4714_, new_n4339_ );
and  ( new_n4716_, new_n4465_, new_n4330_ );
and  ( new_n4717_, new_n4468_, new_n4323_ );
or   ( new_n4718_, new_n4717_, new_n4716_ );
and  ( new_n4719_, new_n4718_, new_n4473_ );
or   ( new_n4720_, new_n4719_, new_n4715_ );
or   ( new_n4721_, new_n4454_, new_n4305_ );
and  ( new_n4722_, new_n4721_, new_n4312_ );
and  ( new_n4723_, new_n4453_, new_n4066_ );
and  ( new_n4724_, new_n4303_, new_n3903_ );
or   ( new_n4725_, new_n4724_, new_n4723_ );
and  ( new_n4726_, new_n4725_, new_n4458_ );
or   ( new_n4727_, new_n4726_, new_n4722_ );
and  ( new_n4728_, new_n4727_, new_n4720_ );
or   ( new_n4729_, new_n4727_, new_n4720_ );
or   ( new_n4730_, new_n4424_, new_n4238_ );
and  ( new_n4731_, new_n4730_, new_n4270_ );
and  ( new_n4732_, new_n4410_, new_n4199_ );
and  ( new_n4733_, new_n4423_, new_n4237_ );
or   ( new_n4734_, new_n4733_, new_n4732_ );
and  ( new_n4735_, new_n4734_, new_n4438_ );
or   ( new_n4736_, new_n4735_, new_n4731_ );
and  ( new_n4737_, new_n4736_, new_n4729_ );
or   ( new_n4738_, new_n4737_, new_n4728_ );
and  ( new_n4739_, new_n4738_, new_n4713_ );
or   ( new_n4740_, new_n4738_, new_n4713_ );
or   ( new_n4741_, new_n4049_, new_n3867_ );
and  ( new_n4742_, new_n4741_, new_n3899_ );
and  ( new_n4743_, new_n4035_, new_n3866_ );
and  ( new_n4744_, new_n4048_, new_n3835_ );
or   ( new_n4745_, new_n4744_, new_n4743_ );
and  ( new_n4746_, new_n4745_, new_n4063_ );
or   ( new_n4747_, new_n4746_, new_n4742_ );
and  ( new_n4748_, new_n4747_, new_n4740_ );
or   ( new_n4749_, new_n4748_, new_n4739_ );
and  ( new_n4750_, new_n4749_, new_n4528_ );
or   ( new_n4751_, new_n4749_, new_n4528_ );
or   ( new_n4752_, new_n4085_, new_n3941_ );
and  ( new_n4753_, new_n4752_, new_n3967_ );
and  ( new_n4754_, new_n4065_, new_n3940_ );
and  ( new_n4755_, new_n4084_, new_n3901_ );
or   ( new_n4756_, new_n4755_, new_n4754_ );
and  ( new_n4757_, new_n4756_, new_n4099_ );
or   ( new_n4758_, new_n4757_, new_n4753_ );
and  ( new_n4759_, new_n4758_, new_n4751_ );
or   ( new_n4760_, new_n4759_, new_n4750_ );
or   ( new_n4761_, new_n4760_, new_n4513_ );
and  ( new_n4762_, new_n4761_, new_n4506_ );
or   ( new_n4763_, new_n4761_, new_n4506_ );
and  ( new_n4764_, new_n4760_, new_n4513_ );
and  ( new_n4765_, new_n4511_, new_n4363_ );
and  ( new_n4766_, new_n4507_, new_n4502_ );
or   ( new_n4767_, new_n4766_, new_n4765_ );
and  ( new_n4768_, new_n4518_, new_n4166_ );
and  ( new_n4769_, new_n4514_, new_n4488_ );
or   ( new_n4770_, new_n4769_, new_n4768_ );
and  ( new_n4771_, new_n4525_, new_n4341_ );
and  ( new_n4772_, new_n4521_, new_n4475_ );
or   ( new_n4773_, new_n4772_, new_n4771_ );
and  ( new_n4774_, new_n4773_, new_n4770_ );
and  ( new_n4775_, new_n4544_, new_n4400_ );
and  ( new_n4776_, new_n4536_, new_n4215_ );
or   ( new_n4777_, new_n4776_, new_n4775_ );
and  ( new_n4778_, new_n4553_, new_n3695_ );
and  ( new_n4779_, new_n4549_, new_n3548_ );
or   ( new_n4780_, new_n4779_, new_n4778_ );
and  ( new_n4781_, new_n4780_, new_n4777_ );
or   ( new_n4782_, new_n4780_, new_n4777_ );
and  ( new_n4783_, new_n4564_, new_n3004_ );
and  ( new_n4784_, new_n4560_, new_n2868_ );
or   ( new_n4785_, new_n4784_, new_n4783_ );
and  ( new_n4786_, new_n4785_, new_n4782_ );
or   ( new_n4787_, new_n4786_, new_n4781_ );
and  ( new_n4788_, new_n4575_, new_n2334_ );
and  ( new_n4789_, new_n4571_, new_n2168_ );
or   ( new_n4790_, new_n4789_, new_n4788_ );
and  ( new_n4791_, new_n4584_, new_n1824_ );
and  ( new_n4792_, new_n4580_, new_n1717_ );
or   ( new_n4793_, new_n4792_, new_n4791_ );
and  ( new_n4794_, new_n4793_, new_n4790_ );
or   ( new_n4795_, new_n4793_, new_n4790_ );
and  ( new_n4796_, new_n4595_, new_n1355_ );
and  ( new_n4797_, new_n4591_, new_n1267_ );
or   ( new_n4798_, new_n4797_, new_n4796_ );
and  ( new_n4799_, new_n4798_, new_n4795_ );
or   ( new_n4800_, new_n4799_, new_n4794_ );
and  ( new_n4801_, new_n4800_, new_n4787_ );
or   ( new_n4802_, new_n4800_, new_n4787_ );
and  ( new_n4803_, new_n4608_, new_n913_ );
and  ( new_n4804_, new_n4604_, new_n938_ );
or   ( new_n4805_, new_n4804_, new_n4803_ );
and  ( new_n4806_, new_n4617_, new_n428_ );
and  ( new_n4807_, new_n4613_, new_n457_ );
or   ( new_n4808_, new_n4807_, new_n4806_ );
and  ( new_n4809_, new_n4808_, new_n4805_ );
or   ( new_n4810_, new_n4808_, new_n4805_ );
and  ( new_n4811_, new_n4628_, new_n505_ );
and  ( new_n4812_, new_n4624_, new_n533_ );
or   ( new_n4813_, new_n4812_, new_n4811_ );
and  ( new_n4814_, new_n4813_, new_n4810_ );
or   ( new_n4815_, new_n4814_, new_n4809_ );
and  ( new_n4816_, new_n4815_, new_n4802_ );
or   ( new_n4817_, new_n4816_, new_n4801_ );
and  ( new_n4818_, new_n4643_, new_n842_ );
and  ( new_n4819_, new_n4639_, new_n866_ );
or   ( new_n4820_, new_n4819_, new_n4818_ );
and  ( new_n4821_, new_n720_, RI2b1c4342e098_90 );
or   ( new_n4822_, new_n4821_, new_n4820_ );
and  ( new_n4823_, new_n4653_, new_n590_ );
and  ( new_n4824_, new_n4649_, new_n619_ );
or   ( new_n4825_, new_n4824_, new_n4823_ );
and  ( new_n4826_, new_n4662_, new_n734_ );
and  ( new_n4827_, new_n4658_, new_n762_ );
or   ( new_n4828_, new_n4827_, new_n4826_ );
and  ( new_n4829_, new_n4828_, new_n4825_ );
or   ( new_n4830_, new_n4828_, new_n4825_ );
and  ( new_n4831_, new_n4673_, new_n785_ );
and  ( new_n4832_, new_n4669_, new_n813_ );
or   ( new_n4833_, new_n4832_, new_n4831_ );
and  ( new_n4834_, new_n4833_, new_n4830_ );
or   ( new_n4835_, new_n4834_, new_n4829_ );
and  ( new_n4836_, new_n4835_, new_n4822_ );
or   ( new_n4837_, new_n4835_, new_n4822_ );
and  ( new_n4838_, new_n4686_, new_n842_ );
and  ( new_n4839_, new_n4682_, new_n866_ );
or   ( new_n4840_, new_n4839_, new_n4838_ );
and  ( new_n4841_, new_n4840_, new_n4837_ );
or   ( new_n4842_, new_n4841_, new_n4836_ );
and  ( new_n4843_, new_n4842_, new_n4817_ );
or   ( new_n4844_, new_n4842_, new_n4817_ );
and  ( new_n4845_, new_n720_, RI2b1c4342e020_89 );
and  ( new_n4846_, new_n4698_, new_n4301_ );
and  ( new_n4847_, new_n4694_, new_n4451_ );
or   ( new_n4848_, new_n4847_, new_n4846_ );
and  ( new_n4849_, new_n4848_, new_n4845_ );
or   ( new_n4850_, new_n4848_, new_n4845_ );
and  ( new_n4851_, new_n4707_, new_n4268_ );
and  ( new_n4852_, new_n4703_, new_n4436_ );
or   ( new_n4853_, new_n4852_, new_n4851_ );
and  ( new_n4854_, new_n4853_, new_n4850_ );
or   ( new_n4855_, new_n4854_, new_n4849_ );
and  ( new_n4856_, new_n4855_, new_n4844_ );
or   ( new_n4857_, new_n4856_, new_n4843_ );
and  ( new_n4858_, new_n4718_, new_n4339_ );
and  ( new_n4859_, new_n4714_, new_n4473_ );
or   ( new_n4860_, new_n4859_, new_n4858_ );
and  ( new_n4861_, new_n4725_, new_n4312_ );
and  ( new_n4862_, new_n4721_, new_n4458_ );
or   ( new_n4863_, new_n4862_, new_n4861_ );
and  ( new_n4864_, new_n4863_, new_n4860_ );
or   ( new_n4865_, new_n4863_, new_n4860_ );
and  ( new_n4866_, new_n4734_, new_n4270_ );
and  ( new_n4867_, new_n4730_, new_n4438_ );
or   ( new_n4868_, new_n4867_, new_n4866_ );
and  ( new_n4869_, new_n4868_, new_n4865_ );
or   ( new_n4870_, new_n4869_, new_n4864_ );
and  ( new_n4871_, new_n4870_, new_n4857_ );
or   ( new_n4872_, new_n4870_, new_n4857_ );
and  ( new_n4873_, new_n4745_, new_n3899_ );
and  ( new_n4874_, new_n4741_, new_n4063_ );
or   ( new_n4875_, new_n4874_, new_n4873_ );
and  ( new_n4876_, new_n4875_, new_n4872_ );
or   ( new_n4877_, new_n4876_, new_n4871_ );
and  ( new_n4878_, new_n4877_, new_n4774_ );
or   ( new_n4879_, new_n4877_, new_n4774_ );
and  ( new_n4880_, new_n4756_, new_n3967_ );
and  ( new_n4881_, new_n4752_, new_n4099_ );
or   ( new_n4882_, new_n4881_, new_n4880_ );
and  ( new_n4883_, new_n4882_, new_n4879_ );
or   ( new_n4884_, new_n4883_, new_n4878_ );
and  ( new_n4885_, new_n4884_, new_n4767_ );
or   ( new_n4886_, new_n4885_, new_n4764_ );
or   ( new_n4887_, new_n4491_, new_n4344_ );
and  ( new_n4888_, new_n4887_, new_n4352_ );
and  ( new_n4889_, new_n4477_, new_n4168_ );
and  ( new_n4890_, new_n4490_, new_n4343_ );
or   ( new_n4891_, new_n4890_, new_n4889_ );
and  ( new_n4892_, new_n4891_, new_n4495_ );
or   ( new_n4893_, new_n4892_, new_n4888_ );
and  ( new_n4894_, new_n4527_, new_n4520_ );
or   ( new_n4895_, new_n4894_, new_n4774_ );
or   ( new_n4896_, new_n4417_, new_n4187_ );
and  ( new_n4897_, new_n4896_, new_n4197_ );
and  ( new_n4898_, new_n4413_, new_n4186_ );
and  ( new_n4899_, new_n4416_, new_n4177_ );
or   ( new_n4900_, new_n4899_, new_n4898_ );
and  ( new_n4901_, new_n4900_, new_n4421_ );
or   ( new_n4902_, new_n4901_, new_n4897_ );
or   ( new_n4903_, new_n4404_, new_n4225_ );
and  ( new_n4904_, new_n4903_, new_n4235_ );
and  ( new_n4905_, new_n4400_, new_n4224_ );
and  ( new_n4906_, new_n4403_, new_n4215_ );
or   ( new_n4907_, new_n4906_, new_n4905_ );
and  ( new_n4908_, new_n4907_, new_n4408_ );
or   ( new_n4909_, new_n4908_, new_n4904_ );
and  ( new_n4910_, new_n4909_, new_n4902_ );
or   ( new_n4911_, new_n4909_, new_n4902_ );
or   ( new_n4912_, new_n4849_, new_n4701_ );
and  ( new_n4913_, new_n4912_, new_n4709_ );
and  ( new_n4914_, new_n4845_, new_n4700_ );
and  ( new_n4915_, new_n4848_, new_n4693_ );
or   ( new_n4916_, new_n4915_, new_n4914_ );
and  ( new_n4917_, new_n4916_, new_n4853_ );
or   ( new_n4918_, new_n4917_, new_n4913_ );
and  ( new_n4919_, new_n4918_, new_n4911_ );
or   ( new_n4920_, new_n4919_, new_n4910_ );
or   ( new_n4921_, new_n524_, new_n2119_ );
or   ( new_n4922_, new_n528_, new_n126_ );
and  ( new_n4923_, new_n4922_, new_n4921_ );
and  ( new_n4924_, new_n4923_, new_n505_ );
and  ( new_n4925_, new_n537_, RI2b1c4342dcd8_82 );
and  ( new_n4926_, new_n522_, RI2b1c4342dc60_81 );
or   ( new_n4927_, new_n4926_, new_n4925_ );
and  ( new_n4928_, new_n4927_, new_n533_ );
or   ( new_n4929_, new_n4928_, new_n4924_ );
or   ( new_n4930_, new_n610_, new_n2541_ );
or   ( new_n4931_, new_n614_, new_n121_ );
and  ( new_n4932_, new_n4931_, new_n4930_ );
and  ( new_n4933_, new_n4932_, new_n590_ );
and  ( new_n4934_, new_n623_, RI2b1c4342ddc8_84 );
and  ( new_n4935_, new_n608_, RI2b1c4342dd50_83 );
or   ( new_n4936_, new_n4935_, new_n4934_ );
and  ( new_n4937_, new_n4936_, new_n619_ );
or   ( new_n4938_, new_n4937_, new_n4933_ );
and  ( new_n4939_, new_n4938_, new_n4929_ );
or   ( new_n4940_, new_n4938_, new_n4929_ );
or   ( new_n4941_, new_n753_, new_n3239_ );
or   ( new_n4942_, new_n757_, new_n2806_ );
and  ( new_n4943_, new_n4942_, new_n4941_ );
and  ( new_n4944_, new_n4943_, new_n734_ );
and  ( new_n4945_, new_n766_, RI2b1c4342deb8_86 );
and  ( new_n4946_, new_n751_, RI2b1c4342de40_85 );
or   ( new_n4947_, new_n4946_, new_n4945_ );
and  ( new_n4948_, new_n4947_, new_n762_ );
or   ( new_n4949_, new_n4948_, new_n4944_ );
and  ( new_n4950_, new_n4949_, new_n4940_ );
or   ( new_n4951_, new_n4950_, new_n4939_ );
or   ( new_n4952_, new_n804_, new_n3902_ );
or   ( new_n4953_, new_n808_, new_n3924_ );
and  ( new_n4954_, new_n4953_, new_n4952_ );
and  ( new_n4955_, new_n4954_, new_n785_ );
and  ( new_n4956_, new_n817_, RI2b1c4342dfa8_88 );
and  ( new_n4957_, new_n802_, RI2b1c4342df30_87 );
or   ( new_n4958_, new_n4957_, new_n4956_ );
and  ( new_n4959_, new_n4958_, new_n813_ );
or   ( new_n4960_, new_n4959_, new_n4955_ );
or   ( new_n4961_, new_n857_, new_n4635_ );
or   ( new_n4962_, new_n861_, new_n132_ );
and  ( new_n4963_, new_n4962_, new_n4961_ );
and  ( new_n4964_, new_n4963_, new_n842_ );
and  ( new_n4965_, new_n870_, RI2b1c4342e098_90 );
and  ( new_n4966_, new_n855_, RI2b1c4342e020_89 );
or   ( new_n4967_, new_n4966_, new_n4965_ );
and  ( new_n4968_, new_n4967_, new_n866_ );
or   ( new_n4969_, new_n4968_, new_n4964_ );
and  ( new_n4970_, new_n4969_, new_n4960_ );
or   ( new_n4971_, new_n4969_, new_n4960_ );
or   ( new_n4972_, new_n841_, new_n117_ );
and  ( new_n4973_, new_n4972_, new_n4971_ );
or   ( new_n4974_, new_n4973_, new_n4970_ );
and  ( new_n4975_, new_n4974_, new_n4951_ );
or   ( new_n4976_, new_n4974_, new_n4951_ );
and  ( new_n4977_, new_n4820_, new_n4636_ );
and  ( new_n4978_, new_n4821_, new_n4645_ );
or   ( new_n4979_, new_n4978_, new_n4977_ );
and  ( new_n4980_, new_n4979_, new_n4976_ );
or   ( new_n4981_, new_n4980_, new_n4975_ );
or   ( new_n4982_, new_n3112_, new_n755_ );
or   ( new_n4983_, new_n3116_, new_n591_ );
and  ( new_n4984_, new_n4983_, new_n4982_ );
and  ( new_n4985_, new_n4984_, new_n3004_ );
and  ( new_n4986_, new_n3120_, RI2b1c4342d738_70 );
and  ( new_n4987_, new_n3110_, RI2b1c4342d6c0_69 );
or   ( new_n4988_, new_n4987_, new_n4986_ );
and  ( new_n4989_, new_n4988_, new_n2868_ );
or   ( new_n4990_, new_n4989_, new_n4985_ );
or   ( new_n4991_, new_n2450_, new_n806_ );
or   ( new_n4992_, new_n2454_, new_n110_ );
and  ( new_n4993_, new_n4992_, new_n4991_ );
and  ( new_n4994_, new_n4993_, new_n2334_ );
and  ( new_n4995_, new_n2458_, RI2b1c4342d828_72 );
and  ( new_n4996_, new_n2448_, RI2b1c4342d7b0_71 );
or   ( new_n4997_, new_n4996_, new_n4995_ );
and  ( new_n4998_, new_n4997_, new_n2168_ );
or   ( new_n4999_, new_n4998_, new_n4994_ );
and  ( new_n5000_, new_n4999_, new_n4990_ );
or   ( new_n5001_, new_n4999_, new_n4990_ );
or   ( new_n5002_, new_n1910_, new_n859_ );
or   ( new_n5003_, new_n1914_, new_n105_ );
and  ( new_n5004_, new_n5003_, new_n5002_ );
and  ( new_n5005_, new_n5004_, new_n1824_ );
and  ( new_n5006_, new_n1918_, RI2b1c4342d918_74 );
and  ( new_n5007_, new_n1908_, RI2b1c4342d8a0_73 );
or   ( new_n5008_, new_n5007_, new_n5006_ );
and  ( new_n5009_, new_n5008_, new_n1717_ );
or   ( new_n5010_, new_n5009_, new_n5005_ );
and  ( new_n5011_, new_n5010_, new_n5001_ );
or   ( new_n5012_, new_n5011_, new_n5000_ );
xor  ( new_n5013_, new_n325_, new_n200_ );
and  ( new_n5014_, new_n5013_, new_n342_ );
xor  ( new_n5015_, RI2b1c4342c400_29, RI2b1c4342d300_61 );
and  ( new_n5016_, new_n5015_, new_n218_ );
and  ( new_n5017_, new_n5016_, new_n138_ );
or   ( new_n5018_, new_n5017_, new_n201_ );
or   ( new_n5019_, new_n5018_, new_n5014_ );
xor  ( new_n5020_, new_n322_, new_n195_ );
and  ( new_n5021_, new_n5020_, new_n344_ );
xor  ( new_n5022_, RI2b1c4342c388_28, RI2b1c4342d288_60 );
and  ( new_n5023_, new_n5022_, new_n220_ );
and  ( new_n5024_, new_n5023_, new_n138_ );
or   ( new_n5025_, new_n5024_, new_n196_ );
or   ( new_n5026_, new_n5025_, new_n5021_ );
or   ( new_n5027_, new_n5026_, new_n5019_ );
and  ( new_n5028_, new_n5027_, new_n4394_ );
or   ( new_n5029_, new_n4535_, new_n526_ );
or   ( new_n5030_, new_n4539_, new_n99_ );
and  ( new_n5031_, new_n5030_, new_n5029_ );
and  ( new_n5032_, new_n5031_, new_n4400_ );
and  ( new_n5033_, new_n4543_, RI2b1c4342d558_66 );
and  ( new_n5034_, new_n4533_, RI2b1c4342d4e0_65 );
or   ( new_n5035_, new_n5034_, new_n5033_ );
and  ( new_n5036_, new_n5035_, new_n4215_ );
or   ( new_n5037_, new_n5036_, new_n5032_ );
and  ( new_n5038_, new_n5037_, new_n5028_ );
or   ( new_n5039_, new_n5037_, new_n5028_ );
or   ( new_n5040_, new_n3802_, new_n612_ );
or   ( new_n5041_, new_n3806_, new_n112_ );
and  ( new_n5042_, new_n5041_, new_n5040_ );
and  ( new_n5043_, new_n5042_, new_n3695_ );
and  ( new_n5044_, new_n3810_, RI2b1c4342d648_68 );
and  ( new_n5045_, new_n3800_, RI2b1c4342d5d0_67 );
or   ( new_n5046_, new_n5045_, new_n5044_ );
and  ( new_n5047_, new_n5046_, new_n3548_ );
or   ( new_n5048_, new_n5047_, new_n5043_ );
and  ( new_n5049_, new_n5048_, new_n5039_ );
or   ( new_n5050_, new_n5049_, new_n5038_ );
and  ( new_n5051_, new_n5050_, new_n5012_ );
or   ( new_n5052_, new_n5050_, new_n5012_ );
or   ( new_n5053_, new_n1425_, new_n886_ );
or   ( new_n5054_, new_n1429_, new_n843_ );
and  ( new_n5055_, new_n5054_, new_n5053_ );
and  ( new_n5056_, new_n5055_, new_n1355_ );
and  ( new_n5057_, new_n1433_, RI2b1c4342da08_76 );
and  ( new_n5058_, new_n1423_, RI2b1c4342d990_75 );
or   ( new_n5059_, new_n5058_, new_n5057_ );
and  ( new_n5060_, new_n5059_, new_n1267_ );
or   ( new_n5061_, new_n5060_, new_n5056_ );
or   ( new_n5062_, new_n934_, new_n1002_ );
or   ( new_n5063_, new_n940_, new_n1004_ );
and  ( new_n5064_, new_n5063_, new_n5062_ );
and  ( new_n5065_, new_n5064_, new_n913_ );
and  ( new_n5066_, new_n944_, RI2b1c4342daf8_78 );
and  ( new_n5067_, new_n932_, RI2b1c4342da80_77 );
or   ( new_n5068_, new_n5067_, new_n5066_ );
and  ( new_n5069_, new_n5068_, new_n938_ );
or   ( new_n5070_, new_n5069_, new_n5065_ );
and  ( new_n5071_, new_n5070_, new_n5061_ );
or   ( new_n5072_, new_n5070_, new_n5061_ );
or   ( new_n5073_, new_n453_, new_n1511_ );
or   ( new_n5074_, new_n459_, new_n1310_ );
and  ( new_n5075_, new_n5074_, new_n5073_ );
and  ( new_n5076_, new_n5075_, new_n428_ );
and  ( new_n5077_, new_n463_, RI2b1c4342dbe8_80 );
and  ( new_n5078_, new_n451_, RI2b1c4342db70_79 );
or   ( new_n5079_, new_n5078_, new_n5077_ );
and  ( new_n5080_, new_n5079_, new_n457_ );
or   ( new_n5081_, new_n5080_, new_n5076_ );
and  ( new_n5082_, new_n5081_, new_n5072_ );
or   ( new_n5083_, new_n5082_, new_n5071_ );
and  ( new_n5084_, new_n5083_, new_n5052_ );
or   ( new_n5085_, new_n5084_, new_n5051_ );
and  ( new_n5086_, new_n5085_, new_n4981_ );
or   ( new_n5087_, new_n5085_, new_n4981_ );
or   ( new_n5088_, new_n4829_, new_n4665_ );
and  ( new_n5089_, new_n5088_, new_n4675_ );
and  ( new_n5090_, new_n4825_, new_n4664_ );
and  ( new_n5091_, new_n4828_, new_n4655_ );
or   ( new_n5092_, new_n5091_, new_n5090_ );
and  ( new_n5093_, new_n5092_, new_n4833_ );
or   ( new_n5094_, new_n5093_, new_n5089_ );
or   ( new_n5095_, new_n4809_, new_n4620_ );
and  ( new_n5096_, new_n5095_, new_n4630_ );
and  ( new_n5097_, new_n4805_, new_n4619_ );
and  ( new_n5098_, new_n4808_, new_n4610_ );
or   ( new_n5099_, new_n5098_, new_n5097_ );
and  ( new_n5100_, new_n5099_, new_n4813_ );
or   ( new_n5101_, new_n5100_, new_n5096_ );
and  ( new_n5102_, new_n5101_, new_n5094_ );
or   ( new_n5103_, new_n5101_, new_n5094_ );
or   ( new_n5104_, new_n4794_, new_n4587_ );
and  ( new_n5105_, new_n5104_, new_n4597_ );
and  ( new_n5106_, new_n4790_, new_n4586_ );
and  ( new_n5107_, new_n4793_, new_n4577_ );
or   ( new_n5108_, new_n5107_, new_n5106_ );
and  ( new_n5109_, new_n5108_, new_n4798_ );
or   ( new_n5110_, new_n5109_, new_n5105_ );
and  ( new_n5111_, new_n5110_, new_n5103_ );
or   ( new_n5112_, new_n5111_, new_n5102_ );
and  ( new_n5113_, new_n5112_, new_n5087_ );
or   ( new_n5114_, new_n5113_, new_n5086_ );
and  ( new_n5115_, new_n5114_, new_n4920_ );
or   ( new_n5116_, new_n5114_, new_n4920_ );
or   ( new_n5117_, new_n4864_, new_n4728_ );
and  ( new_n5118_, new_n5117_, new_n4736_ );
and  ( new_n5119_, new_n4860_, new_n4727_ );
and  ( new_n5120_, new_n4863_, new_n4720_ );
or   ( new_n5121_, new_n5120_, new_n5119_ );
and  ( new_n5122_, new_n5121_, new_n4868_ );
or   ( new_n5123_, new_n5122_, new_n5118_ );
and  ( new_n5124_, new_n5123_, new_n5116_ );
or   ( new_n5125_, new_n5124_, new_n5115_ );
and  ( new_n5126_, new_n5125_, new_n4895_ );
or   ( new_n5127_, new_n5125_, new_n4895_ );
or   ( new_n5128_, new_n4871_, new_n4739_ );
and  ( new_n5129_, new_n5128_, new_n4747_ );
and  ( new_n5130_, new_n4857_, new_n4738_ );
and  ( new_n5131_, new_n4870_, new_n4713_ );
or   ( new_n5132_, new_n5131_, new_n5130_ );
and  ( new_n5133_, new_n5132_, new_n4875_ );
or   ( new_n5134_, new_n5133_, new_n5129_ );
and  ( new_n5135_, new_n5134_, new_n5127_ );
or   ( new_n5136_, new_n5135_, new_n5126_ );
and  ( new_n5137_, new_n5136_, new_n4893_ );
or   ( new_n5138_, new_n5136_, new_n4893_ );
or   ( new_n5139_, new_n4878_, new_n4750_ );
and  ( new_n5140_, new_n5139_, new_n4758_ );
and  ( new_n5141_, new_n4877_, new_n4528_ );
and  ( new_n5142_, new_n4774_, new_n4749_ );
or   ( new_n5143_, new_n5142_, new_n5141_ );
and  ( new_n5144_, new_n5143_, new_n4882_ );
or   ( new_n5145_, new_n5144_, new_n5140_ );
and  ( new_n5146_, new_n5145_, new_n5138_ );
or   ( new_n5147_, new_n5146_, new_n5137_ );
or   ( new_n5148_, new_n5147_, new_n4886_ );
and  ( new_n5149_, new_n5148_, new_n4763_ );
or   ( new_n5150_, new_n5149_, new_n4762_ );
and  ( new_n5151_, new_n5147_, new_n4886_ );
or   ( new_n5152_, new_n5151_, new_n4762_ );
and  ( new_n5153_, new_n4891_, new_n4352_ );
and  ( new_n5154_, new_n4887_, new_n4495_ );
or   ( new_n5155_, new_n5154_, new_n5153_ );
and  ( new_n5156_, new_n4770_, new_n4527_ );
and  ( new_n5157_, new_n4773_, new_n4520_ );
or   ( new_n5158_, new_n5157_, new_n5156_ );
and  ( new_n5159_, new_n4900_, new_n4197_ );
and  ( new_n5160_, new_n4896_, new_n4421_ );
or   ( new_n5161_, new_n5160_, new_n5159_ );
and  ( new_n5162_, new_n4907_, new_n4235_ );
and  ( new_n5163_, new_n4903_, new_n4408_ );
or   ( new_n5164_, new_n5163_, new_n5162_ );
and  ( new_n5165_, new_n5164_, new_n5161_ );
or   ( new_n5166_, new_n5164_, new_n5161_ );
and  ( new_n5167_, new_n4916_, new_n4709_ );
and  ( new_n5168_, new_n4912_, new_n4853_ );
or   ( new_n5169_, new_n5168_, new_n5167_ );
and  ( new_n5170_, new_n5169_, new_n5166_ );
or   ( new_n5171_, new_n5170_, new_n5165_ );
not  ( new_n5172_, new_n218_ );
nor  ( new_n5173_, new_n5015_, new_n5172_ );
and  ( new_n5174_, new_n5015_, new_n342_ );
or   ( new_n5175_, new_n5174_, new_n5173_ );
and  ( new_n5176_, new_n5175_, new_n325_ );
nor  ( new_n5177_, new_n5022_, new_n221_ );
and  ( new_n5178_, new_n5022_, new_n344_ );
or   ( new_n5179_, new_n5178_, new_n5177_ );
and  ( new_n5180_, new_n5179_, new_n322_ );
and  ( new_n5181_, new_n5180_, new_n5176_ );
or   ( new_n5182_, new_n5181_, new_n4206_ );
and  ( new_n5183_, new_n5035_, new_n4400_ );
and  ( new_n5184_, new_n5031_, new_n4215_ );
or   ( new_n5185_, new_n5184_, new_n5183_ );
and  ( new_n5186_, new_n5185_, new_n5182_ );
or   ( new_n5187_, new_n5185_, new_n5182_ );
and  ( new_n5188_, new_n5046_, new_n3695_ );
and  ( new_n5189_, new_n5042_, new_n3548_ );
or   ( new_n5190_, new_n5189_, new_n5188_ );
and  ( new_n5191_, new_n5190_, new_n5187_ );
or   ( new_n5192_, new_n5191_, new_n5186_ );
and  ( new_n5193_, new_n4988_, new_n3004_ );
and  ( new_n5194_, new_n4984_, new_n2868_ );
or   ( new_n5195_, new_n5194_, new_n5193_ );
and  ( new_n5196_, new_n4997_, new_n2334_ );
and  ( new_n5197_, new_n4993_, new_n2168_ );
or   ( new_n5198_, new_n5197_, new_n5196_ );
and  ( new_n5199_, new_n5198_, new_n5195_ );
or   ( new_n5200_, new_n5198_, new_n5195_ );
and  ( new_n5201_, new_n5008_, new_n1824_ );
and  ( new_n5202_, new_n5004_, new_n1717_ );
or   ( new_n5203_, new_n5202_, new_n5201_ );
and  ( new_n5204_, new_n5203_, new_n5200_ );
or   ( new_n5205_, new_n5204_, new_n5199_ );
and  ( new_n5206_, new_n5205_, new_n5192_ );
or   ( new_n5207_, new_n5205_, new_n5192_ );
and  ( new_n5208_, new_n5059_, new_n1355_ );
and  ( new_n5209_, new_n5055_, new_n1267_ );
or   ( new_n5210_, new_n5209_, new_n5208_ );
and  ( new_n5211_, new_n5068_, new_n913_ );
and  ( new_n5212_, new_n5064_, new_n938_ );
or   ( new_n5213_, new_n5212_, new_n5211_ );
and  ( new_n5214_, new_n5213_, new_n5210_ );
or   ( new_n5215_, new_n5213_, new_n5210_ );
and  ( new_n5216_, new_n5079_, new_n428_ );
and  ( new_n5217_, new_n5075_, new_n457_ );
or   ( new_n5218_, new_n5217_, new_n5216_ );
and  ( new_n5219_, new_n5218_, new_n5215_ );
or   ( new_n5220_, new_n5219_, new_n5214_ );
and  ( new_n5221_, new_n5220_, new_n5207_ );
or   ( new_n5222_, new_n5221_, new_n5206_ );
and  ( new_n5223_, new_n4927_, new_n505_ );
and  ( new_n5224_, new_n4923_, new_n533_ );
or   ( new_n5225_, new_n5224_, new_n5223_ );
and  ( new_n5226_, new_n4936_, new_n590_ );
and  ( new_n5227_, new_n4932_, new_n619_ );
or   ( new_n5228_, new_n5227_, new_n5226_ );
and  ( new_n5229_, new_n5228_, new_n5225_ );
or   ( new_n5230_, new_n5228_, new_n5225_ );
and  ( new_n5231_, new_n4947_, new_n734_ );
and  ( new_n5232_, new_n4943_, new_n762_ );
or   ( new_n5233_, new_n5232_, new_n5231_ );
and  ( new_n5234_, new_n5233_, new_n5230_ );
or   ( new_n5235_, new_n5234_, new_n5229_ );
and  ( new_n5236_, new_n4958_, new_n785_ );
and  ( new_n5237_, new_n4954_, new_n813_ );
or   ( new_n5238_, new_n5237_, new_n5236_ );
and  ( new_n5239_, new_n4967_, new_n842_ );
and  ( new_n5240_, new_n4963_, new_n866_ );
or   ( new_n5241_, new_n5240_, new_n5239_ );
or   ( new_n5242_, new_n5241_, new_n5238_ );
and  ( new_n5243_, new_n5241_, new_n5238_ );
and  ( new_n5244_, new_n720_, RI2b1c4342e110_91 );
or   ( new_n5245_, new_n5244_, new_n5243_ );
and  ( new_n5246_, new_n5245_, new_n5242_ );
or   ( new_n5247_, new_n5246_, new_n5235_ );
and  ( new_n5248_, new_n5246_, new_n5235_ );
and  ( new_n5249_, new_n4821_, new_n4820_ );
or   ( new_n5250_, new_n5249_, new_n4646_ );
or   ( new_n5251_, new_n5250_, new_n5248_ );
and  ( new_n5252_, new_n5251_, new_n5247_ );
or   ( new_n5253_, new_n5252_, new_n5222_ );
and  ( new_n5254_, new_n5252_, new_n5222_ );
and  ( new_n5255_, new_n5092_, new_n4675_ );
and  ( new_n5256_, new_n5088_, new_n4833_ );
or   ( new_n5257_, new_n5256_, new_n5255_ );
and  ( new_n5258_, new_n5099_, new_n4630_ );
and  ( new_n5259_, new_n5095_, new_n4813_ );
or   ( new_n5260_, new_n5259_, new_n5258_ );
and  ( new_n5261_, new_n5260_, new_n5257_ );
or   ( new_n5262_, new_n5260_, new_n5257_ );
and  ( new_n5263_, new_n5108_, new_n4597_ );
and  ( new_n5264_, new_n5104_, new_n4798_ );
or   ( new_n5265_, new_n5264_, new_n5263_ );
and  ( new_n5266_, new_n5265_, new_n5262_ );
or   ( new_n5267_, new_n5266_, new_n5261_ );
or   ( new_n5268_, new_n5267_, new_n5254_ );
and  ( new_n5269_, new_n5268_, new_n5253_ );
or   ( new_n5270_, new_n5269_, new_n5171_ );
and  ( new_n5271_, new_n5269_, new_n5171_ );
and  ( new_n5272_, new_n5121_, new_n4736_ );
and  ( new_n5273_, new_n5117_, new_n4868_ );
or   ( new_n5274_, new_n5273_, new_n5272_ );
or   ( new_n5275_, new_n5274_, new_n5271_ );
and  ( new_n5276_, new_n5275_, new_n5270_ );
or   ( new_n5277_, new_n5276_, new_n5158_ );
and  ( new_n5278_, new_n5276_, new_n5158_ );
and  ( new_n5279_, new_n5132_, new_n4747_ );
and  ( new_n5280_, new_n5128_, new_n4875_ );
or   ( new_n5281_, new_n5280_, new_n5279_ );
or   ( new_n5282_, new_n5281_, new_n5278_ );
and  ( new_n5283_, new_n5282_, new_n5277_ );
and  ( new_n5284_, new_n5283_, new_n5155_ );
or   ( new_n5285_, new_n5284_, new_n5137_ );
and  ( new_n5286_, new_n5285_, new_n5145_ );
and  ( new_n5287_, new_n5283_, new_n4893_ );
and  ( new_n5288_, new_n5155_, new_n5136_ );
or   ( new_n5289_, new_n5288_, new_n5287_ );
and  ( new_n5290_, new_n5143_, new_n4758_ );
and  ( new_n5291_, new_n5139_, new_n4882_ );
or   ( new_n5292_, new_n5291_, new_n5290_ );
and  ( new_n5293_, new_n5292_, new_n5289_ );
or   ( new_n5294_, new_n5293_, new_n5286_ );
or   ( new_n5295_, new_n5278_, new_n5126_ );
and  ( new_n5296_, new_n5295_, new_n5134_ );
and  ( new_n5297_, new_n5276_, new_n4895_ );
and  ( new_n5298_, new_n5158_, new_n5125_ );
or   ( new_n5299_, new_n5298_, new_n5297_ );
and  ( new_n5300_, new_n5299_, new_n5281_ );
or   ( new_n5301_, new_n5300_, new_n5296_ );
and  ( new_n5302_, new_n5180_, new_n4394_ );
and  ( new_n5303_, new_n5026_, new_n4206_ );
and  ( new_n5304_, new_n5180_, new_n5019_ );
and  ( new_n5305_, new_n5176_, new_n5026_ );
or   ( new_n5306_, new_n5305_, new_n5304_ );
or   ( new_n5307_, new_n5306_, new_n5303_ );
or   ( new_n5308_, new_n5307_, new_n5302_ );
or   ( new_n5309_, new_n5308_, new_n99_ );
and  ( new_n5310_, new_n5309_, new_n5182_ );
and  ( new_n5311_, new_n5026_, new_n5019_ );
or   ( new_n5312_, new_n5311_, new_n5181_ );
and  ( new_n5313_, new_n5026_, new_n4394_ );
and  ( new_n5314_, new_n5180_, new_n4206_ );
or   ( new_n5315_, new_n5314_, new_n5313_ );
and  ( new_n5316_, new_n5315_, new_n5312_ );
and  ( new_n5317_, new_n5316_, RI2b1c4342d4e0_65 );
and  ( new_n5318_, new_n5317_, new_n5028_ );
or   ( new_n5319_, new_n5318_, new_n5310_ );
or   ( new_n5320_, new_n4535_, new_n112_ );
or   ( new_n5321_, new_n4539_, new_n526_ );
and  ( new_n5322_, new_n5321_, new_n5320_ );
and  ( new_n5323_, new_n5322_, new_n4400_ );
and  ( new_n5324_, new_n4543_, RI2b1c4342d5d0_67 );
and  ( new_n5325_, new_n4533_, RI2b1c4342d558_66 );
or   ( new_n5326_, new_n5325_, new_n5324_ );
and  ( new_n5327_, new_n5326_, new_n4215_ );
or   ( new_n5328_, new_n5327_, new_n5323_ );
and  ( new_n5329_, new_n5328_, new_n5319_ );
or   ( new_n5330_, new_n5328_, new_n5319_ );
or   ( new_n5331_, new_n3802_, new_n591_ );
or   ( new_n5332_, new_n3806_, new_n612_ );
and  ( new_n5333_, new_n5332_, new_n5331_ );
and  ( new_n5334_, new_n5333_, new_n3695_ );
and  ( new_n5335_, new_n3810_, RI2b1c4342d6c0_69 );
and  ( new_n5336_, new_n3800_, RI2b1c4342d648_68 );
or   ( new_n5337_, new_n5336_, new_n5335_ );
and  ( new_n5338_, new_n5337_, new_n3548_ );
or   ( new_n5339_, new_n5338_, new_n5334_ );
and  ( new_n5340_, new_n5339_, new_n5330_ );
or   ( new_n5341_, new_n5340_, new_n5329_ );
or   ( new_n5342_, new_n3112_, new_n110_ );
or   ( new_n5343_, new_n3116_, new_n755_ );
and  ( new_n5344_, new_n5343_, new_n5342_ );
and  ( new_n5345_, new_n5344_, new_n3004_ );
and  ( new_n5346_, new_n3120_, RI2b1c4342d7b0_71 );
and  ( new_n5347_, new_n3110_, RI2b1c4342d738_70 );
or   ( new_n5348_, new_n5347_, new_n5346_ );
and  ( new_n5349_, new_n5348_, new_n2868_ );
or   ( new_n5350_, new_n5349_, new_n5345_ );
or   ( new_n5351_, new_n2450_, new_n105_ );
or   ( new_n5352_, new_n2454_, new_n806_ );
and  ( new_n5353_, new_n5352_, new_n5351_ );
and  ( new_n5354_, new_n5353_, new_n2334_ );
and  ( new_n5355_, new_n2458_, RI2b1c4342d8a0_73 );
and  ( new_n5356_, new_n2448_, RI2b1c4342d828_72 );
or   ( new_n5357_, new_n5356_, new_n5355_ );
and  ( new_n5358_, new_n5357_, new_n2168_ );
or   ( new_n5359_, new_n5358_, new_n5354_ );
and  ( new_n5360_, new_n5359_, new_n5350_ );
or   ( new_n5361_, new_n5359_, new_n5350_ );
or   ( new_n5362_, new_n1910_, new_n843_ );
or   ( new_n5363_, new_n1914_, new_n859_ );
and  ( new_n5364_, new_n5363_, new_n5362_ );
and  ( new_n5365_, new_n5364_, new_n1824_ );
and  ( new_n5366_, new_n1918_, RI2b1c4342d990_75 );
and  ( new_n5367_, new_n1908_, RI2b1c4342d918_74 );
or   ( new_n5368_, new_n5367_, new_n5366_ );
and  ( new_n5369_, new_n5368_, new_n1717_ );
or   ( new_n5370_, new_n5369_, new_n5365_ );
and  ( new_n5371_, new_n5370_, new_n5361_ );
or   ( new_n5372_, new_n5371_, new_n5360_ );
and  ( new_n5373_, new_n5372_, new_n5341_ );
or   ( new_n5374_, new_n5372_, new_n5341_ );
or   ( new_n5375_, new_n1425_, new_n1004_ );
or   ( new_n5376_, new_n1429_, new_n886_ );
and  ( new_n5377_, new_n5376_, new_n5375_ );
and  ( new_n5378_, new_n5377_, new_n1355_ );
and  ( new_n5379_, new_n1433_, RI2b1c4342da80_77 );
and  ( new_n5380_, new_n1423_, RI2b1c4342da08_76 );
or   ( new_n5381_, new_n5380_, new_n5379_ );
and  ( new_n5382_, new_n5381_, new_n1267_ );
or   ( new_n5383_, new_n5382_, new_n5378_ );
or   ( new_n5384_, new_n934_, new_n1310_ );
or   ( new_n5385_, new_n940_, new_n1002_ );
and  ( new_n5386_, new_n5385_, new_n5384_ );
and  ( new_n5387_, new_n5386_, new_n913_ );
and  ( new_n5388_, new_n944_, RI2b1c4342db70_79 );
and  ( new_n5389_, new_n932_, RI2b1c4342daf8_78 );
or   ( new_n5390_, new_n5389_, new_n5388_ );
and  ( new_n5391_, new_n5390_, new_n938_ );
or   ( new_n5392_, new_n5391_, new_n5387_ );
and  ( new_n5393_, new_n5392_, new_n5383_ );
or   ( new_n5394_, new_n5392_, new_n5383_ );
or   ( new_n5395_, new_n453_, new_n126_ );
or   ( new_n5396_, new_n459_, new_n1511_ );
and  ( new_n5397_, new_n5396_, new_n5395_ );
and  ( new_n5398_, new_n5397_, new_n428_ );
and  ( new_n5399_, new_n463_, RI2b1c4342dc60_81 );
and  ( new_n5400_, new_n451_, RI2b1c4342dbe8_80 );
or   ( new_n5401_, new_n5400_, new_n5399_ );
and  ( new_n5402_, new_n5401_, new_n457_ );
or   ( new_n5403_, new_n5402_, new_n5398_ );
and  ( new_n5404_, new_n5403_, new_n5394_ );
or   ( new_n5405_, new_n5404_, new_n5393_ );
and  ( new_n5406_, new_n5405_, new_n5374_ );
or   ( new_n5407_, new_n5406_, new_n5373_ );
or   ( new_n5408_, new_n524_, new_n121_ );
or   ( new_n5409_, new_n528_, new_n2119_ );
and  ( new_n5410_, new_n5409_, new_n5408_ );
and  ( new_n5411_, new_n5410_, new_n505_ );
and  ( new_n5412_, new_n537_, RI2b1c4342dd50_83 );
and  ( new_n5413_, new_n522_, RI2b1c4342dcd8_82 );
or   ( new_n5414_, new_n5413_, new_n5412_ );
and  ( new_n5415_, new_n5414_, new_n533_ );
or   ( new_n5416_, new_n5415_, new_n5411_ );
or   ( new_n5417_, new_n610_, new_n2806_ );
or   ( new_n5418_, new_n614_, new_n2541_ );
and  ( new_n5419_, new_n5418_, new_n5417_ );
and  ( new_n5420_, new_n5419_, new_n590_ );
and  ( new_n5421_, new_n623_, RI2b1c4342de40_85 );
and  ( new_n5422_, new_n608_, RI2b1c4342ddc8_84 );
or   ( new_n5423_, new_n5422_, new_n5421_ );
and  ( new_n5424_, new_n5423_, new_n619_ );
or   ( new_n5425_, new_n5424_, new_n5420_ );
and  ( new_n5426_, new_n5425_, new_n5416_ );
or   ( new_n5427_, new_n5425_, new_n5416_ );
or   ( new_n5428_, new_n753_, new_n3924_ );
or   ( new_n5429_, new_n757_, new_n3239_ );
and  ( new_n5430_, new_n5429_, new_n5428_ );
and  ( new_n5431_, new_n5430_, new_n734_ );
and  ( new_n5432_, new_n766_, RI2b1c4342df30_87 );
and  ( new_n5433_, new_n751_, RI2b1c4342deb8_86 );
or   ( new_n5434_, new_n5433_, new_n5432_ );
and  ( new_n5435_, new_n5434_, new_n762_ );
or   ( new_n5436_, new_n5435_, new_n5431_ );
and  ( new_n5437_, new_n5436_, new_n5427_ );
or   ( new_n5438_, new_n5437_, new_n5426_ );
or   ( new_n5439_, new_n804_, new_n132_ );
or   ( new_n5440_, new_n808_, new_n3902_ );
and  ( new_n5441_, new_n5440_, new_n5439_ );
and  ( new_n5442_, new_n5441_, new_n785_ );
and  ( new_n5443_, new_n817_, RI2b1c4342e020_89 );
and  ( new_n5444_, new_n802_, RI2b1c4342dfa8_88 );
or   ( new_n5445_, new_n5444_, new_n5443_ );
and  ( new_n5446_, new_n5445_, new_n813_ );
or   ( new_n5447_, new_n5446_, new_n5442_ );
or   ( new_n5448_, new_n857_, new_n117_ );
or   ( new_n5449_, new_n861_, new_n4635_ );
and  ( new_n5450_, new_n5449_, new_n5448_ );
and  ( new_n5451_, new_n5450_, new_n842_ );
and  ( new_n5452_, new_n870_, RI2b1c4342e110_91 );
and  ( new_n5453_, new_n855_, RI2b1c4342e098_90 );
or   ( new_n5454_, new_n5453_, new_n5452_ );
and  ( new_n5455_, new_n5454_, new_n866_ );
or   ( new_n5456_, new_n5455_, new_n5451_ );
and  ( new_n5457_, new_n5456_, new_n5447_ );
or   ( new_n5458_, new_n5456_, new_n5447_ );
not  ( new_n5459_, RI2b1c4342e188_92 );
or   ( new_n5460_, new_n841_, new_n5459_ );
and  ( new_n5461_, new_n5460_, new_n5458_ );
or   ( new_n5462_, new_n5461_, new_n5457_ );
and  ( new_n5463_, new_n5462_, new_n5438_ );
or   ( new_n5464_, new_n5462_, new_n5438_ );
or   ( new_n5465_, new_n5243_, new_n4970_ );
and  ( new_n5466_, new_n5465_, new_n4972_ );
and  ( new_n5467_, new_n5238_, new_n4969_ );
and  ( new_n5468_, new_n5241_, new_n4960_ );
or   ( new_n5469_, new_n5468_, new_n5467_ );
and  ( new_n5470_, new_n5469_, new_n5244_ );
or   ( new_n5471_, new_n5470_, new_n5466_ );
and  ( new_n5472_, new_n5471_, new_n5464_ );
or   ( new_n5473_, new_n5472_, new_n5463_ );
and  ( new_n5474_, new_n5473_, new_n5407_ );
or   ( new_n5475_, new_n5473_, new_n5407_ );
or   ( new_n5476_, new_n5229_, new_n4939_ );
and  ( new_n5477_, new_n5476_, new_n4949_ );
and  ( new_n5478_, new_n5225_, new_n4938_ );
and  ( new_n5479_, new_n5228_, new_n4929_ );
or   ( new_n5480_, new_n5479_, new_n5478_ );
and  ( new_n5481_, new_n5480_, new_n5233_ );
or   ( new_n5482_, new_n5481_, new_n5477_ );
or   ( new_n5483_, new_n5214_, new_n5071_ );
and  ( new_n5484_, new_n5483_, new_n5081_ );
and  ( new_n5485_, new_n5210_, new_n5070_ );
and  ( new_n5486_, new_n5213_, new_n5061_ );
or   ( new_n5487_, new_n5486_, new_n5485_ );
and  ( new_n5488_, new_n5487_, new_n5218_ );
or   ( new_n5489_, new_n5488_, new_n5484_ );
and  ( new_n5490_, new_n5489_, new_n5482_ );
or   ( new_n5491_, new_n5489_, new_n5482_ );
or   ( new_n5492_, new_n5199_, new_n5000_ );
and  ( new_n5493_, new_n5492_, new_n5010_ );
and  ( new_n5494_, new_n5195_, new_n4999_ );
and  ( new_n5495_, new_n5198_, new_n4990_ );
or   ( new_n5496_, new_n5495_, new_n5494_ );
and  ( new_n5497_, new_n5496_, new_n5203_ );
or   ( new_n5498_, new_n5497_, new_n5493_ );
and  ( new_n5499_, new_n5498_, new_n5491_ );
or   ( new_n5500_, new_n5499_, new_n5490_ );
and  ( new_n5501_, new_n5500_, new_n5475_ );
or   ( new_n5502_, new_n5501_, new_n5474_ );
or   ( new_n5503_, new_n4781_, new_n4556_ );
and  ( new_n5504_, new_n5503_, new_n4566_ );
and  ( new_n5505_, new_n4777_, new_n4555_ );
and  ( new_n5506_, new_n4780_, new_n4546_ );
or   ( new_n5507_, new_n5506_, new_n5505_ );
and  ( new_n5508_, new_n5507_, new_n4785_ );
or   ( new_n5509_, new_n5508_, new_n5504_ );
or   ( new_n5510_, new_n5261_, new_n5102_ );
and  ( new_n5511_, new_n5510_, new_n5110_ );
and  ( new_n5512_, new_n5257_, new_n5101_ );
and  ( new_n5513_, new_n5260_, new_n5094_ );
or   ( new_n5514_, new_n5513_, new_n5512_ );
and  ( new_n5515_, new_n5514_, new_n5265_ );
or   ( new_n5516_, new_n5515_, new_n5511_ );
and  ( new_n5517_, new_n5516_, new_n5509_ );
or   ( new_n5518_, new_n5516_, new_n5509_ );
or   ( new_n5519_, new_n5248_, new_n4975_ );
and  ( new_n5520_, new_n5519_, new_n4979_ );
and  ( new_n5521_, new_n5235_, new_n4974_ );
and  ( new_n5522_, new_n5246_, new_n4951_ );
or   ( new_n5523_, new_n5522_, new_n5521_ );
and  ( new_n5524_, new_n5523_, new_n5250_ );
or   ( new_n5525_, new_n5524_, new_n5520_ );
and  ( new_n5526_, new_n5525_, new_n5518_ );
or   ( new_n5527_, new_n5526_, new_n5517_ );
and  ( new_n5528_, new_n5527_, new_n5502_ );
or   ( new_n5529_, new_n5527_, new_n5502_ );
or   ( new_n5530_, new_n4836_, new_n4678_ );
and  ( new_n5531_, new_n5530_, new_n4688_ );
and  ( new_n5532_, new_n4835_, new_n4646_ );
and  ( new_n5533_, new_n4822_, new_n4677_ );
or   ( new_n5534_, new_n5533_, new_n5532_ );
and  ( new_n5535_, new_n5534_, new_n4840_ );
or   ( new_n5536_, new_n5535_, new_n5531_ );
and  ( new_n5537_, new_n5536_, new_n5529_ );
or   ( new_n5538_, new_n5537_, new_n5528_ );
or   ( new_n5539_, new_n4801_, new_n4600_ );
and  ( new_n5540_, new_n5539_, new_n4632_ );
and  ( new_n5541_, new_n4787_, new_n4599_ );
and  ( new_n5542_, new_n4800_, new_n4568_ );
or   ( new_n5543_, new_n5542_, new_n5541_ );
and  ( new_n5544_, new_n5543_, new_n4815_ );
or   ( new_n5545_, new_n5544_, new_n5540_ );
or   ( new_n5546_, new_n5165_, new_n4910_ );
and  ( new_n5547_, new_n5546_, new_n4918_ );
and  ( new_n5548_, new_n5161_, new_n4909_ );
and  ( new_n5549_, new_n5164_, new_n4902_ );
or   ( new_n5550_, new_n5549_, new_n5548_ );
and  ( new_n5551_, new_n5550_, new_n5169_ );
or   ( new_n5552_, new_n5551_, new_n5547_ );
and  ( new_n5553_, new_n5552_, new_n5545_ );
or   ( new_n5554_, new_n5552_, new_n5545_ );
or   ( new_n5555_, new_n5254_, new_n5086_ );
and  ( new_n5556_, new_n5555_, new_n5112_ );
and  ( new_n5557_, new_n5222_, new_n4981_ );
and  ( new_n5558_, new_n5252_, new_n5085_ );
or   ( new_n5559_, new_n5558_, new_n5557_ );
and  ( new_n5560_, new_n5559_, new_n5267_ );
or   ( new_n5561_, new_n5560_, new_n5556_ );
and  ( new_n5562_, new_n5561_, new_n5554_ );
or   ( new_n5563_, new_n5562_, new_n5553_ );
and  ( new_n5564_, new_n5563_, new_n5538_ );
or   ( new_n5565_, new_n5563_, new_n5538_ );
or   ( new_n5566_, new_n4843_, new_n4691_ );
and  ( new_n5567_, new_n5566_, new_n4711_ );
and  ( new_n5568_, new_n4817_, new_n4690_ );
and  ( new_n5569_, new_n4842_, new_n4634_ );
or   ( new_n5570_, new_n5569_, new_n5568_ );
and  ( new_n5571_, new_n5570_, new_n4855_ );
or   ( new_n5572_, new_n5571_, new_n5567_ );
and  ( new_n5573_, new_n5572_, new_n5565_ );
or   ( new_n5574_, new_n5573_, new_n5564_ );
or   ( new_n5575_, new_n5574_, new_n5301_ );
and  ( new_n5576_, new_n5575_, new_n5294_ );
or   ( new_n5577_, new_n5575_, new_n5294_ );
and  ( new_n5578_, new_n5574_, new_n5301_ );
and  ( new_n5579_, new_n5299_, new_n5134_ );
and  ( new_n5580_, new_n5295_, new_n5281_ );
or   ( new_n5581_, new_n5580_, new_n5579_ );
and  ( new_n5582_, new_n5543_, new_n4632_ );
and  ( new_n5583_, new_n5539_, new_n4815_ );
or   ( new_n5584_, new_n5583_, new_n5582_ );
and  ( new_n5585_, new_n5550_, new_n4918_ );
and  ( new_n5586_, new_n5546_, new_n5169_ );
or   ( new_n5587_, new_n5586_, new_n5585_ );
and  ( new_n5588_, new_n5587_, new_n5584_ );
or   ( new_n5589_, new_n5587_, new_n5584_ );
and  ( new_n5590_, new_n5559_, new_n5112_ );
and  ( new_n5591_, new_n5555_, new_n5267_ );
or   ( new_n5592_, new_n5591_, new_n5590_ );
and  ( new_n5593_, new_n5592_, new_n5589_ );
or   ( new_n5594_, new_n5593_, new_n5588_ );
and  ( new_n5595_, new_n5507_, new_n4566_ );
and  ( new_n5596_, new_n5503_, new_n4785_ );
or   ( new_n5597_, new_n5596_, new_n5595_ );
and  ( new_n5598_, new_n5514_, new_n5110_ );
and  ( new_n5599_, new_n5510_, new_n5265_ );
or   ( new_n5600_, new_n5599_, new_n5598_ );
and  ( new_n5601_, new_n5600_, new_n5597_ );
or   ( new_n5602_, new_n5600_, new_n5597_ );
and  ( new_n5603_, new_n5523_, new_n4979_ );
and  ( new_n5604_, new_n5519_, new_n5250_ );
or   ( new_n5605_, new_n5604_, new_n5603_ );
and  ( new_n5606_, new_n5605_, new_n5602_ );
or   ( new_n5607_, new_n5606_, new_n5601_ );
and  ( new_n5608_, new_n5317_, new_n5182_ );
and  ( new_n5609_, new_n5309_, new_n5028_ );
or   ( new_n5610_, new_n5609_, new_n5608_ );
and  ( new_n5611_, new_n5326_, new_n4400_ );
and  ( new_n5612_, new_n5322_, new_n4215_ );
or   ( new_n5613_, new_n5612_, new_n5611_ );
and  ( new_n5614_, new_n5613_, new_n5610_ );
or   ( new_n5615_, new_n5613_, new_n5610_ );
and  ( new_n5616_, new_n5337_, new_n3695_ );
and  ( new_n5617_, new_n5333_, new_n3548_ );
or   ( new_n5618_, new_n5617_, new_n5616_ );
and  ( new_n5619_, new_n5618_, new_n5615_ );
or   ( new_n5620_, new_n5619_, new_n5614_ );
and  ( new_n5621_, new_n5348_, new_n3004_ );
and  ( new_n5622_, new_n5344_, new_n2868_ );
or   ( new_n5623_, new_n5622_, new_n5621_ );
and  ( new_n5624_, new_n5357_, new_n2334_ );
and  ( new_n5625_, new_n5353_, new_n2168_ );
or   ( new_n5626_, new_n5625_, new_n5624_ );
and  ( new_n5627_, new_n5626_, new_n5623_ );
or   ( new_n5628_, new_n5626_, new_n5623_ );
and  ( new_n5629_, new_n5368_, new_n1824_ );
and  ( new_n5630_, new_n5364_, new_n1717_ );
or   ( new_n5631_, new_n5630_, new_n5629_ );
and  ( new_n5632_, new_n5631_, new_n5628_ );
or   ( new_n5633_, new_n5632_, new_n5627_ );
and  ( new_n5634_, new_n5633_, new_n5620_ );
or   ( new_n5635_, new_n5633_, new_n5620_ );
and  ( new_n5636_, new_n5381_, new_n1355_ );
and  ( new_n5637_, new_n5377_, new_n1267_ );
or   ( new_n5638_, new_n5637_, new_n5636_ );
and  ( new_n5639_, new_n5390_, new_n913_ );
and  ( new_n5640_, new_n5386_, new_n938_ );
or   ( new_n5641_, new_n5640_, new_n5639_ );
and  ( new_n5642_, new_n5641_, new_n5638_ );
or   ( new_n5643_, new_n5641_, new_n5638_ );
and  ( new_n5644_, new_n5401_, new_n428_ );
and  ( new_n5645_, new_n5397_, new_n457_ );
or   ( new_n5646_, new_n5645_, new_n5644_ );
and  ( new_n5647_, new_n5646_, new_n5643_ );
or   ( new_n5648_, new_n5647_, new_n5642_ );
and  ( new_n5649_, new_n5648_, new_n5635_ );
or   ( new_n5650_, new_n5649_, new_n5634_ );
and  ( new_n5651_, new_n5414_, new_n505_ );
and  ( new_n5652_, new_n5410_, new_n533_ );
or   ( new_n5653_, new_n5652_, new_n5651_ );
and  ( new_n5654_, new_n5423_, new_n590_ );
and  ( new_n5655_, new_n5419_, new_n619_ );
or   ( new_n5656_, new_n5655_, new_n5654_ );
and  ( new_n5657_, new_n5656_, new_n5653_ );
or   ( new_n5658_, new_n5656_, new_n5653_ );
and  ( new_n5659_, new_n5434_, new_n734_ );
and  ( new_n5660_, new_n5430_, new_n762_ );
or   ( new_n5661_, new_n5660_, new_n5659_ );
and  ( new_n5662_, new_n5661_, new_n5658_ );
or   ( new_n5663_, new_n5662_, new_n5657_ );
and  ( new_n5664_, new_n5445_, new_n785_ );
and  ( new_n5665_, new_n5441_, new_n813_ );
or   ( new_n5666_, new_n5665_, new_n5664_ );
and  ( new_n5667_, new_n5454_, new_n842_ );
and  ( new_n5668_, new_n5450_, new_n866_ );
or   ( new_n5669_, new_n5668_, new_n5667_ );
or   ( new_n5670_, new_n5669_, new_n5666_ );
and  ( new_n5671_, new_n5669_, new_n5666_ );
and  ( new_n5672_, new_n720_, RI2b1c4342e188_92 );
or   ( new_n5673_, new_n5672_, new_n5671_ );
and  ( new_n5674_, new_n5673_, new_n5670_ );
or   ( new_n5675_, new_n5674_, new_n5663_ );
and  ( new_n5676_, new_n5674_, new_n5663_ );
and  ( new_n5677_, new_n5469_, new_n4972_ );
and  ( new_n5678_, new_n5465_, new_n5244_ );
or   ( new_n5679_, new_n5678_, new_n5677_ );
or   ( new_n5680_, new_n5679_, new_n5676_ );
and  ( new_n5681_, new_n5680_, new_n5675_ );
or   ( new_n5682_, new_n5681_, new_n5650_ );
and  ( new_n5683_, new_n5681_, new_n5650_ );
and  ( new_n5684_, new_n5480_, new_n4949_ );
and  ( new_n5685_, new_n5476_, new_n5233_ );
or   ( new_n5686_, new_n5685_, new_n5684_ );
and  ( new_n5687_, new_n5487_, new_n5081_ );
and  ( new_n5688_, new_n5483_, new_n5218_ );
or   ( new_n5689_, new_n5688_, new_n5687_ );
and  ( new_n5690_, new_n5689_, new_n5686_ );
or   ( new_n5691_, new_n5689_, new_n5686_ );
and  ( new_n5692_, new_n5496_, new_n5010_ );
and  ( new_n5693_, new_n5492_, new_n5203_ );
or   ( new_n5694_, new_n5693_, new_n5692_ );
and  ( new_n5695_, new_n5694_, new_n5691_ );
or   ( new_n5696_, new_n5695_, new_n5690_ );
or   ( new_n5697_, new_n5696_, new_n5683_ );
and  ( new_n5698_, new_n5697_, new_n5682_ );
or   ( new_n5699_, new_n5698_, new_n5607_ );
and  ( new_n5700_, new_n5698_, new_n5607_ );
and  ( new_n5701_, new_n5534_, new_n4688_ );
and  ( new_n5702_, new_n5530_, new_n4840_ );
or   ( new_n5703_, new_n5702_, new_n5701_ );
or   ( new_n5704_, new_n5703_, new_n5700_ );
and  ( new_n5705_, new_n5704_, new_n5699_ );
or   ( new_n5706_, new_n5705_, new_n5594_ );
and  ( new_n5707_, new_n5705_, new_n5594_ );
and  ( new_n5708_, new_n5570_, new_n4711_ );
and  ( new_n5709_, new_n5566_, new_n4855_ );
or   ( new_n5710_, new_n5709_, new_n5708_ );
or   ( new_n5711_, new_n5710_, new_n5707_ );
and  ( new_n5712_, new_n5711_, new_n5706_ );
and  ( new_n5713_, new_n5712_, new_n5581_ );
or   ( new_n5714_, new_n5713_, new_n5578_ );
or   ( new_n5715_, new_n5271_, new_n5115_ );
and  ( new_n5716_, new_n5715_, new_n5123_ );
and  ( new_n5717_, new_n5269_, new_n4920_ );
and  ( new_n5718_, new_n5171_, new_n5114_ );
or   ( new_n5719_, new_n5718_, new_n5717_ );
and  ( new_n5720_, new_n5719_, new_n5274_ );
or   ( new_n5721_, new_n5720_, new_n5716_ );
or   ( new_n5722_, new_n5588_, new_n5553_ );
and  ( new_n5723_, new_n5722_, new_n5561_ );
and  ( new_n5724_, new_n5584_, new_n5552_ );
and  ( new_n5725_, new_n5587_, new_n5545_ );
or   ( new_n5726_, new_n5725_, new_n5724_ );
and  ( new_n5727_, new_n5726_, new_n5592_ );
or   ( new_n5728_, new_n5727_, new_n5723_ );
or   ( new_n5729_, new_n5186_, new_n5038_ );
and  ( new_n5730_, new_n5729_, new_n5048_ );
and  ( new_n5731_, new_n5182_, new_n5037_ );
and  ( new_n5732_, new_n5185_, new_n5028_ );
or   ( new_n5733_, new_n5732_, new_n5731_ );
and  ( new_n5734_, new_n5733_, new_n5190_ );
or   ( new_n5735_, new_n5734_, new_n5730_ );
or   ( new_n5736_, new_n5690_, new_n5490_ );
and  ( new_n5737_, new_n5736_, new_n5498_ );
and  ( new_n5738_, new_n5686_, new_n5489_ );
and  ( new_n5739_, new_n5689_, new_n5482_ );
or   ( new_n5740_, new_n5739_, new_n5738_ );
and  ( new_n5741_, new_n5740_, new_n5694_ );
or   ( new_n5742_, new_n5741_, new_n5737_ );
and  ( new_n5743_, new_n5742_, new_n5735_ );
or   ( new_n5744_, new_n5742_, new_n5735_ );
or   ( new_n5745_, new_n5676_, new_n5463_ );
and  ( new_n5746_, new_n5745_, new_n5471_ );
and  ( new_n5747_, new_n5663_, new_n5462_ );
and  ( new_n5748_, new_n5674_, new_n5438_ );
or   ( new_n5749_, new_n5748_, new_n5747_ );
and  ( new_n5750_, new_n5749_, new_n5679_ );
or   ( new_n5751_, new_n5750_, new_n5746_ );
and  ( new_n5752_, new_n5751_, new_n5744_ );
or   ( new_n5753_, new_n5752_, new_n5743_ );
or   ( new_n5754_, new_n753_, new_n3902_ );
or   ( new_n5755_, new_n757_, new_n3924_ );
and  ( new_n5756_, new_n5755_, new_n5754_ );
and  ( new_n5757_, new_n5756_, new_n734_ );
and  ( new_n5758_, new_n766_, RI2b1c4342dfa8_88 );
and  ( new_n5759_, new_n751_, RI2b1c4342df30_87 );
or   ( new_n5760_, new_n5759_, new_n5758_ );
and  ( new_n5761_, new_n5760_, new_n762_ );
or   ( new_n5762_, new_n5761_, new_n5757_ );
or   ( new_n5763_, new_n804_, new_n4635_ );
or   ( new_n5764_, new_n808_, new_n132_ );
and  ( new_n5765_, new_n5764_, new_n5763_ );
and  ( new_n5766_, new_n5765_, new_n785_ );
and  ( new_n5767_, new_n817_, RI2b1c4342e098_90 );
and  ( new_n5768_, new_n802_, RI2b1c4342e020_89 );
or   ( new_n5769_, new_n5768_, new_n5767_ );
and  ( new_n5770_, new_n5769_, new_n813_ );
or   ( new_n5771_, new_n5770_, new_n5766_ );
and  ( new_n5772_, new_n5771_, new_n5762_ );
or   ( new_n5773_, new_n5771_, new_n5762_ );
or   ( new_n5774_, new_n857_, new_n5459_ );
or   ( new_n5775_, new_n861_, new_n117_ );
and  ( new_n5776_, new_n5775_, new_n5774_ );
and  ( new_n5777_, new_n5776_, new_n842_ );
and  ( new_n5778_, new_n870_, RI2b1c4342e188_92 );
and  ( new_n5779_, new_n855_, RI2b1c4342e110_91 );
or   ( new_n5780_, new_n5779_, new_n5778_ );
and  ( new_n5781_, new_n5780_, new_n866_ );
or   ( new_n5782_, new_n5781_, new_n5777_ );
and  ( new_n5783_, new_n5782_, new_n5773_ );
or   ( new_n5784_, new_n5783_, new_n5772_ );
or   ( new_n5785_, new_n453_, new_n2119_ );
or   ( new_n5786_, new_n459_, new_n126_ );
and  ( new_n5787_, new_n5786_, new_n5785_ );
and  ( new_n5788_, new_n5787_, new_n428_ );
and  ( new_n5789_, new_n463_, RI2b1c4342dcd8_82 );
and  ( new_n5790_, new_n451_, RI2b1c4342dc60_81 );
or   ( new_n5791_, new_n5790_, new_n5789_ );
and  ( new_n5792_, new_n5791_, new_n457_ );
or   ( new_n5793_, new_n5792_, new_n5788_ );
or   ( new_n5794_, new_n524_, new_n2541_ );
or   ( new_n5795_, new_n528_, new_n121_ );
and  ( new_n5796_, new_n5795_, new_n5794_ );
and  ( new_n5797_, new_n5796_, new_n505_ );
and  ( new_n5798_, new_n537_, RI2b1c4342ddc8_84 );
and  ( new_n5799_, new_n522_, RI2b1c4342dd50_83 );
or   ( new_n5800_, new_n5799_, new_n5798_ );
and  ( new_n5801_, new_n5800_, new_n533_ );
or   ( new_n5802_, new_n5801_, new_n5797_ );
and  ( new_n5803_, new_n5802_, new_n5793_ );
or   ( new_n5804_, new_n5802_, new_n5793_ );
or   ( new_n5805_, new_n610_, new_n3239_ );
or   ( new_n5806_, new_n614_, new_n2806_ );
and  ( new_n5807_, new_n5806_, new_n5805_ );
and  ( new_n5808_, new_n5807_, new_n590_ );
and  ( new_n5809_, new_n623_, RI2b1c4342deb8_86 );
and  ( new_n5810_, new_n608_, RI2b1c4342de40_85 );
or   ( new_n5811_, new_n5810_, new_n5809_ );
and  ( new_n5812_, new_n5811_, new_n619_ );
or   ( new_n5813_, new_n5812_, new_n5808_ );
and  ( new_n5814_, new_n5813_, new_n5804_ );
or   ( new_n5815_, new_n5814_, new_n5803_ );
and  ( new_n5816_, new_n5815_, new_n5784_ );
or   ( new_n5817_, new_n3802_, new_n755_ );
or   ( new_n5818_, new_n3806_, new_n591_ );
and  ( new_n5819_, new_n5818_, new_n5817_ );
and  ( new_n5820_, new_n5819_, new_n3695_ );
and  ( new_n5821_, new_n3810_, RI2b1c4342d738_70 );
and  ( new_n5822_, new_n3800_, RI2b1c4342d6c0_69 );
or   ( new_n5823_, new_n5822_, new_n5821_ );
and  ( new_n5824_, new_n5823_, new_n3548_ );
or   ( new_n5825_, new_n5824_, new_n5820_ );
or   ( new_n5826_, new_n3112_, new_n806_ );
or   ( new_n5827_, new_n3116_, new_n110_ );
and  ( new_n5828_, new_n5827_, new_n5826_ );
and  ( new_n5829_, new_n5828_, new_n3004_ );
and  ( new_n5830_, new_n3120_, RI2b1c4342d828_72 );
and  ( new_n5831_, new_n3110_, RI2b1c4342d7b0_71 );
or   ( new_n5832_, new_n5831_, new_n5830_ );
and  ( new_n5833_, new_n5832_, new_n2868_ );
or   ( new_n5834_, new_n5833_, new_n5829_ );
and  ( new_n5835_, new_n5834_, new_n5825_ );
or   ( new_n5836_, new_n5834_, new_n5825_ );
or   ( new_n5837_, new_n2450_, new_n859_ );
or   ( new_n5838_, new_n2454_, new_n105_ );
and  ( new_n5839_, new_n5838_, new_n5837_ );
and  ( new_n5840_, new_n5839_, new_n2334_ );
and  ( new_n5841_, new_n2458_, RI2b1c4342d918_74 );
and  ( new_n5842_, new_n2448_, RI2b1c4342d8a0_73 );
or   ( new_n5843_, new_n5842_, new_n5841_ );
and  ( new_n5844_, new_n5843_, new_n2168_ );
or   ( new_n5845_, new_n5844_, new_n5840_ );
and  ( new_n5846_, new_n5845_, new_n5836_ );
or   ( new_n5847_, new_n5846_, new_n5835_ );
xor  ( new_n5848_, new_n335_, new_n208_ );
not  ( new_n5849_, RI2b1c4342d468_64 );
not  ( new_n5850_, RI2b1c4342c568_32 );
and  ( new_n5851_, new_n138_, new_n5850_ );
or   ( new_n5852_, new_n5851_, new_n5849_ );
and  ( new_n5853_, new_n5852_, new_n5848_ );
or   ( new_n5854_, new_n5853_, new_n209_ );
and  ( new_n5855_, new_n138_, RI2b1c4342c568_32 );
and  ( new_n5856_, new_n5855_, RI2b1c4342d468_64 );
and  ( new_n5857_, new_n5856_, new_n208_ );
or   ( new_n5858_, new_n5857_, new_n5854_ );
xor  ( new_n5859_, new_n332_, new_n204_ );
and  ( new_n5860_, new_n5859_, new_n340_ );
xor  ( new_n5861_, RI2b1c4342c478_30, RI2b1c4342d378_62 );
and  ( new_n5862_, new_n5861_, new_n216_ );
and  ( new_n5863_, new_n5862_, new_n138_ );
or   ( new_n5864_, new_n5863_, new_n205_ );
or   ( new_n5865_, new_n5864_, new_n5860_ );
or   ( new_n5866_, new_n5865_, new_n5858_ );
and  ( new_n5867_, new_n5866_, new_n5176_ );
or   ( new_n5868_, new_n5308_, new_n526_ );
or   ( new_n5869_, new_n5312_, new_n99_ );
and  ( new_n5870_, new_n5869_, new_n5868_ );
and  ( new_n5871_, new_n5870_, new_n5182_ );
and  ( new_n5872_, new_n5316_, RI2b1c4342d558_66 );
and  ( new_n5873_, new_n5306_, RI2b1c4342d4e0_65 );
or   ( new_n5874_, new_n5873_, new_n5872_ );
and  ( new_n5875_, new_n5874_, new_n5028_ );
or   ( new_n5876_, new_n5875_, new_n5871_ );
and  ( new_n5877_, new_n5876_, new_n5867_ );
or   ( new_n5878_, new_n5876_, new_n5867_ );
or   ( new_n5879_, new_n4535_, new_n612_ );
or   ( new_n5880_, new_n4539_, new_n112_ );
and  ( new_n5881_, new_n5880_, new_n5879_ );
and  ( new_n5882_, new_n5881_, new_n4400_ );
and  ( new_n5883_, new_n4543_, RI2b1c4342d648_68 );
and  ( new_n5884_, new_n4533_, RI2b1c4342d5d0_67 );
or   ( new_n5885_, new_n5884_, new_n5883_ );
and  ( new_n5886_, new_n5885_, new_n4215_ );
or   ( new_n5887_, new_n5886_, new_n5882_ );
and  ( new_n5888_, new_n5887_, new_n5878_ );
or   ( new_n5889_, new_n5888_, new_n5877_ );
and  ( new_n5890_, new_n5889_, new_n5847_ );
or   ( new_n5891_, new_n5889_, new_n5847_ );
or   ( new_n5892_, new_n1910_, new_n886_ );
or   ( new_n5893_, new_n1914_, new_n843_ );
and  ( new_n5894_, new_n5893_, new_n5892_ );
and  ( new_n5895_, new_n5894_, new_n1824_ );
and  ( new_n5896_, new_n1918_, RI2b1c4342da08_76 );
and  ( new_n5897_, new_n1908_, RI2b1c4342d990_75 );
or   ( new_n5898_, new_n5897_, new_n5896_ );
and  ( new_n5899_, new_n5898_, new_n1717_ );
or   ( new_n5900_, new_n5899_, new_n5895_ );
or   ( new_n5901_, new_n1425_, new_n1002_ );
or   ( new_n5902_, new_n1429_, new_n1004_ );
and  ( new_n5903_, new_n5902_, new_n5901_ );
and  ( new_n5904_, new_n5903_, new_n1355_ );
and  ( new_n5905_, new_n1433_, RI2b1c4342daf8_78 );
and  ( new_n5906_, new_n1423_, RI2b1c4342da80_77 );
or   ( new_n5907_, new_n5906_, new_n5905_ );
and  ( new_n5908_, new_n5907_, new_n1267_ );
or   ( new_n5909_, new_n5908_, new_n5904_ );
and  ( new_n5910_, new_n5909_, new_n5900_ );
or   ( new_n5911_, new_n5909_, new_n5900_ );
or   ( new_n5912_, new_n934_, new_n1511_ );
or   ( new_n5913_, new_n940_, new_n1310_ );
and  ( new_n5914_, new_n5913_, new_n5912_ );
and  ( new_n5915_, new_n5914_, new_n913_ );
and  ( new_n5916_, new_n944_, RI2b1c4342dbe8_80 );
and  ( new_n5917_, new_n932_, RI2b1c4342db70_79 );
or   ( new_n5918_, new_n5917_, new_n5916_ );
and  ( new_n5919_, new_n5918_, new_n938_ );
or   ( new_n5920_, new_n5919_, new_n5915_ );
and  ( new_n5921_, new_n5920_, new_n5911_ );
or   ( new_n5922_, new_n5921_, new_n5910_ );
and  ( new_n5923_, new_n5922_, new_n5891_ );
or   ( new_n5924_, new_n5923_, new_n5890_ );
and  ( new_n5925_, new_n5924_, new_n5816_ );
or   ( new_n5926_, new_n5924_, new_n5816_ );
or   ( new_n5927_, new_n5671_, new_n5457_ );
and  ( new_n5928_, new_n5927_, new_n5460_ );
and  ( new_n5929_, new_n5666_, new_n5456_ );
and  ( new_n5930_, new_n5669_, new_n5447_ );
or   ( new_n5931_, new_n5930_, new_n5929_ );
and  ( new_n5932_, new_n5931_, new_n5672_ );
or   ( new_n5933_, new_n5932_, new_n5928_ );
or   ( new_n5934_, new_n5657_, new_n5426_ );
and  ( new_n5935_, new_n5934_, new_n5436_ );
and  ( new_n5936_, new_n5653_, new_n5425_ );
and  ( new_n5937_, new_n5656_, new_n5416_ );
or   ( new_n5938_, new_n5937_, new_n5936_ );
and  ( new_n5939_, new_n5938_, new_n5661_ );
or   ( new_n5940_, new_n5939_, new_n5935_ );
and  ( new_n5941_, new_n5940_, new_n5933_ );
or   ( new_n5942_, new_n5940_, new_n5933_ );
or   ( new_n5943_, new_n5642_, new_n5393_ );
and  ( new_n5944_, new_n5943_, new_n5403_ );
and  ( new_n5945_, new_n5638_, new_n5392_ );
and  ( new_n5946_, new_n5641_, new_n5383_ );
or   ( new_n5947_, new_n5946_, new_n5945_ );
and  ( new_n5948_, new_n5947_, new_n5646_ );
or   ( new_n5949_, new_n5948_, new_n5944_ );
and  ( new_n5950_, new_n5949_, new_n5942_ );
or   ( new_n5951_, new_n5950_, new_n5941_ );
and  ( new_n5952_, new_n5951_, new_n5926_ );
or   ( new_n5953_, new_n5952_, new_n5925_ );
and  ( new_n5954_, new_n5953_, new_n5753_ );
or   ( new_n5955_, new_n5953_, new_n5753_ );
or   ( new_n5956_, new_n5206_, new_n5051_ );
and  ( new_n5957_, new_n5956_, new_n5083_ );
and  ( new_n5958_, new_n5192_, new_n5012_ );
and  ( new_n5959_, new_n5205_, new_n5050_ );
or   ( new_n5960_, new_n5959_, new_n5958_ );
and  ( new_n5961_, new_n5960_, new_n5220_ );
or   ( new_n5962_, new_n5961_, new_n5957_ );
and  ( new_n5963_, new_n5962_, new_n5955_ );
or   ( new_n5964_, new_n5963_, new_n5954_ );
and  ( new_n5965_, new_n5964_, new_n5728_ );
or   ( new_n5966_, new_n5964_, new_n5728_ );
or   ( new_n5967_, new_n5700_, new_n5528_ );
and  ( new_n5968_, new_n5967_, new_n5536_ );
and  ( new_n5969_, new_n5698_, new_n5527_ );
and  ( new_n5970_, new_n5607_, new_n5502_ );
or   ( new_n5971_, new_n5970_, new_n5969_ );
and  ( new_n5972_, new_n5971_, new_n5703_ );
or   ( new_n5973_, new_n5972_, new_n5968_ );
and  ( new_n5974_, new_n5973_, new_n5966_ );
or   ( new_n5975_, new_n5974_, new_n5965_ );
and  ( new_n5976_, new_n5975_, new_n5721_ );
or   ( new_n5977_, new_n5975_, new_n5721_ );
or   ( new_n5978_, new_n5707_, new_n5564_ );
and  ( new_n5979_, new_n5978_, new_n5572_ );
and  ( new_n5980_, new_n5705_, new_n5563_ );
and  ( new_n5981_, new_n5594_, new_n5538_ );
or   ( new_n5982_, new_n5981_, new_n5980_ );
and  ( new_n5983_, new_n5982_, new_n5710_ );
or   ( new_n5984_, new_n5983_, new_n5979_ );
and  ( new_n5985_, new_n5984_, new_n5977_ );
or   ( new_n5986_, new_n5985_, new_n5976_ );
or   ( new_n5987_, new_n5986_, new_n5714_ );
and  ( new_n5988_, new_n5987_, new_n5577_ );
or   ( new_n5989_, new_n5988_, new_n5576_ );
or   ( new_n5990_, new_n5989_, new_n5152_ );
and  ( new_n5991_, new_n5990_, new_n5150_ );
and  ( new_n5992_, new_n5986_, new_n5714_ );
or   ( new_n5993_, new_n5992_, new_n5576_ );
or   ( new_n5994_, new_n5993_, new_n5152_ );
and  ( new_n5995_, new_n5719_, new_n5123_ );
and  ( new_n5996_, new_n5715_, new_n5274_ );
or   ( new_n5997_, new_n5996_, new_n5995_ );
and  ( new_n5998_, new_n5726_, new_n5561_ );
and  ( new_n5999_, new_n5722_, new_n5592_ );
or   ( new_n6000_, new_n5999_, new_n5998_ );
and  ( new_n6001_, new_n5791_, new_n428_ );
and  ( new_n6002_, new_n5787_, new_n457_ );
or   ( new_n6003_, new_n6002_, new_n6001_ );
and  ( new_n6004_, new_n5800_, new_n505_ );
and  ( new_n6005_, new_n5796_, new_n533_ );
or   ( new_n6006_, new_n6005_, new_n6004_ );
and  ( new_n6007_, new_n6006_, new_n6003_ );
or   ( new_n6008_, new_n6006_, new_n6003_ );
and  ( new_n6009_, new_n5811_, new_n590_ );
and  ( new_n6010_, new_n5807_, new_n619_ );
or   ( new_n6011_, new_n6010_, new_n6009_ );
and  ( new_n6012_, new_n6011_, new_n6008_ );
or   ( new_n6013_, new_n6012_, new_n6007_ );
and  ( new_n6014_, new_n5760_, new_n734_ );
and  ( new_n6015_, new_n5756_, new_n762_ );
or   ( new_n6016_, new_n6015_, new_n6014_ );
and  ( new_n6017_, new_n5769_, new_n785_ );
and  ( new_n6018_, new_n5765_, new_n813_ );
or   ( new_n6019_, new_n6018_, new_n6017_ );
and  ( new_n6020_, new_n6019_, new_n6016_ );
or   ( new_n6021_, new_n6019_, new_n6016_ );
and  ( new_n6022_, new_n5780_, new_n842_ );
and  ( new_n6023_, new_n5776_, new_n866_ );
or   ( new_n6024_, new_n6023_, new_n6022_ );
and  ( new_n6025_, new_n6024_, new_n6021_ );
or   ( new_n6026_, new_n6025_, new_n6020_ );
or   ( new_n6027_, new_n6026_, new_n6013_ );
not  ( new_n6028_, new_n216_ );
nor  ( new_n6029_, new_n5861_, new_n6028_ );
and  ( new_n6030_, new_n5861_, new_n340_ );
or   ( new_n6031_, new_n6030_, new_n6029_ );
and  ( new_n6032_, new_n6031_, new_n332_ );
xor  ( new_n6033_, RI2b1c4342c4f0_31, RI2b1c4342d3f0_63 );
nor  ( new_n6034_, new_n6033_, new_n214_ );
and  ( new_n6035_, new_n214_, new_n208_ );
or   ( new_n6036_, new_n6035_, new_n6034_ );
and  ( new_n6037_, new_n6036_, new_n335_ );
and  ( new_n6038_, new_n6037_, new_n6032_ );
or   ( new_n6039_, new_n6038_, new_n5019_ );
and  ( new_n6040_, new_n5874_, new_n5182_ );
and  ( new_n6041_, new_n5870_, new_n5028_ );
or   ( new_n6042_, new_n6041_, new_n6040_ );
and  ( new_n6043_, new_n6042_, new_n6039_ );
or   ( new_n6044_, new_n6042_, new_n6039_ );
and  ( new_n6045_, new_n5885_, new_n4400_ );
and  ( new_n6046_, new_n5881_, new_n4215_ );
or   ( new_n6047_, new_n6046_, new_n6045_ );
and  ( new_n6048_, new_n6047_, new_n6044_ );
or   ( new_n6049_, new_n6048_, new_n6043_ );
and  ( new_n6050_, new_n5823_, new_n3695_ );
and  ( new_n6051_, new_n5819_, new_n3548_ );
or   ( new_n6052_, new_n6051_, new_n6050_ );
and  ( new_n6053_, new_n5832_, new_n3004_ );
and  ( new_n6054_, new_n5828_, new_n2868_ );
or   ( new_n6055_, new_n6054_, new_n6053_ );
and  ( new_n6056_, new_n6055_, new_n6052_ );
or   ( new_n6057_, new_n6055_, new_n6052_ );
and  ( new_n6058_, new_n5843_, new_n2334_ );
and  ( new_n6059_, new_n5839_, new_n2168_ );
or   ( new_n6060_, new_n6059_, new_n6058_ );
and  ( new_n6061_, new_n6060_, new_n6057_ );
or   ( new_n6062_, new_n6061_, new_n6056_ );
and  ( new_n6063_, new_n6062_, new_n6049_ );
or   ( new_n6064_, new_n6062_, new_n6049_ );
and  ( new_n6065_, new_n5898_, new_n1824_ );
and  ( new_n6066_, new_n5894_, new_n1717_ );
or   ( new_n6067_, new_n6066_, new_n6065_ );
and  ( new_n6068_, new_n5907_, new_n1355_ );
and  ( new_n6069_, new_n5903_, new_n1267_ );
or   ( new_n6070_, new_n6069_, new_n6068_ );
and  ( new_n6071_, new_n6070_, new_n6067_ );
or   ( new_n6072_, new_n6070_, new_n6067_ );
and  ( new_n6073_, new_n5918_, new_n913_ );
and  ( new_n6074_, new_n5914_, new_n938_ );
or   ( new_n6075_, new_n6074_, new_n6073_ );
and  ( new_n6076_, new_n6075_, new_n6072_ );
or   ( new_n6077_, new_n6076_, new_n6071_ );
and  ( new_n6078_, new_n6077_, new_n6064_ );
or   ( new_n6079_, new_n6078_, new_n6063_ );
and  ( new_n6080_, new_n6079_, new_n6027_ );
or   ( new_n6081_, new_n6079_, new_n6027_ );
and  ( new_n6082_, new_n5931_, new_n5460_ );
and  ( new_n6083_, new_n5927_, new_n5672_ );
or   ( new_n6084_, new_n6083_, new_n6082_ );
and  ( new_n6085_, new_n5938_, new_n5436_ );
and  ( new_n6086_, new_n5934_, new_n5661_ );
or   ( new_n6087_, new_n6086_, new_n6085_ );
and  ( new_n6088_, new_n6087_, new_n6084_ );
or   ( new_n6089_, new_n6087_, new_n6084_ );
and  ( new_n6090_, new_n5947_, new_n5403_ );
and  ( new_n6091_, new_n5943_, new_n5646_ );
or   ( new_n6092_, new_n6091_, new_n6090_ );
and  ( new_n6093_, new_n6092_, new_n6089_ );
or   ( new_n6094_, new_n6093_, new_n6088_ );
and  ( new_n6095_, new_n6094_, new_n6081_ );
or   ( new_n6096_, new_n6095_, new_n6080_ );
and  ( new_n6097_, new_n5733_, new_n5048_ );
and  ( new_n6098_, new_n5729_, new_n5190_ );
or   ( new_n6099_, new_n6098_, new_n6097_ );
and  ( new_n6100_, new_n5740_, new_n5498_ );
and  ( new_n6101_, new_n5736_, new_n5694_ );
or   ( new_n6102_, new_n6101_, new_n6100_ );
and  ( new_n6103_, new_n6102_, new_n6099_ );
or   ( new_n6104_, new_n6102_, new_n6099_ );
and  ( new_n6105_, new_n5749_, new_n5471_ );
and  ( new_n6106_, new_n5745_, new_n5679_ );
or   ( new_n6107_, new_n6106_, new_n6105_ );
and  ( new_n6108_, new_n6107_, new_n6104_ );
or   ( new_n6109_, new_n6108_, new_n6103_ );
and  ( new_n6110_, new_n6109_, new_n6096_ );
or   ( new_n6111_, new_n6109_, new_n6096_ );
and  ( new_n6112_, new_n5960_, new_n5083_ );
and  ( new_n6113_, new_n5956_, new_n5220_ );
or   ( new_n6114_, new_n6113_, new_n6112_ );
and  ( new_n6115_, new_n6114_, new_n6111_ );
or   ( new_n6116_, new_n6115_, new_n6110_ );
and  ( new_n6117_, new_n6116_, new_n6000_ );
or   ( new_n6118_, new_n6116_, new_n6000_ );
and  ( new_n6119_, new_n5971_, new_n5536_ );
and  ( new_n6120_, new_n5967_, new_n5703_ );
or   ( new_n6121_, new_n6120_, new_n6119_ );
and  ( new_n6122_, new_n6121_, new_n6118_ );
or   ( new_n6123_, new_n6122_, new_n6117_ );
and  ( new_n6124_, new_n6123_, new_n5997_ );
or   ( new_n6125_, new_n6124_, new_n5976_ );
and  ( new_n6126_, new_n6125_, new_n5984_ );
and  ( new_n6127_, new_n6123_, new_n5721_ );
and  ( new_n6128_, new_n5997_, new_n5975_ );
or   ( new_n6129_, new_n6128_, new_n6127_ );
and  ( new_n6130_, new_n5982_, new_n5572_ );
and  ( new_n6131_, new_n5978_, new_n5710_ );
or   ( new_n6132_, new_n6131_, new_n6130_ );
and  ( new_n6133_, new_n6132_, new_n6129_ );
or   ( new_n6134_, new_n6133_, new_n6126_ );
or   ( new_n6135_, new_n5683_, new_n5474_ );
and  ( new_n6136_, new_n6135_, new_n5500_ );
and  ( new_n6137_, new_n5650_, new_n5473_ );
and  ( new_n6138_, new_n5681_, new_n5407_ );
or   ( new_n6139_, new_n6138_, new_n6137_ );
and  ( new_n6140_, new_n6139_, new_n5696_ );
or   ( new_n6141_, new_n6140_, new_n6136_ );
or   ( new_n6142_, new_n6110_, new_n5954_ );
and  ( new_n6143_, new_n6142_, new_n5962_ );
and  ( new_n6144_, new_n6096_, new_n5753_ );
and  ( new_n6145_, new_n6109_, new_n5953_ );
or   ( new_n6146_, new_n6145_, new_n6144_ );
and  ( new_n6147_, new_n6146_, new_n6114_ );
or   ( new_n6148_, new_n6147_, new_n6143_ );
or   ( new_n6149_, new_n6148_, new_n6141_ );
and  ( new_n6150_, new_n6032_, new_n5176_ );
and  ( new_n6151_, new_n5865_, new_n5019_ );
and  ( new_n6152_, new_n6032_, new_n5858_ );
and  ( new_n6153_, new_n6037_, new_n5865_ );
or   ( new_n6154_, new_n6153_, new_n6152_ );
or   ( new_n6155_, new_n6154_, new_n6151_ );
or   ( new_n6156_, new_n6155_, new_n6150_ );
or   ( new_n6157_, new_n6156_, new_n99_ );
and  ( new_n6158_, new_n6157_, new_n6039_ );
and  ( new_n6159_, new_n5865_, new_n5858_ );
or   ( new_n6160_, new_n6159_, new_n6038_ );
and  ( new_n6161_, new_n5865_, new_n5176_ );
and  ( new_n6162_, new_n6032_, new_n5019_ );
or   ( new_n6163_, new_n6162_, new_n6161_ );
and  ( new_n6164_, new_n6163_, new_n6160_ );
and  ( new_n6165_, new_n6164_, RI2b1c4342d4e0_65 );
and  ( new_n6166_, new_n6165_, new_n5867_ );
or   ( new_n6167_, new_n6166_, new_n6158_ );
or   ( new_n6168_, new_n5308_, new_n112_ );
or   ( new_n6169_, new_n5312_, new_n526_ );
and  ( new_n6170_, new_n6169_, new_n6168_ );
and  ( new_n6171_, new_n6170_, new_n5182_ );
and  ( new_n6172_, new_n5316_, RI2b1c4342d5d0_67 );
and  ( new_n6173_, new_n5306_, RI2b1c4342d558_66 );
or   ( new_n6174_, new_n6173_, new_n6172_ );
and  ( new_n6175_, new_n6174_, new_n5028_ );
or   ( new_n6176_, new_n6175_, new_n6171_ );
and  ( new_n6177_, new_n6176_, new_n6167_ );
or   ( new_n6178_, new_n6176_, new_n6167_ );
or   ( new_n6179_, new_n4535_, new_n591_ );
or   ( new_n6180_, new_n4539_, new_n612_ );
and  ( new_n6181_, new_n6180_, new_n6179_ );
and  ( new_n6182_, new_n6181_, new_n4400_ );
and  ( new_n6183_, new_n4543_, RI2b1c4342d6c0_69 );
and  ( new_n6184_, new_n4533_, RI2b1c4342d648_68 );
or   ( new_n6185_, new_n6184_, new_n6183_ );
and  ( new_n6186_, new_n6185_, new_n4215_ );
or   ( new_n6187_, new_n6186_, new_n6182_ );
and  ( new_n6188_, new_n6187_, new_n6178_ );
or   ( new_n6189_, new_n6188_, new_n6177_ );
or   ( new_n6190_, new_n3802_, new_n110_ );
or   ( new_n6191_, new_n3806_, new_n755_ );
and  ( new_n6192_, new_n6191_, new_n6190_ );
and  ( new_n6193_, new_n6192_, new_n3695_ );
and  ( new_n6194_, new_n3810_, RI2b1c4342d7b0_71 );
and  ( new_n6195_, new_n3800_, RI2b1c4342d738_70 );
or   ( new_n6196_, new_n6195_, new_n6194_ );
and  ( new_n6197_, new_n6196_, new_n3548_ );
or   ( new_n6198_, new_n6197_, new_n6193_ );
or   ( new_n6199_, new_n3112_, new_n105_ );
or   ( new_n6200_, new_n3116_, new_n806_ );
and  ( new_n6201_, new_n6200_, new_n6199_ );
and  ( new_n6202_, new_n6201_, new_n3004_ );
and  ( new_n6203_, new_n3120_, RI2b1c4342d8a0_73 );
and  ( new_n6204_, new_n3110_, RI2b1c4342d828_72 );
or   ( new_n6205_, new_n6204_, new_n6203_ );
and  ( new_n6206_, new_n6205_, new_n2868_ );
or   ( new_n6207_, new_n6206_, new_n6202_ );
and  ( new_n6208_, new_n6207_, new_n6198_ );
or   ( new_n6209_, new_n6207_, new_n6198_ );
or   ( new_n6210_, new_n2450_, new_n843_ );
or   ( new_n6211_, new_n2454_, new_n859_ );
and  ( new_n6212_, new_n6211_, new_n6210_ );
and  ( new_n6213_, new_n6212_, new_n2334_ );
and  ( new_n6214_, new_n2458_, RI2b1c4342d990_75 );
and  ( new_n6215_, new_n2448_, RI2b1c4342d918_74 );
or   ( new_n6216_, new_n6215_, new_n6214_ );
and  ( new_n6217_, new_n6216_, new_n2168_ );
or   ( new_n6218_, new_n6217_, new_n6213_ );
and  ( new_n6219_, new_n6218_, new_n6209_ );
or   ( new_n6220_, new_n6219_, new_n6208_ );
and  ( new_n6221_, new_n6220_, new_n6189_ );
or   ( new_n6222_, new_n6220_, new_n6189_ );
or   ( new_n6223_, new_n1910_, new_n1004_ );
or   ( new_n6224_, new_n1914_, new_n886_ );
and  ( new_n6225_, new_n6224_, new_n6223_ );
and  ( new_n6226_, new_n6225_, new_n1824_ );
and  ( new_n6227_, new_n1918_, RI2b1c4342da80_77 );
and  ( new_n6228_, new_n1908_, RI2b1c4342da08_76 );
or   ( new_n6229_, new_n6228_, new_n6227_ );
and  ( new_n6230_, new_n6229_, new_n1717_ );
or   ( new_n6231_, new_n6230_, new_n6226_ );
or   ( new_n6232_, new_n1425_, new_n1310_ );
or   ( new_n6233_, new_n1429_, new_n1002_ );
and  ( new_n6234_, new_n6233_, new_n6232_ );
and  ( new_n6235_, new_n6234_, new_n1355_ );
and  ( new_n6236_, new_n1433_, RI2b1c4342db70_79 );
and  ( new_n6237_, new_n1423_, RI2b1c4342daf8_78 );
or   ( new_n6238_, new_n6237_, new_n6236_ );
and  ( new_n6239_, new_n6238_, new_n1267_ );
or   ( new_n6240_, new_n6239_, new_n6235_ );
and  ( new_n6241_, new_n6240_, new_n6231_ );
or   ( new_n6242_, new_n6240_, new_n6231_ );
or   ( new_n6243_, new_n934_, new_n126_ );
or   ( new_n6244_, new_n940_, new_n1511_ );
and  ( new_n6245_, new_n6244_, new_n6243_ );
and  ( new_n6246_, new_n6245_, new_n913_ );
and  ( new_n6247_, new_n944_, RI2b1c4342dc60_81 );
and  ( new_n6248_, new_n932_, RI2b1c4342dbe8_80 );
or   ( new_n6249_, new_n6248_, new_n6247_ );
and  ( new_n6250_, new_n6249_, new_n938_ );
or   ( new_n6251_, new_n6250_, new_n6246_ );
and  ( new_n6252_, new_n6251_, new_n6242_ );
or   ( new_n6253_, new_n6252_, new_n6241_ );
and  ( new_n6254_, new_n6253_, new_n6222_ );
or   ( new_n6255_, new_n6254_, new_n6221_ );
or   ( new_n6256_, new_n453_, new_n121_ );
or   ( new_n6257_, new_n459_, new_n2119_ );
and  ( new_n6258_, new_n6257_, new_n6256_ );
and  ( new_n6259_, new_n6258_, new_n428_ );
and  ( new_n6260_, new_n463_, RI2b1c4342dd50_83 );
and  ( new_n6261_, new_n451_, RI2b1c4342dcd8_82 );
or   ( new_n6262_, new_n6261_, new_n6260_ );
and  ( new_n6263_, new_n6262_, new_n457_ );
or   ( new_n6264_, new_n6263_, new_n6259_ );
or   ( new_n6265_, new_n524_, new_n2806_ );
or   ( new_n6266_, new_n528_, new_n2541_ );
and  ( new_n6267_, new_n6266_, new_n6265_ );
and  ( new_n6268_, new_n6267_, new_n505_ );
and  ( new_n6269_, new_n537_, RI2b1c4342de40_85 );
and  ( new_n6270_, new_n522_, RI2b1c4342ddc8_84 );
or   ( new_n6271_, new_n6270_, new_n6269_ );
and  ( new_n6272_, new_n6271_, new_n533_ );
or   ( new_n6273_, new_n6272_, new_n6268_ );
and  ( new_n6274_, new_n6273_, new_n6264_ );
or   ( new_n6275_, new_n6273_, new_n6264_ );
or   ( new_n6276_, new_n610_, new_n3924_ );
or   ( new_n6277_, new_n614_, new_n3239_ );
and  ( new_n6278_, new_n6277_, new_n6276_ );
and  ( new_n6279_, new_n6278_, new_n590_ );
and  ( new_n6280_, new_n623_, RI2b1c4342df30_87 );
and  ( new_n6281_, new_n608_, RI2b1c4342deb8_86 );
or   ( new_n6282_, new_n6281_, new_n6280_ );
and  ( new_n6283_, new_n6282_, new_n619_ );
or   ( new_n6284_, new_n6283_, new_n6279_ );
and  ( new_n6285_, new_n6284_, new_n6275_ );
or   ( new_n6286_, new_n6285_, new_n6274_ );
or   ( new_n6287_, new_n753_, new_n132_ );
or   ( new_n6288_, new_n757_, new_n3902_ );
and  ( new_n6289_, new_n6288_, new_n6287_ );
and  ( new_n6290_, new_n6289_, new_n734_ );
and  ( new_n6291_, new_n766_, RI2b1c4342e020_89 );
and  ( new_n6292_, new_n751_, RI2b1c4342dfa8_88 );
or   ( new_n6293_, new_n6292_, new_n6291_ );
and  ( new_n6294_, new_n6293_, new_n762_ );
or   ( new_n6295_, new_n6294_, new_n6290_ );
or   ( new_n6296_, new_n804_, new_n117_ );
or   ( new_n6297_, new_n808_, new_n4635_ );
and  ( new_n6298_, new_n6297_, new_n6296_ );
and  ( new_n6299_, new_n6298_, new_n785_ );
and  ( new_n6300_, new_n817_, RI2b1c4342e110_91 );
and  ( new_n6301_, new_n802_, RI2b1c4342e098_90 );
or   ( new_n6302_, new_n6301_, new_n6300_ );
and  ( new_n6303_, new_n6302_, new_n813_ );
or   ( new_n6304_, new_n6303_, new_n6299_ );
and  ( new_n6305_, new_n6304_, new_n6295_ );
or   ( new_n6306_, new_n6304_, new_n6295_ );
not  ( new_n6307_, RI2b1c4342e200_93 );
or   ( new_n6308_, new_n857_, new_n6307_ );
or   ( new_n6309_, new_n861_, new_n5459_ );
and  ( new_n6310_, new_n6309_, new_n6308_ );
and  ( new_n6311_, new_n6310_, new_n842_ );
and  ( new_n6312_, new_n870_, RI2b1c4342e200_93 );
and  ( new_n6313_, new_n855_, RI2b1c4342e188_92 );
or   ( new_n6314_, new_n6313_, new_n6312_ );
and  ( new_n6315_, new_n6314_, new_n866_ );
or   ( new_n6316_, new_n6315_, new_n6311_ );
and  ( new_n6317_, new_n6316_, new_n6306_ );
or   ( new_n6318_, new_n6317_, new_n6305_ );
and  ( new_n6319_, new_n6318_, new_n6286_ );
or   ( new_n6320_, new_n6318_, new_n6286_ );
not  ( new_n6321_, RI2b1c4342e278_94 );
or   ( new_n6322_, new_n841_, new_n6321_ );
and  ( new_n6323_, new_n6322_, new_n6320_ );
or   ( new_n6324_, new_n6323_, new_n6319_ );
and  ( new_n6325_, new_n6324_, new_n6255_ );
or   ( new_n6326_, new_n6324_, new_n6255_ );
or   ( new_n6327_, new_n841_, new_n6307_ );
or   ( new_n6328_, new_n6020_, new_n5772_ );
and  ( new_n6329_, new_n6328_, new_n5782_ );
and  ( new_n6330_, new_n6016_, new_n5771_ );
and  ( new_n6331_, new_n6019_, new_n5762_ );
or   ( new_n6332_, new_n6331_, new_n6330_ );
and  ( new_n6333_, new_n6332_, new_n6024_ );
or   ( new_n6334_, new_n6333_, new_n6329_ );
and  ( new_n6335_, new_n6334_, new_n6327_ );
or   ( new_n6336_, new_n6334_, new_n6327_ );
or   ( new_n6337_, new_n6007_, new_n5803_ );
and  ( new_n6338_, new_n6337_, new_n5813_ );
and  ( new_n6339_, new_n6003_, new_n5802_ );
and  ( new_n6340_, new_n6006_, new_n5793_ );
or   ( new_n6341_, new_n6340_, new_n6339_ );
and  ( new_n6342_, new_n6341_, new_n6011_ );
or   ( new_n6343_, new_n6342_, new_n6338_ );
and  ( new_n6344_, new_n6343_, new_n6336_ );
or   ( new_n6345_, new_n6344_, new_n6335_ );
and  ( new_n6346_, new_n6345_, new_n6326_ );
or   ( new_n6347_, new_n6346_, new_n6325_ );
or   ( new_n6348_, new_n5627_, new_n5360_ );
and  ( new_n6349_, new_n6348_, new_n5370_ );
and  ( new_n6350_, new_n5623_, new_n5359_ );
and  ( new_n6351_, new_n5626_, new_n5350_ );
or   ( new_n6352_, new_n6351_, new_n6350_ );
and  ( new_n6353_, new_n6352_, new_n5631_ );
or   ( new_n6354_, new_n6353_, new_n6349_ );
or   ( new_n6355_, new_n6071_, new_n5910_ );
and  ( new_n6356_, new_n6355_, new_n5920_ );
and  ( new_n6357_, new_n6067_, new_n5909_ );
and  ( new_n6358_, new_n6070_, new_n5900_ );
or   ( new_n6359_, new_n6358_, new_n6357_ );
and  ( new_n6360_, new_n6359_, new_n6075_ );
or   ( new_n6361_, new_n6360_, new_n6356_ );
or   ( new_n6362_, new_n6056_, new_n5835_ );
and  ( new_n6363_, new_n6362_, new_n5845_ );
and  ( new_n6364_, new_n6052_, new_n5834_ );
and  ( new_n6365_, new_n6055_, new_n5825_ );
or   ( new_n6366_, new_n6365_, new_n6364_ );
and  ( new_n6367_, new_n6366_, new_n6060_ );
or   ( new_n6368_, new_n6367_, new_n6363_ );
and  ( new_n6369_, new_n6368_, new_n6361_ );
or   ( new_n6370_, new_n6368_, new_n6361_ );
or   ( new_n6371_, new_n6043_, new_n5877_ );
and  ( new_n6372_, new_n6371_, new_n5887_ );
and  ( new_n6373_, new_n6039_, new_n5876_ );
and  ( new_n6374_, new_n6042_, new_n5867_ );
or   ( new_n6375_, new_n6374_, new_n6373_ );
and  ( new_n6376_, new_n6375_, new_n6047_ );
or   ( new_n6377_, new_n6376_, new_n6372_ );
and  ( new_n6378_, new_n6377_, new_n6370_ );
or   ( new_n6379_, new_n6378_, new_n6369_ );
and  ( new_n6380_, new_n6379_, new_n6354_ );
or   ( new_n6381_, new_n6379_, new_n6354_ );
or   ( new_n6382_, new_n5614_, new_n5329_ );
and  ( new_n6383_, new_n6382_, new_n5339_ );
and  ( new_n6384_, new_n5610_, new_n5328_ );
and  ( new_n6385_, new_n5613_, new_n5319_ );
or   ( new_n6386_, new_n6385_, new_n6384_ );
and  ( new_n6387_, new_n6386_, new_n5618_ );
or   ( new_n6388_, new_n6387_, new_n6383_ );
and  ( new_n6389_, new_n6388_, new_n6381_ );
or   ( new_n6390_, new_n6389_, new_n6380_ );
and  ( new_n6391_, new_n6390_, new_n6347_ );
or   ( new_n6392_, new_n6390_, new_n6347_ );
or   ( new_n6393_, new_n6088_, new_n5941_ );
and  ( new_n6394_, new_n6393_, new_n5949_ );
and  ( new_n6395_, new_n6084_, new_n5940_ );
and  ( new_n6396_, new_n6087_, new_n5933_ );
or   ( new_n6397_, new_n6396_, new_n6395_ );
and  ( new_n6398_, new_n6397_, new_n6092_ );
or   ( new_n6399_, new_n6398_, new_n6394_ );
and  ( new_n6400_, new_n6013_, new_n5784_ );
and  ( new_n6401_, new_n6026_, new_n5815_ );
or   ( new_n6402_, new_n6401_, new_n6400_ );
and  ( new_n6403_, new_n6402_, new_n6399_ );
or   ( new_n6404_, new_n6402_, new_n6399_ );
or   ( new_n6405_, new_n6063_, new_n5890_ );
and  ( new_n6406_, new_n6405_, new_n5922_ );
and  ( new_n6407_, new_n6049_, new_n5847_ );
and  ( new_n6408_, new_n6062_, new_n5889_ );
or   ( new_n6409_, new_n6408_, new_n6407_ );
and  ( new_n6410_, new_n6409_, new_n6077_ );
or   ( new_n6411_, new_n6410_, new_n6406_ );
and  ( new_n6412_, new_n6411_, new_n6404_ );
or   ( new_n6413_, new_n6412_, new_n6403_ );
and  ( new_n6414_, new_n6413_, new_n6392_ );
or   ( new_n6415_, new_n6414_, new_n6391_ );
or   ( new_n6416_, new_n5634_, new_n5373_ );
and  ( new_n6417_, new_n6416_, new_n5405_ );
and  ( new_n6418_, new_n5620_, new_n5372_ );
and  ( new_n6419_, new_n5633_, new_n5341_ );
or   ( new_n6420_, new_n6419_, new_n6418_ );
and  ( new_n6421_, new_n6420_, new_n5648_ );
or   ( new_n6422_, new_n6421_, new_n6417_ );
or   ( new_n6423_, new_n6103_, new_n5743_ );
and  ( new_n6424_, new_n6423_, new_n5751_ );
and  ( new_n6425_, new_n6099_, new_n5742_ );
and  ( new_n6426_, new_n6102_, new_n5735_ );
or   ( new_n6427_, new_n6426_, new_n6425_ );
and  ( new_n6428_, new_n6427_, new_n6107_ );
or   ( new_n6429_, new_n6428_, new_n6424_ );
and  ( new_n6430_, new_n6429_, new_n6422_ );
or   ( new_n6431_, new_n6429_, new_n6422_ );
or   ( new_n6432_, new_n6080_, new_n5925_ );
and  ( new_n6433_, new_n6432_, new_n5951_ );
and  ( new_n6434_, new_n6079_, new_n5816_ );
and  ( new_n6435_, new_n6027_, new_n5924_ );
or   ( new_n6436_, new_n6435_, new_n6434_ );
and  ( new_n6437_, new_n6436_, new_n6094_ );
or   ( new_n6438_, new_n6437_, new_n6433_ );
and  ( new_n6439_, new_n6438_, new_n6431_ );
or   ( new_n6440_, new_n6439_, new_n6430_ );
and  ( new_n6441_, new_n6440_, new_n6415_ );
or   ( new_n6442_, new_n6440_, new_n6415_ );
or   ( new_n6443_, new_n5601_, new_n5517_ );
and  ( new_n6444_, new_n6443_, new_n5525_ );
and  ( new_n6445_, new_n5597_, new_n5516_ );
and  ( new_n6446_, new_n5600_, new_n5509_ );
or   ( new_n6447_, new_n6446_, new_n6445_ );
and  ( new_n6448_, new_n6447_, new_n5605_ );
or   ( new_n6449_, new_n6448_, new_n6444_ );
and  ( new_n6450_, new_n6449_, new_n6442_ );
or   ( new_n6451_, new_n6450_, new_n6441_ );
and  ( new_n6452_, new_n6451_, new_n6149_ );
or   ( new_n6453_, new_n6451_, new_n6149_ );
or   ( new_n6454_, new_n6117_, new_n5965_ );
and  ( new_n6455_, new_n6454_, new_n5973_ );
and  ( new_n6456_, new_n6116_, new_n5728_ );
and  ( new_n6457_, new_n6000_, new_n5964_ );
or   ( new_n6458_, new_n6457_, new_n6456_ );
and  ( new_n6459_, new_n6458_, new_n6121_ );
or   ( new_n6460_, new_n6459_, new_n6455_ );
and  ( new_n6461_, new_n6460_, new_n6453_ );
or   ( new_n6462_, new_n6461_, new_n6452_ );
and  ( new_n6463_, new_n6462_, new_n6134_ );
or   ( new_n6464_, new_n6462_, new_n6134_ );
and  ( new_n6465_, new_n6139_, new_n5500_ );
and  ( new_n6466_, new_n6135_, new_n5696_ );
or   ( new_n6467_, new_n6466_, new_n6465_ );
and  ( new_n6468_, new_n6146_, new_n5962_ );
and  ( new_n6469_, new_n6142_, new_n6114_ );
or   ( new_n6470_, new_n6469_, new_n6468_ );
and  ( new_n6471_, new_n6470_, new_n6467_ );
and  ( new_n6472_, new_n6420_, new_n5405_ );
and  ( new_n6473_, new_n6416_, new_n5648_ );
or   ( new_n6474_, new_n6473_, new_n6472_ );
and  ( new_n6475_, new_n6427_, new_n5751_ );
and  ( new_n6476_, new_n6423_, new_n6107_ );
or   ( new_n6477_, new_n6476_, new_n6475_ );
and  ( new_n6478_, new_n6477_, new_n6474_ );
or   ( new_n6479_, new_n6477_, new_n6474_ );
and  ( new_n6480_, new_n6436_, new_n5951_ );
and  ( new_n6481_, new_n6432_, new_n6094_ );
or   ( new_n6482_, new_n6481_, new_n6480_ );
and  ( new_n6483_, new_n6482_, new_n6479_ );
or   ( new_n6484_, new_n6483_, new_n6478_ );
and  ( new_n6485_, new_n6352_, new_n5370_ );
and  ( new_n6486_, new_n6348_, new_n5631_ );
or   ( new_n6487_, new_n6486_, new_n6485_ );
and  ( new_n6488_, new_n6359_, new_n5920_ );
and  ( new_n6489_, new_n6355_, new_n6075_ );
or   ( new_n6490_, new_n6489_, new_n6488_ );
and  ( new_n6491_, new_n6366_, new_n5845_ );
and  ( new_n6492_, new_n6362_, new_n6060_ );
or   ( new_n6493_, new_n6492_, new_n6491_ );
and  ( new_n6494_, new_n6493_, new_n6490_ );
or   ( new_n6495_, new_n6493_, new_n6490_ );
and  ( new_n6496_, new_n6375_, new_n5887_ );
and  ( new_n6497_, new_n6371_, new_n6047_ );
or   ( new_n6498_, new_n6497_, new_n6496_ );
and  ( new_n6499_, new_n6498_, new_n6495_ );
or   ( new_n6500_, new_n6499_, new_n6494_ );
and  ( new_n6501_, new_n6500_, new_n6487_ );
or   ( new_n6502_, new_n6500_, new_n6487_ );
and  ( new_n6503_, new_n6386_, new_n5339_ );
and  ( new_n6504_, new_n6382_, new_n5618_ );
or   ( new_n6505_, new_n6504_, new_n6503_ );
and  ( new_n6506_, new_n6505_, new_n6502_ );
or   ( new_n6507_, new_n6506_, new_n6501_ );
and  ( new_n6508_, new_n6165_, new_n6039_ );
and  ( new_n6509_, new_n6157_, new_n5867_ );
or   ( new_n6510_, new_n6509_, new_n6508_ );
and  ( new_n6511_, new_n6174_, new_n5182_ );
and  ( new_n6512_, new_n6170_, new_n5028_ );
or   ( new_n6513_, new_n6512_, new_n6511_ );
and  ( new_n6514_, new_n6513_, new_n6510_ );
or   ( new_n6515_, new_n6513_, new_n6510_ );
and  ( new_n6516_, new_n6185_, new_n4400_ );
and  ( new_n6517_, new_n6181_, new_n4215_ );
or   ( new_n6518_, new_n6517_, new_n6516_ );
and  ( new_n6519_, new_n6518_, new_n6515_ );
or   ( new_n6520_, new_n6519_, new_n6514_ );
and  ( new_n6521_, new_n6196_, new_n3695_ );
and  ( new_n6522_, new_n6192_, new_n3548_ );
or   ( new_n6523_, new_n6522_, new_n6521_ );
and  ( new_n6524_, new_n6205_, new_n3004_ );
and  ( new_n6525_, new_n6201_, new_n2868_ );
or   ( new_n6526_, new_n6525_, new_n6524_ );
and  ( new_n6527_, new_n6526_, new_n6523_ );
or   ( new_n6528_, new_n6526_, new_n6523_ );
and  ( new_n6529_, new_n6216_, new_n2334_ );
and  ( new_n6530_, new_n6212_, new_n2168_ );
or   ( new_n6531_, new_n6530_, new_n6529_ );
and  ( new_n6532_, new_n6531_, new_n6528_ );
or   ( new_n6533_, new_n6532_, new_n6527_ );
and  ( new_n6534_, new_n6533_, new_n6520_ );
or   ( new_n6535_, new_n6533_, new_n6520_ );
and  ( new_n6536_, new_n6229_, new_n1824_ );
and  ( new_n6537_, new_n6225_, new_n1717_ );
or   ( new_n6538_, new_n6537_, new_n6536_ );
and  ( new_n6539_, new_n6238_, new_n1355_ );
and  ( new_n6540_, new_n6234_, new_n1267_ );
or   ( new_n6541_, new_n6540_, new_n6539_ );
and  ( new_n6542_, new_n6541_, new_n6538_ );
or   ( new_n6543_, new_n6541_, new_n6538_ );
and  ( new_n6544_, new_n6249_, new_n913_ );
and  ( new_n6545_, new_n6245_, new_n938_ );
or   ( new_n6546_, new_n6545_, new_n6544_ );
and  ( new_n6547_, new_n6546_, new_n6543_ );
or   ( new_n6548_, new_n6547_, new_n6542_ );
and  ( new_n6549_, new_n6548_, new_n6535_ );
or   ( new_n6550_, new_n6549_, new_n6534_ );
and  ( new_n6551_, new_n6262_, new_n428_ );
and  ( new_n6552_, new_n6258_, new_n457_ );
or   ( new_n6553_, new_n6552_, new_n6551_ );
and  ( new_n6554_, new_n6271_, new_n505_ );
and  ( new_n6555_, new_n6267_, new_n533_ );
or   ( new_n6556_, new_n6555_, new_n6554_ );
and  ( new_n6557_, new_n6556_, new_n6553_ );
or   ( new_n6558_, new_n6556_, new_n6553_ );
and  ( new_n6559_, new_n6282_, new_n590_ );
and  ( new_n6560_, new_n6278_, new_n619_ );
or   ( new_n6561_, new_n6560_, new_n6559_ );
and  ( new_n6562_, new_n6561_, new_n6558_ );
or   ( new_n6563_, new_n6562_, new_n6557_ );
and  ( new_n6564_, new_n6293_, new_n734_ );
and  ( new_n6565_, new_n6289_, new_n762_ );
or   ( new_n6566_, new_n6565_, new_n6564_ );
and  ( new_n6567_, new_n6302_, new_n785_ );
and  ( new_n6568_, new_n6298_, new_n813_ );
or   ( new_n6569_, new_n6568_, new_n6567_ );
and  ( new_n6570_, new_n6569_, new_n6566_ );
or   ( new_n6571_, new_n6569_, new_n6566_ );
and  ( new_n6572_, new_n6314_, new_n842_ );
and  ( new_n6573_, new_n6310_, new_n866_ );
or   ( new_n6574_, new_n6573_, new_n6572_ );
and  ( new_n6575_, new_n6574_, new_n6571_ );
or   ( new_n6576_, new_n6575_, new_n6570_ );
or   ( new_n6577_, new_n6576_, new_n6563_ );
and  ( new_n6578_, new_n6576_, new_n6563_ );
and  ( new_n6579_, new_n720_, RI2b1c4342e278_94 );
or   ( new_n6580_, new_n6579_, new_n6578_ );
and  ( new_n6581_, new_n6580_, new_n6577_ );
or   ( new_n6582_, new_n6581_, new_n6550_ );
and  ( new_n6583_, new_n6581_, new_n6550_ );
and  ( new_n6584_, new_n720_, RI2b1c4342e200_93 );
and  ( new_n6585_, new_n6332_, new_n5782_ );
and  ( new_n6586_, new_n6328_, new_n6024_ );
or   ( new_n6587_, new_n6586_, new_n6585_ );
and  ( new_n6588_, new_n6587_, new_n6584_ );
or   ( new_n6589_, new_n6587_, new_n6584_ );
and  ( new_n6590_, new_n6341_, new_n5813_ );
and  ( new_n6591_, new_n6337_, new_n6011_ );
or   ( new_n6592_, new_n6591_, new_n6590_ );
and  ( new_n6593_, new_n6592_, new_n6589_ );
or   ( new_n6594_, new_n6593_, new_n6588_ );
or   ( new_n6595_, new_n6594_, new_n6583_ );
and  ( new_n6596_, new_n6595_, new_n6582_ );
or   ( new_n6597_, new_n6596_, new_n6507_ );
and  ( new_n6598_, new_n6596_, new_n6507_ );
and  ( new_n6599_, new_n6397_, new_n5949_ );
and  ( new_n6600_, new_n6393_, new_n6092_ );
or   ( new_n6601_, new_n6600_, new_n6599_ );
and  ( new_n6602_, new_n6026_, new_n6013_ );
or   ( new_n6603_, new_n6602_, new_n5816_ );
and  ( new_n6604_, new_n6603_, new_n6601_ );
or   ( new_n6605_, new_n6603_, new_n6601_ );
and  ( new_n6606_, new_n6409_, new_n5922_ );
and  ( new_n6607_, new_n6405_, new_n6077_ );
or   ( new_n6608_, new_n6607_, new_n6606_ );
and  ( new_n6609_, new_n6608_, new_n6605_ );
or   ( new_n6610_, new_n6609_, new_n6604_ );
or   ( new_n6611_, new_n6610_, new_n6598_ );
and  ( new_n6612_, new_n6611_, new_n6597_ );
or   ( new_n6613_, new_n6612_, new_n6484_ );
and  ( new_n6614_, new_n6612_, new_n6484_ );
and  ( new_n6615_, new_n6447_, new_n5525_ );
and  ( new_n6616_, new_n6443_, new_n5605_ );
or   ( new_n6617_, new_n6616_, new_n6615_ );
or   ( new_n6618_, new_n6617_, new_n6614_ );
and  ( new_n6619_, new_n6618_, new_n6613_ );
and  ( new_n6620_, new_n6619_, new_n6471_ );
or   ( new_n6621_, new_n6620_, new_n6452_ );
and  ( new_n6622_, new_n6621_, new_n6460_ );
and  ( new_n6623_, new_n6619_, new_n6149_ );
and  ( new_n6624_, new_n6471_, new_n6451_ );
or   ( new_n6625_, new_n6624_, new_n6623_ );
and  ( new_n6626_, new_n6458_, new_n5973_ );
and  ( new_n6627_, new_n6454_, new_n6121_ );
or   ( new_n6628_, new_n6627_, new_n6626_ );
and  ( new_n6629_, new_n6628_, new_n6625_ );
or   ( new_n6630_, new_n6629_, new_n6622_ );
and  ( new_n6631_, new_n6148_, new_n6141_ );
or   ( new_n6632_, new_n6631_, new_n6471_ );
or   ( new_n6633_, new_n6478_, new_n6430_ );
and  ( new_n6634_, new_n6633_, new_n6438_ );
and  ( new_n6635_, new_n6474_, new_n6429_ );
and  ( new_n6636_, new_n6477_, new_n6422_ );
or   ( new_n6637_, new_n6636_, new_n6635_ );
and  ( new_n6638_, new_n6637_, new_n6482_ );
or   ( new_n6639_, new_n6638_, new_n6634_ );
or   ( new_n6640_, new_n934_, new_n2119_ );
or   ( new_n6641_, new_n940_, new_n126_ );
and  ( new_n6642_, new_n6641_, new_n6640_ );
and  ( new_n6643_, new_n6642_, new_n913_ );
and  ( new_n6644_, new_n944_, RI2b1c4342dcd8_82 );
and  ( new_n6645_, new_n932_, RI2b1c4342dc60_81 );
or   ( new_n6646_, new_n6645_, new_n6644_ );
and  ( new_n6647_, new_n6646_, new_n938_ );
or   ( new_n6648_, new_n6647_, new_n6643_ );
or   ( new_n6649_, new_n453_, new_n2541_ );
or   ( new_n6650_, new_n459_, new_n121_ );
and  ( new_n6651_, new_n6650_, new_n6649_ );
and  ( new_n6652_, new_n6651_, new_n428_ );
and  ( new_n6653_, new_n463_, RI2b1c4342ddc8_84 );
and  ( new_n6654_, new_n451_, RI2b1c4342dd50_83 );
or   ( new_n6655_, new_n6654_, new_n6653_ );
and  ( new_n6656_, new_n6655_, new_n457_ );
or   ( new_n6657_, new_n6656_, new_n6652_ );
and  ( new_n6658_, new_n6657_, new_n6648_ );
or   ( new_n6659_, new_n6657_, new_n6648_ );
or   ( new_n6660_, new_n524_, new_n3239_ );
or   ( new_n6661_, new_n528_, new_n2806_ );
and  ( new_n6662_, new_n6661_, new_n6660_ );
and  ( new_n6663_, new_n6662_, new_n505_ );
and  ( new_n6664_, new_n537_, RI2b1c4342deb8_86 );
and  ( new_n6665_, new_n522_, RI2b1c4342de40_85 );
or   ( new_n6666_, new_n6665_, new_n6664_ );
and  ( new_n6667_, new_n6666_, new_n533_ );
or   ( new_n6668_, new_n6667_, new_n6663_ );
and  ( new_n6669_, new_n6668_, new_n6659_ );
or   ( new_n6670_, new_n6669_, new_n6658_ );
or   ( new_n6671_, new_n610_, new_n3902_ );
or   ( new_n6672_, new_n614_, new_n3924_ );
and  ( new_n6673_, new_n6672_, new_n6671_ );
and  ( new_n6674_, new_n6673_, new_n590_ );
and  ( new_n6675_, new_n623_, RI2b1c4342dfa8_88 );
and  ( new_n6676_, new_n608_, RI2b1c4342df30_87 );
or   ( new_n6677_, new_n6676_, new_n6675_ );
and  ( new_n6678_, new_n6677_, new_n619_ );
or   ( new_n6679_, new_n6678_, new_n6674_ );
or   ( new_n6680_, new_n753_, new_n4635_ );
or   ( new_n6681_, new_n757_, new_n132_ );
and  ( new_n6682_, new_n6681_, new_n6680_ );
and  ( new_n6683_, new_n6682_, new_n734_ );
and  ( new_n6684_, new_n766_, RI2b1c4342e098_90 );
and  ( new_n6685_, new_n751_, RI2b1c4342e020_89 );
or   ( new_n6686_, new_n6685_, new_n6684_ );
and  ( new_n6687_, new_n6686_, new_n762_ );
or   ( new_n6688_, new_n6687_, new_n6683_ );
and  ( new_n6689_, new_n6688_, new_n6679_ );
or   ( new_n6690_, new_n6688_, new_n6679_ );
or   ( new_n6691_, new_n804_, new_n5459_ );
or   ( new_n6692_, new_n808_, new_n117_ );
and  ( new_n6693_, new_n6692_, new_n6691_ );
and  ( new_n6694_, new_n6693_, new_n785_ );
and  ( new_n6695_, new_n817_, RI2b1c4342e188_92 );
and  ( new_n6696_, new_n802_, RI2b1c4342e110_91 );
or   ( new_n6697_, new_n6696_, new_n6695_ );
and  ( new_n6698_, new_n6697_, new_n813_ );
or   ( new_n6699_, new_n6698_, new_n6694_ );
and  ( new_n6700_, new_n6699_, new_n6690_ );
or   ( new_n6701_, new_n6700_, new_n6689_ );
and  ( new_n6702_, new_n6701_, new_n6670_ );
or   ( new_n6703_, new_n6701_, new_n6670_ );
or   ( new_n6704_, new_n841_, new_n124_ );
or   ( new_n6705_, new_n857_, new_n6321_ );
or   ( new_n6706_, new_n861_, new_n6307_ );
and  ( new_n6707_, new_n6706_, new_n6705_ );
and  ( new_n6708_, new_n6707_, new_n842_ );
and  ( new_n6709_, new_n870_, RI2b1c4342e278_94 );
and  ( new_n6710_, new_n855_, RI2b1c4342e200_93 );
or   ( new_n6711_, new_n6710_, new_n6709_ );
and  ( new_n6712_, new_n6711_, new_n866_ );
or   ( new_n6713_, new_n6712_, new_n6708_ );
and  ( new_n6714_, new_n6713_, new_n6704_ );
and  ( new_n6715_, new_n6714_, new_n6703_ );
or   ( new_n6716_, new_n6715_, new_n6702_ );
or   ( new_n6717_, new_n4535_, new_n755_ );
or   ( new_n6718_, new_n4539_, new_n591_ );
and  ( new_n6719_, new_n6718_, new_n6717_ );
and  ( new_n6720_, new_n6719_, new_n4400_ );
and  ( new_n6721_, new_n4543_, RI2b1c4342d738_70 );
and  ( new_n6722_, new_n4533_, RI2b1c4342d6c0_69 );
or   ( new_n6723_, new_n6722_, new_n6721_ );
and  ( new_n6724_, new_n6723_, new_n4215_ );
or   ( new_n6725_, new_n6724_, new_n6720_ );
or   ( new_n6726_, new_n3802_, new_n806_ );
or   ( new_n6727_, new_n3806_, new_n110_ );
and  ( new_n6728_, new_n6727_, new_n6726_ );
and  ( new_n6729_, new_n6728_, new_n3695_ );
and  ( new_n6730_, new_n3810_, RI2b1c4342d828_72 );
and  ( new_n6731_, new_n3800_, RI2b1c4342d7b0_71 );
or   ( new_n6732_, new_n6731_, new_n6730_ );
and  ( new_n6733_, new_n6732_, new_n3548_ );
or   ( new_n6734_, new_n6733_, new_n6729_ );
and  ( new_n6735_, new_n6734_, new_n6725_ );
or   ( new_n6736_, new_n6734_, new_n6725_ );
or   ( new_n6737_, new_n3112_, new_n859_ );
or   ( new_n6738_, new_n3116_, new_n105_ );
and  ( new_n6739_, new_n6738_, new_n6737_ );
and  ( new_n6740_, new_n6739_, new_n3004_ );
and  ( new_n6741_, new_n3120_, RI2b1c4342d918_74 );
and  ( new_n6742_, new_n3110_, RI2b1c4342d8a0_73 );
or   ( new_n6743_, new_n6742_, new_n6741_ );
and  ( new_n6744_, new_n6743_, new_n2868_ );
or   ( new_n6745_, new_n6744_, new_n6740_ );
and  ( new_n6746_, new_n6745_, new_n6736_ );
or   ( new_n6747_, new_n6746_, new_n6735_ );
or   ( new_n6748_, new_n6156_, new_n526_ );
or   ( new_n6749_, new_n6160_, new_n99_ );
and  ( new_n6750_, new_n6749_, new_n6748_ );
and  ( new_n6751_, new_n6750_, new_n6039_ );
and  ( new_n6752_, new_n6164_, RI2b1c4342d558_66 );
and  ( new_n6753_, new_n6154_, RI2b1c4342d4e0_65 );
or   ( new_n6754_, new_n6753_, new_n6752_ );
and  ( new_n6755_, new_n6754_, new_n5867_ );
or   ( new_n6756_, new_n6755_, new_n6751_ );
and  ( new_n6757_, new_n6756_, new_n6037_ );
or   ( new_n6758_, new_n6756_, new_n6037_ );
or   ( new_n6759_, new_n5308_, new_n612_ );
or   ( new_n6760_, new_n5312_, new_n112_ );
and  ( new_n6761_, new_n6760_, new_n6759_ );
and  ( new_n6762_, new_n6761_, new_n5182_ );
and  ( new_n6763_, new_n5316_, RI2b1c4342d648_68 );
and  ( new_n6764_, new_n5306_, RI2b1c4342d5d0_67 );
or   ( new_n6765_, new_n6764_, new_n6763_ );
and  ( new_n6766_, new_n6765_, new_n5028_ );
or   ( new_n6767_, new_n6766_, new_n6762_ );
and  ( new_n6768_, new_n6767_, new_n6758_ );
or   ( new_n6769_, new_n6768_, new_n6757_ );
and  ( new_n6770_, new_n6769_, new_n6747_ );
or   ( new_n6771_, new_n6769_, new_n6747_ );
or   ( new_n6772_, new_n2450_, new_n886_ );
or   ( new_n6773_, new_n2454_, new_n843_ );
and  ( new_n6774_, new_n6773_, new_n6772_ );
and  ( new_n6775_, new_n6774_, new_n2334_ );
and  ( new_n6776_, new_n2458_, RI2b1c4342da08_76 );
and  ( new_n6777_, new_n2448_, RI2b1c4342d990_75 );
or   ( new_n6778_, new_n6777_, new_n6776_ );
and  ( new_n6779_, new_n6778_, new_n2168_ );
or   ( new_n6780_, new_n6779_, new_n6775_ );
or   ( new_n6781_, new_n1910_, new_n1002_ );
or   ( new_n6782_, new_n1914_, new_n1004_ );
and  ( new_n6783_, new_n6782_, new_n6781_ );
and  ( new_n6784_, new_n6783_, new_n1824_ );
and  ( new_n6785_, new_n1918_, RI2b1c4342daf8_78 );
and  ( new_n6786_, new_n1908_, RI2b1c4342da80_77 );
or   ( new_n6787_, new_n6786_, new_n6785_ );
and  ( new_n6788_, new_n6787_, new_n1717_ );
or   ( new_n6789_, new_n6788_, new_n6784_ );
and  ( new_n6790_, new_n6789_, new_n6780_ );
or   ( new_n6791_, new_n6789_, new_n6780_ );
or   ( new_n6792_, new_n1425_, new_n1511_ );
or   ( new_n6793_, new_n1429_, new_n1310_ );
and  ( new_n6794_, new_n6793_, new_n6792_ );
and  ( new_n6795_, new_n6794_, new_n1355_ );
and  ( new_n6796_, new_n1433_, RI2b1c4342dbe8_80 );
and  ( new_n6797_, new_n1423_, RI2b1c4342db70_79 );
or   ( new_n6798_, new_n6797_, new_n6796_ );
and  ( new_n6799_, new_n6798_, new_n1267_ );
or   ( new_n6800_, new_n6799_, new_n6795_ );
and  ( new_n6801_, new_n6800_, new_n6791_ );
or   ( new_n6802_, new_n6801_, new_n6790_ );
and  ( new_n6803_, new_n6802_, new_n6771_ );
or   ( new_n6804_, new_n6803_, new_n6770_ );
and  ( new_n6805_, new_n6804_, new_n6716_ );
or   ( new_n6806_, new_n6804_, new_n6716_ );
or   ( new_n6807_, new_n6570_, new_n6305_ );
and  ( new_n6808_, new_n6807_, new_n6316_ );
and  ( new_n6809_, new_n6566_, new_n6304_ );
and  ( new_n6810_, new_n6569_, new_n6295_ );
or   ( new_n6811_, new_n6810_, new_n6809_ );
and  ( new_n6812_, new_n6811_, new_n6574_ );
or   ( new_n6813_, new_n6812_, new_n6808_ );
and  ( new_n6814_, new_n6813_, new_n6579_ );
or   ( new_n6815_, new_n6813_, new_n6579_ );
or   ( new_n6816_, new_n6557_, new_n6274_ );
and  ( new_n6817_, new_n6816_, new_n6284_ );
and  ( new_n6818_, new_n6553_, new_n6273_ );
and  ( new_n6819_, new_n6556_, new_n6264_ );
or   ( new_n6820_, new_n6819_, new_n6818_ );
and  ( new_n6821_, new_n6820_, new_n6561_ );
or   ( new_n6822_, new_n6821_, new_n6817_ );
and  ( new_n6823_, new_n6822_, new_n6815_ );
or   ( new_n6824_, new_n6823_, new_n6814_ );
and  ( new_n6825_, new_n6824_, new_n6806_ );
or   ( new_n6826_, new_n6825_, new_n6805_ );
or   ( new_n6827_, new_n6494_, new_n6369_ );
and  ( new_n6828_, new_n6827_, new_n6377_ );
and  ( new_n6829_, new_n6490_, new_n6368_ );
and  ( new_n6830_, new_n6493_, new_n6361_ );
or   ( new_n6831_, new_n6830_, new_n6829_ );
and  ( new_n6832_, new_n6831_, new_n6498_ );
or   ( new_n6833_, new_n6832_, new_n6828_ );
or   ( new_n6834_, new_n6542_, new_n6241_ );
and  ( new_n6835_, new_n6834_, new_n6251_ );
and  ( new_n6836_, new_n6538_, new_n6240_ );
and  ( new_n6837_, new_n6541_, new_n6231_ );
or   ( new_n6838_, new_n6837_, new_n6836_ );
and  ( new_n6839_, new_n6838_, new_n6546_ );
or   ( new_n6840_, new_n6839_, new_n6835_ );
or   ( new_n6841_, new_n6527_, new_n6208_ );
and  ( new_n6842_, new_n6841_, new_n6218_ );
and  ( new_n6843_, new_n6523_, new_n6207_ );
and  ( new_n6844_, new_n6526_, new_n6198_ );
or   ( new_n6845_, new_n6844_, new_n6843_ );
and  ( new_n6846_, new_n6845_, new_n6531_ );
or   ( new_n6847_, new_n6846_, new_n6842_ );
and  ( new_n6848_, new_n6847_, new_n6840_ );
or   ( new_n6849_, new_n6847_, new_n6840_ );
or   ( new_n6850_, new_n6514_, new_n6177_ );
and  ( new_n6851_, new_n6850_, new_n6187_ );
and  ( new_n6852_, new_n6510_, new_n6176_ );
and  ( new_n6853_, new_n6513_, new_n6167_ );
or   ( new_n6854_, new_n6853_, new_n6852_ );
and  ( new_n6855_, new_n6854_, new_n6518_ );
or   ( new_n6856_, new_n6855_, new_n6851_ );
and  ( new_n6857_, new_n6856_, new_n6849_ );
or   ( new_n6858_, new_n6857_, new_n6848_ );
and  ( new_n6859_, new_n6858_, new_n6833_ );
or   ( new_n6860_, new_n6858_, new_n6833_ );
or   ( new_n6861_, new_n6588_, new_n6335_ );
and  ( new_n6862_, new_n6861_, new_n6343_ );
and  ( new_n6863_, new_n6584_, new_n6334_ );
and  ( new_n6864_, new_n6587_, new_n6327_ );
or   ( new_n6865_, new_n6864_, new_n6863_ );
and  ( new_n6866_, new_n6865_, new_n6592_ );
or   ( new_n6867_, new_n6866_, new_n6862_ );
and  ( new_n6868_, new_n6867_, new_n6860_ );
or   ( new_n6869_, new_n6868_, new_n6859_ );
and  ( new_n6870_, new_n6869_, new_n6826_ );
or   ( new_n6871_, new_n6869_, new_n6826_ );
or   ( new_n6872_, new_n6604_, new_n6403_ );
and  ( new_n6873_, new_n6872_, new_n6411_ );
and  ( new_n6874_, new_n6601_, new_n6402_ );
and  ( new_n6875_, new_n6603_, new_n6399_ );
or   ( new_n6876_, new_n6875_, new_n6874_ );
and  ( new_n6877_, new_n6876_, new_n6608_ );
or   ( new_n6878_, new_n6877_, new_n6873_ );
and  ( new_n6879_, new_n6878_, new_n6871_ );
or   ( new_n6880_, new_n6879_, new_n6870_ );
and  ( new_n6881_, new_n6880_, new_n6639_ );
or   ( new_n6882_, new_n6880_, new_n6639_ );
or   ( new_n6883_, new_n6598_, new_n6391_ );
and  ( new_n6884_, new_n6883_, new_n6413_ );
and  ( new_n6885_, new_n6596_, new_n6390_ );
and  ( new_n6886_, new_n6507_, new_n6347_ );
or   ( new_n6887_, new_n6886_, new_n6885_ );
and  ( new_n6888_, new_n6887_, new_n6610_ );
or   ( new_n6889_, new_n6888_, new_n6884_ );
and  ( new_n6890_, new_n6889_, new_n6882_ );
or   ( new_n6891_, new_n6890_, new_n6881_ );
and  ( new_n6892_, new_n6891_, new_n6632_ );
or   ( new_n6893_, new_n6891_, new_n6632_ );
or   ( new_n6894_, new_n6614_, new_n6441_ );
and  ( new_n6895_, new_n6894_, new_n6449_ );
and  ( new_n6896_, new_n6612_, new_n6440_ );
and  ( new_n6897_, new_n6484_, new_n6415_ );
or   ( new_n6898_, new_n6897_, new_n6896_ );
and  ( new_n6899_, new_n6898_, new_n6617_ );
or   ( new_n6900_, new_n6899_, new_n6895_ );
and  ( new_n6901_, new_n6900_, new_n6893_ );
or   ( new_n6902_, new_n6901_, new_n6892_ );
or   ( new_n6903_, new_n6902_, new_n6630_ );
and  ( new_n6904_, new_n6903_, new_n6464_ );
or   ( new_n6905_, new_n6904_, new_n6463_ );
and  ( new_n6906_, new_n6902_, new_n6630_ );
or   ( new_n6907_, new_n6906_, new_n6463_ );
and  ( new_n6908_, new_n6467_, new_n6148_ );
and  ( new_n6909_, new_n6470_, new_n6141_ );
or   ( new_n6910_, new_n6909_, new_n6908_ );
and  ( new_n6911_, new_n6637_, new_n6438_ );
and  ( new_n6912_, new_n6633_, new_n6482_ );
or   ( new_n6913_, new_n6912_, new_n6911_ );
and  ( new_n6914_, new_n6754_, new_n6039_ );
and  ( new_n6915_, new_n6750_, new_n5867_ );
or   ( new_n6916_, new_n6915_, new_n6914_ );
and  ( new_n6917_, new_n6916_, new_n5858_ );
or   ( new_n6918_, new_n6916_, new_n5858_ );
and  ( new_n6919_, new_n6765_, new_n5182_ );
and  ( new_n6920_, new_n6761_, new_n5028_ );
or   ( new_n6921_, new_n6920_, new_n6919_ );
and  ( new_n6922_, new_n6921_, new_n6918_ );
or   ( new_n6923_, new_n6922_, new_n6917_ );
and  ( new_n6924_, new_n6723_, new_n4400_ );
and  ( new_n6925_, new_n6719_, new_n4215_ );
or   ( new_n6926_, new_n6925_, new_n6924_ );
and  ( new_n6927_, new_n6732_, new_n3695_ );
and  ( new_n6928_, new_n6728_, new_n3548_ );
or   ( new_n6929_, new_n6928_, new_n6927_ );
and  ( new_n6930_, new_n6929_, new_n6926_ );
or   ( new_n6931_, new_n6929_, new_n6926_ );
and  ( new_n6932_, new_n6743_, new_n3004_ );
and  ( new_n6933_, new_n6739_, new_n2868_ );
or   ( new_n6934_, new_n6933_, new_n6932_ );
and  ( new_n6935_, new_n6934_, new_n6931_ );
or   ( new_n6936_, new_n6935_, new_n6930_ );
and  ( new_n6937_, new_n6936_, new_n6923_ );
or   ( new_n6938_, new_n6936_, new_n6923_ );
and  ( new_n6939_, new_n6778_, new_n2334_ );
and  ( new_n6940_, new_n6774_, new_n2168_ );
or   ( new_n6941_, new_n6940_, new_n6939_ );
and  ( new_n6942_, new_n6787_, new_n1824_ );
and  ( new_n6943_, new_n6783_, new_n1717_ );
or   ( new_n6944_, new_n6943_, new_n6942_ );
and  ( new_n6945_, new_n6944_, new_n6941_ );
or   ( new_n6946_, new_n6944_, new_n6941_ );
and  ( new_n6947_, new_n6798_, new_n1355_ );
and  ( new_n6948_, new_n6794_, new_n1267_ );
or   ( new_n6949_, new_n6948_, new_n6947_ );
and  ( new_n6950_, new_n6949_, new_n6946_ );
or   ( new_n6951_, new_n6950_, new_n6945_ );
and  ( new_n6952_, new_n6951_, new_n6938_ );
or   ( new_n6953_, new_n6952_, new_n6937_ );
and  ( new_n6954_, new_n6646_, new_n913_ );
and  ( new_n6955_, new_n6642_, new_n938_ );
or   ( new_n6956_, new_n6955_, new_n6954_ );
and  ( new_n6957_, new_n6655_, new_n428_ );
and  ( new_n6958_, new_n6651_, new_n457_ );
or   ( new_n6959_, new_n6958_, new_n6957_ );
and  ( new_n6960_, new_n6959_, new_n6956_ );
or   ( new_n6961_, new_n6959_, new_n6956_ );
and  ( new_n6962_, new_n6666_, new_n505_ );
and  ( new_n6963_, new_n6662_, new_n533_ );
or   ( new_n6964_, new_n6963_, new_n6962_ );
and  ( new_n6965_, new_n6964_, new_n6961_ );
or   ( new_n6966_, new_n6965_, new_n6960_ );
and  ( new_n6967_, new_n6677_, new_n590_ );
and  ( new_n6968_, new_n6673_, new_n619_ );
or   ( new_n6969_, new_n6968_, new_n6967_ );
and  ( new_n6970_, new_n6686_, new_n734_ );
and  ( new_n6971_, new_n6682_, new_n762_ );
or   ( new_n6972_, new_n6971_, new_n6970_ );
and  ( new_n6973_, new_n6972_, new_n6969_ );
or   ( new_n6974_, new_n6972_, new_n6969_ );
and  ( new_n6975_, new_n6697_, new_n785_ );
and  ( new_n6976_, new_n6693_, new_n813_ );
or   ( new_n6977_, new_n6976_, new_n6975_ );
and  ( new_n6978_, new_n6977_, new_n6974_ );
or   ( new_n6979_, new_n6978_, new_n6973_ );
and  ( new_n6980_, new_n6979_, new_n6966_ );
or   ( new_n6981_, new_n6979_, new_n6966_ );
and  ( new_n6982_, new_n6711_, new_n842_ );
and  ( new_n6983_, new_n6707_, new_n866_ );
or   ( new_n6984_, new_n6983_, new_n6982_ );
and  ( new_n6985_, new_n720_, RI2b1c4342e2f0_95 );
or   ( new_n6986_, new_n6985_, new_n6984_ );
and  ( new_n6987_, new_n6986_, new_n6981_ );
or   ( new_n6988_, new_n6987_, new_n6980_ );
and  ( new_n6989_, new_n6988_, new_n6953_ );
or   ( new_n6990_, new_n6988_, new_n6953_ );
and  ( new_n6991_, new_n6811_, new_n6316_ );
and  ( new_n6992_, new_n6807_, new_n6574_ );
or   ( new_n6993_, new_n6992_, new_n6991_ );
and  ( new_n6994_, new_n6993_, new_n6322_ );
or   ( new_n6995_, new_n6993_, new_n6322_ );
and  ( new_n6996_, new_n6820_, new_n6284_ );
and  ( new_n6997_, new_n6816_, new_n6561_ );
or   ( new_n6998_, new_n6997_, new_n6996_ );
and  ( new_n6999_, new_n6998_, new_n6995_ );
or   ( new_n7000_, new_n6999_, new_n6994_ );
and  ( new_n7001_, new_n7000_, new_n6990_ );
or   ( new_n7002_, new_n7001_, new_n6989_ );
and  ( new_n7003_, new_n6831_, new_n6377_ );
and  ( new_n7004_, new_n6827_, new_n6498_ );
or   ( new_n7005_, new_n7004_, new_n7003_ );
and  ( new_n7006_, new_n6838_, new_n6251_ );
and  ( new_n7007_, new_n6834_, new_n6546_ );
or   ( new_n7008_, new_n7007_, new_n7006_ );
and  ( new_n7009_, new_n6845_, new_n6218_ );
and  ( new_n7010_, new_n6841_, new_n6531_ );
or   ( new_n7011_, new_n7010_, new_n7009_ );
and  ( new_n7012_, new_n7011_, new_n7008_ );
or   ( new_n7013_, new_n7011_, new_n7008_ );
and  ( new_n7014_, new_n6854_, new_n6187_ );
and  ( new_n7015_, new_n6850_, new_n6518_ );
or   ( new_n7016_, new_n7015_, new_n7014_ );
and  ( new_n7017_, new_n7016_, new_n7013_ );
or   ( new_n7018_, new_n7017_, new_n7012_ );
and  ( new_n7019_, new_n7018_, new_n7005_ );
or   ( new_n7020_, new_n7018_, new_n7005_ );
and  ( new_n7021_, new_n6865_, new_n6343_ );
and  ( new_n7022_, new_n6861_, new_n6592_ );
or   ( new_n7023_, new_n7022_, new_n7021_ );
and  ( new_n7024_, new_n7023_, new_n7020_ );
or   ( new_n7025_, new_n7024_, new_n7019_ );
and  ( new_n7026_, new_n7025_, new_n7002_ );
and  ( new_n7027_, new_n6876_, new_n6411_ );
and  ( new_n7028_, new_n6872_, new_n6608_ );
or   ( new_n7029_, new_n7028_, new_n7027_ );
or   ( new_n7030_, new_n7025_, new_n7002_ );
and  ( new_n7031_, new_n7030_, new_n7029_ );
or   ( new_n7032_, new_n7031_, new_n7026_ );
and  ( new_n7033_, new_n7032_, new_n6913_ );
and  ( new_n7034_, new_n6887_, new_n6413_ );
and  ( new_n7035_, new_n6883_, new_n6610_ );
or   ( new_n7036_, new_n7035_, new_n7034_ );
or   ( new_n7037_, new_n7032_, new_n6913_ );
and  ( new_n7038_, new_n7037_, new_n7036_ );
or   ( new_n7039_, new_n7038_, new_n7033_ );
and  ( new_n7040_, new_n7039_, new_n6910_ );
or   ( new_n7041_, new_n7040_, new_n6892_ );
and  ( new_n7042_, new_n7041_, new_n6900_ );
and  ( new_n7043_, new_n7039_, new_n6632_ );
and  ( new_n7044_, new_n6910_, new_n6891_ );
or   ( new_n7045_, new_n7044_, new_n7043_ );
and  ( new_n7046_, new_n6898_, new_n6449_ );
and  ( new_n7047_, new_n6894_, new_n6617_ );
or   ( new_n7048_, new_n7047_, new_n7046_ );
and  ( new_n7049_, new_n7048_, new_n7045_ );
or   ( new_n7050_, new_n7049_, new_n7042_ );
or   ( new_n7051_, new_n6583_, new_n6325_ );
and  ( new_n7052_, new_n7051_, new_n6345_ );
and  ( new_n7053_, new_n6550_, new_n6324_ );
and  ( new_n7054_, new_n6581_, new_n6255_ );
or   ( new_n7055_, new_n7054_, new_n7053_ );
and  ( new_n7056_, new_n7055_, new_n6594_ );
or   ( new_n7057_, new_n7056_, new_n7052_ );
or   ( new_n7058_, new_n7026_, new_n6870_ );
and  ( new_n7059_, new_n7058_, new_n6878_ );
and  ( new_n7060_, new_n7002_, new_n6869_ );
and  ( new_n7061_, new_n7025_, new_n6826_ );
or   ( new_n7062_, new_n7061_, new_n7060_ );
and  ( new_n7063_, new_n7062_, new_n7029_ );
or   ( new_n7064_, new_n7063_, new_n7059_ );
or   ( new_n7065_, new_n7064_, new_n7057_ );
xor  ( new_n7066_, RI2b1c4342d0a8_56, new_n173_ );
xor  ( new_n7067_, RI2b1c4342cec8_52, new_n157_ );
xor  ( new_n7068_, new_n7067_, new_n7066_ );
xor  ( new_n7069_, new_n7068_, new_n5850_ );
xor  ( new_n7070_, RI2b1c4342d198_58, RI2b1c4342d120_57 );
xor  ( new_n7071_, RI2b1c4342d378_62, RI2b1c4342d300_61 );
xor  ( new_n7072_, new_n7071_, new_n7070_ );
xor  ( new_n7073_, RI2b1c4342cce8_48, RI2b1c4342cc70_47 );
xor  ( new_n7074_, RI2b1c4342c658_34, new_n670_ );
xor  ( new_n7075_, RI2b1c4342c838_38, RI2b1c4342c7c0_37 );
xor  ( new_n7076_, new_n7075_, new_n7074_ );
xor  ( new_n7077_, new_n7076_, new_n7073_ );
xor  ( new_n7078_, RI2b1c4342cb08_44, RI2b1c4342ca90_43 );
xor  ( new_n7079_, RI2b1c4342ca18_42, new_n482_ );
xor  ( new_n7080_, RI2b1c4342cbf8_46, RI2b1c4342cb80_45 );
xor  ( new_n7081_, new_n7080_, new_n7079_ );
xor  ( new_n7082_, new_n7081_, new_n7078_ );
xor  ( new_n7083_, RI2b1c4342c928_40, new_n567_ );
xor  ( new_n7084_, RI2b1c4342c748_36, new_n659_ );
xor  ( new_n7085_, new_n7084_, new_n7083_ );
xor  ( new_n7086_, new_n7085_, new_n7082_ );
xor  ( new_n7087_, new_n7086_, new_n7077_ );
xor  ( new_n7088_, RI2b1c4342d288_60, new_n191_ );
xor  ( new_n7089_, new_n7088_, new_n7087_ );
xor  ( new_n7090_, new_n7089_, new_n7072_ );
xor  ( new_n7091_, RI2b1c4342d468_64, new_n208_ );
xor  ( new_n7092_, RI2b1c4342cdd8_50, new_n150_ );
xor  ( new_n7093_, RI2b1c4342cfb8_54, RI2b1c4342cf40_53 );
xor  ( new_n7094_, new_n7093_, new_n7092_ );
xor  ( new_n7095_, new_n7094_, new_n7091_ );
xor  ( new_n7096_, new_n7095_, new_n7090_ );
xor  ( new_n7097_, new_n7096_, new_n7069_ );
xor  ( new_n7098_, new_n5855_, RI2b1c4342d468_64 );
nand ( new_n7099_, new_n7098_, new_n7097_ );
and  ( new_n7100_, new_n7099_, new_n5858_ );
and  ( new_n7101_, new_n5850_, new_n5849_ );
not  ( new_n7102_, new_n7101_ );
and  ( new_n7103_, new_n7102_, new_n338_ );
and  ( new_n7104_, new_n7103_, new_n7097_ );
or   ( new_n7105_, new_n7104_, new_n7100_ );
or   ( new_n7106_, new_n7105_, new_n99_ );
and  ( new_n7107_, new_n7106_, new_n5858_ );
and  ( new_n7108_, new_n7104_, new_n5858_ );
or   ( new_n7109_, new_n7108_, new_n6037_ );
and  ( new_n7110_, new_n7109_, new_n7099_ );
and  ( new_n7111_, new_n7110_, RI2b1c4342d4e0_65 );
and  ( new_n7112_, new_n7111_, new_n6037_ );
or   ( new_n7113_, new_n7112_, new_n7107_ );
or   ( new_n7114_, new_n6156_, new_n112_ );
or   ( new_n7115_, new_n6160_, new_n526_ );
and  ( new_n7116_, new_n7115_, new_n7114_ );
and  ( new_n7117_, new_n7116_, new_n6039_ );
and  ( new_n7118_, new_n6164_, RI2b1c4342d5d0_67 );
and  ( new_n7119_, new_n6154_, RI2b1c4342d558_66 );
or   ( new_n7120_, new_n7119_, new_n7118_ );
and  ( new_n7121_, new_n7120_, new_n5867_ );
or   ( new_n7122_, new_n7121_, new_n7117_ );
or   ( new_n7123_, new_n7122_, new_n7113_ );
or   ( new_n7124_, new_n5308_, new_n591_ );
or   ( new_n7125_, new_n5312_, new_n612_ );
and  ( new_n7126_, new_n7125_, new_n7124_ );
and  ( new_n7127_, new_n7126_, new_n5182_ );
and  ( new_n7128_, new_n5316_, RI2b1c4342d6c0_69 );
and  ( new_n7129_, new_n5306_, RI2b1c4342d648_68 );
or   ( new_n7130_, new_n7129_, new_n7128_ );
and  ( new_n7131_, new_n7130_, new_n5028_ );
or   ( new_n7132_, new_n7131_, new_n7127_ );
or   ( new_n7133_, new_n4535_, new_n110_ );
or   ( new_n7134_, new_n4539_, new_n755_ );
and  ( new_n7135_, new_n7134_, new_n7133_ );
and  ( new_n7136_, new_n7135_, new_n4400_ );
and  ( new_n7137_, new_n4543_, RI2b1c4342d7b0_71 );
and  ( new_n7138_, new_n4533_, RI2b1c4342d738_70 );
or   ( new_n7139_, new_n7138_, new_n7137_ );
and  ( new_n7140_, new_n7139_, new_n4215_ );
or   ( new_n7141_, new_n7140_, new_n7136_ );
and  ( new_n7142_, new_n7141_, new_n7132_ );
or   ( new_n7143_, new_n7141_, new_n7132_ );
or   ( new_n7144_, new_n3802_, new_n105_ );
or   ( new_n7145_, new_n3806_, new_n806_ );
and  ( new_n7146_, new_n7145_, new_n7144_ );
and  ( new_n7147_, new_n7146_, new_n3695_ );
and  ( new_n7148_, new_n3810_, RI2b1c4342d8a0_73 );
and  ( new_n7149_, new_n3800_, RI2b1c4342d828_72 );
or   ( new_n7150_, new_n7149_, new_n7148_ );
and  ( new_n7151_, new_n7150_, new_n3548_ );
or   ( new_n7152_, new_n7151_, new_n7147_ );
and  ( new_n7153_, new_n7152_, new_n7143_ );
or   ( new_n7154_, new_n7153_, new_n7142_ );
and  ( new_n7155_, new_n7154_, new_n7123_ );
or   ( new_n7156_, new_n7154_, new_n7123_ );
or   ( new_n7157_, new_n3112_, new_n843_ );
or   ( new_n7158_, new_n3116_, new_n859_ );
and  ( new_n7159_, new_n7158_, new_n7157_ );
and  ( new_n7160_, new_n7159_, new_n3004_ );
and  ( new_n7161_, new_n3120_, RI2b1c4342d990_75 );
and  ( new_n7162_, new_n3110_, RI2b1c4342d918_74 );
or   ( new_n7163_, new_n7162_, new_n7161_ );
and  ( new_n7164_, new_n7163_, new_n2868_ );
or   ( new_n7165_, new_n7164_, new_n7160_ );
or   ( new_n7166_, new_n2450_, new_n1004_ );
or   ( new_n7167_, new_n2454_, new_n886_ );
and  ( new_n7168_, new_n7167_, new_n7166_ );
and  ( new_n7169_, new_n7168_, new_n2334_ );
and  ( new_n7170_, new_n2458_, RI2b1c4342da80_77 );
and  ( new_n7171_, new_n2448_, RI2b1c4342da08_76 );
or   ( new_n7172_, new_n7171_, new_n7170_ );
and  ( new_n7173_, new_n7172_, new_n2168_ );
or   ( new_n7174_, new_n7173_, new_n7169_ );
and  ( new_n7175_, new_n7174_, new_n7165_ );
or   ( new_n7176_, new_n7174_, new_n7165_ );
or   ( new_n7177_, new_n1910_, new_n1310_ );
or   ( new_n7178_, new_n1914_, new_n1002_ );
and  ( new_n7179_, new_n7178_, new_n7177_ );
and  ( new_n7180_, new_n7179_, new_n1824_ );
and  ( new_n7181_, new_n1918_, RI2b1c4342db70_79 );
and  ( new_n7182_, new_n1908_, RI2b1c4342daf8_78 );
or   ( new_n7183_, new_n7182_, new_n7181_ );
and  ( new_n7184_, new_n7183_, new_n1717_ );
or   ( new_n7185_, new_n7184_, new_n7180_ );
and  ( new_n7186_, new_n7185_, new_n7176_ );
or   ( new_n7187_, new_n7186_, new_n7175_ );
and  ( new_n7188_, new_n7187_, new_n7156_ );
or   ( new_n7189_, new_n7188_, new_n7155_ );
or   ( new_n7190_, new_n1425_, new_n126_ );
or   ( new_n7191_, new_n1429_, new_n1511_ );
and  ( new_n7192_, new_n7191_, new_n7190_ );
and  ( new_n7193_, new_n7192_, new_n1355_ );
and  ( new_n7194_, new_n1433_, RI2b1c4342dc60_81 );
and  ( new_n7195_, new_n1423_, RI2b1c4342dbe8_80 );
or   ( new_n7196_, new_n7195_, new_n7194_ );
and  ( new_n7197_, new_n7196_, new_n1267_ );
or   ( new_n7198_, new_n7197_, new_n7193_ );
or   ( new_n7199_, new_n934_, new_n121_ );
or   ( new_n7200_, new_n940_, new_n2119_ );
and  ( new_n7201_, new_n7200_, new_n7199_ );
and  ( new_n7202_, new_n7201_, new_n913_ );
and  ( new_n7203_, new_n944_, RI2b1c4342dd50_83 );
and  ( new_n7204_, new_n932_, RI2b1c4342dcd8_82 );
or   ( new_n7205_, new_n7204_, new_n7203_ );
and  ( new_n7206_, new_n7205_, new_n938_ );
or   ( new_n7207_, new_n7206_, new_n7202_ );
and  ( new_n7208_, new_n7207_, new_n7198_ );
or   ( new_n7209_, new_n7207_, new_n7198_ );
or   ( new_n7210_, new_n453_, new_n2806_ );
or   ( new_n7211_, new_n459_, new_n2541_ );
and  ( new_n7212_, new_n7211_, new_n7210_ );
and  ( new_n7213_, new_n7212_, new_n428_ );
and  ( new_n7214_, new_n463_, RI2b1c4342de40_85 );
and  ( new_n7215_, new_n451_, RI2b1c4342ddc8_84 );
or   ( new_n7216_, new_n7215_, new_n7214_ );
and  ( new_n7217_, new_n7216_, new_n457_ );
or   ( new_n7218_, new_n7217_, new_n7213_ );
and  ( new_n7219_, new_n7218_, new_n7209_ );
or   ( new_n7220_, new_n7219_, new_n7208_ );
or   ( new_n7221_, new_n524_, new_n3924_ );
or   ( new_n7222_, new_n528_, new_n3239_ );
and  ( new_n7223_, new_n7222_, new_n7221_ );
and  ( new_n7224_, new_n7223_, new_n505_ );
and  ( new_n7225_, new_n537_, RI2b1c4342df30_87 );
and  ( new_n7226_, new_n522_, RI2b1c4342deb8_86 );
or   ( new_n7227_, new_n7226_, new_n7225_ );
and  ( new_n7228_, new_n7227_, new_n533_ );
or   ( new_n7229_, new_n7228_, new_n7224_ );
or   ( new_n7230_, new_n610_, new_n132_ );
or   ( new_n7231_, new_n614_, new_n3902_ );
and  ( new_n7232_, new_n7231_, new_n7230_ );
and  ( new_n7233_, new_n7232_, new_n590_ );
and  ( new_n7234_, new_n623_, RI2b1c4342e020_89 );
and  ( new_n7235_, new_n608_, RI2b1c4342dfa8_88 );
or   ( new_n7236_, new_n7235_, new_n7234_ );
and  ( new_n7237_, new_n7236_, new_n619_ );
or   ( new_n7238_, new_n7237_, new_n7233_ );
and  ( new_n7239_, new_n7238_, new_n7229_ );
or   ( new_n7240_, new_n7238_, new_n7229_ );
or   ( new_n7241_, new_n753_, new_n117_ );
or   ( new_n7242_, new_n757_, new_n4635_ );
and  ( new_n7243_, new_n7242_, new_n7241_ );
and  ( new_n7244_, new_n7243_, new_n734_ );
and  ( new_n7245_, new_n766_, RI2b1c4342e110_91 );
and  ( new_n7246_, new_n751_, RI2b1c4342e098_90 );
or   ( new_n7247_, new_n7246_, new_n7245_ );
and  ( new_n7248_, new_n7247_, new_n762_ );
or   ( new_n7249_, new_n7248_, new_n7244_ );
and  ( new_n7250_, new_n7249_, new_n7240_ );
or   ( new_n7251_, new_n7250_, new_n7239_ );
and  ( new_n7252_, new_n7251_, new_n7220_ );
or   ( new_n7253_, new_n7251_, new_n7220_ );
or   ( new_n7254_, new_n804_, new_n6307_ );
or   ( new_n7255_, new_n808_, new_n5459_ );
and  ( new_n7256_, new_n7255_, new_n7254_ );
and  ( new_n7257_, new_n7256_, new_n785_ );
and  ( new_n7258_, new_n817_, RI2b1c4342e200_93 );
and  ( new_n7259_, new_n802_, RI2b1c4342e188_92 );
or   ( new_n7260_, new_n7259_, new_n7258_ );
and  ( new_n7261_, new_n7260_, new_n813_ );
or   ( new_n7262_, new_n7261_, new_n7257_ );
or   ( new_n7263_, new_n857_, new_n124_ );
or   ( new_n7264_, new_n861_, new_n6321_ );
and  ( new_n7265_, new_n7264_, new_n7263_ );
and  ( new_n7266_, new_n7265_, new_n842_ );
and  ( new_n7267_, new_n870_, RI2b1c4342e2f0_95 );
and  ( new_n7268_, new_n855_, RI2b1c4342e278_94 );
or   ( new_n7269_, new_n7268_, new_n7267_ );
and  ( new_n7270_, new_n7269_, new_n866_ );
or   ( new_n7271_, new_n7270_, new_n7266_ );
and  ( new_n7272_, new_n7271_, new_n7262_ );
or   ( new_n7273_, new_n7271_, new_n7262_ );
not  ( new_n7274_, RI2b1c4342e368_96 );
or   ( new_n7275_, new_n841_, new_n7274_ );
and  ( new_n7276_, new_n7275_, new_n7273_ );
or   ( new_n7277_, new_n7276_, new_n7272_ );
and  ( new_n7278_, new_n7277_, new_n7253_ );
or   ( new_n7279_, new_n7278_, new_n7252_ );
and  ( new_n7280_, new_n7279_, new_n7189_ );
or   ( new_n7281_, new_n7279_, new_n7189_ );
and  ( new_n7282_, new_n6984_, new_n6704_ );
and  ( new_n7283_, new_n6985_, new_n6713_ );
or   ( new_n7284_, new_n7283_, new_n7282_ );
or   ( new_n7285_, new_n6973_, new_n6689_ );
and  ( new_n7286_, new_n7285_, new_n6699_ );
and  ( new_n7287_, new_n6969_, new_n6688_ );
and  ( new_n7288_, new_n6972_, new_n6679_ );
or   ( new_n7289_, new_n7288_, new_n7287_ );
and  ( new_n7290_, new_n7289_, new_n6977_ );
or   ( new_n7291_, new_n7290_, new_n7286_ );
and  ( new_n7292_, new_n7291_, new_n7284_ );
or   ( new_n7293_, new_n7291_, new_n7284_ );
or   ( new_n7294_, new_n6960_, new_n6658_ );
and  ( new_n7295_, new_n7294_, new_n6668_ );
and  ( new_n7296_, new_n6956_, new_n6657_ );
and  ( new_n7297_, new_n6959_, new_n6648_ );
or   ( new_n7298_, new_n7297_, new_n7296_ );
and  ( new_n7299_, new_n7298_, new_n6964_ );
or   ( new_n7300_, new_n7299_, new_n7295_ );
and  ( new_n7301_, new_n7300_, new_n7293_ );
or   ( new_n7302_, new_n7301_, new_n7292_ );
and  ( new_n7303_, new_n7302_, new_n7281_ );
or   ( new_n7304_, new_n7303_, new_n7280_ );
or   ( new_n7305_, new_n7012_, new_n6848_ );
and  ( new_n7306_, new_n7305_, new_n6856_ );
and  ( new_n7307_, new_n7008_, new_n6847_ );
and  ( new_n7308_, new_n7011_, new_n6840_ );
or   ( new_n7309_, new_n7308_, new_n7307_ );
and  ( new_n7310_, new_n7309_, new_n7016_ );
or   ( new_n7311_, new_n7310_, new_n7306_ );
or   ( new_n7312_, new_n6945_, new_n6790_ );
and  ( new_n7313_, new_n7312_, new_n6800_ );
and  ( new_n7314_, new_n6941_, new_n6789_ );
and  ( new_n7315_, new_n6944_, new_n6780_ );
or   ( new_n7316_, new_n7315_, new_n7314_ );
and  ( new_n7317_, new_n7316_, new_n6949_ );
or   ( new_n7318_, new_n7317_, new_n7313_ );
or   ( new_n7319_, new_n6930_, new_n6735_ );
and  ( new_n7320_, new_n7319_, new_n6745_ );
and  ( new_n7321_, new_n6926_, new_n6734_ );
and  ( new_n7322_, new_n6929_, new_n6725_ );
or   ( new_n7323_, new_n7322_, new_n7321_ );
and  ( new_n7324_, new_n7323_, new_n6934_ );
or   ( new_n7325_, new_n7324_, new_n7320_ );
and  ( new_n7326_, new_n7325_, new_n7318_ );
or   ( new_n7327_, new_n7325_, new_n7318_ );
or   ( new_n7328_, new_n6917_, new_n6757_ );
and  ( new_n7329_, new_n7328_, new_n6767_ );
and  ( new_n7330_, new_n6756_, new_n5858_ );
and  ( new_n7331_, new_n6916_, new_n6037_ );
or   ( new_n7332_, new_n7331_, new_n7330_ );
and  ( new_n7333_, new_n7332_, new_n6921_ );
or   ( new_n7334_, new_n7333_, new_n7329_ );
and  ( new_n7335_, new_n7334_, new_n7327_ );
or   ( new_n7336_, new_n7335_, new_n7326_ );
and  ( new_n7337_, new_n7336_, new_n7311_ );
or   ( new_n7338_, new_n7336_, new_n7311_ );
or   ( new_n7339_, new_n6994_, new_n6814_ );
and  ( new_n7340_, new_n7339_, new_n6822_ );
and  ( new_n7341_, new_n6813_, new_n6322_ );
and  ( new_n7342_, new_n6993_, new_n6579_ );
or   ( new_n7343_, new_n7342_, new_n7341_ );
and  ( new_n7344_, new_n7343_, new_n6998_ );
or   ( new_n7345_, new_n7344_, new_n7340_ );
and  ( new_n7346_, new_n7345_, new_n7338_ );
or   ( new_n7347_, new_n7346_, new_n7337_ );
and  ( new_n7348_, new_n7347_, new_n7304_ );
or   ( new_n7349_, new_n7347_, new_n7304_ );
or   ( new_n7350_, new_n6578_, new_n6319_ );
and  ( new_n7351_, new_n7350_, new_n6322_ );
and  ( new_n7352_, new_n6563_, new_n6318_ );
and  ( new_n7353_, new_n6576_, new_n6286_ );
or   ( new_n7354_, new_n7353_, new_n7352_ );
and  ( new_n7355_, new_n7354_, new_n6579_ );
or   ( new_n7356_, new_n7355_, new_n7351_ );
and  ( new_n7357_, new_n7356_, new_n7349_ );
or   ( new_n7358_, new_n7357_, new_n7348_ );
or   ( new_n7359_, new_n6534_, new_n6221_ );
and  ( new_n7360_, new_n7359_, new_n6253_ );
and  ( new_n7361_, new_n6520_, new_n6220_ );
and  ( new_n7362_, new_n6533_, new_n6189_ );
or   ( new_n7363_, new_n7362_, new_n7361_ );
and  ( new_n7364_, new_n7363_, new_n6548_ );
or   ( new_n7365_, new_n7364_, new_n7360_ );
or   ( new_n7366_, new_n7019_, new_n6859_ );
and  ( new_n7367_, new_n7366_, new_n6867_ );
and  ( new_n7368_, new_n7018_, new_n6833_ );
and  ( new_n7369_, new_n7005_, new_n6858_ );
or   ( new_n7370_, new_n7369_, new_n7368_ );
and  ( new_n7371_, new_n7370_, new_n7023_ );
or   ( new_n7372_, new_n7371_, new_n7367_ );
and  ( new_n7373_, new_n7372_, new_n7365_ );
or   ( new_n7374_, new_n7372_, new_n7365_ );
or   ( new_n7375_, new_n6989_, new_n6805_ );
and  ( new_n7376_, new_n7375_, new_n6824_ );
and  ( new_n7377_, new_n6953_, new_n6716_ );
and  ( new_n7378_, new_n6988_, new_n6804_ );
or   ( new_n7379_, new_n7378_, new_n7377_ );
and  ( new_n7380_, new_n7379_, new_n7000_ );
or   ( new_n7381_, new_n7380_, new_n7376_ );
and  ( new_n7382_, new_n7381_, new_n7374_ );
or   ( new_n7383_, new_n7382_, new_n7373_ );
and  ( new_n7384_, new_n7383_, new_n7358_ );
or   ( new_n7385_, new_n7383_, new_n7358_ );
or   ( new_n7386_, new_n6501_, new_n6380_ );
and  ( new_n7387_, new_n7386_, new_n6388_ );
and  ( new_n7388_, new_n6500_, new_n6354_ );
and  ( new_n7389_, new_n6487_, new_n6379_ );
or   ( new_n7390_, new_n7389_, new_n7388_ );
and  ( new_n7391_, new_n7390_, new_n6505_ );
or   ( new_n7392_, new_n7391_, new_n7387_ );
and  ( new_n7393_, new_n7392_, new_n7385_ );
or   ( new_n7394_, new_n7393_, new_n7384_ );
and  ( new_n7395_, new_n7394_, new_n7065_ );
or   ( new_n7396_, new_n7033_, new_n6881_ );
and  ( new_n7397_, new_n7396_, new_n6889_ );
and  ( new_n7398_, new_n7032_, new_n6639_ );
and  ( new_n7399_, new_n6913_, new_n6880_ );
or   ( new_n7400_, new_n7399_, new_n7398_ );
and  ( new_n7401_, new_n7400_, new_n7036_ );
or   ( new_n7402_, new_n7401_, new_n7397_ );
or   ( new_n7403_, new_n7394_, new_n7065_ );
and  ( new_n7404_, new_n7403_, new_n7402_ );
or   ( new_n7405_, new_n7404_, new_n7395_ );
and  ( new_n7406_, new_n7405_, new_n7050_ );
or   ( new_n7407_, new_n7405_, new_n7050_ );
and  ( new_n7408_, new_n7055_, new_n6345_ );
and  ( new_n7409_, new_n7051_, new_n6594_ );
or   ( new_n7410_, new_n7409_, new_n7408_ );
and  ( new_n7411_, new_n7062_, new_n6878_ );
and  ( new_n7412_, new_n7058_, new_n7029_ );
or   ( new_n7413_, new_n7412_, new_n7411_ );
and  ( new_n7414_, new_n7413_, new_n7410_ );
and  ( new_n7415_, new_n7363_, new_n6253_ );
and  ( new_n7416_, new_n7359_, new_n6548_ );
or   ( new_n7417_, new_n7416_, new_n7415_ );
and  ( new_n7418_, new_n7370_, new_n6867_ );
and  ( new_n7419_, new_n7366_, new_n7023_ );
or   ( new_n7420_, new_n7419_, new_n7418_ );
and  ( new_n7421_, new_n7420_, new_n7417_ );
or   ( new_n7422_, new_n7420_, new_n7417_ );
and  ( new_n7423_, new_n7379_, new_n6824_ );
and  ( new_n7424_, new_n7375_, new_n7000_ );
or   ( new_n7425_, new_n7424_, new_n7423_ );
and  ( new_n7426_, new_n7425_, new_n7422_ );
or   ( new_n7427_, new_n7426_, new_n7421_ );
and  ( new_n7428_, new_n7309_, new_n6856_ );
and  ( new_n7429_, new_n7305_, new_n7016_ );
or   ( new_n7430_, new_n7429_, new_n7428_ );
and  ( new_n7431_, new_n7316_, new_n6800_ );
and  ( new_n7432_, new_n7312_, new_n6949_ );
or   ( new_n7433_, new_n7432_, new_n7431_ );
and  ( new_n7434_, new_n7323_, new_n6745_ );
and  ( new_n7435_, new_n7319_, new_n6934_ );
or   ( new_n7436_, new_n7435_, new_n7434_ );
and  ( new_n7437_, new_n7436_, new_n7433_ );
or   ( new_n7438_, new_n7436_, new_n7433_ );
and  ( new_n7439_, new_n7332_, new_n6767_ );
and  ( new_n7440_, new_n7328_, new_n6921_ );
or   ( new_n7441_, new_n7440_, new_n7439_ );
and  ( new_n7442_, new_n7441_, new_n7438_ );
or   ( new_n7443_, new_n7442_, new_n7437_ );
and  ( new_n7444_, new_n7443_, new_n7430_ );
or   ( new_n7445_, new_n7443_, new_n7430_ );
and  ( new_n7446_, new_n7343_, new_n6822_ );
and  ( new_n7447_, new_n7339_, new_n6998_ );
or   ( new_n7448_, new_n7447_, new_n7446_ );
and  ( new_n7449_, new_n7448_, new_n7445_ );
or   ( new_n7450_, new_n7449_, new_n7444_ );
and  ( new_n7451_, new_n7111_, new_n5858_ );
and  ( new_n7452_, new_n7106_, new_n6037_ );
or   ( new_n7453_, new_n7452_, new_n7451_ );
and  ( new_n7454_, new_n7120_, new_n6039_ );
and  ( new_n7455_, new_n7116_, new_n5867_ );
or   ( new_n7456_, new_n7455_, new_n7454_ );
and  ( new_n7457_, new_n7456_, new_n7453_ );
and  ( new_n7458_, new_n7130_, new_n5182_ );
and  ( new_n7459_, new_n7126_, new_n5028_ );
or   ( new_n7460_, new_n7459_, new_n7458_ );
and  ( new_n7461_, new_n7139_, new_n4400_ );
and  ( new_n7462_, new_n7135_, new_n4215_ );
or   ( new_n7463_, new_n7462_, new_n7461_ );
and  ( new_n7464_, new_n7463_, new_n7460_ );
or   ( new_n7465_, new_n7463_, new_n7460_ );
and  ( new_n7466_, new_n7150_, new_n3695_ );
and  ( new_n7467_, new_n7146_, new_n3548_ );
or   ( new_n7468_, new_n7467_, new_n7466_ );
and  ( new_n7469_, new_n7468_, new_n7465_ );
or   ( new_n7470_, new_n7469_, new_n7464_ );
and  ( new_n7471_, new_n7470_, new_n7457_ );
or   ( new_n7472_, new_n7470_, new_n7457_ );
and  ( new_n7473_, new_n7163_, new_n3004_ );
and  ( new_n7474_, new_n7159_, new_n2868_ );
or   ( new_n7475_, new_n7474_, new_n7473_ );
and  ( new_n7476_, new_n7172_, new_n2334_ );
and  ( new_n7477_, new_n7168_, new_n2168_ );
or   ( new_n7478_, new_n7477_, new_n7476_ );
and  ( new_n7479_, new_n7478_, new_n7475_ );
or   ( new_n7480_, new_n7478_, new_n7475_ );
and  ( new_n7481_, new_n7183_, new_n1824_ );
and  ( new_n7482_, new_n7179_, new_n1717_ );
or   ( new_n7483_, new_n7482_, new_n7481_ );
and  ( new_n7484_, new_n7483_, new_n7480_ );
or   ( new_n7485_, new_n7484_, new_n7479_ );
and  ( new_n7486_, new_n7485_, new_n7472_ );
or   ( new_n7487_, new_n7486_, new_n7471_ );
and  ( new_n7488_, new_n7196_, new_n1355_ );
and  ( new_n7489_, new_n7192_, new_n1267_ );
or   ( new_n7490_, new_n7489_, new_n7488_ );
and  ( new_n7491_, new_n7205_, new_n913_ );
and  ( new_n7492_, new_n7201_, new_n938_ );
or   ( new_n7493_, new_n7492_, new_n7491_ );
and  ( new_n7494_, new_n7493_, new_n7490_ );
or   ( new_n7495_, new_n7493_, new_n7490_ );
and  ( new_n7496_, new_n7216_, new_n428_ );
and  ( new_n7497_, new_n7212_, new_n457_ );
or   ( new_n7498_, new_n7497_, new_n7496_ );
and  ( new_n7499_, new_n7498_, new_n7495_ );
or   ( new_n7500_, new_n7499_, new_n7494_ );
and  ( new_n7501_, new_n7227_, new_n505_ );
and  ( new_n7502_, new_n7223_, new_n533_ );
or   ( new_n7503_, new_n7502_, new_n7501_ );
and  ( new_n7504_, new_n7236_, new_n590_ );
and  ( new_n7505_, new_n7232_, new_n619_ );
or   ( new_n7506_, new_n7505_, new_n7504_ );
and  ( new_n7507_, new_n7506_, new_n7503_ );
or   ( new_n7508_, new_n7506_, new_n7503_ );
and  ( new_n7509_, new_n7247_, new_n734_ );
and  ( new_n7510_, new_n7243_, new_n762_ );
or   ( new_n7511_, new_n7510_, new_n7509_ );
and  ( new_n7512_, new_n7511_, new_n7508_ );
or   ( new_n7513_, new_n7512_, new_n7507_ );
or   ( new_n7514_, new_n7513_, new_n7500_ );
and  ( new_n7515_, new_n7513_, new_n7500_ );
and  ( new_n7516_, new_n7260_, new_n785_ );
and  ( new_n7517_, new_n7256_, new_n813_ );
or   ( new_n7518_, new_n7517_, new_n7516_ );
and  ( new_n7519_, new_n7269_, new_n842_ );
and  ( new_n7520_, new_n7265_, new_n866_ );
or   ( new_n7521_, new_n7520_, new_n7519_ );
or   ( new_n7522_, new_n7521_, new_n7518_ );
and  ( new_n7523_, new_n7521_, new_n7518_ );
and  ( new_n7524_, new_n720_, RI2b1c4342e368_96 );
or   ( new_n7525_, new_n7524_, new_n7523_ );
and  ( new_n7526_, new_n7525_, new_n7522_ );
or   ( new_n7527_, new_n7526_, new_n7515_ );
and  ( new_n7528_, new_n7527_, new_n7514_ );
or   ( new_n7529_, new_n7528_, new_n7487_ );
and  ( new_n7530_, new_n7528_, new_n7487_ );
and  ( new_n7531_, new_n6985_, new_n6984_ );
or   ( new_n7532_, new_n7531_, new_n6714_ );
and  ( new_n7533_, new_n7289_, new_n6699_ );
and  ( new_n7534_, new_n7285_, new_n6977_ );
or   ( new_n7535_, new_n7534_, new_n7533_ );
and  ( new_n7536_, new_n7535_, new_n7532_ );
or   ( new_n7537_, new_n7535_, new_n7532_ );
and  ( new_n7538_, new_n7298_, new_n6668_ );
and  ( new_n7539_, new_n7294_, new_n6964_ );
or   ( new_n7540_, new_n7539_, new_n7538_ );
and  ( new_n7541_, new_n7540_, new_n7537_ );
or   ( new_n7542_, new_n7541_, new_n7536_ );
or   ( new_n7543_, new_n7542_, new_n7530_ );
and  ( new_n7544_, new_n7543_, new_n7529_ );
or   ( new_n7545_, new_n7544_, new_n7450_ );
and  ( new_n7546_, new_n7544_, new_n7450_ );
and  ( new_n7547_, new_n7354_, new_n6322_ );
and  ( new_n7548_, new_n7350_, new_n6579_ );
or   ( new_n7549_, new_n7548_, new_n7547_ );
or   ( new_n7550_, new_n7549_, new_n7546_ );
and  ( new_n7551_, new_n7550_, new_n7545_ );
or   ( new_n7552_, new_n7551_, new_n7427_ );
and  ( new_n7553_, new_n7551_, new_n7427_ );
and  ( new_n7554_, new_n7390_, new_n6388_ );
and  ( new_n7555_, new_n7386_, new_n6505_ );
or   ( new_n7556_, new_n7555_, new_n7554_ );
or   ( new_n7557_, new_n7556_, new_n7553_ );
and  ( new_n7558_, new_n7557_, new_n7552_ );
and  ( new_n7559_, new_n7558_, new_n7414_ );
or   ( new_n7560_, new_n7559_, new_n7395_ );
and  ( new_n7561_, new_n7560_, new_n7402_ );
and  ( new_n7562_, new_n7558_, new_n7065_ );
and  ( new_n7563_, new_n7414_, new_n7394_ );
or   ( new_n7564_, new_n7563_, new_n7562_ );
and  ( new_n7565_, new_n7400_, new_n6889_ );
and  ( new_n7566_, new_n7396_, new_n7036_ );
or   ( new_n7567_, new_n7566_, new_n7565_ );
and  ( new_n7568_, new_n7567_, new_n7564_ );
or   ( new_n7569_, new_n7568_, new_n7561_ );
and  ( new_n7570_, new_n7064_, new_n7057_ );
or   ( new_n7571_, new_n7570_, new_n7414_ );
or   ( new_n7572_, new_n6937_, new_n6770_ );
and  ( new_n7573_, new_n7572_, new_n6802_ );
and  ( new_n7574_, new_n6923_, new_n6747_ );
and  ( new_n7575_, new_n6936_, new_n6769_ );
or   ( new_n7576_, new_n7575_, new_n7574_ );
and  ( new_n7577_, new_n7576_, new_n6951_ );
or   ( new_n7578_, new_n7577_, new_n7573_ );
or   ( new_n7579_, new_n7444_, new_n7337_ );
and  ( new_n7580_, new_n7579_, new_n7345_ );
and  ( new_n7581_, new_n7443_, new_n7311_ );
and  ( new_n7582_, new_n7430_, new_n7336_ );
or   ( new_n7583_, new_n7582_, new_n7581_ );
and  ( new_n7584_, new_n7583_, new_n7448_ );
or   ( new_n7585_, new_n7584_, new_n7580_ );
and  ( new_n7586_, new_n7585_, new_n7578_ );
or   ( new_n7587_, new_n7585_, new_n7578_ );
or   ( new_n7588_, new_n7530_, new_n7280_ );
and  ( new_n7589_, new_n7588_, new_n7302_ );
and  ( new_n7590_, new_n7487_, new_n7279_ );
and  ( new_n7591_, new_n7528_, new_n7189_ );
or   ( new_n7592_, new_n7591_, new_n7590_ );
and  ( new_n7593_, new_n7592_, new_n7542_ );
or   ( new_n7594_, new_n7593_, new_n7589_ );
and  ( new_n7595_, new_n7594_, new_n7587_ );
or   ( new_n7596_, new_n7595_, new_n7586_ );
or   ( new_n7597_, new_n7105_, new_n526_ );
or   ( new_n7598_, new_n7099_, new_n99_ );
and  ( new_n7599_, new_n7598_, new_n7597_ );
and  ( new_n7600_, new_n7599_, new_n5858_ );
and  ( new_n7601_, new_n7104_, RI2b1c4342d4e0_65 );
and  ( new_n7602_, new_n7110_, RI2b1c4342d558_66 );
or   ( new_n7603_, new_n7602_, new_n7601_ );
and  ( new_n7604_, new_n7603_, new_n6037_ );
or   ( new_n7605_, new_n7604_, new_n7600_ );
or   ( new_n7606_, new_n6156_, new_n612_ );
or   ( new_n7607_, new_n6160_, new_n112_ );
and  ( new_n7608_, new_n7607_, new_n7606_ );
and  ( new_n7609_, new_n7608_, new_n6039_ );
and  ( new_n7610_, new_n6164_, RI2b1c4342d648_68 );
and  ( new_n7611_, new_n6154_, RI2b1c4342d5d0_67 );
or   ( new_n7612_, new_n7611_, new_n7610_ );
and  ( new_n7613_, new_n7612_, new_n5867_ );
or   ( new_n7614_, new_n7613_, new_n7609_ );
and  ( new_n7615_, new_n7614_, new_n7605_ );
or   ( new_n7616_, new_n7614_, new_n7605_ );
or   ( new_n7617_, new_n5308_, new_n755_ );
or   ( new_n7618_, new_n5312_, new_n591_ );
and  ( new_n7619_, new_n7618_, new_n7617_ );
and  ( new_n7620_, new_n7619_, new_n5182_ );
and  ( new_n7621_, new_n5316_, RI2b1c4342d738_70 );
and  ( new_n7622_, new_n5306_, RI2b1c4342d6c0_69 );
or   ( new_n7623_, new_n7622_, new_n7621_ );
and  ( new_n7624_, new_n7623_, new_n5028_ );
or   ( new_n7625_, new_n7624_, new_n7620_ );
and  ( new_n7626_, new_n7625_, new_n7616_ );
or   ( new_n7627_, new_n7626_, new_n7615_ );
or   ( new_n7628_, new_n4535_, new_n806_ );
or   ( new_n7629_, new_n4539_, new_n110_ );
and  ( new_n7630_, new_n7629_, new_n7628_ );
and  ( new_n7631_, new_n7630_, new_n4400_ );
and  ( new_n7632_, new_n4543_, RI2b1c4342d828_72 );
and  ( new_n7633_, new_n4533_, RI2b1c4342d7b0_71 );
or   ( new_n7634_, new_n7633_, new_n7632_ );
and  ( new_n7635_, new_n7634_, new_n4215_ );
or   ( new_n7636_, new_n7635_, new_n7631_ );
or   ( new_n7637_, new_n3802_, new_n859_ );
or   ( new_n7638_, new_n3806_, new_n105_ );
and  ( new_n7639_, new_n7638_, new_n7637_ );
and  ( new_n7640_, new_n7639_, new_n3695_ );
and  ( new_n7641_, new_n3810_, RI2b1c4342d918_74 );
and  ( new_n7642_, new_n3800_, RI2b1c4342d8a0_73 );
or   ( new_n7643_, new_n7642_, new_n7641_ );
and  ( new_n7644_, new_n7643_, new_n3548_ );
or   ( new_n7645_, new_n7644_, new_n7640_ );
and  ( new_n7646_, new_n7645_, new_n7636_ );
or   ( new_n7647_, new_n7645_, new_n7636_ );
or   ( new_n7648_, new_n3112_, new_n886_ );
or   ( new_n7649_, new_n3116_, new_n843_ );
and  ( new_n7650_, new_n7649_, new_n7648_ );
and  ( new_n7651_, new_n7650_, new_n3004_ );
and  ( new_n7652_, new_n3120_, RI2b1c4342da08_76 );
and  ( new_n7653_, new_n3110_, RI2b1c4342d990_75 );
or   ( new_n7654_, new_n7653_, new_n7652_ );
and  ( new_n7655_, new_n7654_, new_n2868_ );
or   ( new_n7656_, new_n7655_, new_n7651_ );
and  ( new_n7657_, new_n7656_, new_n7647_ );
or   ( new_n7658_, new_n7657_, new_n7646_ );
and  ( new_n7659_, new_n7658_, new_n7627_ );
or   ( new_n7660_, new_n7658_, new_n7627_ );
or   ( new_n7661_, new_n2450_, new_n1002_ );
or   ( new_n7662_, new_n2454_, new_n1004_ );
and  ( new_n7663_, new_n7662_, new_n7661_ );
and  ( new_n7664_, new_n7663_, new_n2334_ );
and  ( new_n7665_, new_n2458_, RI2b1c4342daf8_78 );
and  ( new_n7666_, new_n2448_, RI2b1c4342da80_77 );
or   ( new_n7667_, new_n7666_, new_n7665_ );
and  ( new_n7668_, new_n7667_, new_n2168_ );
or   ( new_n7669_, new_n7668_, new_n7664_ );
or   ( new_n7670_, new_n1910_, new_n1511_ );
or   ( new_n7671_, new_n1914_, new_n1310_ );
and  ( new_n7672_, new_n7671_, new_n7670_ );
and  ( new_n7673_, new_n7672_, new_n1824_ );
and  ( new_n7674_, new_n1918_, RI2b1c4342dbe8_80 );
and  ( new_n7675_, new_n1908_, RI2b1c4342db70_79 );
or   ( new_n7676_, new_n7675_, new_n7674_ );
and  ( new_n7677_, new_n7676_, new_n1717_ );
or   ( new_n7678_, new_n7677_, new_n7673_ );
and  ( new_n7679_, new_n7678_, new_n7669_ );
or   ( new_n7680_, new_n7678_, new_n7669_ );
or   ( new_n7681_, new_n1425_, new_n2119_ );
or   ( new_n7682_, new_n1429_, new_n126_ );
and  ( new_n7683_, new_n7682_, new_n7681_ );
and  ( new_n7684_, new_n7683_, new_n1355_ );
and  ( new_n7685_, new_n1433_, RI2b1c4342dcd8_82 );
and  ( new_n7686_, new_n1423_, RI2b1c4342dc60_81 );
or   ( new_n7687_, new_n7686_, new_n7685_ );
and  ( new_n7688_, new_n7687_, new_n1267_ );
or   ( new_n7689_, new_n7688_, new_n7684_ );
and  ( new_n7690_, new_n7689_, new_n7680_ );
or   ( new_n7691_, new_n7690_, new_n7679_ );
and  ( new_n7692_, new_n7691_, new_n7660_ );
or   ( new_n7693_, new_n7692_, new_n7659_ );
or   ( new_n7694_, new_n934_, new_n2541_ );
or   ( new_n7695_, new_n940_, new_n121_ );
and  ( new_n7696_, new_n7695_, new_n7694_ );
and  ( new_n7697_, new_n7696_, new_n913_ );
and  ( new_n7698_, new_n944_, RI2b1c4342ddc8_84 );
and  ( new_n7699_, new_n932_, RI2b1c4342dd50_83 );
or   ( new_n7700_, new_n7699_, new_n7698_ );
and  ( new_n7701_, new_n7700_, new_n938_ );
or   ( new_n7702_, new_n7701_, new_n7697_ );
or   ( new_n7703_, new_n453_, new_n3239_ );
or   ( new_n7704_, new_n459_, new_n2806_ );
and  ( new_n7705_, new_n7704_, new_n7703_ );
and  ( new_n7706_, new_n7705_, new_n428_ );
and  ( new_n7707_, new_n463_, RI2b1c4342deb8_86 );
and  ( new_n7708_, new_n451_, RI2b1c4342de40_85 );
or   ( new_n7709_, new_n7708_, new_n7707_ );
and  ( new_n7710_, new_n7709_, new_n457_ );
or   ( new_n7711_, new_n7710_, new_n7706_ );
and  ( new_n7712_, new_n7711_, new_n7702_ );
or   ( new_n7713_, new_n7711_, new_n7702_ );
or   ( new_n7714_, new_n524_, new_n3902_ );
or   ( new_n7715_, new_n528_, new_n3924_ );
and  ( new_n7716_, new_n7715_, new_n7714_ );
and  ( new_n7717_, new_n7716_, new_n505_ );
and  ( new_n7718_, new_n537_, RI2b1c4342dfa8_88 );
and  ( new_n7719_, new_n522_, RI2b1c4342df30_87 );
or   ( new_n7720_, new_n7719_, new_n7718_ );
and  ( new_n7721_, new_n7720_, new_n533_ );
or   ( new_n7722_, new_n7721_, new_n7717_ );
and  ( new_n7723_, new_n7722_, new_n7713_ );
or   ( new_n7724_, new_n7723_, new_n7712_ );
or   ( new_n7725_, new_n610_, new_n4635_ );
or   ( new_n7726_, new_n614_, new_n132_ );
and  ( new_n7727_, new_n7726_, new_n7725_ );
and  ( new_n7728_, new_n7727_, new_n590_ );
and  ( new_n7729_, new_n623_, RI2b1c4342e098_90 );
and  ( new_n7730_, new_n608_, RI2b1c4342e020_89 );
or   ( new_n7731_, new_n7730_, new_n7729_ );
and  ( new_n7732_, new_n7731_, new_n619_ );
or   ( new_n7733_, new_n7732_, new_n7728_ );
or   ( new_n7734_, new_n753_, new_n5459_ );
or   ( new_n7735_, new_n757_, new_n117_ );
and  ( new_n7736_, new_n7735_, new_n7734_ );
and  ( new_n7737_, new_n7736_, new_n734_ );
and  ( new_n7738_, new_n766_, RI2b1c4342e188_92 );
and  ( new_n7739_, new_n751_, RI2b1c4342e110_91 );
or   ( new_n7740_, new_n7739_, new_n7738_ );
and  ( new_n7741_, new_n7740_, new_n762_ );
or   ( new_n7742_, new_n7741_, new_n7737_ );
and  ( new_n7743_, new_n7742_, new_n7733_ );
or   ( new_n7744_, new_n7742_, new_n7733_ );
or   ( new_n7745_, new_n804_, new_n6321_ );
or   ( new_n7746_, new_n808_, new_n6307_ );
and  ( new_n7747_, new_n7746_, new_n7745_ );
and  ( new_n7748_, new_n7747_, new_n785_ );
and  ( new_n7749_, new_n817_, RI2b1c4342e278_94 );
and  ( new_n7750_, new_n802_, RI2b1c4342e200_93 );
or   ( new_n7751_, new_n7750_, new_n7749_ );
and  ( new_n7752_, new_n7751_, new_n813_ );
or   ( new_n7753_, new_n7752_, new_n7748_ );
and  ( new_n7754_, new_n7753_, new_n7744_ );
or   ( new_n7755_, new_n7754_, new_n7743_ );
and  ( new_n7756_, new_n7755_, new_n7724_ );
or   ( new_n7757_, new_n7755_, new_n7724_ );
or   ( new_n7758_, new_n7523_, new_n7272_ );
and  ( new_n7759_, new_n7758_, new_n7275_ );
and  ( new_n7760_, new_n7518_, new_n7271_ );
and  ( new_n7761_, new_n7521_, new_n7262_ );
or   ( new_n7762_, new_n7761_, new_n7760_ );
and  ( new_n7763_, new_n7762_, new_n7524_ );
or   ( new_n7764_, new_n7763_, new_n7759_ );
and  ( new_n7765_, new_n7764_, new_n7757_ );
or   ( new_n7766_, new_n7765_, new_n7756_ );
and  ( new_n7767_, new_n7766_, new_n7693_ );
or   ( new_n7768_, new_n7766_, new_n7693_ );
or   ( new_n7769_, new_n7507_, new_n7239_ );
and  ( new_n7770_, new_n7769_, new_n7249_ );
and  ( new_n7771_, new_n7503_, new_n7238_ );
and  ( new_n7772_, new_n7506_, new_n7229_ );
or   ( new_n7773_, new_n7772_, new_n7771_ );
and  ( new_n7774_, new_n7773_, new_n7511_ );
or   ( new_n7775_, new_n7774_, new_n7770_ );
or   ( new_n7776_, new_n7494_, new_n7208_ );
and  ( new_n7777_, new_n7776_, new_n7218_ );
and  ( new_n7778_, new_n7490_, new_n7207_ );
and  ( new_n7779_, new_n7493_, new_n7198_ );
or   ( new_n7780_, new_n7779_, new_n7778_ );
and  ( new_n7781_, new_n7780_, new_n7498_ );
or   ( new_n7782_, new_n7781_, new_n7777_ );
and  ( new_n7783_, new_n7782_, new_n7775_ );
or   ( new_n7784_, new_n7782_, new_n7775_ );
or   ( new_n7785_, new_n7479_, new_n7175_ );
and  ( new_n7786_, new_n7785_, new_n7185_ );
and  ( new_n7787_, new_n7475_, new_n7174_ );
and  ( new_n7788_, new_n7478_, new_n7165_ );
or   ( new_n7789_, new_n7788_, new_n7787_ );
and  ( new_n7790_, new_n7789_, new_n7483_ );
or   ( new_n7791_, new_n7790_, new_n7786_ );
and  ( new_n7792_, new_n7791_, new_n7784_ );
or   ( new_n7793_, new_n7792_, new_n7783_ );
and  ( new_n7794_, new_n7793_, new_n7768_ );
or   ( new_n7795_, new_n7794_, new_n7767_ );
or   ( new_n7796_, new_n7437_, new_n7326_ );
and  ( new_n7797_, new_n7796_, new_n7334_ );
and  ( new_n7798_, new_n7433_, new_n7325_ );
and  ( new_n7799_, new_n7436_, new_n7318_ );
or   ( new_n7800_, new_n7799_, new_n7798_ );
and  ( new_n7801_, new_n7800_, new_n7441_ );
or   ( new_n7802_, new_n7801_, new_n7797_ );
or   ( new_n7803_, new_n7536_, new_n7292_ );
and  ( new_n7804_, new_n7803_, new_n7300_ );
and  ( new_n7805_, new_n7532_, new_n7291_ );
and  ( new_n7806_, new_n7535_, new_n7284_ );
or   ( new_n7807_, new_n7806_, new_n7805_ );
and  ( new_n7808_, new_n7807_, new_n7540_ );
or   ( new_n7809_, new_n7808_, new_n7804_ );
and  ( new_n7810_, new_n7809_, new_n7802_ );
or   ( new_n7811_, new_n7809_, new_n7802_ );
or   ( new_n7812_, new_n7515_, new_n7252_ );
and  ( new_n7813_, new_n7812_, new_n7277_ );
and  ( new_n7814_, new_n7500_, new_n7251_ );
and  ( new_n7815_, new_n7513_, new_n7220_ );
or   ( new_n7816_, new_n7815_, new_n7814_ );
and  ( new_n7817_, new_n7816_, new_n7526_ );
or   ( new_n7818_, new_n7817_, new_n7813_ );
and  ( new_n7819_, new_n7818_, new_n7811_ );
or   ( new_n7820_, new_n7819_, new_n7810_ );
and  ( new_n7821_, new_n7820_, new_n7795_ );
or   ( new_n7822_, new_n7820_, new_n7795_ );
or   ( new_n7823_, new_n6980_, new_n6702_ );
and  ( new_n7824_, new_n7823_, new_n6714_ );
and  ( new_n7825_, new_n6966_, new_n6701_ );
and  ( new_n7826_, new_n6979_, new_n6670_ );
or   ( new_n7827_, new_n7826_, new_n7825_ );
and  ( new_n7828_, new_n7827_, new_n6986_ );
or   ( new_n7829_, new_n7828_, new_n7824_ );
and  ( new_n7830_, new_n7829_, new_n7822_ );
or   ( new_n7831_, new_n7830_, new_n7821_ );
and  ( new_n7832_, new_n7831_, new_n7596_ );
or   ( new_n7833_, new_n7831_, new_n7596_ );
or   ( new_n7834_, new_n7421_, new_n7373_ );
and  ( new_n7835_, new_n7834_, new_n7381_ );
and  ( new_n7836_, new_n7417_, new_n7372_ );
and  ( new_n7837_, new_n7420_, new_n7365_ );
or   ( new_n7838_, new_n7837_, new_n7836_ );
and  ( new_n7839_, new_n7838_, new_n7425_ );
or   ( new_n7840_, new_n7839_, new_n7835_ );
and  ( new_n7841_, new_n7840_, new_n7833_ );
or   ( new_n7842_, new_n7841_, new_n7832_ );
and  ( new_n7843_, new_n7842_, new_n7571_ );
or   ( new_n7844_, new_n7842_, new_n7571_ );
or   ( new_n7845_, new_n7553_, new_n7384_ );
and  ( new_n7846_, new_n7845_, new_n7392_ );
and  ( new_n7847_, new_n7551_, new_n7383_ );
and  ( new_n7848_, new_n7427_, new_n7358_ );
or   ( new_n7849_, new_n7848_, new_n7847_ );
and  ( new_n7850_, new_n7849_, new_n7556_ );
or   ( new_n7851_, new_n7850_, new_n7846_ );
and  ( new_n7852_, new_n7851_, new_n7844_ );
or   ( new_n7853_, new_n7852_, new_n7843_ );
or   ( new_n7854_, new_n7853_, new_n7569_ );
and  ( new_n7855_, new_n7854_, new_n7407_ );
or   ( new_n7856_, new_n7855_, new_n7406_ );
or   ( new_n7857_, new_n7856_, new_n6907_ );
and  ( new_n7858_, new_n7857_, new_n6905_ );
or   ( new_n7859_, new_n7858_, new_n5994_ );
and  ( new_n7860_, new_n7859_, new_n5991_ );
and  ( new_n7861_, new_n7410_, new_n7064_ );
and  ( new_n7862_, new_n7413_, new_n7057_ );
or   ( new_n7863_, new_n7862_, new_n7861_ );
and  ( new_n7864_, new_n7603_, new_n5858_ );
and  ( new_n7865_, new_n7599_, new_n6037_ );
or   ( new_n7866_, new_n7865_, new_n7864_ );
and  ( new_n7867_, new_n7612_, new_n6039_ );
and  ( new_n7868_, new_n7608_, new_n5867_ );
or   ( new_n7869_, new_n7868_, new_n7867_ );
and  ( new_n7870_, new_n7869_, new_n7866_ );
or   ( new_n7871_, new_n7869_, new_n7866_ );
and  ( new_n7872_, new_n7623_, new_n5182_ );
and  ( new_n7873_, new_n7619_, new_n5028_ );
or   ( new_n7874_, new_n7873_, new_n7872_ );
and  ( new_n7875_, new_n7874_, new_n7871_ );
or   ( new_n7876_, new_n7875_, new_n7870_ );
and  ( new_n7877_, new_n7634_, new_n4400_ );
and  ( new_n7878_, new_n7630_, new_n4215_ );
or   ( new_n7879_, new_n7878_, new_n7877_ );
and  ( new_n7880_, new_n7643_, new_n3695_ );
and  ( new_n7881_, new_n7639_, new_n3548_ );
or   ( new_n7882_, new_n7881_, new_n7880_ );
and  ( new_n7883_, new_n7882_, new_n7879_ );
or   ( new_n7884_, new_n7882_, new_n7879_ );
and  ( new_n7885_, new_n7654_, new_n3004_ );
and  ( new_n7886_, new_n7650_, new_n2868_ );
or   ( new_n7887_, new_n7886_, new_n7885_ );
and  ( new_n7888_, new_n7887_, new_n7884_ );
or   ( new_n7889_, new_n7888_, new_n7883_ );
and  ( new_n7890_, new_n7889_, new_n7876_ );
or   ( new_n7891_, new_n7889_, new_n7876_ );
and  ( new_n7892_, new_n7667_, new_n2334_ );
and  ( new_n7893_, new_n7663_, new_n2168_ );
or   ( new_n7894_, new_n7893_, new_n7892_ );
and  ( new_n7895_, new_n7676_, new_n1824_ );
and  ( new_n7896_, new_n7672_, new_n1717_ );
or   ( new_n7897_, new_n7896_, new_n7895_ );
and  ( new_n7898_, new_n7897_, new_n7894_ );
or   ( new_n7899_, new_n7897_, new_n7894_ );
and  ( new_n7900_, new_n7687_, new_n1355_ );
and  ( new_n7901_, new_n7683_, new_n1267_ );
or   ( new_n7902_, new_n7901_, new_n7900_ );
and  ( new_n7903_, new_n7902_, new_n7899_ );
or   ( new_n7904_, new_n7903_, new_n7898_ );
and  ( new_n7905_, new_n7904_, new_n7891_ );
or   ( new_n7906_, new_n7905_, new_n7890_ );
and  ( new_n7907_, new_n7700_, new_n913_ );
and  ( new_n7908_, new_n7696_, new_n938_ );
or   ( new_n7909_, new_n7908_, new_n7907_ );
and  ( new_n7910_, new_n7709_, new_n428_ );
and  ( new_n7911_, new_n7705_, new_n457_ );
or   ( new_n7912_, new_n7911_, new_n7910_ );
and  ( new_n7913_, new_n7912_, new_n7909_ );
or   ( new_n7914_, new_n7912_, new_n7909_ );
and  ( new_n7915_, new_n7720_, new_n505_ );
and  ( new_n7916_, new_n7716_, new_n533_ );
or   ( new_n7917_, new_n7916_, new_n7915_ );
and  ( new_n7918_, new_n7917_, new_n7914_ );
or   ( new_n7919_, new_n7918_, new_n7913_ );
and  ( new_n7920_, new_n7731_, new_n590_ );
and  ( new_n7921_, new_n7727_, new_n619_ );
or   ( new_n7922_, new_n7921_, new_n7920_ );
and  ( new_n7923_, new_n7740_, new_n734_ );
and  ( new_n7924_, new_n7736_, new_n762_ );
or   ( new_n7925_, new_n7924_, new_n7923_ );
and  ( new_n7926_, new_n7925_, new_n7922_ );
or   ( new_n7927_, new_n7925_, new_n7922_ );
and  ( new_n7928_, new_n7751_, new_n785_ );
and  ( new_n7929_, new_n7747_, new_n813_ );
or   ( new_n7930_, new_n7929_, new_n7928_ );
and  ( new_n7931_, new_n7930_, new_n7927_ );
or   ( new_n7932_, new_n7931_, new_n7926_ );
and  ( new_n7933_, new_n7932_, new_n7919_ );
or   ( new_n7934_, new_n7932_, new_n7919_ );
and  ( new_n7935_, new_n7762_, new_n7275_ );
and  ( new_n7936_, new_n7758_, new_n7524_ );
or   ( new_n7937_, new_n7936_, new_n7935_ );
and  ( new_n7938_, new_n7937_, new_n7934_ );
or   ( new_n7939_, new_n7938_, new_n7933_ );
and  ( new_n7940_, new_n7939_, new_n7906_ );
or   ( new_n7941_, new_n7939_, new_n7906_ );
and  ( new_n7942_, new_n7773_, new_n7249_ );
and  ( new_n7943_, new_n7769_, new_n7511_ );
or   ( new_n7944_, new_n7943_, new_n7942_ );
and  ( new_n7945_, new_n7780_, new_n7218_ );
and  ( new_n7946_, new_n7776_, new_n7498_ );
or   ( new_n7947_, new_n7946_, new_n7945_ );
and  ( new_n7948_, new_n7947_, new_n7944_ );
or   ( new_n7949_, new_n7947_, new_n7944_ );
and  ( new_n7950_, new_n7789_, new_n7185_ );
and  ( new_n7951_, new_n7785_, new_n7483_ );
or   ( new_n7952_, new_n7951_, new_n7950_ );
and  ( new_n7953_, new_n7952_, new_n7949_ );
or   ( new_n7954_, new_n7953_, new_n7948_ );
and  ( new_n7955_, new_n7954_, new_n7941_ );
or   ( new_n7956_, new_n7955_, new_n7940_ );
and  ( new_n7957_, new_n7800_, new_n7334_ );
and  ( new_n7958_, new_n7796_, new_n7441_ );
or   ( new_n7959_, new_n7958_, new_n7957_ );
and  ( new_n7960_, new_n7807_, new_n7300_ );
and  ( new_n7961_, new_n7803_, new_n7540_ );
or   ( new_n7962_, new_n7961_, new_n7960_ );
and  ( new_n7963_, new_n7962_, new_n7959_ );
or   ( new_n7964_, new_n7962_, new_n7959_ );
and  ( new_n7965_, new_n7816_, new_n7277_ );
and  ( new_n7966_, new_n7812_, new_n7526_ );
or   ( new_n7967_, new_n7966_, new_n7965_ );
and  ( new_n7968_, new_n7967_, new_n7964_ );
or   ( new_n7969_, new_n7968_, new_n7963_ );
and  ( new_n7970_, new_n7969_, new_n7956_ );
or   ( new_n7971_, new_n7969_, new_n7956_ );
and  ( new_n7972_, new_n7827_, new_n6714_ );
and  ( new_n7973_, new_n7823_, new_n6986_ );
or   ( new_n7974_, new_n7973_, new_n7972_ );
and  ( new_n7975_, new_n7974_, new_n7971_ );
or   ( new_n7976_, new_n7975_, new_n7970_ );
and  ( new_n7977_, new_n7576_, new_n6802_ );
and  ( new_n7978_, new_n7572_, new_n6951_ );
or   ( new_n7979_, new_n7978_, new_n7977_ );
and  ( new_n7980_, new_n7583_, new_n7345_ );
and  ( new_n7981_, new_n7579_, new_n7448_ );
or   ( new_n7982_, new_n7981_, new_n7980_ );
and  ( new_n7983_, new_n7982_, new_n7979_ );
or   ( new_n7984_, new_n7982_, new_n7979_ );
and  ( new_n7985_, new_n7592_, new_n7302_ );
and  ( new_n7986_, new_n7588_, new_n7542_ );
or   ( new_n7987_, new_n7986_, new_n7985_ );
and  ( new_n7988_, new_n7987_, new_n7984_ );
or   ( new_n7989_, new_n7988_, new_n7983_ );
and  ( new_n7990_, new_n7989_, new_n7976_ );
or   ( new_n7991_, new_n7989_, new_n7976_ );
and  ( new_n7992_, new_n7838_, new_n7381_ );
and  ( new_n7993_, new_n7834_, new_n7425_ );
or   ( new_n7994_, new_n7993_, new_n7992_ );
and  ( new_n7995_, new_n7994_, new_n7991_ );
or   ( new_n7996_, new_n7995_, new_n7990_ );
and  ( new_n7997_, new_n7996_, new_n7863_ );
or   ( new_n7998_, new_n7997_, new_n7843_ );
and  ( new_n7999_, new_n7998_, new_n7851_ );
and  ( new_n8000_, new_n7996_, new_n7571_ );
and  ( new_n8001_, new_n7863_, new_n7842_ );
or   ( new_n8002_, new_n8001_, new_n8000_ );
and  ( new_n8003_, new_n7849_, new_n7392_ );
and  ( new_n8004_, new_n7845_, new_n7556_ );
or   ( new_n8005_, new_n8004_, new_n8003_ );
and  ( new_n8006_, new_n8005_, new_n8002_ );
or   ( new_n8007_, new_n8006_, new_n7999_ );
or   ( new_n8008_, new_n7546_, new_n7348_ );
and  ( new_n8009_, new_n8008_, new_n7356_ );
and  ( new_n8010_, new_n7544_, new_n7347_ );
and  ( new_n8011_, new_n7450_, new_n7304_ );
or   ( new_n8012_, new_n8011_, new_n8010_ );
and  ( new_n8013_, new_n8012_, new_n7549_ );
or   ( new_n8014_, new_n8013_, new_n8009_ );
or   ( new_n8015_, new_n7471_, new_n7155_ );
and  ( new_n8016_, new_n8015_, new_n7187_ );
and  ( new_n8017_, new_n7457_, new_n7154_ );
and  ( new_n8018_, new_n7470_, new_n7123_ );
or   ( new_n8019_, new_n8018_, new_n8017_ );
and  ( new_n8020_, new_n8019_, new_n7485_ );
or   ( new_n8021_, new_n8020_, new_n8016_ );
or   ( new_n8022_, new_n7963_, new_n7810_ );
and  ( new_n8023_, new_n8022_, new_n7818_ );
and  ( new_n8024_, new_n7959_, new_n7809_ );
and  ( new_n8025_, new_n7962_, new_n7802_ );
or   ( new_n8026_, new_n8025_, new_n8024_ );
and  ( new_n8027_, new_n8026_, new_n7967_ );
or   ( new_n8028_, new_n8027_, new_n8023_ );
and  ( new_n8029_, new_n8028_, new_n8021_ );
or   ( new_n8030_, new_n8028_, new_n8021_ );
or   ( new_n8031_, new_n7940_, new_n7767_ );
and  ( new_n8032_, new_n8031_, new_n7793_ );
and  ( new_n8033_, new_n7906_, new_n7766_ );
and  ( new_n8034_, new_n7939_, new_n7693_ );
or   ( new_n8035_, new_n8034_, new_n8033_ );
and  ( new_n8036_, new_n8035_, new_n7954_ );
or   ( new_n8037_, new_n8036_, new_n8032_ );
and  ( new_n8038_, new_n8037_, new_n8030_ );
or   ( new_n8039_, new_n8038_, new_n8029_ );
or   ( new_n8040_, new_n7464_, new_n7142_ );
and  ( new_n8041_, new_n8040_, new_n7152_ );
and  ( new_n8042_, new_n7460_, new_n7141_ );
and  ( new_n8043_, new_n7463_, new_n7132_ );
or   ( new_n8044_, new_n8043_, new_n8042_ );
and  ( new_n8045_, new_n8044_, new_n7468_ );
or   ( new_n8046_, new_n8045_, new_n8041_ );
and  ( new_n8047_, new_n7122_, new_n7113_ );
or   ( new_n8048_, new_n8047_, new_n7457_ );
and  ( new_n8049_, new_n8048_, new_n8046_ );
or   ( new_n8050_, new_n8048_, new_n8046_ );
or   ( new_n8051_, new_n7948_, new_n7783_ );
and  ( new_n8052_, new_n8051_, new_n7791_ );
and  ( new_n8053_, new_n7944_, new_n7782_ );
and  ( new_n8054_, new_n7947_, new_n7775_ );
or   ( new_n8055_, new_n8054_, new_n8053_ );
and  ( new_n8056_, new_n8055_, new_n7952_ );
or   ( new_n8057_, new_n8056_, new_n8052_ );
and  ( new_n8058_, new_n8057_, new_n8050_ );
or   ( new_n8059_, new_n8058_, new_n8049_ );
or   ( new_n8060_, new_n1425_, new_n121_ );
or   ( new_n8061_, new_n1429_, new_n2119_ );
and  ( new_n8062_, new_n8061_, new_n8060_ );
and  ( new_n8063_, new_n8062_, new_n1355_ );
and  ( new_n8064_, new_n1433_, RI2b1c4342dd50_83 );
and  ( new_n8065_, new_n1423_, RI2b1c4342dcd8_82 );
or   ( new_n8066_, new_n8065_, new_n8064_ );
and  ( new_n8067_, new_n8066_, new_n1267_ );
or   ( new_n8068_, new_n8067_, new_n8063_ );
or   ( new_n8069_, new_n934_, new_n2806_ );
or   ( new_n8070_, new_n940_, new_n2541_ );
and  ( new_n8071_, new_n8070_, new_n8069_ );
and  ( new_n8072_, new_n8071_, new_n913_ );
and  ( new_n8073_, new_n944_, RI2b1c4342de40_85 );
and  ( new_n8074_, new_n932_, RI2b1c4342ddc8_84 );
or   ( new_n8075_, new_n8074_, new_n8073_ );
and  ( new_n8076_, new_n8075_, new_n938_ );
or   ( new_n8077_, new_n8076_, new_n8072_ );
and  ( new_n8078_, new_n8077_, new_n8068_ );
or   ( new_n8079_, new_n8077_, new_n8068_ );
or   ( new_n8080_, new_n453_, new_n3924_ );
or   ( new_n8081_, new_n459_, new_n3239_ );
and  ( new_n8082_, new_n8081_, new_n8080_ );
and  ( new_n8083_, new_n8082_, new_n428_ );
and  ( new_n8084_, new_n463_, RI2b1c4342df30_87 );
and  ( new_n8085_, new_n451_, RI2b1c4342deb8_86 );
or   ( new_n8086_, new_n8085_, new_n8084_ );
and  ( new_n8087_, new_n8086_, new_n457_ );
or   ( new_n8088_, new_n8087_, new_n8083_ );
and  ( new_n8089_, new_n8088_, new_n8079_ );
or   ( new_n8090_, new_n8089_, new_n8078_ );
or   ( new_n8091_, new_n524_, new_n132_ );
or   ( new_n8092_, new_n528_, new_n3902_ );
and  ( new_n8093_, new_n8092_, new_n8091_ );
and  ( new_n8094_, new_n8093_, new_n505_ );
and  ( new_n8095_, new_n537_, RI2b1c4342e020_89 );
and  ( new_n8096_, new_n522_, RI2b1c4342dfa8_88 );
or   ( new_n8097_, new_n8096_, new_n8095_ );
and  ( new_n8098_, new_n8097_, new_n533_ );
or   ( new_n8099_, new_n8098_, new_n8094_ );
or   ( new_n8100_, new_n610_, new_n117_ );
or   ( new_n8101_, new_n614_, new_n4635_ );
and  ( new_n8102_, new_n8101_, new_n8100_ );
and  ( new_n8103_, new_n8102_, new_n590_ );
and  ( new_n8104_, new_n623_, RI2b1c4342e110_91 );
and  ( new_n8105_, new_n608_, RI2b1c4342e098_90 );
or   ( new_n8106_, new_n8105_, new_n8104_ );
and  ( new_n8107_, new_n8106_, new_n619_ );
or   ( new_n8108_, new_n8107_, new_n8103_ );
and  ( new_n8109_, new_n8108_, new_n8099_ );
or   ( new_n8110_, new_n8108_, new_n8099_ );
or   ( new_n8111_, new_n753_, new_n6307_ );
or   ( new_n8112_, new_n757_, new_n5459_ );
and  ( new_n8113_, new_n8112_, new_n8111_ );
and  ( new_n8114_, new_n8113_, new_n734_ );
and  ( new_n8115_, new_n766_, RI2b1c4342e200_93 );
and  ( new_n8116_, new_n751_, RI2b1c4342e188_92 );
or   ( new_n8117_, new_n8116_, new_n8115_ );
and  ( new_n8118_, new_n8117_, new_n762_ );
or   ( new_n8119_, new_n8118_, new_n8114_ );
and  ( new_n8120_, new_n8119_, new_n8110_ );
or   ( new_n8121_, new_n8120_, new_n8109_ );
and  ( new_n8122_, new_n8121_, new_n8090_ );
or   ( new_n8123_, new_n8121_, new_n8090_ );
or   ( new_n8124_, new_n857_, new_n7274_ );
or   ( new_n8125_, new_n861_, new_n124_ );
and  ( new_n8126_, new_n8125_, new_n8124_ );
and  ( new_n8127_, new_n8126_, new_n842_ );
and  ( new_n8128_, new_n870_, RI2b1c4342e368_96 );
and  ( new_n8129_, new_n855_, RI2b1c4342e2f0_95 );
or   ( new_n8130_, new_n8129_, new_n8128_ );
and  ( new_n8131_, new_n8130_, new_n866_ );
or   ( new_n8132_, new_n8131_, new_n8127_ );
and  ( new_n8133_, new_n8132_, new_n8123_ );
or   ( new_n8134_, new_n8133_, new_n8122_ );
or   ( new_n8135_, new_n5308_, new_n110_ );
or   ( new_n8136_, new_n5312_, new_n755_ );
and  ( new_n8137_, new_n8136_, new_n8135_ );
and  ( new_n8138_, new_n8137_, new_n5182_ );
and  ( new_n8139_, new_n5316_, RI2b1c4342d7b0_71 );
and  ( new_n8140_, new_n5306_, RI2b1c4342d738_70 );
or   ( new_n8141_, new_n8140_, new_n8139_ );
and  ( new_n8142_, new_n8141_, new_n5028_ );
or   ( new_n8143_, new_n8142_, new_n8138_ );
or   ( new_n8144_, new_n4535_, new_n105_ );
or   ( new_n8145_, new_n4539_, new_n806_ );
and  ( new_n8146_, new_n8145_, new_n8144_ );
and  ( new_n8147_, new_n8146_, new_n4400_ );
and  ( new_n8148_, new_n4543_, RI2b1c4342d8a0_73 );
and  ( new_n8149_, new_n4533_, RI2b1c4342d828_72 );
or   ( new_n8150_, new_n8149_, new_n8148_ );
and  ( new_n8151_, new_n8150_, new_n4215_ );
or   ( new_n8152_, new_n8151_, new_n8147_ );
and  ( new_n8153_, new_n8152_, new_n8143_ );
or   ( new_n8154_, new_n8152_, new_n8143_ );
or   ( new_n8155_, new_n3802_, new_n843_ );
or   ( new_n8156_, new_n3806_, new_n859_ );
and  ( new_n8157_, new_n8156_, new_n8155_ );
and  ( new_n8158_, new_n8157_, new_n3695_ );
and  ( new_n8159_, new_n3810_, RI2b1c4342d990_75 );
and  ( new_n8160_, new_n3800_, RI2b1c4342d918_74 );
or   ( new_n8161_, new_n8160_, new_n8159_ );
and  ( new_n8162_, new_n8161_, new_n3548_ );
or   ( new_n8163_, new_n8162_, new_n8158_ );
and  ( new_n8164_, new_n8163_, new_n8154_ );
or   ( new_n8165_, new_n8164_, new_n8153_ );
or   ( new_n8166_, new_n7105_, new_n112_ );
or   ( new_n8167_, new_n7099_, new_n526_ );
and  ( new_n8168_, new_n8167_, new_n8166_ );
and  ( new_n8169_, new_n8168_, new_n5858_ );
and  ( new_n8170_, new_n7104_, RI2b1c4342d558_66 );
and  ( new_n8171_, new_n7110_, RI2b1c4342d5d0_67 );
or   ( new_n8172_, new_n8171_, new_n8170_ );
and  ( new_n8173_, new_n8172_, new_n6037_ );
or   ( new_n8174_, new_n8173_, new_n8169_ );
and  ( new_n8175_, new_n8174_, new_n842_ );
or   ( new_n8176_, new_n8174_, new_n842_ );
or   ( new_n8177_, new_n6156_, new_n591_ );
or   ( new_n8178_, new_n6160_, new_n612_ );
and  ( new_n8179_, new_n8178_, new_n8177_ );
and  ( new_n8180_, new_n8179_, new_n6039_ );
and  ( new_n8181_, new_n6164_, RI2b1c4342d6c0_69 );
and  ( new_n8182_, new_n6154_, RI2b1c4342d648_68 );
or   ( new_n8183_, new_n8182_, new_n8181_ );
and  ( new_n8184_, new_n8183_, new_n5867_ );
or   ( new_n8185_, new_n8184_, new_n8180_ );
and  ( new_n8186_, new_n8185_, new_n8176_ );
or   ( new_n8187_, new_n8186_, new_n8175_ );
and  ( new_n8188_, new_n8187_, new_n8165_ );
or   ( new_n8189_, new_n8187_, new_n8165_ );
or   ( new_n8190_, new_n3112_, new_n1004_ );
or   ( new_n8191_, new_n3116_, new_n886_ );
and  ( new_n8192_, new_n8191_, new_n8190_ );
and  ( new_n8193_, new_n8192_, new_n3004_ );
and  ( new_n8194_, new_n3120_, RI2b1c4342da80_77 );
and  ( new_n8195_, new_n3110_, RI2b1c4342da08_76 );
or   ( new_n8196_, new_n8195_, new_n8194_ );
and  ( new_n8197_, new_n8196_, new_n2868_ );
or   ( new_n8198_, new_n8197_, new_n8193_ );
or   ( new_n8199_, new_n2450_, new_n1310_ );
or   ( new_n8200_, new_n2454_, new_n1002_ );
and  ( new_n8201_, new_n8200_, new_n8199_ );
and  ( new_n8202_, new_n8201_, new_n2334_ );
and  ( new_n8203_, new_n2458_, RI2b1c4342db70_79 );
and  ( new_n8204_, new_n2448_, RI2b1c4342daf8_78 );
or   ( new_n8205_, new_n8204_, new_n8203_ );
and  ( new_n8206_, new_n8205_, new_n2168_ );
or   ( new_n8207_, new_n8206_, new_n8202_ );
and  ( new_n8208_, new_n8207_, new_n8198_ );
or   ( new_n8209_, new_n8207_, new_n8198_ );
or   ( new_n8210_, new_n1910_, new_n126_ );
or   ( new_n8211_, new_n1914_, new_n1511_ );
and  ( new_n8212_, new_n8211_, new_n8210_ );
and  ( new_n8213_, new_n8212_, new_n1824_ );
and  ( new_n8214_, new_n1918_, RI2b1c4342dc60_81 );
and  ( new_n8215_, new_n1908_, RI2b1c4342dbe8_80 );
or   ( new_n8216_, new_n8215_, new_n8214_ );
and  ( new_n8217_, new_n8216_, new_n1717_ );
or   ( new_n8218_, new_n8217_, new_n8213_ );
and  ( new_n8219_, new_n8218_, new_n8209_ );
or   ( new_n8220_, new_n8219_, new_n8208_ );
and  ( new_n8221_, new_n8220_, new_n8189_ );
or   ( new_n8222_, new_n8221_, new_n8188_ );
and  ( new_n8223_, new_n8222_, new_n8134_ );
or   ( new_n8224_, new_n8222_, new_n8134_ );
or   ( new_n8225_, new_n7926_, new_n7743_ );
and  ( new_n8226_, new_n8225_, new_n7753_ );
and  ( new_n8227_, new_n7922_, new_n7742_ );
and  ( new_n8228_, new_n7925_, new_n7733_ );
or   ( new_n8229_, new_n8228_, new_n8227_ );
and  ( new_n8230_, new_n8229_, new_n7930_ );
or   ( new_n8231_, new_n8230_, new_n8226_ );
or   ( new_n8232_, new_n7913_, new_n7712_ );
and  ( new_n8233_, new_n8232_, new_n7722_ );
and  ( new_n8234_, new_n7909_, new_n7711_ );
and  ( new_n8235_, new_n7912_, new_n7702_ );
or   ( new_n8236_, new_n8235_, new_n8234_ );
and  ( new_n8237_, new_n8236_, new_n7917_ );
or   ( new_n8238_, new_n8237_, new_n8233_ );
and  ( new_n8239_, new_n8238_, new_n8231_ );
or   ( new_n8240_, new_n8238_, new_n8231_ );
or   ( new_n8241_, new_n7898_, new_n7679_ );
and  ( new_n8242_, new_n8241_, new_n7689_ );
and  ( new_n8243_, new_n7894_, new_n7678_ );
and  ( new_n8244_, new_n7897_, new_n7669_ );
or   ( new_n8245_, new_n8244_, new_n8243_ );
and  ( new_n8246_, new_n8245_, new_n7902_ );
or   ( new_n8247_, new_n8246_, new_n8242_ );
and  ( new_n8248_, new_n8247_, new_n8240_ );
or   ( new_n8249_, new_n8248_, new_n8239_ );
and  ( new_n8250_, new_n8249_, new_n8224_ );
or   ( new_n8251_, new_n8250_, new_n8223_ );
and  ( new_n8252_, new_n8251_, new_n8059_ );
or   ( new_n8253_, new_n8251_, new_n8059_ );
or   ( new_n8254_, new_n7933_, new_n7756_ );
and  ( new_n8255_, new_n8254_, new_n7764_ );
and  ( new_n8256_, new_n7919_, new_n7755_ );
and  ( new_n8257_, new_n7932_, new_n7724_ );
or   ( new_n8258_, new_n8257_, new_n8256_ );
and  ( new_n8259_, new_n8258_, new_n7937_ );
or   ( new_n8260_, new_n8259_, new_n8255_ );
or   ( new_n8261_, new_n7890_, new_n7659_ );
and  ( new_n8262_, new_n8261_, new_n7691_ );
and  ( new_n8263_, new_n7876_, new_n7658_ );
and  ( new_n8264_, new_n7889_, new_n7627_ );
or   ( new_n8265_, new_n8264_, new_n8263_ );
and  ( new_n8266_, new_n8265_, new_n7904_ );
or   ( new_n8267_, new_n8266_, new_n8262_ );
or   ( new_n8268_, new_n8267_, new_n8260_ );
and  ( new_n8269_, new_n8268_, new_n8253_ );
or   ( new_n8270_, new_n8269_, new_n8252_ );
and  ( new_n8271_, new_n8270_, new_n8039_ );
or   ( new_n8272_, new_n8270_, new_n8039_ );
or   ( new_n8273_, new_n7983_, new_n7586_ );
and  ( new_n8274_, new_n8273_, new_n7594_ );
and  ( new_n8275_, new_n7979_, new_n7585_ );
and  ( new_n8276_, new_n7982_, new_n7578_ );
or   ( new_n8277_, new_n8276_, new_n8275_ );
and  ( new_n8278_, new_n8277_, new_n7987_ );
or   ( new_n8279_, new_n8278_, new_n8274_ );
and  ( new_n8280_, new_n8279_, new_n8272_ );
or   ( new_n8281_, new_n8280_, new_n8271_ );
and  ( new_n8282_, new_n8281_, new_n8014_ );
or   ( new_n8283_, new_n8281_, new_n8014_ );
or   ( new_n8284_, new_n7990_, new_n7832_ );
and  ( new_n8285_, new_n8284_, new_n7840_ );
and  ( new_n8286_, new_n7976_, new_n7596_ );
and  ( new_n8287_, new_n7989_, new_n7831_ );
or   ( new_n8288_, new_n8287_, new_n8286_ );
and  ( new_n8289_, new_n8288_, new_n7994_ );
or   ( new_n8290_, new_n8289_, new_n8285_ );
and  ( new_n8291_, new_n8290_, new_n8283_ );
or   ( new_n8292_, new_n8291_, new_n8282_ );
and  ( new_n8293_, new_n8292_, new_n8007_ );
or   ( new_n8294_, new_n8292_, new_n8007_ );
and  ( new_n8295_, new_n8012_, new_n7356_ );
and  ( new_n8296_, new_n8008_, new_n7549_ );
or   ( new_n8297_, new_n8296_, new_n8295_ );
and  ( new_n8298_, new_n8019_, new_n7187_ );
and  ( new_n8299_, new_n8015_, new_n7485_ );
or   ( new_n8300_, new_n8299_, new_n8298_ );
and  ( new_n8301_, new_n8026_, new_n7818_ );
and  ( new_n8302_, new_n8022_, new_n7967_ );
or   ( new_n8303_, new_n8302_, new_n8301_ );
and  ( new_n8304_, new_n8303_, new_n8300_ );
or   ( new_n8305_, new_n8303_, new_n8300_ );
and  ( new_n8306_, new_n8035_, new_n7793_ );
and  ( new_n8307_, new_n8031_, new_n7954_ );
or   ( new_n8308_, new_n8307_, new_n8306_ );
and  ( new_n8309_, new_n8308_, new_n8305_ );
or   ( new_n8310_, new_n8309_, new_n8304_ );
and  ( new_n8311_, new_n8044_, new_n7152_ );
and  ( new_n8312_, new_n8040_, new_n7468_ );
or   ( new_n8313_, new_n8312_, new_n8311_ );
and  ( new_n8314_, new_n7453_, new_n7122_ );
and  ( new_n8315_, new_n7456_, new_n7113_ );
or   ( new_n8316_, new_n8315_, new_n8314_ );
and  ( new_n8317_, new_n8316_, new_n8313_ );
or   ( new_n8318_, new_n8316_, new_n8313_ );
and  ( new_n8319_, new_n8055_, new_n7791_ );
and  ( new_n8320_, new_n8051_, new_n7952_ );
or   ( new_n8321_, new_n8320_, new_n8319_ );
and  ( new_n8322_, new_n8321_, new_n8318_ );
or   ( new_n8323_, new_n8322_, new_n8317_ );
and  ( new_n8324_, new_n8066_, new_n1355_ );
and  ( new_n8325_, new_n8062_, new_n1267_ );
or   ( new_n8326_, new_n8325_, new_n8324_ );
and  ( new_n8327_, new_n8075_, new_n913_ );
and  ( new_n8328_, new_n8071_, new_n938_ );
or   ( new_n8329_, new_n8328_, new_n8327_ );
and  ( new_n8330_, new_n8329_, new_n8326_ );
or   ( new_n8331_, new_n8329_, new_n8326_ );
and  ( new_n8332_, new_n8086_, new_n428_ );
and  ( new_n8333_, new_n8082_, new_n457_ );
or   ( new_n8334_, new_n8333_, new_n8332_ );
and  ( new_n8335_, new_n8334_, new_n8331_ );
or   ( new_n8336_, new_n8335_, new_n8330_ );
and  ( new_n8337_, new_n8097_, new_n505_ );
and  ( new_n8338_, new_n8093_, new_n533_ );
or   ( new_n8339_, new_n8338_, new_n8337_ );
and  ( new_n8340_, new_n8106_, new_n590_ );
and  ( new_n8341_, new_n8102_, new_n619_ );
or   ( new_n8342_, new_n8341_, new_n8340_ );
and  ( new_n8343_, new_n8342_, new_n8339_ );
or   ( new_n8344_, new_n8342_, new_n8339_ );
and  ( new_n8345_, new_n8117_, new_n734_ );
and  ( new_n8346_, new_n8113_, new_n762_ );
or   ( new_n8347_, new_n8346_, new_n8345_ );
and  ( new_n8348_, new_n8347_, new_n8344_ );
or   ( new_n8349_, new_n8348_, new_n8343_ );
and  ( new_n8350_, new_n8349_, new_n8336_ );
or   ( new_n8351_, new_n8349_, new_n8336_ );
and  ( new_n8352_, new_n8130_, new_n842_ );
and  ( new_n8353_, new_n8126_, new_n866_ );
or   ( new_n8354_, new_n8353_, new_n8352_ );
and  ( new_n8355_, new_n8354_, new_n8351_ );
or   ( new_n8356_, new_n8355_, new_n8350_ );
and  ( new_n8357_, new_n8141_, new_n5182_ );
and  ( new_n8358_, new_n8137_, new_n5028_ );
or   ( new_n8359_, new_n8358_, new_n8357_ );
and  ( new_n8360_, new_n8150_, new_n4400_ );
and  ( new_n8361_, new_n8146_, new_n4215_ );
or   ( new_n8362_, new_n8361_, new_n8360_ );
and  ( new_n8363_, new_n8362_, new_n8359_ );
or   ( new_n8364_, new_n8362_, new_n8359_ );
and  ( new_n8365_, new_n8161_, new_n3695_ );
and  ( new_n8366_, new_n8157_, new_n3548_ );
or   ( new_n8367_, new_n8366_, new_n8365_ );
and  ( new_n8368_, new_n8367_, new_n8364_ );
or   ( new_n8369_, new_n8368_, new_n8363_ );
and  ( new_n8370_, new_n8172_, new_n5858_ );
and  ( new_n8371_, new_n8168_, new_n6037_ );
or   ( new_n8372_, new_n8371_, new_n8370_ );
or   ( new_n8373_, new_n8372_, new_n866_ );
and  ( new_n8374_, new_n8372_, new_n866_ );
and  ( new_n8375_, new_n8183_, new_n6039_ );
and  ( new_n8376_, new_n8179_, new_n5867_ );
or   ( new_n8377_, new_n8376_, new_n8375_ );
or   ( new_n8378_, new_n8377_, new_n8374_ );
and  ( new_n8379_, new_n8378_, new_n8373_ );
or   ( new_n8380_, new_n8379_, new_n8369_ );
and  ( new_n8381_, new_n8379_, new_n8369_ );
and  ( new_n8382_, new_n8196_, new_n3004_ );
and  ( new_n8383_, new_n8192_, new_n2868_ );
or   ( new_n8384_, new_n8383_, new_n8382_ );
and  ( new_n8385_, new_n8205_, new_n2334_ );
and  ( new_n8386_, new_n8201_, new_n2168_ );
or   ( new_n8387_, new_n8386_, new_n8385_ );
and  ( new_n8388_, new_n8387_, new_n8384_ );
or   ( new_n8389_, new_n8387_, new_n8384_ );
and  ( new_n8390_, new_n8216_, new_n1824_ );
and  ( new_n8391_, new_n8212_, new_n1717_ );
or   ( new_n8392_, new_n8391_, new_n8390_ );
and  ( new_n8393_, new_n8392_, new_n8389_ );
or   ( new_n8394_, new_n8393_, new_n8388_ );
or   ( new_n8395_, new_n8394_, new_n8381_ );
and  ( new_n8396_, new_n8395_, new_n8380_ );
or   ( new_n8397_, new_n8396_, new_n8356_ );
and  ( new_n8398_, new_n8396_, new_n8356_ );
and  ( new_n8399_, new_n8229_, new_n7753_ );
and  ( new_n8400_, new_n8225_, new_n7930_ );
or   ( new_n8401_, new_n8400_, new_n8399_ );
and  ( new_n8402_, new_n8236_, new_n7722_ );
and  ( new_n8403_, new_n8232_, new_n7917_ );
or   ( new_n8404_, new_n8403_, new_n8402_ );
and  ( new_n8405_, new_n8404_, new_n8401_ );
or   ( new_n8406_, new_n8404_, new_n8401_ );
and  ( new_n8407_, new_n8245_, new_n7689_ );
and  ( new_n8408_, new_n8241_, new_n7902_ );
or   ( new_n8409_, new_n8408_, new_n8407_ );
and  ( new_n8410_, new_n8409_, new_n8406_ );
or   ( new_n8411_, new_n8410_, new_n8405_ );
or   ( new_n8412_, new_n8411_, new_n8398_ );
and  ( new_n8413_, new_n8412_, new_n8397_ );
or   ( new_n8414_, new_n8413_, new_n8323_ );
and  ( new_n8415_, new_n8413_, new_n8323_ );
and  ( new_n8416_, new_n8258_, new_n7764_ );
and  ( new_n8417_, new_n8254_, new_n7937_ );
or   ( new_n8418_, new_n8417_, new_n8416_ );
and  ( new_n8419_, new_n8265_, new_n7691_ );
and  ( new_n8420_, new_n8261_, new_n7904_ );
or   ( new_n8421_, new_n8420_, new_n8419_ );
and  ( new_n8422_, new_n8421_, new_n8418_ );
or   ( new_n8423_, new_n8422_, new_n8415_ );
and  ( new_n8424_, new_n8423_, new_n8414_ );
or   ( new_n8425_, new_n8424_, new_n8310_ );
and  ( new_n8426_, new_n8424_, new_n8310_ );
and  ( new_n8427_, new_n8277_, new_n7594_ );
and  ( new_n8428_, new_n8273_, new_n7987_ );
or   ( new_n8429_, new_n8428_, new_n8427_ );
or   ( new_n8430_, new_n8429_, new_n8426_ );
and  ( new_n8431_, new_n8430_, new_n8425_ );
and  ( new_n8432_, new_n8431_, new_n8297_ );
or   ( new_n8433_, new_n8432_, new_n8282_ );
and  ( new_n8434_, new_n8433_, new_n8290_ );
and  ( new_n8435_, new_n8431_, new_n8014_ );
and  ( new_n8436_, new_n8297_, new_n8281_ );
or   ( new_n8437_, new_n8436_, new_n8435_ );
and  ( new_n8438_, new_n8288_, new_n7840_ );
and  ( new_n8439_, new_n8284_, new_n7994_ );
or   ( new_n8440_, new_n8439_, new_n8438_ );
and  ( new_n8441_, new_n8440_, new_n8437_ );
or   ( new_n8442_, new_n8441_, new_n8434_ );
or   ( new_n8443_, new_n7970_, new_n7821_ );
and  ( new_n8444_, new_n8443_, new_n7829_ );
and  ( new_n8445_, new_n7956_, new_n7820_ );
and  ( new_n8446_, new_n7969_, new_n7795_ );
or   ( new_n8447_, new_n8446_, new_n8445_ );
and  ( new_n8448_, new_n8447_, new_n7974_ );
or   ( new_n8449_, new_n8448_, new_n8444_ );
or   ( new_n8450_, new_n6156_, new_n755_ );
or   ( new_n8451_, new_n6160_, new_n591_ );
and  ( new_n8452_, new_n8451_, new_n8450_ );
and  ( new_n8453_, new_n8452_, new_n6039_ );
and  ( new_n8454_, new_n6164_, RI2b1c4342d738_70 );
and  ( new_n8455_, new_n6154_, RI2b1c4342d6c0_69 );
or   ( new_n8456_, new_n8455_, new_n8454_ );
and  ( new_n8457_, new_n8456_, new_n5867_ );
or   ( new_n8458_, new_n8457_, new_n8453_ );
or   ( new_n8459_, new_n7105_, new_n612_ );
or   ( new_n8460_, new_n7099_, new_n112_ );
and  ( new_n8461_, new_n8460_, new_n8459_ );
and  ( new_n8462_, new_n8461_, new_n5858_ );
and  ( new_n8463_, new_n7104_, RI2b1c4342d5d0_67 );
and  ( new_n8464_, new_n7110_, RI2b1c4342d648_68 );
or   ( new_n8465_, new_n8464_, new_n8463_ );
and  ( new_n8466_, new_n8465_, new_n6037_ );
or   ( new_n8467_, new_n8466_, new_n8462_ );
and  ( new_n8468_, new_n8467_, new_n8458_ );
or   ( new_n8469_, new_n8467_, new_n8458_ );
or   ( new_n8470_, new_n5308_, new_n806_ );
or   ( new_n8471_, new_n5312_, new_n110_ );
and  ( new_n8472_, new_n8471_, new_n8470_ );
and  ( new_n8473_, new_n8472_, new_n5182_ );
and  ( new_n8474_, new_n5316_, RI2b1c4342d828_72 );
and  ( new_n8475_, new_n5306_, RI2b1c4342d7b0_71 );
or   ( new_n8476_, new_n8475_, new_n8474_ );
and  ( new_n8477_, new_n8476_, new_n5028_ );
or   ( new_n8478_, new_n8477_, new_n8473_ );
and  ( new_n8479_, new_n8478_, new_n8469_ );
or   ( new_n8480_, new_n8479_, new_n8468_ );
or   ( new_n8481_, new_n4535_, new_n859_ );
or   ( new_n8482_, new_n4539_, new_n105_ );
and  ( new_n8483_, new_n8482_, new_n8481_ );
and  ( new_n8484_, new_n8483_, new_n4400_ );
and  ( new_n8485_, new_n4543_, RI2b1c4342d918_74 );
and  ( new_n8486_, new_n4533_, RI2b1c4342d8a0_73 );
or   ( new_n8487_, new_n8486_, new_n8485_ );
and  ( new_n8488_, new_n8487_, new_n4215_ );
or   ( new_n8489_, new_n8488_, new_n8484_ );
or   ( new_n8490_, new_n3802_, new_n886_ );
or   ( new_n8491_, new_n3806_, new_n843_ );
and  ( new_n8492_, new_n8491_, new_n8490_ );
and  ( new_n8493_, new_n8492_, new_n3695_ );
and  ( new_n8494_, new_n3810_, RI2b1c4342da08_76 );
and  ( new_n8495_, new_n3800_, RI2b1c4342d990_75 );
or   ( new_n8496_, new_n8495_, new_n8494_ );
and  ( new_n8497_, new_n8496_, new_n3548_ );
or   ( new_n8498_, new_n8497_, new_n8493_ );
and  ( new_n8499_, new_n8498_, new_n8489_ );
or   ( new_n8500_, new_n8498_, new_n8489_ );
or   ( new_n8501_, new_n3112_, new_n1002_ );
or   ( new_n8502_, new_n3116_, new_n1004_ );
and  ( new_n8503_, new_n8502_, new_n8501_ );
and  ( new_n8504_, new_n8503_, new_n3004_ );
and  ( new_n8505_, new_n3120_, RI2b1c4342daf8_78 );
and  ( new_n8506_, new_n3110_, RI2b1c4342da80_77 );
or   ( new_n8507_, new_n8506_, new_n8505_ );
and  ( new_n8508_, new_n8507_, new_n2868_ );
or   ( new_n8509_, new_n8508_, new_n8504_ );
and  ( new_n8510_, new_n8509_, new_n8500_ );
or   ( new_n8511_, new_n8510_, new_n8499_ );
and  ( new_n8512_, new_n8511_, new_n8480_ );
or   ( new_n8513_, new_n8511_, new_n8480_ );
or   ( new_n8514_, new_n2450_, new_n1511_ );
or   ( new_n8515_, new_n2454_, new_n1310_ );
and  ( new_n8516_, new_n8515_, new_n8514_ );
and  ( new_n8517_, new_n8516_, new_n2334_ );
and  ( new_n8518_, new_n2458_, RI2b1c4342dbe8_80 );
and  ( new_n8519_, new_n2448_, RI2b1c4342db70_79 );
or   ( new_n8520_, new_n8519_, new_n8518_ );
and  ( new_n8521_, new_n8520_, new_n2168_ );
or   ( new_n8522_, new_n8521_, new_n8517_ );
or   ( new_n8523_, new_n1910_, new_n2119_ );
or   ( new_n8524_, new_n1914_, new_n126_ );
and  ( new_n8525_, new_n8524_, new_n8523_ );
and  ( new_n8526_, new_n8525_, new_n1824_ );
and  ( new_n8527_, new_n1918_, RI2b1c4342dcd8_82 );
and  ( new_n8528_, new_n1908_, RI2b1c4342dc60_81 );
or   ( new_n8529_, new_n8528_, new_n8527_ );
and  ( new_n8530_, new_n8529_, new_n1717_ );
or   ( new_n8531_, new_n8530_, new_n8526_ );
and  ( new_n8532_, new_n8531_, new_n8522_ );
or   ( new_n8533_, new_n8531_, new_n8522_ );
or   ( new_n8534_, new_n1425_, new_n2541_ );
or   ( new_n8535_, new_n1429_, new_n121_ );
and  ( new_n8536_, new_n8535_, new_n8534_ );
and  ( new_n8537_, new_n8536_, new_n1355_ );
and  ( new_n8538_, new_n1433_, RI2b1c4342ddc8_84 );
and  ( new_n8539_, new_n1423_, RI2b1c4342dd50_83 );
or   ( new_n8540_, new_n8539_, new_n8538_ );
and  ( new_n8541_, new_n8540_, new_n1267_ );
or   ( new_n8542_, new_n8541_, new_n8537_ );
and  ( new_n8543_, new_n8542_, new_n8533_ );
or   ( new_n8544_, new_n8543_, new_n8532_ );
and  ( new_n8545_, new_n8544_, new_n8513_ );
or   ( new_n8546_, new_n8545_, new_n8512_ );
or   ( new_n8547_, new_n934_, new_n3239_ );
or   ( new_n8548_, new_n940_, new_n2806_ );
and  ( new_n8549_, new_n8548_, new_n8547_ );
and  ( new_n8550_, new_n8549_, new_n913_ );
and  ( new_n8551_, new_n944_, RI2b1c4342deb8_86 );
and  ( new_n8552_, new_n932_, RI2b1c4342de40_85 );
or   ( new_n8553_, new_n8552_, new_n8551_ );
and  ( new_n8554_, new_n8553_, new_n938_ );
or   ( new_n8555_, new_n8554_, new_n8550_ );
or   ( new_n8556_, new_n453_, new_n3902_ );
or   ( new_n8557_, new_n459_, new_n3924_ );
and  ( new_n8558_, new_n8557_, new_n8556_ );
and  ( new_n8559_, new_n8558_, new_n428_ );
and  ( new_n8560_, new_n463_, RI2b1c4342dfa8_88 );
and  ( new_n8561_, new_n451_, RI2b1c4342df30_87 );
or   ( new_n8562_, new_n8561_, new_n8560_ );
and  ( new_n8563_, new_n8562_, new_n457_ );
or   ( new_n8564_, new_n8563_, new_n8559_ );
and  ( new_n8565_, new_n8564_, new_n8555_ );
or   ( new_n8566_, new_n8564_, new_n8555_ );
or   ( new_n8567_, new_n524_, new_n4635_ );
or   ( new_n8568_, new_n528_, new_n132_ );
and  ( new_n8569_, new_n8568_, new_n8567_ );
and  ( new_n8570_, new_n8569_, new_n505_ );
and  ( new_n8571_, new_n537_, RI2b1c4342e098_90 );
and  ( new_n8572_, new_n522_, RI2b1c4342e020_89 );
or   ( new_n8573_, new_n8572_, new_n8571_ );
and  ( new_n8574_, new_n8573_, new_n533_ );
or   ( new_n8575_, new_n8574_, new_n8570_ );
and  ( new_n8576_, new_n8575_, new_n8566_ );
or   ( new_n8577_, new_n8576_, new_n8565_ );
or   ( new_n8578_, new_n610_, new_n5459_ );
or   ( new_n8579_, new_n614_, new_n117_ );
and  ( new_n8580_, new_n8579_, new_n8578_ );
and  ( new_n8581_, new_n8580_, new_n590_ );
and  ( new_n8582_, new_n623_, RI2b1c4342e188_92 );
and  ( new_n8583_, new_n608_, RI2b1c4342e110_91 );
or   ( new_n8584_, new_n8583_, new_n8582_ );
and  ( new_n8585_, new_n8584_, new_n619_ );
or   ( new_n8586_, new_n8585_, new_n8581_ );
or   ( new_n8587_, new_n753_, new_n6321_ );
or   ( new_n8588_, new_n757_, new_n6307_ );
and  ( new_n8589_, new_n8588_, new_n8587_ );
and  ( new_n8590_, new_n8589_, new_n734_ );
and  ( new_n8591_, new_n766_, RI2b1c4342e278_94 );
and  ( new_n8592_, new_n751_, RI2b1c4342e200_93 );
or   ( new_n8593_, new_n8592_, new_n8591_ );
and  ( new_n8594_, new_n8593_, new_n762_ );
or   ( new_n8595_, new_n8594_, new_n8590_ );
and  ( new_n8596_, new_n8595_, new_n8586_ );
or   ( new_n8597_, new_n8595_, new_n8586_ );
or   ( new_n8598_, new_n804_, new_n7274_ );
or   ( new_n8599_, new_n808_, new_n124_ );
and  ( new_n8600_, new_n8599_, new_n8598_ );
and  ( new_n8601_, new_n8600_, new_n785_ );
and  ( new_n8602_, new_n817_, RI2b1c4342e368_96 );
and  ( new_n8603_, new_n802_, RI2b1c4342e2f0_95 );
or   ( new_n8604_, new_n8603_, new_n8602_ );
and  ( new_n8605_, new_n8604_, new_n813_ );
or   ( new_n8606_, new_n8605_, new_n8601_ );
and  ( new_n8607_, new_n8606_, new_n8597_ );
or   ( new_n8608_, new_n8607_, new_n8596_ );
and  ( new_n8609_, new_n8608_, new_n8577_ );
or   ( new_n8610_, new_n8608_, new_n8577_ );
or   ( new_n8611_, new_n804_, new_n124_ );
or   ( new_n8612_, new_n808_, new_n6321_ );
and  ( new_n8613_, new_n8612_, new_n8611_ );
and  ( new_n8614_, new_n8613_, new_n785_ );
and  ( new_n8615_, new_n817_, RI2b1c4342e2f0_95 );
and  ( new_n8616_, new_n802_, RI2b1c4342e278_94 );
or   ( new_n8617_, new_n8616_, new_n8615_ );
and  ( new_n8618_, new_n8617_, new_n813_ );
or   ( new_n8619_, new_n8618_, new_n8614_ );
and  ( new_n8620_, new_n8619_, new_n8610_ );
or   ( new_n8621_, new_n8620_, new_n8609_ );
and  ( new_n8622_, new_n8621_, new_n8546_ );
or   ( new_n8623_, new_n8621_, new_n8546_ );
or   ( new_n8624_, new_n861_, new_n7274_ );
and  ( new_n8625_, new_n8624_, new_n842_ );
and  ( new_n8626_, new_n855_, RI2b1c4342e368_96 );
and  ( new_n8627_, new_n8626_, new_n866_ );
or   ( new_n8628_, new_n8627_, new_n8625_ );
or   ( new_n8629_, new_n8343_, new_n8109_ );
and  ( new_n8630_, new_n8629_, new_n8119_ );
and  ( new_n8631_, new_n8339_, new_n8108_ );
and  ( new_n8632_, new_n8342_, new_n8099_ );
or   ( new_n8633_, new_n8632_, new_n8631_ );
and  ( new_n8634_, new_n8633_, new_n8347_ );
or   ( new_n8635_, new_n8634_, new_n8630_ );
and  ( new_n8636_, new_n8635_, new_n8628_ );
or   ( new_n8637_, new_n8635_, new_n8628_ );
or   ( new_n8638_, new_n8330_, new_n8078_ );
and  ( new_n8639_, new_n8638_, new_n8088_ );
and  ( new_n8640_, new_n8326_, new_n8077_ );
and  ( new_n8641_, new_n8329_, new_n8068_ );
or   ( new_n8642_, new_n8641_, new_n8640_ );
and  ( new_n8643_, new_n8642_, new_n8334_ );
or   ( new_n8644_, new_n8643_, new_n8639_ );
and  ( new_n8645_, new_n8644_, new_n8637_ );
or   ( new_n8646_, new_n8645_, new_n8636_ );
and  ( new_n8647_, new_n8646_, new_n8623_ );
or   ( new_n8648_, new_n8647_, new_n8622_ );
or   ( new_n8649_, new_n7883_, new_n7646_ );
and  ( new_n8650_, new_n8649_, new_n7656_ );
and  ( new_n8651_, new_n7879_, new_n7645_ );
and  ( new_n8652_, new_n7882_, new_n7636_ );
or   ( new_n8653_, new_n8652_, new_n8651_ );
and  ( new_n8654_, new_n8653_, new_n7887_ );
or   ( new_n8655_, new_n8654_, new_n8650_ );
or   ( new_n8656_, new_n8388_, new_n8208_ );
and  ( new_n8657_, new_n8656_, new_n8218_ );
and  ( new_n8658_, new_n8384_, new_n8207_ );
and  ( new_n8659_, new_n8387_, new_n8198_ );
or   ( new_n8660_, new_n8659_, new_n8658_ );
and  ( new_n8661_, new_n8660_, new_n8392_ );
or   ( new_n8662_, new_n8661_, new_n8657_ );
or   ( new_n8663_, new_n8363_, new_n8153_ );
and  ( new_n8664_, new_n8663_, new_n8163_ );
and  ( new_n8665_, new_n8359_, new_n8152_ );
and  ( new_n8666_, new_n8362_, new_n8143_ );
or   ( new_n8667_, new_n8666_, new_n8665_ );
and  ( new_n8668_, new_n8667_, new_n8367_ );
or   ( new_n8669_, new_n8668_, new_n8664_ );
and  ( new_n8670_, new_n8669_, new_n8662_ );
or   ( new_n8671_, new_n8669_, new_n8662_ );
or   ( new_n8672_, new_n8374_, new_n8175_ );
and  ( new_n8673_, new_n8672_, new_n8185_ );
and  ( new_n8674_, new_n8174_, new_n866_ );
and  ( new_n8675_, new_n8372_, new_n842_ );
or   ( new_n8676_, new_n8675_, new_n8674_ );
and  ( new_n8677_, new_n8676_, new_n8377_ );
or   ( new_n8678_, new_n8677_, new_n8673_ );
and  ( new_n8679_, new_n8678_, new_n8671_ );
or   ( new_n8680_, new_n8679_, new_n8670_ );
and  ( new_n8681_, new_n8680_, new_n8655_ );
or   ( new_n8682_, new_n8680_, new_n8655_ );
or   ( new_n8683_, new_n7870_, new_n7615_ );
and  ( new_n8684_, new_n8683_, new_n7625_ );
and  ( new_n8685_, new_n7866_, new_n7614_ );
and  ( new_n8686_, new_n7869_, new_n7605_ );
or   ( new_n8687_, new_n8686_, new_n8685_ );
and  ( new_n8688_, new_n8687_, new_n7874_ );
or   ( new_n8689_, new_n8688_, new_n8684_ );
and  ( new_n8690_, new_n8689_, new_n8682_ );
or   ( new_n8691_, new_n8690_, new_n8681_ );
and  ( new_n8692_, new_n8691_, new_n8648_ );
or   ( new_n8693_, new_n8691_, new_n8648_ );
or   ( new_n8694_, new_n8405_, new_n8239_ );
and  ( new_n8695_, new_n8694_, new_n8247_ );
and  ( new_n8696_, new_n8401_, new_n8238_ );
and  ( new_n8697_, new_n8404_, new_n8231_ );
or   ( new_n8698_, new_n8697_, new_n8696_ );
and  ( new_n8699_, new_n8698_, new_n8409_ );
or   ( new_n8700_, new_n8699_, new_n8695_ );
or   ( new_n8701_, new_n8350_, new_n8122_ );
and  ( new_n8702_, new_n8701_, new_n8132_ );
and  ( new_n8703_, new_n8336_, new_n8121_ );
and  ( new_n8704_, new_n8349_, new_n8090_ );
or   ( new_n8705_, new_n8704_, new_n8703_ );
and  ( new_n8706_, new_n8705_, new_n8354_ );
or   ( new_n8707_, new_n8706_, new_n8702_ );
and  ( new_n8708_, new_n8707_, new_n8700_ );
or   ( new_n8709_, new_n8707_, new_n8700_ );
or   ( new_n8710_, new_n8381_, new_n8188_ );
and  ( new_n8711_, new_n8710_, new_n8220_ );
and  ( new_n8712_, new_n8379_, new_n8165_ );
and  ( new_n8713_, new_n8369_, new_n8187_ );
or   ( new_n8714_, new_n8713_, new_n8712_ );
and  ( new_n8715_, new_n8714_, new_n8394_ );
or   ( new_n8716_, new_n8715_, new_n8711_ );
and  ( new_n8717_, new_n8716_, new_n8709_ );
or   ( new_n8718_, new_n8717_, new_n8708_ );
and  ( new_n8719_, new_n8718_, new_n8693_ );
or   ( new_n8720_, new_n8719_, new_n8692_ );
and  ( new_n8721_, new_n8267_, new_n8260_ );
or   ( new_n8722_, new_n8721_, new_n8422_ );
or   ( new_n8723_, new_n8317_, new_n8049_ );
and  ( new_n8724_, new_n8723_, new_n8057_ );
and  ( new_n8725_, new_n8313_, new_n8048_ );
and  ( new_n8726_, new_n8316_, new_n8046_ );
or   ( new_n8727_, new_n8726_, new_n8725_ );
and  ( new_n8728_, new_n8727_, new_n8321_ );
or   ( new_n8729_, new_n8728_, new_n8724_ );
and  ( new_n8730_, new_n8729_, new_n8722_ );
or   ( new_n8731_, new_n8729_, new_n8722_ );
or   ( new_n8732_, new_n8398_, new_n8223_ );
and  ( new_n8733_, new_n8732_, new_n8249_ );
and  ( new_n8734_, new_n8396_, new_n8134_ );
and  ( new_n8735_, new_n8356_, new_n8222_ );
or   ( new_n8736_, new_n8735_, new_n8734_ );
and  ( new_n8737_, new_n8736_, new_n8411_ );
or   ( new_n8738_, new_n8737_, new_n8733_ );
and  ( new_n8739_, new_n8738_, new_n8731_ );
or   ( new_n8740_, new_n8739_, new_n8730_ );
and  ( new_n8741_, new_n8740_, new_n8720_ );
or   ( new_n8742_, new_n8740_, new_n8720_ );
or   ( new_n8743_, new_n8304_, new_n8029_ );
and  ( new_n8744_, new_n8743_, new_n8037_ );
and  ( new_n8745_, new_n8300_, new_n8028_ );
and  ( new_n8746_, new_n8303_, new_n8021_ );
or   ( new_n8747_, new_n8746_, new_n8745_ );
and  ( new_n8748_, new_n8747_, new_n8308_ );
or   ( new_n8749_, new_n8748_, new_n8744_ );
and  ( new_n8750_, new_n8749_, new_n8742_ );
or   ( new_n8751_, new_n8750_, new_n8741_ );
and  ( new_n8752_, new_n8751_, new_n8449_ );
or   ( new_n8753_, new_n8751_, new_n8449_ );
or   ( new_n8754_, new_n8426_, new_n8271_ );
and  ( new_n8755_, new_n8754_, new_n8279_ );
and  ( new_n8756_, new_n8424_, new_n8039_ );
and  ( new_n8757_, new_n8310_, new_n8270_ );
or   ( new_n8758_, new_n8757_, new_n8756_ );
and  ( new_n8759_, new_n8758_, new_n8429_ );
or   ( new_n8760_, new_n8759_, new_n8755_ );
and  ( new_n8761_, new_n8760_, new_n8753_ );
or   ( new_n8762_, new_n8761_, new_n8752_ );
or   ( new_n8763_, new_n8762_, new_n8442_ );
and  ( new_n8764_, new_n8763_, new_n8294_ );
or   ( new_n8765_, new_n8764_, new_n8293_ );
and  ( new_n8766_, new_n8762_, new_n8442_ );
or   ( new_n8767_, new_n8766_, new_n8293_ );
and  ( new_n8768_, new_n8447_, new_n7829_ );
and  ( new_n8769_, new_n8443_, new_n7974_ );
or   ( new_n8770_, new_n8769_, new_n8768_ );
and  ( new_n8771_, new_n8465_, new_n5858_ );
and  ( new_n8772_, new_n8461_, new_n6037_ );
or   ( new_n8773_, new_n8772_, new_n8771_ );
and  ( new_n8774_, new_n8456_, new_n6039_ );
and  ( new_n8775_, new_n8452_, new_n5867_ );
or   ( new_n8776_, new_n8775_, new_n8774_ );
and  ( new_n8777_, new_n8776_, new_n8773_ );
or   ( new_n8778_, new_n8776_, new_n8773_ );
and  ( new_n8779_, new_n8476_, new_n5182_ );
and  ( new_n8780_, new_n8472_, new_n5028_ );
or   ( new_n8781_, new_n8780_, new_n8779_ );
and  ( new_n8782_, new_n8781_, new_n8778_ );
or   ( new_n8783_, new_n8782_, new_n8777_ );
and  ( new_n8784_, new_n8487_, new_n4400_ );
and  ( new_n8785_, new_n8483_, new_n4215_ );
or   ( new_n8786_, new_n8785_, new_n8784_ );
and  ( new_n8787_, new_n8496_, new_n3695_ );
and  ( new_n8788_, new_n8492_, new_n3548_ );
or   ( new_n8789_, new_n8788_, new_n8787_ );
and  ( new_n8790_, new_n8789_, new_n8786_ );
or   ( new_n8791_, new_n8789_, new_n8786_ );
and  ( new_n8792_, new_n8507_, new_n3004_ );
and  ( new_n8793_, new_n8503_, new_n2868_ );
or   ( new_n8794_, new_n8793_, new_n8792_ );
and  ( new_n8795_, new_n8794_, new_n8791_ );
or   ( new_n8796_, new_n8795_, new_n8790_ );
and  ( new_n8797_, new_n8796_, new_n8783_ );
or   ( new_n8798_, new_n8796_, new_n8783_ );
and  ( new_n8799_, new_n8520_, new_n2334_ );
and  ( new_n8800_, new_n8516_, new_n2168_ );
or   ( new_n8801_, new_n8800_, new_n8799_ );
and  ( new_n8802_, new_n8529_, new_n1824_ );
and  ( new_n8803_, new_n8525_, new_n1717_ );
or   ( new_n8804_, new_n8803_, new_n8802_ );
and  ( new_n8805_, new_n8804_, new_n8801_ );
or   ( new_n8806_, new_n8804_, new_n8801_ );
and  ( new_n8807_, new_n8540_, new_n1355_ );
and  ( new_n8808_, new_n8536_, new_n1267_ );
or   ( new_n8809_, new_n8808_, new_n8807_ );
and  ( new_n8810_, new_n8809_, new_n8806_ );
or   ( new_n8811_, new_n8810_, new_n8805_ );
and  ( new_n8812_, new_n8811_, new_n8798_ );
or   ( new_n8813_, new_n8812_, new_n8797_ );
and  ( new_n8814_, new_n8553_, new_n913_ );
and  ( new_n8815_, new_n8549_, new_n938_ );
or   ( new_n8816_, new_n8815_, new_n8814_ );
and  ( new_n8817_, new_n8562_, new_n428_ );
and  ( new_n8818_, new_n8558_, new_n457_ );
or   ( new_n8819_, new_n8818_, new_n8817_ );
and  ( new_n8820_, new_n8819_, new_n8816_ );
or   ( new_n8821_, new_n8819_, new_n8816_ );
and  ( new_n8822_, new_n8573_, new_n505_ );
and  ( new_n8823_, new_n8569_, new_n533_ );
or   ( new_n8824_, new_n8823_, new_n8822_ );
and  ( new_n8825_, new_n8824_, new_n8821_ );
or   ( new_n8826_, new_n8825_, new_n8820_ );
and  ( new_n8827_, new_n8584_, new_n590_ );
and  ( new_n8828_, new_n8580_, new_n619_ );
or   ( new_n8829_, new_n8828_, new_n8827_ );
and  ( new_n8830_, new_n8593_, new_n734_ );
and  ( new_n8831_, new_n8589_, new_n762_ );
or   ( new_n8832_, new_n8831_, new_n8830_ );
and  ( new_n8833_, new_n8832_, new_n8829_ );
or   ( new_n8834_, new_n8832_, new_n8829_ );
and  ( new_n8835_, new_n8604_, new_n785_ );
and  ( new_n8836_, new_n8600_, new_n813_ );
or   ( new_n8837_, new_n8836_, new_n8835_ );
and  ( new_n8838_, new_n8837_, new_n8834_ );
or   ( new_n8839_, new_n8838_, new_n8833_ );
and  ( new_n8840_, new_n8839_, new_n8826_ );
or   ( new_n8841_, new_n8839_, new_n8826_ );
and  ( new_n8842_, new_n8617_, new_n785_ );
and  ( new_n8843_, new_n8613_, new_n813_ );
or   ( new_n8844_, new_n8843_, new_n8842_ );
and  ( new_n8845_, new_n8844_, new_n8841_ );
or   ( new_n8846_, new_n8845_, new_n8840_ );
and  ( new_n8847_, new_n8846_, new_n8813_ );
or   ( new_n8848_, new_n8846_, new_n8813_ );
and  ( new_n8849_, new_n8626_, new_n842_ );
and  ( new_n8850_, new_n8624_, new_n866_ );
or   ( new_n8851_, new_n8850_, new_n8849_ );
and  ( new_n8852_, new_n8633_, new_n8119_ );
and  ( new_n8853_, new_n8629_, new_n8347_ );
or   ( new_n8854_, new_n8853_, new_n8852_ );
and  ( new_n8855_, new_n8854_, new_n8851_ );
or   ( new_n8856_, new_n8854_, new_n8851_ );
and  ( new_n8857_, new_n8642_, new_n8088_ );
and  ( new_n8858_, new_n8638_, new_n8334_ );
or   ( new_n8859_, new_n8858_, new_n8857_ );
and  ( new_n8860_, new_n8859_, new_n8856_ );
or   ( new_n8861_, new_n8860_, new_n8855_ );
and  ( new_n8862_, new_n8861_, new_n8848_ );
or   ( new_n8863_, new_n8862_, new_n8847_ );
and  ( new_n8864_, new_n8653_, new_n7656_ );
and  ( new_n8865_, new_n8649_, new_n7887_ );
or   ( new_n8866_, new_n8865_, new_n8864_ );
and  ( new_n8867_, new_n8660_, new_n8218_ );
and  ( new_n8868_, new_n8656_, new_n8392_ );
or   ( new_n8869_, new_n8868_, new_n8867_ );
and  ( new_n8870_, new_n8667_, new_n8163_ );
and  ( new_n8871_, new_n8663_, new_n8367_ );
or   ( new_n8872_, new_n8871_, new_n8870_ );
and  ( new_n8873_, new_n8872_, new_n8869_ );
or   ( new_n8874_, new_n8872_, new_n8869_ );
and  ( new_n8875_, new_n8676_, new_n8185_ );
and  ( new_n8876_, new_n8672_, new_n8377_ );
or   ( new_n8877_, new_n8876_, new_n8875_ );
and  ( new_n8878_, new_n8877_, new_n8874_ );
or   ( new_n8879_, new_n8878_, new_n8873_ );
and  ( new_n8880_, new_n8879_, new_n8866_ );
or   ( new_n8881_, new_n8879_, new_n8866_ );
and  ( new_n8882_, new_n8687_, new_n7625_ );
and  ( new_n8883_, new_n8683_, new_n7874_ );
or   ( new_n8884_, new_n8883_, new_n8882_ );
and  ( new_n8885_, new_n8884_, new_n8881_ );
or   ( new_n8886_, new_n8885_, new_n8880_ );
and  ( new_n8887_, new_n8886_, new_n8863_ );
or   ( new_n8888_, new_n8886_, new_n8863_ );
and  ( new_n8889_, new_n8698_, new_n8247_ );
and  ( new_n8890_, new_n8694_, new_n8409_ );
or   ( new_n8891_, new_n8890_, new_n8889_ );
and  ( new_n8892_, new_n8705_, new_n8132_ );
and  ( new_n8893_, new_n8701_, new_n8354_ );
or   ( new_n8894_, new_n8893_, new_n8892_ );
and  ( new_n8895_, new_n8894_, new_n8891_ );
or   ( new_n8896_, new_n8894_, new_n8891_ );
and  ( new_n8897_, new_n8714_, new_n8220_ );
and  ( new_n8898_, new_n8710_, new_n8394_ );
or   ( new_n8899_, new_n8898_, new_n8897_ );
and  ( new_n8900_, new_n8899_, new_n8896_ );
or   ( new_n8901_, new_n8900_, new_n8895_ );
and  ( new_n8902_, new_n8901_, new_n8888_ );
or   ( new_n8903_, new_n8902_, new_n8887_ );
and  ( new_n8904_, new_n8418_, new_n8267_ );
and  ( new_n8905_, new_n8421_, new_n8260_ );
or   ( new_n8906_, new_n8905_, new_n8904_ );
and  ( new_n8907_, new_n8727_, new_n8057_ );
and  ( new_n8908_, new_n8723_, new_n8321_ );
or   ( new_n8909_, new_n8908_, new_n8907_ );
and  ( new_n8910_, new_n8909_, new_n8906_ );
or   ( new_n8911_, new_n8909_, new_n8906_ );
and  ( new_n8912_, new_n8736_, new_n8249_ );
and  ( new_n8913_, new_n8732_, new_n8411_ );
or   ( new_n8914_, new_n8913_, new_n8912_ );
and  ( new_n8915_, new_n8914_, new_n8911_ );
or   ( new_n8916_, new_n8915_, new_n8910_ );
and  ( new_n8917_, new_n8916_, new_n8903_ );
or   ( new_n8918_, new_n8916_, new_n8903_ );
and  ( new_n8919_, new_n8747_, new_n8037_ );
and  ( new_n8920_, new_n8743_, new_n8308_ );
or   ( new_n8921_, new_n8920_, new_n8919_ );
and  ( new_n8922_, new_n8921_, new_n8918_ );
or   ( new_n8923_, new_n8922_, new_n8917_ );
and  ( new_n8924_, new_n8923_, new_n8770_ );
or   ( new_n8925_, new_n8924_, new_n8752_ );
and  ( new_n8926_, new_n8925_, new_n8760_ );
and  ( new_n8927_, new_n8923_, new_n8449_ );
and  ( new_n8928_, new_n8770_, new_n8751_ );
or   ( new_n8929_, new_n8928_, new_n8927_ );
and  ( new_n8930_, new_n8758_, new_n8279_ );
and  ( new_n8931_, new_n8754_, new_n8429_ );
or   ( new_n8932_, new_n8931_, new_n8930_ );
and  ( new_n8933_, new_n8932_, new_n8929_ );
or   ( new_n8934_, new_n8933_, new_n8926_ );
or   ( new_n8935_, new_n8415_, new_n8252_ );
and  ( new_n8936_, new_n8935_, new_n8268_ );
and  ( new_n8937_, new_n8413_, new_n8059_ );
and  ( new_n8938_, new_n8323_, new_n8251_ );
or   ( new_n8939_, new_n8938_, new_n8937_ );
and  ( new_n8940_, new_n8939_, new_n8422_ );
or   ( new_n8941_, new_n8940_, new_n8936_ );
or   ( new_n8942_, new_n8880_, new_n8681_ );
and  ( new_n8943_, new_n8942_, new_n8689_ );
and  ( new_n8944_, new_n8879_, new_n8655_ );
and  ( new_n8945_, new_n8866_, new_n8680_ );
or   ( new_n8946_, new_n8945_, new_n8944_ );
and  ( new_n8947_, new_n8946_, new_n8884_ );
or   ( new_n8948_, new_n8947_, new_n8943_ );
or   ( new_n8949_, new_n8847_, new_n8622_ );
and  ( new_n8950_, new_n8949_, new_n8646_ );
and  ( new_n8951_, new_n8813_, new_n8621_ );
and  ( new_n8952_, new_n8846_, new_n8546_ );
or   ( new_n8953_, new_n8952_, new_n8951_ );
and  ( new_n8954_, new_n8953_, new_n8861_ );
or   ( new_n8955_, new_n8954_, new_n8950_ );
or   ( new_n8956_, new_n8955_, new_n8948_ );
or   ( new_n8957_, new_n8873_, new_n8670_ );
and  ( new_n8958_, new_n8957_, new_n8678_ );
and  ( new_n8959_, new_n8869_, new_n8669_ );
and  ( new_n8960_, new_n8872_, new_n8662_ );
or   ( new_n8961_, new_n8960_, new_n8959_ );
and  ( new_n8962_, new_n8961_, new_n8877_ );
or   ( new_n8963_, new_n8962_, new_n8958_ );
or   ( new_n8964_, new_n8855_, new_n8636_ );
and  ( new_n8965_, new_n8964_, new_n8644_ );
and  ( new_n8966_, new_n8851_, new_n8635_ );
and  ( new_n8967_, new_n8854_, new_n8628_ );
or   ( new_n8968_, new_n8967_, new_n8966_ );
and  ( new_n8969_, new_n8968_, new_n8859_ );
or   ( new_n8970_, new_n8969_, new_n8965_ );
and  ( new_n8971_, new_n8970_, new_n8963_ );
or   ( new_n8972_, new_n8970_, new_n8963_ );
or   ( new_n8973_, new_n8840_, new_n8609_ );
and  ( new_n8974_, new_n8973_, new_n8619_ );
and  ( new_n8975_, new_n8826_, new_n8608_ );
and  ( new_n8976_, new_n8839_, new_n8577_ );
or   ( new_n8977_, new_n8976_, new_n8975_ );
and  ( new_n8978_, new_n8977_, new_n8844_ );
or   ( new_n8979_, new_n8978_, new_n8974_ );
and  ( new_n8980_, new_n8979_, new_n8972_ );
or   ( new_n8981_, new_n8980_, new_n8971_ );
or   ( new_n8982_, new_n934_, new_n3924_ );
or   ( new_n8983_, new_n940_, new_n3239_ );
and  ( new_n8984_, new_n8983_, new_n8982_ );
and  ( new_n8985_, new_n8984_, new_n913_ );
and  ( new_n8986_, new_n944_, RI2b1c4342df30_87 );
and  ( new_n8987_, new_n932_, RI2b1c4342deb8_86 );
or   ( new_n8988_, new_n8987_, new_n8986_ );
and  ( new_n8989_, new_n8988_, new_n938_ );
or   ( new_n8990_, new_n8989_, new_n8985_ );
or   ( new_n8991_, new_n1425_, new_n2806_ );
or   ( new_n8992_, new_n1429_, new_n2541_ );
and  ( new_n8993_, new_n8992_, new_n8991_ );
and  ( new_n8994_, new_n8993_, new_n1355_ );
and  ( new_n8995_, new_n1433_, RI2b1c4342de40_85 );
and  ( new_n8996_, new_n1423_, RI2b1c4342ddc8_84 );
or   ( new_n8997_, new_n8996_, new_n8995_ );
and  ( new_n8998_, new_n8997_, new_n1267_ );
or   ( new_n8999_, new_n8998_, new_n8994_ );
and  ( new_n9000_, new_n8999_, new_n8990_ );
or   ( new_n9001_, new_n8999_, new_n8990_ );
or   ( new_n9002_, new_n453_, new_n132_ );
or   ( new_n9003_, new_n459_, new_n3902_ );
and  ( new_n9004_, new_n9003_, new_n9002_ );
and  ( new_n9005_, new_n9004_, new_n428_ );
and  ( new_n9006_, new_n463_, RI2b1c4342e020_89 );
and  ( new_n9007_, new_n451_, RI2b1c4342dfa8_88 );
or   ( new_n9008_, new_n9007_, new_n9006_ );
and  ( new_n9009_, new_n9008_, new_n457_ );
or   ( new_n9010_, new_n9009_, new_n9005_ );
and  ( new_n9011_, new_n9010_, new_n9001_ );
or   ( new_n9012_, new_n9011_, new_n9000_ );
or   ( new_n9013_, new_n524_, new_n117_ );
or   ( new_n9014_, new_n528_, new_n4635_ );
and  ( new_n9015_, new_n9014_, new_n9013_ );
and  ( new_n9016_, new_n9015_, new_n505_ );
and  ( new_n9017_, new_n537_, RI2b1c4342e110_91 );
and  ( new_n9018_, new_n522_, RI2b1c4342e098_90 );
or   ( new_n9019_, new_n9018_, new_n9017_ );
and  ( new_n9020_, new_n9019_, new_n533_ );
or   ( new_n9021_, new_n9020_, new_n9016_ );
or   ( new_n9022_, new_n610_, new_n6307_ );
or   ( new_n9023_, new_n614_, new_n5459_ );
and  ( new_n9024_, new_n9023_, new_n9022_ );
and  ( new_n9025_, new_n9024_, new_n590_ );
and  ( new_n9026_, new_n623_, RI2b1c4342e200_93 );
and  ( new_n9027_, new_n608_, RI2b1c4342e188_92 );
or   ( new_n9028_, new_n9027_, new_n9026_ );
and  ( new_n9029_, new_n9028_, new_n619_ );
or   ( new_n9030_, new_n9029_, new_n9025_ );
and  ( new_n9031_, new_n9030_, new_n9021_ );
or   ( new_n9032_, new_n9030_, new_n9021_ );
or   ( new_n9033_, new_n753_, new_n124_ );
or   ( new_n9034_, new_n757_, new_n6321_ );
and  ( new_n9035_, new_n9034_, new_n9033_ );
and  ( new_n9036_, new_n9035_, new_n734_ );
and  ( new_n9037_, new_n766_, RI2b1c4342e2f0_95 );
and  ( new_n9038_, new_n751_, RI2b1c4342e278_94 );
or   ( new_n9039_, new_n9038_, new_n9037_ );
and  ( new_n9040_, new_n9039_, new_n762_ );
or   ( new_n9041_, new_n9040_, new_n9036_ );
and  ( new_n9042_, new_n9041_, new_n9032_ );
or   ( new_n9043_, new_n9042_, new_n9031_ );
and  ( new_n9044_, new_n9043_, new_n9012_ );
or   ( new_n9045_, new_n9043_, new_n9012_ );
or   ( new_n9046_, new_n8833_, new_n8596_ );
and  ( new_n9047_, new_n9046_, new_n8606_ );
and  ( new_n9048_, new_n8829_, new_n8595_ );
and  ( new_n9049_, new_n8832_, new_n8586_ );
or   ( new_n9050_, new_n9049_, new_n9048_ );
and  ( new_n9051_, new_n9050_, new_n8837_ );
or   ( new_n9052_, new_n9051_, new_n9047_ );
and  ( new_n9053_, new_n9052_, new_n9045_ );
or   ( new_n9054_, new_n9053_, new_n9044_ );
or   ( new_n9055_, new_n5308_, new_n105_ );
or   ( new_n9056_, new_n5312_, new_n806_ );
and  ( new_n9057_, new_n9056_, new_n9055_ );
and  ( new_n9058_, new_n9057_, new_n5182_ );
and  ( new_n9059_, new_n5316_, RI2b1c4342d8a0_73 );
and  ( new_n9060_, new_n5306_, RI2b1c4342d828_72 );
or   ( new_n9061_, new_n9060_, new_n9059_ );
and  ( new_n9062_, new_n9061_, new_n5028_ );
or   ( new_n9063_, new_n9062_, new_n9058_ );
or   ( new_n9064_, new_n4535_, new_n843_ );
or   ( new_n9065_, new_n4539_, new_n859_ );
and  ( new_n9066_, new_n9065_, new_n9064_ );
and  ( new_n9067_, new_n9066_, new_n4400_ );
and  ( new_n9068_, new_n4543_, RI2b1c4342d990_75 );
and  ( new_n9069_, new_n4533_, RI2b1c4342d918_74 );
or   ( new_n9070_, new_n9069_, new_n9068_ );
and  ( new_n9071_, new_n9070_, new_n4215_ );
or   ( new_n9072_, new_n9071_, new_n9067_ );
and  ( new_n9073_, new_n9072_, new_n9063_ );
or   ( new_n9074_, new_n9072_, new_n9063_ );
or   ( new_n9075_, new_n3802_, new_n1004_ );
or   ( new_n9076_, new_n3806_, new_n886_ );
and  ( new_n9077_, new_n9076_, new_n9075_ );
and  ( new_n9078_, new_n9077_, new_n3695_ );
and  ( new_n9079_, new_n3810_, RI2b1c4342da80_77 );
and  ( new_n9080_, new_n3800_, RI2b1c4342da08_76 );
or   ( new_n9081_, new_n9080_, new_n9079_ );
and  ( new_n9082_, new_n9081_, new_n3548_ );
or   ( new_n9083_, new_n9082_, new_n9078_ );
and  ( new_n9084_, new_n9083_, new_n9074_ );
or   ( new_n9085_, new_n9084_, new_n9073_ );
or   ( new_n9086_, new_n7105_, new_n591_ );
or   ( new_n9087_, new_n7099_, new_n612_ );
and  ( new_n9088_, new_n9087_, new_n9086_ );
and  ( new_n9089_, new_n9088_, new_n5858_ );
and  ( new_n9090_, new_n7104_, RI2b1c4342d648_68 );
and  ( new_n9091_, new_n7110_, RI2b1c4342d6c0_69 );
or   ( new_n9092_, new_n9091_, new_n9090_ );
and  ( new_n9093_, new_n9092_, new_n6037_ );
or   ( new_n9094_, new_n9093_, new_n9089_ );
and  ( new_n9095_, new_n9094_, new_n785_ );
or   ( new_n9096_, new_n9094_, new_n785_ );
or   ( new_n9097_, new_n6156_, new_n110_ );
or   ( new_n9098_, new_n6160_, new_n755_ );
and  ( new_n9099_, new_n9098_, new_n9097_ );
and  ( new_n9100_, new_n9099_, new_n6039_ );
and  ( new_n9101_, new_n6164_, RI2b1c4342d7b0_71 );
and  ( new_n9102_, new_n6154_, RI2b1c4342d738_70 );
or   ( new_n9103_, new_n9102_, new_n9101_ );
and  ( new_n9104_, new_n9103_, new_n5867_ );
or   ( new_n9105_, new_n9104_, new_n9100_ );
and  ( new_n9106_, new_n9105_, new_n9096_ );
or   ( new_n9107_, new_n9106_, new_n9095_ );
and  ( new_n9108_, new_n9107_, new_n9085_ );
or   ( new_n9109_, new_n9107_, new_n9085_ );
or   ( new_n9110_, new_n3112_, new_n1310_ );
or   ( new_n9111_, new_n3116_, new_n1002_ );
and  ( new_n9112_, new_n9111_, new_n9110_ );
and  ( new_n9113_, new_n9112_, new_n3004_ );
and  ( new_n9114_, new_n3120_, RI2b1c4342db70_79 );
and  ( new_n9115_, new_n3110_, RI2b1c4342daf8_78 );
or   ( new_n9116_, new_n9115_, new_n9114_ );
and  ( new_n9117_, new_n9116_, new_n2868_ );
or   ( new_n9118_, new_n9117_, new_n9113_ );
or   ( new_n9119_, new_n2450_, new_n126_ );
or   ( new_n9120_, new_n2454_, new_n1511_ );
and  ( new_n9121_, new_n9120_, new_n9119_ );
and  ( new_n9122_, new_n9121_, new_n2334_ );
and  ( new_n9123_, new_n2458_, RI2b1c4342dc60_81 );
and  ( new_n9124_, new_n2448_, RI2b1c4342dbe8_80 );
or   ( new_n9125_, new_n9124_, new_n9123_ );
and  ( new_n9126_, new_n9125_, new_n2168_ );
or   ( new_n9127_, new_n9126_, new_n9122_ );
and  ( new_n9128_, new_n9127_, new_n9118_ );
or   ( new_n9129_, new_n9127_, new_n9118_ );
or   ( new_n9130_, new_n1910_, new_n121_ );
or   ( new_n9131_, new_n1914_, new_n2119_ );
and  ( new_n9132_, new_n9131_, new_n9130_ );
and  ( new_n9133_, new_n9132_, new_n1824_ );
and  ( new_n9134_, new_n1918_, RI2b1c4342dd50_83 );
and  ( new_n9135_, new_n1908_, RI2b1c4342dcd8_82 );
or   ( new_n9136_, new_n9135_, new_n9134_ );
and  ( new_n9137_, new_n9136_, new_n1717_ );
or   ( new_n9138_, new_n9137_, new_n9133_ );
and  ( new_n9139_, new_n9138_, new_n9129_ );
or   ( new_n9140_, new_n9139_, new_n9128_ );
and  ( new_n9141_, new_n9140_, new_n9109_ );
or   ( new_n9142_, new_n9141_, new_n9108_ );
and  ( new_n9143_, new_n9142_, new_n9054_ );
or   ( new_n9144_, new_n9142_, new_n9054_ );
or   ( new_n9145_, new_n8820_, new_n8565_ );
and  ( new_n9146_, new_n9145_, new_n8575_ );
and  ( new_n9147_, new_n8816_, new_n8564_ );
and  ( new_n9148_, new_n8819_, new_n8555_ );
or   ( new_n9149_, new_n9148_, new_n9147_ );
and  ( new_n9150_, new_n9149_, new_n8824_ );
or   ( new_n9151_, new_n9150_, new_n9146_ );
or   ( new_n9152_, new_n8805_, new_n8532_ );
and  ( new_n9153_, new_n9152_, new_n8542_ );
and  ( new_n9154_, new_n8801_, new_n8531_ );
and  ( new_n9155_, new_n8804_, new_n8522_ );
or   ( new_n9156_, new_n9155_, new_n9154_ );
and  ( new_n9157_, new_n9156_, new_n8809_ );
or   ( new_n9158_, new_n9157_, new_n9153_ );
and  ( new_n9159_, new_n9158_, new_n9151_ );
or   ( new_n9160_, new_n9158_, new_n9151_ );
or   ( new_n9161_, new_n8790_, new_n8499_ );
and  ( new_n9162_, new_n9161_, new_n8509_ );
and  ( new_n9163_, new_n8786_, new_n8498_ );
and  ( new_n9164_, new_n8789_, new_n8489_ );
or   ( new_n9165_, new_n9164_, new_n9163_ );
and  ( new_n9166_, new_n9165_, new_n8794_ );
or   ( new_n9167_, new_n9166_, new_n9162_ );
and  ( new_n9168_, new_n9167_, new_n9160_ );
or   ( new_n9169_, new_n9168_, new_n9159_ );
and  ( new_n9170_, new_n9169_, new_n9144_ );
or   ( new_n9171_, new_n9170_, new_n9143_ );
and  ( new_n9172_, new_n9171_, new_n8981_ );
or   ( new_n9173_, new_n9171_, new_n8981_ );
or   ( new_n9174_, new_n8895_, new_n8708_ );
and  ( new_n9175_, new_n9174_, new_n8716_ );
and  ( new_n9176_, new_n8891_, new_n8707_ );
and  ( new_n9177_, new_n8894_, new_n8700_ );
or   ( new_n9178_, new_n9177_, new_n9176_ );
and  ( new_n9179_, new_n9178_, new_n8899_ );
or   ( new_n9180_, new_n9179_, new_n9175_ );
and  ( new_n9181_, new_n9180_, new_n9173_ );
or   ( new_n9182_, new_n9181_, new_n9172_ );
and  ( new_n9183_, new_n9182_, new_n8956_ );
or   ( new_n9184_, new_n9182_, new_n8956_ );
or   ( new_n9185_, new_n8910_, new_n8730_ );
and  ( new_n9186_, new_n9185_, new_n8738_ );
and  ( new_n9187_, new_n8906_, new_n8729_ );
and  ( new_n9188_, new_n8909_, new_n8722_ );
or   ( new_n9189_, new_n9188_, new_n9187_ );
and  ( new_n9190_, new_n9189_, new_n8914_ );
or   ( new_n9191_, new_n9190_, new_n9186_ );
and  ( new_n9192_, new_n9191_, new_n9184_ );
or   ( new_n9193_, new_n9192_, new_n9183_ );
and  ( new_n9194_, new_n9193_, new_n8941_ );
or   ( new_n9195_, new_n9193_, new_n8941_ );
or   ( new_n9196_, new_n8917_, new_n8741_ );
and  ( new_n9197_, new_n9196_, new_n8749_ );
and  ( new_n9198_, new_n8903_, new_n8740_ );
and  ( new_n9199_, new_n8916_, new_n8720_ );
or   ( new_n9200_, new_n9199_, new_n9198_ );
and  ( new_n9201_, new_n9200_, new_n8921_ );
or   ( new_n9202_, new_n9201_, new_n9197_ );
and  ( new_n9203_, new_n9202_, new_n9195_ );
or   ( new_n9204_, new_n9203_, new_n9194_ );
and  ( new_n9205_, new_n9204_, new_n8934_ );
or   ( new_n9206_, new_n9204_, new_n8934_ );
and  ( new_n9207_, new_n8939_, new_n8268_ );
and  ( new_n9208_, new_n8935_, new_n8422_ );
or   ( new_n9209_, new_n9208_, new_n9207_ );
and  ( new_n9210_, new_n8946_, new_n8689_ );
and  ( new_n9211_, new_n8942_, new_n8884_ );
or   ( new_n9212_, new_n9211_, new_n9210_ );
and  ( new_n9213_, new_n8953_, new_n8646_ );
and  ( new_n9214_, new_n8949_, new_n8861_ );
or   ( new_n9215_, new_n9214_, new_n9213_ );
and  ( new_n9216_, new_n9215_, new_n9212_ );
and  ( new_n9217_, new_n8961_, new_n8678_ );
and  ( new_n9218_, new_n8957_, new_n8877_ );
or   ( new_n9219_, new_n9218_, new_n9217_ );
and  ( new_n9220_, new_n8968_, new_n8644_ );
and  ( new_n9221_, new_n8964_, new_n8859_ );
or   ( new_n9222_, new_n9221_, new_n9220_ );
and  ( new_n9223_, new_n9222_, new_n9219_ );
or   ( new_n9224_, new_n9222_, new_n9219_ );
and  ( new_n9225_, new_n8977_, new_n8619_ );
and  ( new_n9226_, new_n8973_, new_n8844_ );
or   ( new_n9227_, new_n9226_, new_n9225_ );
and  ( new_n9228_, new_n9227_, new_n9224_ );
or   ( new_n9229_, new_n9228_, new_n9223_ );
and  ( new_n9230_, new_n8997_, new_n1355_ );
and  ( new_n9231_, new_n8993_, new_n1267_ );
or   ( new_n9232_, new_n9231_, new_n9230_ );
and  ( new_n9233_, new_n8988_, new_n913_ );
and  ( new_n9234_, new_n8984_, new_n938_ );
or   ( new_n9235_, new_n9234_, new_n9233_ );
and  ( new_n9236_, new_n9235_, new_n9232_ );
or   ( new_n9237_, new_n9235_, new_n9232_ );
and  ( new_n9238_, new_n9008_, new_n428_ );
and  ( new_n9239_, new_n9004_, new_n457_ );
or   ( new_n9240_, new_n9239_, new_n9238_ );
and  ( new_n9241_, new_n9240_, new_n9237_ );
or   ( new_n9242_, new_n9241_, new_n9236_ );
and  ( new_n9243_, new_n9019_, new_n505_ );
and  ( new_n9244_, new_n9015_, new_n533_ );
or   ( new_n9245_, new_n9244_, new_n9243_ );
and  ( new_n9246_, new_n9028_, new_n590_ );
and  ( new_n9247_, new_n9024_, new_n619_ );
or   ( new_n9248_, new_n9247_, new_n9246_ );
and  ( new_n9249_, new_n9248_, new_n9245_ );
or   ( new_n9250_, new_n9248_, new_n9245_ );
and  ( new_n9251_, new_n9039_, new_n734_ );
and  ( new_n9252_, new_n9035_, new_n762_ );
or   ( new_n9253_, new_n9252_, new_n9251_ );
and  ( new_n9254_, new_n9253_, new_n9250_ );
or   ( new_n9255_, new_n9254_, new_n9249_ );
and  ( new_n9256_, new_n9255_, new_n9242_ );
or   ( new_n9257_, new_n9255_, new_n9242_ );
and  ( new_n9258_, new_n9050_, new_n8606_ );
and  ( new_n9259_, new_n9046_, new_n8837_ );
or   ( new_n9260_, new_n9259_, new_n9258_ );
and  ( new_n9261_, new_n9260_, new_n9257_ );
or   ( new_n9262_, new_n9261_, new_n9256_ );
and  ( new_n9263_, new_n9061_, new_n5182_ );
and  ( new_n9264_, new_n9057_, new_n5028_ );
or   ( new_n9265_, new_n9264_, new_n9263_ );
and  ( new_n9266_, new_n9070_, new_n4400_ );
and  ( new_n9267_, new_n9066_, new_n4215_ );
or   ( new_n9268_, new_n9267_, new_n9266_ );
and  ( new_n9269_, new_n9268_, new_n9265_ );
or   ( new_n9270_, new_n9268_, new_n9265_ );
and  ( new_n9271_, new_n9081_, new_n3695_ );
and  ( new_n9272_, new_n9077_, new_n3548_ );
or   ( new_n9273_, new_n9272_, new_n9271_ );
and  ( new_n9274_, new_n9273_, new_n9270_ );
or   ( new_n9275_, new_n9274_, new_n9269_ );
and  ( new_n9276_, new_n9092_, new_n5858_ );
and  ( new_n9277_, new_n9088_, new_n6037_ );
or   ( new_n9278_, new_n9277_, new_n9276_ );
or   ( new_n9279_, new_n9278_, new_n813_ );
and  ( new_n9280_, new_n9278_, new_n813_ );
and  ( new_n9281_, new_n9103_, new_n6039_ );
and  ( new_n9282_, new_n9099_, new_n5867_ );
or   ( new_n9283_, new_n9282_, new_n9281_ );
or   ( new_n9284_, new_n9283_, new_n9280_ );
and  ( new_n9285_, new_n9284_, new_n9279_ );
or   ( new_n9286_, new_n9285_, new_n9275_ );
and  ( new_n9287_, new_n9285_, new_n9275_ );
and  ( new_n9288_, new_n9116_, new_n3004_ );
and  ( new_n9289_, new_n9112_, new_n2868_ );
or   ( new_n9290_, new_n9289_, new_n9288_ );
and  ( new_n9291_, new_n9125_, new_n2334_ );
and  ( new_n9292_, new_n9121_, new_n2168_ );
or   ( new_n9293_, new_n9292_, new_n9291_ );
and  ( new_n9294_, new_n9293_, new_n9290_ );
or   ( new_n9295_, new_n9293_, new_n9290_ );
and  ( new_n9296_, new_n9136_, new_n1824_ );
and  ( new_n9297_, new_n9132_, new_n1717_ );
or   ( new_n9298_, new_n9297_, new_n9296_ );
and  ( new_n9299_, new_n9298_, new_n9295_ );
or   ( new_n9300_, new_n9299_, new_n9294_ );
or   ( new_n9301_, new_n9300_, new_n9287_ );
and  ( new_n9302_, new_n9301_, new_n9286_ );
or   ( new_n9303_, new_n9302_, new_n9262_ );
and  ( new_n9304_, new_n9302_, new_n9262_ );
and  ( new_n9305_, new_n9149_, new_n8575_ );
and  ( new_n9306_, new_n9145_, new_n8824_ );
or   ( new_n9307_, new_n9306_, new_n9305_ );
and  ( new_n9308_, new_n9156_, new_n8542_ );
and  ( new_n9309_, new_n9152_, new_n8809_ );
or   ( new_n9310_, new_n9309_, new_n9308_ );
and  ( new_n9311_, new_n9310_, new_n9307_ );
or   ( new_n9312_, new_n9310_, new_n9307_ );
and  ( new_n9313_, new_n9165_, new_n8509_ );
and  ( new_n9314_, new_n9161_, new_n8794_ );
or   ( new_n9315_, new_n9314_, new_n9313_ );
and  ( new_n9316_, new_n9315_, new_n9312_ );
or   ( new_n9317_, new_n9316_, new_n9311_ );
or   ( new_n9318_, new_n9317_, new_n9304_ );
and  ( new_n9319_, new_n9318_, new_n9303_ );
or   ( new_n9320_, new_n9319_, new_n9229_ );
and  ( new_n9321_, new_n9319_, new_n9229_ );
and  ( new_n9322_, new_n9178_, new_n8716_ );
and  ( new_n9323_, new_n9174_, new_n8899_ );
or   ( new_n9324_, new_n9323_, new_n9322_ );
or   ( new_n9325_, new_n9324_, new_n9321_ );
and  ( new_n9326_, new_n9325_, new_n9320_ );
or   ( new_n9327_, new_n9326_, new_n9216_ );
and  ( new_n9328_, new_n9326_, new_n9216_ );
and  ( new_n9329_, new_n9189_, new_n8738_ );
and  ( new_n9330_, new_n9185_, new_n8914_ );
or   ( new_n9331_, new_n9330_, new_n9329_ );
or   ( new_n9332_, new_n9331_, new_n9328_ );
and  ( new_n9333_, new_n9332_, new_n9327_ );
and  ( new_n9334_, new_n9333_, new_n9209_ );
or   ( new_n9335_, new_n9334_, new_n9194_ );
and  ( new_n9336_, new_n9335_, new_n9202_ );
and  ( new_n9337_, new_n9333_, new_n8941_ );
and  ( new_n9338_, new_n9209_, new_n9193_ );
or   ( new_n9339_, new_n9338_, new_n9337_ );
and  ( new_n9340_, new_n9200_, new_n8749_ );
and  ( new_n9341_, new_n9196_, new_n8921_ );
or   ( new_n9342_, new_n9341_, new_n9340_ );
and  ( new_n9343_, new_n9342_, new_n9339_ );
or   ( new_n9344_, new_n9343_, new_n9336_ );
or   ( new_n9345_, new_n8887_, new_n8692_ );
and  ( new_n9346_, new_n9345_, new_n8718_ );
and  ( new_n9347_, new_n8863_, new_n8691_ );
and  ( new_n9348_, new_n8886_, new_n8648_ );
or   ( new_n9349_, new_n9348_, new_n9347_ );
and  ( new_n9350_, new_n9349_, new_n8901_ );
or   ( new_n9351_, new_n9350_, new_n9346_ );
and  ( new_n9352_, new_n8955_, new_n8948_ );
or   ( new_n9353_, new_n9352_, new_n9216_ );
or   ( new_n9354_, new_n9311_, new_n9159_ );
and  ( new_n9355_, new_n9354_, new_n9167_ );
and  ( new_n9356_, new_n9307_, new_n9158_ );
and  ( new_n9357_, new_n9310_, new_n9151_ );
or   ( new_n9358_, new_n9357_, new_n9356_ );
and  ( new_n9359_, new_n9358_, new_n9315_ );
or   ( new_n9360_, new_n9359_, new_n9355_ );
or   ( new_n9361_, new_n8777_, new_n8468_ );
and  ( new_n9362_, new_n9361_, new_n8478_ );
and  ( new_n9363_, new_n8773_, new_n8458_ );
and  ( new_n9364_, new_n8776_, new_n8467_ );
or   ( new_n9365_, new_n9364_, new_n9363_ );
and  ( new_n9366_, new_n9365_, new_n8781_ );
or   ( new_n9367_, new_n9366_, new_n9362_ );
and  ( new_n9368_, new_n9367_, new_n9360_ );
or   ( new_n9369_, new_n9367_, new_n9360_ );
or   ( new_n9370_, new_n9256_, new_n9044_ );
and  ( new_n9371_, new_n9370_, new_n9052_ );
and  ( new_n9372_, new_n9242_, new_n9043_ );
and  ( new_n9373_, new_n9255_, new_n9012_ );
or   ( new_n9374_, new_n9373_, new_n9372_ );
and  ( new_n9375_, new_n9374_, new_n9260_ );
or   ( new_n9376_, new_n9375_, new_n9371_ );
and  ( new_n9377_, new_n9376_, new_n9369_ );
or   ( new_n9378_, new_n9377_, new_n9368_ );
or   ( new_n9379_, new_n808_, new_n7274_ );
and  ( new_n9380_, new_n9379_, new_n785_ );
and  ( new_n9381_, new_n802_, RI2b1c4342e368_96 );
and  ( new_n9382_, new_n9381_, new_n813_ );
or   ( new_n9383_, new_n9382_, new_n9380_ );
or   ( new_n9384_, new_n453_, new_n4635_ );
or   ( new_n9385_, new_n459_, new_n132_ );
and  ( new_n9386_, new_n9385_, new_n9384_ );
and  ( new_n9387_, new_n9386_, new_n428_ );
and  ( new_n9388_, new_n463_, RI2b1c4342e098_90 );
and  ( new_n9389_, new_n451_, RI2b1c4342e020_89 );
or   ( new_n9390_, new_n9389_, new_n9388_ );
and  ( new_n9391_, new_n9390_, new_n457_ );
or   ( new_n9392_, new_n9391_, new_n9387_ );
or   ( new_n9393_, new_n934_, new_n3902_ );
or   ( new_n9394_, new_n940_, new_n3924_ );
and  ( new_n9395_, new_n9394_, new_n9393_ );
and  ( new_n9396_, new_n9395_, new_n913_ );
and  ( new_n9397_, new_n944_, RI2b1c4342dfa8_88 );
and  ( new_n9398_, new_n932_, RI2b1c4342df30_87 );
or   ( new_n9399_, new_n9398_, new_n9397_ );
and  ( new_n9400_, new_n9399_, new_n938_ );
or   ( new_n9401_, new_n9400_, new_n9396_ );
and  ( new_n9402_, new_n9401_, new_n9392_ );
or   ( new_n9403_, new_n9401_, new_n9392_ );
or   ( new_n9404_, new_n524_, new_n5459_ );
or   ( new_n9405_, new_n528_, new_n117_ );
and  ( new_n9406_, new_n9405_, new_n9404_ );
and  ( new_n9407_, new_n9406_, new_n505_ );
and  ( new_n9408_, new_n537_, RI2b1c4342e188_92 );
and  ( new_n9409_, new_n522_, RI2b1c4342e110_91 );
or   ( new_n9410_, new_n9409_, new_n9408_ );
and  ( new_n9411_, new_n9410_, new_n533_ );
or   ( new_n9412_, new_n9411_, new_n9407_ );
and  ( new_n9413_, new_n9412_, new_n9403_ );
or   ( new_n9414_, new_n9413_, new_n9402_ );
and  ( new_n9415_, new_n9414_, new_n9383_ );
or   ( new_n9416_, new_n9414_, new_n9383_ );
or   ( new_n9417_, new_n9249_, new_n9031_ );
and  ( new_n9418_, new_n9417_, new_n9041_ );
and  ( new_n9419_, new_n9245_, new_n9030_ );
and  ( new_n9420_, new_n9248_, new_n9021_ );
or   ( new_n9421_, new_n9420_, new_n9419_ );
and  ( new_n9422_, new_n9421_, new_n9253_ );
or   ( new_n9423_, new_n9422_, new_n9418_ );
and  ( new_n9424_, new_n9423_, new_n9416_ );
or   ( new_n9425_, new_n9424_, new_n9415_ );
or   ( new_n9426_, new_n7105_, new_n755_ );
or   ( new_n9427_, new_n7099_, new_n591_ );
and  ( new_n9428_, new_n9427_, new_n9426_ );
and  ( new_n9429_, new_n9428_, new_n5858_ );
and  ( new_n9430_, new_n7104_, RI2b1c4342d6c0_69 );
and  ( new_n9431_, new_n7110_, RI2b1c4342d738_70 );
or   ( new_n9432_, new_n9431_, new_n9430_ );
and  ( new_n9433_, new_n9432_, new_n6037_ );
or   ( new_n9434_, new_n9433_, new_n9429_ );
or   ( new_n9435_, new_n6156_, new_n806_ );
or   ( new_n9436_, new_n6160_, new_n110_ );
and  ( new_n9437_, new_n9436_, new_n9435_ );
and  ( new_n9438_, new_n9437_, new_n6039_ );
and  ( new_n9439_, new_n6164_, RI2b1c4342d828_72 );
and  ( new_n9440_, new_n6154_, RI2b1c4342d7b0_71 );
or   ( new_n9441_, new_n9440_, new_n9439_ );
and  ( new_n9442_, new_n9441_, new_n5867_ );
or   ( new_n9443_, new_n9442_, new_n9438_ );
and  ( new_n9444_, new_n9443_, new_n9434_ );
or   ( new_n9445_, new_n9443_, new_n9434_ );
or   ( new_n9446_, new_n5308_, new_n859_ );
or   ( new_n9447_, new_n5312_, new_n105_ );
and  ( new_n9448_, new_n9447_, new_n9446_ );
and  ( new_n9449_, new_n9448_, new_n5182_ );
and  ( new_n9450_, new_n5316_, RI2b1c4342d918_74 );
and  ( new_n9451_, new_n5306_, RI2b1c4342d8a0_73 );
or   ( new_n9452_, new_n9451_, new_n9450_ );
and  ( new_n9453_, new_n9452_, new_n5028_ );
or   ( new_n9454_, new_n9453_, new_n9449_ );
and  ( new_n9455_, new_n9454_, new_n9445_ );
or   ( new_n9456_, new_n9455_, new_n9444_ );
or   ( new_n9457_, new_n4535_, new_n886_ );
or   ( new_n9458_, new_n4539_, new_n843_ );
and  ( new_n9459_, new_n9458_, new_n9457_ );
and  ( new_n9460_, new_n9459_, new_n4400_ );
and  ( new_n9461_, new_n4543_, RI2b1c4342da08_76 );
and  ( new_n9462_, new_n4533_, RI2b1c4342d990_75 );
or   ( new_n9463_, new_n9462_, new_n9461_ );
and  ( new_n9464_, new_n9463_, new_n4215_ );
or   ( new_n9465_, new_n9464_, new_n9460_ );
or   ( new_n9466_, new_n3802_, new_n1002_ );
or   ( new_n9467_, new_n3806_, new_n1004_ );
and  ( new_n9468_, new_n9467_, new_n9466_ );
and  ( new_n9469_, new_n9468_, new_n3695_ );
and  ( new_n9470_, new_n3810_, RI2b1c4342daf8_78 );
and  ( new_n9471_, new_n3800_, RI2b1c4342da80_77 );
or   ( new_n9472_, new_n9471_, new_n9470_ );
and  ( new_n9473_, new_n9472_, new_n3548_ );
or   ( new_n9474_, new_n9473_, new_n9469_ );
and  ( new_n9475_, new_n9474_, new_n9465_ );
or   ( new_n9476_, new_n9474_, new_n9465_ );
or   ( new_n9477_, new_n3112_, new_n1511_ );
or   ( new_n9478_, new_n3116_, new_n1310_ );
and  ( new_n9479_, new_n9478_, new_n9477_ );
and  ( new_n9480_, new_n9479_, new_n3004_ );
and  ( new_n9481_, new_n3120_, RI2b1c4342dbe8_80 );
and  ( new_n9482_, new_n3110_, RI2b1c4342db70_79 );
or   ( new_n9483_, new_n9482_, new_n9481_ );
and  ( new_n9484_, new_n9483_, new_n2868_ );
or   ( new_n9485_, new_n9484_, new_n9480_ );
and  ( new_n9486_, new_n9485_, new_n9476_ );
or   ( new_n9487_, new_n9486_, new_n9475_ );
and  ( new_n9488_, new_n9487_, new_n9456_ );
or   ( new_n9489_, new_n9487_, new_n9456_ );
or   ( new_n9490_, new_n2450_, new_n2119_ );
or   ( new_n9491_, new_n2454_, new_n126_ );
and  ( new_n9492_, new_n9491_, new_n9490_ );
and  ( new_n9493_, new_n9492_, new_n2334_ );
and  ( new_n9494_, new_n2458_, RI2b1c4342dcd8_82 );
and  ( new_n9495_, new_n2448_, RI2b1c4342dc60_81 );
or   ( new_n9496_, new_n9495_, new_n9494_ );
and  ( new_n9497_, new_n9496_, new_n2168_ );
or   ( new_n9498_, new_n9497_, new_n9493_ );
or   ( new_n9499_, new_n1910_, new_n2541_ );
or   ( new_n9500_, new_n1914_, new_n121_ );
and  ( new_n9501_, new_n9500_, new_n9499_ );
and  ( new_n9502_, new_n9501_, new_n1824_ );
and  ( new_n9503_, new_n1918_, RI2b1c4342ddc8_84 );
and  ( new_n9504_, new_n1908_, RI2b1c4342dd50_83 );
or   ( new_n9505_, new_n9504_, new_n9503_ );
and  ( new_n9506_, new_n9505_, new_n1717_ );
or   ( new_n9507_, new_n9506_, new_n9502_ );
and  ( new_n9508_, new_n9507_, new_n9498_ );
or   ( new_n9509_, new_n9507_, new_n9498_ );
or   ( new_n9510_, new_n1425_, new_n3239_ );
or   ( new_n9511_, new_n1429_, new_n2806_ );
and  ( new_n9512_, new_n9511_, new_n9510_ );
and  ( new_n9513_, new_n9512_, new_n1355_ );
and  ( new_n9514_, new_n1433_, RI2b1c4342deb8_86 );
and  ( new_n9515_, new_n1423_, RI2b1c4342de40_85 );
or   ( new_n9516_, new_n9515_, new_n9514_ );
and  ( new_n9517_, new_n9516_, new_n1267_ );
or   ( new_n9518_, new_n9517_, new_n9513_ );
and  ( new_n9519_, new_n9518_, new_n9509_ );
or   ( new_n9520_, new_n9519_, new_n9508_ );
and  ( new_n9521_, new_n9520_, new_n9489_ );
or   ( new_n9522_, new_n9521_, new_n9488_ );
and  ( new_n9523_, new_n9522_, new_n9425_ );
or   ( new_n9524_, new_n9522_, new_n9425_ );
or   ( new_n9525_, new_n9294_, new_n9128_ );
and  ( new_n9526_, new_n9525_, new_n9138_ );
and  ( new_n9527_, new_n9290_, new_n9127_ );
and  ( new_n9528_, new_n9293_, new_n9118_ );
or   ( new_n9529_, new_n9528_, new_n9527_ );
and  ( new_n9530_, new_n9529_, new_n9298_ );
or   ( new_n9531_, new_n9530_, new_n9526_ );
or   ( new_n9532_, new_n9236_, new_n9000_ );
and  ( new_n9533_, new_n9532_, new_n9010_ );
and  ( new_n9534_, new_n9232_, new_n8990_ );
and  ( new_n9535_, new_n9235_, new_n8999_ );
or   ( new_n9536_, new_n9535_, new_n9534_ );
and  ( new_n9537_, new_n9536_, new_n9240_ );
or   ( new_n9538_, new_n9537_, new_n9533_ );
and  ( new_n9539_, new_n9538_, new_n9531_ );
or   ( new_n9540_, new_n9538_, new_n9531_ );
or   ( new_n9541_, new_n9269_, new_n9073_ );
and  ( new_n9542_, new_n9541_, new_n9083_ );
and  ( new_n9543_, new_n9265_, new_n9072_ );
and  ( new_n9544_, new_n9268_, new_n9063_ );
or   ( new_n9545_, new_n9544_, new_n9543_ );
and  ( new_n9546_, new_n9545_, new_n9273_ );
or   ( new_n9547_, new_n9546_, new_n9542_ );
and  ( new_n9548_, new_n9547_, new_n9540_ );
or   ( new_n9549_, new_n9548_, new_n9539_ );
and  ( new_n9550_, new_n9549_, new_n9524_ );
or   ( new_n9551_, new_n9550_, new_n9523_ );
and  ( new_n9552_, new_n9551_, new_n9378_ );
or   ( new_n9553_, new_n9551_, new_n9378_ );
or   ( new_n9554_, new_n8797_, new_n8512_ );
and  ( new_n9555_, new_n9554_, new_n8544_ );
and  ( new_n9556_, new_n8783_, new_n8511_ );
and  ( new_n9557_, new_n8796_, new_n8480_ );
or   ( new_n9558_, new_n9557_, new_n9556_ );
and  ( new_n9559_, new_n9558_, new_n8811_ );
or   ( new_n9560_, new_n9559_, new_n9555_ );
and  ( new_n9561_, new_n9560_, new_n9553_ );
or   ( new_n9562_, new_n9561_, new_n9552_ );
and  ( new_n9563_, new_n9562_, new_n9353_ );
or   ( new_n9564_, new_n9562_, new_n9353_ );
or   ( new_n9565_, new_n9321_, new_n9172_ );
and  ( new_n9566_, new_n9565_, new_n9180_ );
and  ( new_n9567_, new_n9319_, new_n8981_ );
and  ( new_n9568_, new_n9229_, new_n9171_ );
or   ( new_n9569_, new_n9568_, new_n9567_ );
and  ( new_n9570_, new_n9569_, new_n9324_ );
or   ( new_n9571_, new_n9570_, new_n9566_ );
and  ( new_n9572_, new_n9571_, new_n9564_ );
or   ( new_n9573_, new_n9572_, new_n9563_ );
and  ( new_n9574_, new_n9573_, new_n9351_ );
or   ( new_n9575_, new_n9573_, new_n9351_ );
or   ( new_n9576_, new_n9328_, new_n9183_ );
and  ( new_n9577_, new_n9576_, new_n9191_ );
and  ( new_n9578_, new_n9326_, new_n8956_ );
and  ( new_n9579_, new_n9216_, new_n9182_ );
or   ( new_n9580_, new_n9579_, new_n9578_ );
and  ( new_n9581_, new_n9580_, new_n9331_ );
or   ( new_n9582_, new_n9581_, new_n9577_ );
and  ( new_n9583_, new_n9582_, new_n9575_ );
or   ( new_n9584_, new_n9583_, new_n9574_ );
or   ( new_n9585_, new_n9584_, new_n9344_ );
and  ( new_n9586_, new_n9585_, new_n9206_ );
or   ( new_n9587_, new_n9586_, new_n9205_ );
or   ( new_n9588_, new_n9587_, new_n8767_ );
and  ( new_n9589_, new_n9588_, new_n8765_ );
and  ( new_n9590_, new_n9584_, new_n9344_ );
or   ( new_n9591_, new_n9590_, new_n9205_ );
or   ( new_n9592_, new_n9591_, new_n8767_ );
and  ( new_n9593_, new_n9349_, new_n8718_ );
and  ( new_n9594_, new_n9345_, new_n8901_ );
or   ( new_n9595_, new_n9594_, new_n9593_ );
and  ( new_n9596_, new_n9212_, new_n8955_ );
and  ( new_n9597_, new_n9215_, new_n8948_ );
or   ( new_n9598_, new_n9597_, new_n9596_ );
and  ( new_n9599_, new_n9432_, new_n5858_ );
and  ( new_n9600_, new_n9428_, new_n6037_ );
or   ( new_n9601_, new_n9600_, new_n9599_ );
and  ( new_n9602_, new_n9441_, new_n6039_ );
and  ( new_n9603_, new_n9437_, new_n5867_ );
or   ( new_n9604_, new_n9603_, new_n9602_ );
and  ( new_n9605_, new_n9604_, new_n9601_ );
or   ( new_n9606_, new_n9604_, new_n9601_ );
and  ( new_n9607_, new_n9452_, new_n5182_ );
and  ( new_n9608_, new_n9448_, new_n5028_ );
or   ( new_n9609_, new_n9608_, new_n9607_ );
and  ( new_n9610_, new_n9609_, new_n9606_ );
or   ( new_n9611_, new_n9610_, new_n9605_ );
and  ( new_n9612_, new_n9463_, new_n4400_ );
and  ( new_n9613_, new_n9459_, new_n4215_ );
or   ( new_n9614_, new_n9613_, new_n9612_ );
and  ( new_n9615_, new_n9472_, new_n3695_ );
and  ( new_n9616_, new_n9468_, new_n3548_ );
or   ( new_n9617_, new_n9616_, new_n9615_ );
and  ( new_n9618_, new_n9617_, new_n9614_ );
or   ( new_n9619_, new_n9617_, new_n9614_ );
and  ( new_n9620_, new_n9483_, new_n3004_ );
and  ( new_n9621_, new_n9479_, new_n2868_ );
or   ( new_n9622_, new_n9621_, new_n9620_ );
and  ( new_n9623_, new_n9622_, new_n9619_ );
or   ( new_n9624_, new_n9623_, new_n9618_ );
and  ( new_n9625_, new_n9624_, new_n9611_ );
or   ( new_n9626_, new_n9624_, new_n9611_ );
and  ( new_n9627_, new_n9496_, new_n2334_ );
and  ( new_n9628_, new_n9492_, new_n2168_ );
or   ( new_n9629_, new_n9628_, new_n9627_ );
and  ( new_n9630_, new_n9505_, new_n1824_ );
and  ( new_n9631_, new_n9501_, new_n1717_ );
or   ( new_n9632_, new_n9631_, new_n9630_ );
and  ( new_n9633_, new_n9632_, new_n9629_ );
or   ( new_n9634_, new_n9632_, new_n9629_ );
and  ( new_n9635_, new_n9516_, new_n1355_ );
and  ( new_n9636_, new_n9512_, new_n1267_ );
or   ( new_n9637_, new_n9636_, new_n9635_ );
and  ( new_n9638_, new_n9637_, new_n9634_ );
or   ( new_n9639_, new_n9638_, new_n9633_ );
and  ( new_n9640_, new_n9639_, new_n9626_ );
or   ( new_n9641_, new_n9640_, new_n9625_ );
and  ( new_n9642_, new_n9381_, new_n785_ );
and  ( new_n9643_, new_n9379_, new_n813_ );
or   ( new_n9644_, new_n9643_, new_n9642_ );
and  ( new_n9645_, new_n9399_, new_n913_ );
and  ( new_n9646_, new_n9395_, new_n938_ );
or   ( new_n9647_, new_n9646_, new_n9645_ );
and  ( new_n9648_, new_n9390_, new_n428_ );
and  ( new_n9649_, new_n9386_, new_n457_ );
or   ( new_n9650_, new_n9649_, new_n9648_ );
and  ( new_n9651_, new_n9650_, new_n9647_ );
or   ( new_n9652_, new_n9650_, new_n9647_ );
and  ( new_n9653_, new_n9410_, new_n505_ );
and  ( new_n9654_, new_n9406_, new_n533_ );
or   ( new_n9655_, new_n9654_, new_n9653_ );
and  ( new_n9656_, new_n9655_, new_n9652_ );
or   ( new_n9657_, new_n9656_, new_n9651_ );
and  ( new_n9658_, new_n9657_, new_n9644_ );
or   ( new_n9659_, new_n9657_, new_n9644_ );
and  ( new_n9660_, new_n9421_, new_n9041_ );
and  ( new_n9661_, new_n9417_, new_n9253_ );
or   ( new_n9662_, new_n9661_, new_n9660_ );
and  ( new_n9663_, new_n9662_, new_n9659_ );
or   ( new_n9664_, new_n9663_, new_n9658_ );
and  ( new_n9665_, new_n9664_, new_n9641_ );
or   ( new_n9666_, new_n9664_, new_n9641_ );
and  ( new_n9667_, new_n9536_, new_n9010_ );
and  ( new_n9668_, new_n9532_, new_n9240_ );
or   ( new_n9669_, new_n9668_, new_n9667_ );
and  ( new_n9670_, new_n9529_, new_n9138_ );
and  ( new_n9671_, new_n9525_, new_n9298_ );
or   ( new_n9672_, new_n9671_, new_n9670_ );
and  ( new_n9673_, new_n9672_, new_n9669_ );
or   ( new_n9674_, new_n9672_, new_n9669_ );
and  ( new_n9675_, new_n9545_, new_n9083_ );
and  ( new_n9676_, new_n9541_, new_n9273_ );
or   ( new_n9677_, new_n9676_, new_n9675_ );
and  ( new_n9678_, new_n9677_, new_n9674_ );
or   ( new_n9679_, new_n9678_, new_n9673_ );
and  ( new_n9680_, new_n9679_, new_n9666_ );
or   ( new_n9681_, new_n9680_, new_n9665_ );
and  ( new_n9682_, new_n9365_, new_n8478_ );
and  ( new_n9683_, new_n9361_, new_n8781_ );
or   ( new_n9684_, new_n9683_, new_n9682_ );
and  ( new_n9685_, new_n9358_, new_n9167_ );
and  ( new_n9686_, new_n9354_, new_n9315_ );
or   ( new_n9687_, new_n9686_, new_n9685_ );
and  ( new_n9688_, new_n9687_, new_n9684_ );
or   ( new_n9689_, new_n9687_, new_n9684_ );
and  ( new_n9690_, new_n9374_, new_n9052_ );
and  ( new_n9691_, new_n9370_, new_n9260_ );
or   ( new_n9692_, new_n9691_, new_n9690_ );
and  ( new_n9693_, new_n9692_, new_n9689_ );
or   ( new_n9694_, new_n9693_, new_n9688_ );
and  ( new_n9695_, new_n9694_, new_n9681_ );
or   ( new_n9696_, new_n9694_, new_n9681_ );
and  ( new_n9697_, new_n9558_, new_n8544_ );
and  ( new_n9698_, new_n9554_, new_n8811_ );
or   ( new_n9699_, new_n9698_, new_n9697_ );
and  ( new_n9700_, new_n9699_, new_n9696_ );
or   ( new_n9701_, new_n9700_, new_n9695_ );
and  ( new_n9702_, new_n9701_, new_n9598_ );
or   ( new_n9703_, new_n9701_, new_n9598_ );
and  ( new_n9704_, new_n9569_, new_n9180_ );
and  ( new_n9705_, new_n9565_, new_n9324_ );
or   ( new_n9706_, new_n9705_, new_n9704_ );
and  ( new_n9707_, new_n9706_, new_n9703_ );
or   ( new_n9708_, new_n9707_, new_n9702_ );
and  ( new_n9709_, new_n9708_, new_n9595_ );
or   ( new_n9710_, new_n9709_, new_n9574_ );
and  ( new_n9711_, new_n9710_, new_n9582_ );
and  ( new_n9712_, new_n9708_, new_n9351_ );
and  ( new_n9713_, new_n9595_, new_n9573_ );
or   ( new_n9714_, new_n9713_, new_n9712_ );
and  ( new_n9715_, new_n9580_, new_n9191_ );
and  ( new_n9716_, new_n9576_, new_n9331_ );
or   ( new_n9717_, new_n9716_, new_n9715_ );
and  ( new_n9718_, new_n9717_, new_n9714_ );
or   ( new_n9719_, new_n9718_, new_n9711_ );
or   ( new_n9720_, new_n9304_, new_n9143_ );
and  ( new_n9721_, new_n9720_, new_n9169_ );
and  ( new_n9722_, new_n9302_, new_n9054_ );
and  ( new_n9723_, new_n9262_, new_n9142_ );
or   ( new_n9724_, new_n9723_, new_n9722_ );
and  ( new_n9725_, new_n9724_, new_n9317_ );
or   ( new_n9726_, new_n9725_, new_n9721_ );
or   ( new_n9727_, new_n9695_, new_n9552_ );
and  ( new_n9728_, new_n9727_, new_n9560_ );
and  ( new_n9729_, new_n9681_, new_n9378_ );
and  ( new_n9730_, new_n9694_, new_n9551_ );
or   ( new_n9731_, new_n9730_, new_n9729_ );
and  ( new_n9732_, new_n9731_, new_n9699_ );
or   ( new_n9733_, new_n9732_, new_n9728_ );
or   ( new_n9734_, new_n9733_, new_n9726_ );
or   ( new_n9735_, new_n9688_, new_n9368_ );
and  ( new_n9736_, new_n9735_, new_n9376_ );
and  ( new_n9737_, new_n9684_, new_n9360_ );
and  ( new_n9738_, new_n9687_, new_n9367_ );
or   ( new_n9739_, new_n9738_, new_n9737_ );
and  ( new_n9740_, new_n9739_, new_n9692_ );
or   ( new_n9741_, new_n9740_, new_n9736_ );
or   ( new_n9742_, new_n9665_, new_n9523_ );
and  ( new_n9743_, new_n9742_, new_n9549_ );
and  ( new_n9744_, new_n9641_, new_n9425_ );
and  ( new_n9745_, new_n9664_, new_n9522_ );
or   ( new_n9746_, new_n9745_, new_n9744_ );
and  ( new_n9747_, new_n9746_, new_n9679_ );
or   ( new_n9748_, new_n9747_, new_n9743_ );
or   ( new_n9749_, new_n9748_, new_n9741_ );
or   ( new_n9750_, new_n9280_, new_n9095_ );
and  ( new_n9751_, new_n9750_, new_n9105_ );
and  ( new_n9752_, new_n9094_, new_n813_ );
and  ( new_n9753_, new_n9278_, new_n785_ );
or   ( new_n9754_, new_n9753_, new_n9752_ );
and  ( new_n9755_, new_n9754_, new_n9283_ );
or   ( new_n9756_, new_n9755_, new_n9751_ );
or   ( new_n9757_, new_n9673_, new_n9539_ );
and  ( new_n9758_, new_n9757_, new_n9547_ );
and  ( new_n9759_, new_n9669_, new_n9531_ );
and  ( new_n9760_, new_n9672_, new_n9538_ );
or   ( new_n9761_, new_n9760_, new_n9759_ );
and  ( new_n9762_, new_n9761_, new_n9677_ );
or   ( new_n9763_, new_n9762_, new_n9758_ );
and  ( new_n9764_, new_n9763_, new_n9756_ );
or   ( new_n9765_, new_n9763_, new_n9756_ );
or   ( new_n9766_, new_n9658_, new_n9415_ );
and  ( new_n9767_, new_n9766_, new_n9423_ );
and  ( new_n9768_, new_n9657_, new_n9383_ );
and  ( new_n9769_, new_n9644_, new_n9414_ );
or   ( new_n9770_, new_n9769_, new_n9768_ );
and  ( new_n9771_, new_n9770_, new_n9662_ );
or   ( new_n9772_, new_n9771_, new_n9767_ );
and  ( new_n9773_, new_n9772_, new_n9765_ );
or   ( new_n9774_, new_n9773_, new_n9764_ );
or   ( new_n9775_, new_n1425_, new_n3924_ );
or   ( new_n9776_, new_n1429_, new_n3239_ );
and  ( new_n9777_, new_n9776_, new_n9775_ );
and  ( new_n9778_, new_n9777_, new_n1355_ );
and  ( new_n9779_, new_n1433_, RI2b1c4342df30_87 );
and  ( new_n9780_, new_n1423_, RI2b1c4342deb8_86 );
or   ( new_n9781_, new_n9780_, new_n9779_ );
and  ( new_n9782_, new_n9781_, new_n1267_ );
or   ( new_n9783_, new_n9782_, new_n9778_ );
or   ( new_n9784_, new_n934_, new_n132_ );
or   ( new_n9785_, new_n940_, new_n3902_ );
and  ( new_n9786_, new_n9785_, new_n9784_ );
and  ( new_n9787_, new_n9786_, new_n913_ );
and  ( new_n9788_, new_n944_, RI2b1c4342e020_89 );
and  ( new_n9789_, new_n932_, RI2b1c4342dfa8_88 );
or   ( new_n9790_, new_n9789_, new_n9788_ );
and  ( new_n9791_, new_n9790_, new_n938_ );
or   ( new_n9792_, new_n9791_, new_n9787_ );
and  ( new_n9793_, new_n9792_, new_n9783_ );
or   ( new_n9794_, new_n9792_, new_n9783_ );
or   ( new_n9795_, new_n453_, new_n117_ );
or   ( new_n9796_, new_n459_, new_n4635_ );
and  ( new_n9797_, new_n9796_, new_n9795_ );
and  ( new_n9798_, new_n9797_, new_n428_ );
and  ( new_n9799_, new_n463_, RI2b1c4342e110_91 );
and  ( new_n9800_, new_n451_, RI2b1c4342e098_90 );
or   ( new_n9801_, new_n9800_, new_n9799_ );
and  ( new_n9802_, new_n9801_, new_n457_ );
or   ( new_n9803_, new_n9802_, new_n9798_ );
and  ( new_n9804_, new_n9803_, new_n9794_ );
or   ( new_n9805_, new_n9804_, new_n9793_ );
or   ( new_n9806_, new_n524_, new_n6307_ );
or   ( new_n9807_, new_n528_, new_n5459_ );
and  ( new_n9808_, new_n9807_, new_n9806_ );
and  ( new_n9809_, new_n9808_, new_n505_ );
and  ( new_n9810_, new_n537_, RI2b1c4342e200_93 );
and  ( new_n9811_, new_n522_, RI2b1c4342e188_92 );
or   ( new_n9812_, new_n9811_, new_n9810_ );
and  ( new_n9813_, new_n9812_, new_n533_ );
or   ( new_n9814_, new_n9813_, new_n9809_ );
or   ( new_n9815_, new_n610_, new_n124_ );
or   ( new_n9816_, new_n614_, new_n6321_ );
and  ( new_n9817_, new_n9816_, new_n9815_ );
and  ( new_n9818_, new_n9817_, new_n590_ );
and  ( new_n9819_, new_n623_, RI2b1c4342e2f0_95 );
and  ( new_n9820_, new_n608_, RI2b1c4342e278_94 );
or   ( new_n9821_, new_n9820_, new_n9819_ );
and  ( new_n9822_, new_n9821_, new_n619_ );
or   ( new_n9823_, new_n9822_, new_n9818_ );
and  ( new_n9824_, new_n9823_, new_n9814_ );
or   ( new_n9825_, new_n9823_, new_n9814_ );
or   ( new_n9826_, new_n757_, new_n7274_ );
and  ( new_n9827_, new_n9826_, new_n734_ );
and  ( new_n9828_, new_n751_, RI2b1c4342e368_96 );
and  ( new_n9829_, new_n9828_, new_n762_ );
or   ( new_n9830_, new_n9829_, new_n9827_ );
and  ( new_n9831_, new_n9830_, new_n9825_ );
or   ( new_n9832_, new_n9831_, new_n9824_ );
and  ( new_n9833_, new_n9832_, new_n9805_ );
or   ( new_n9834_, new_n9832_, new_n9805_ );
or   ( new_n9835_, new_n610_, new_n6321_ );
or   ( new_n9836_, new_n614_, new_n6307_ );
and  ( new_n9837_, new_n9836_, new_n9835_ );
and  ( new_n9838_, new_n9837_, new_n590_ );
and  ( new_n9839_, new_n623_, RI2b1c4342e278_94 );
and  ( new_n9840_, new_n608_, RI2b1c4342e200_93 );
or   ( new_n9841_, new_n9840_, new_n9839_ );
and  ( new_n9842_, new_n9841_, new_n619_ );
or   ( new_n9843_, new_n9842_, new_n9838_ );
and  ( new_n9844_, new_n9843_, new_n9834_ );
or   ( new_n9845_, new_n9844_, new_n9833_ );
or   ( new_n9846_, new_n5308_, new_n843_ );
or   ( new_n9847_, new_n5312_, new_n859_ );
and  ( new_n9848_, new_n9847_, new_n9846_ );
and  ( new_n9849_, new_n9848_, new_n5182_ );
and  ( new_n9850_, new_n5316_, RI2b1c4342d990_75 );
and  ( new_n9851_, new_n5306_, RI2b1c4342d918_74 );
or   ( new_n9852_, new_n9851_, new_n9850_ );
and  ( new_n9853_, new_n9852_, new_n5028_ );
or   ( new_n9854_, new_n9853_, new_n9849_ );
or   ( new_n9855_, new_n4535_, new_n1004_ );
or   ( new_n9856_, new_n4539_, new_n886_ );
and  ( new_n9857_, new_n9856_, new_n9855_ );
and  ( new_n9858_, new_n9857_, new_n4400_ );
and  ( new_n9859_, new_n4543_, RI2b1c4342da80_77 );
and  ( new_n9860_, new_n4533_, RI2b1c4342da08_76 );
or   ( new_n9861_, new_n9860_, new_n9859_ );
and  ( new_n9862_, new_n9861_, new_n4215_ );
or   ( new_n9863_, new_n9862_, new_n9858_ );
and  ( new_n9864_, new_n9863_, new_n9854_ );
or   ( new_n9865_, new_n9863_, new_n9854_ );
or   ( new_n9866_, new_n3802_, new_n1310_ );
or   ( new_n9867_, new_n3806_, new_n1002_ );
and  ( new_n9868_, new_n9867_, new_n9866_ );
and  ( new_n9869_, new_n9868_, new_n3695_ );
and  ( new_n9870_, new_n3810_, RI2b1c4342db70_79 );
and  ( new_n9871_, new_n3800_, RI2b1c4342daf8_78 );
or   ( new_n9872_, new_n9871_, new_n9870_ );
and  ( new_n9873_, new_n9872_, new_n3548_ );
or   ( new_n9874_, new_n9873_, new_n9869_ );
and  ( new_n9875_, new_n9874_, new_n9865_ );
or   ( new_n9876_, new_n9875_, new_n9864_ );
or   ( new_n9877_, new_n7105_, new_n110_ );
or   ( new_n9878_, new_n7099_, new_n755_ );
and  ( new_n9879_, new_n9878_, new_n9877_ );
and  ( new_n9880_, new_n9879_, new_n5858_ );
and  ( new_n9881_, new_n7104_, RI2b1c4342d738_70 );
and  ( new_n9882_, new_n7110_, RI2b1c4342d7b0_71 );
or   ( new_n9883_, new_n9882_, new_n9881_ );
and  ( new_n9884_, new_n9883_, new_n6037_ );
or   ( new_n9885_, new_n9884_, new_n9880_ );
and  ( new_n9886_, new_n9885_, new_n734_ );
or   ( new_n9887_, new_n9885_, new_n734_ );
or   ( new_n9888_, new_n6156_, new_n105_ );
or   ( new_n9889_, new_n6160_, new_n806_ );
and  ( new_n9890_, new_n9889_, new_n9888_ );
and  ( new_n9891_, new_n9890_, new_n6039_ );
and  ( new_n9892_, new_n6164_, RI2b1c4342d8a0_73 );
and  ( new_n9893_, new_n6154_, RI2b1c4342d828_72 );
or   ( new_n9894_, new_n9893_, new_n9892_ );
and  ( new_n9895_, new_n9894_, new_n5867_ );
or   ( new_n9896_, new_n9895_, new_n9891_ );
and  ( new_n9897_, new_n9896_, new_n9887_ );
or   ( new_n9898_, new_n9897_, new_n9886_ );
and  ( new_n9899_, new_n9898_, new_n9876_ );
or   ( new_n9900_, new_n9898_, new_n9876_ );
or   ( new_n9901_, new_n3112_, new_n126_ );
or   ( new_n9902_, new_n3116_, new_n1511_ );
and  ( new_n9903_, new_n9902_, new_n9901_ );
and  ( new_n9904_, new_n9903_, new_n3004_ );
and  ( new_n9905_, new_n3120_, RI2b1c4342dc60_81 );
and  ( new_n9906_, new_n3110_, RI2b1c4342dbe8_80 );
or   ( new_n9907_, new_n9906_, new_n9905_ );
and  ( new_n9908_, new_n9907_, new_n2868_ );
or   ( new_n9909_, new_n9908_, new_n9904_ );
or   ( new_n9910_, new_n2450_, new_n121_ );
or   ( new_n9911_, new_n2454_, new_n2119_ );
and  ( new_n9912_, new_n9911_, new_n9910_ );
and  ( new_n9913_, new_n9912_, new_n2334_ );
and  ( new_n9914_, new_n2458_, RI2b1c4342dd50_83 );
and  ( new_n9915_, new_n2448_, RI2b1c4342dcd8_82 );
or   ( new_n9916_, new_n9915_, new_n9914_ );
and  ( new_n9917_, new_n9916_, new_n2168_ );
or   ( new_n9918_, new_n9917_, new_n9913_ );
and  ( new_n9919_, new_n9918_, new_n9909_ );
or   ( new_n9920_, new_n9918_, new_n9909_ );
or   ( new_n9921_, new_n1910_, new_n2806_ );
or   ( new_n9922_, new_n1914_, new_n2541_ );
and  ( new_n9923_, new_n9922_, new_n9921_ );
and  ( new_n9924_, new_n9923_, new_n1824_ );
and  ( new_n9925_, new_n1918_, RI2b1c4342de40_85 );
and  ( new_n9926_, new_n1908_, RI2b1c4342ddc8_84 );
or   ( new_n9927_, new_n9926_, new_n9925_ );
and  ( new_n9928_, new_n9927_, new_n1717_ );
or   ( new_n9929_, new_n9928_, new_n9924_ );
and  ( new_n9930_, new_n9929_, new_n9920_ );
or   ( new_n9931_, new_n9930_, new_n9919_ );
and  ( new_n9932_, new_n9931_, new_n9900_ );
or   ( new_n9933_, new_n9932_, new_n9899_ );
and  ( new_n9934_, new_n9933_, new_n9845_ );
or   ( new_n9935_, new_n9933_, new_n9845_ );
or   ( new_n9936_, new_n753_, new_n7274_ );
or   ( new_n9937_, new_n757_, new_n124_ );
and  ( new_n9938_, new_n9937_, new_n9936_ );
and  ( new_n9939_, new_n9938_, new_n734_ );
and  ( new_n9940_, new_n766_, RI2b1c4342e368_96 );
and  ( new_n9941_, new_n751_, RI2b1c4342e2f0_95 );
or   ( new_n9942_, new_n9941_, new_n9940_ );
and  ( new_n9943_, new_n9942_, new_n762_ );
or   ( new_n9944_, new_n9943_, new_n9939_ );
or   ( new_n9945_, new_n9651_, new_n9402_ );
and  ( new_n9946_, new_n9945_, new_n9412_ );
and  ( new_n9947_, new_n9647_, new_n9392_ );
and  ( new_n9948_, new_n9650_, new_n9401_ );
or   ( new_n9949_, new_n9948_, new_n9947_ );
and  ( new_n9950_, new_n9949_, new_n9655_ );
or   ( new_n9951_, new_n9950_, new_n9946_ );
and  ( new_n9952_, new_n9951_, new_n9944_ );
or   ( new_n9953_, new_n9951_, new_n9944_ );
or   ( new_n9954_, new_n9633_, new_n9508_ );
and  ( new_n9955_, new_n9954_, new_n9518_ );
and  ( new_n9956_, new_n9629_, new_n9507_ );
and  ( new_n9957_, new_n9632_, new_n9498_ );
or   ( new_n9958_, new_n9957_, new_n9956_ );
and  ( new_n9959_, new_n9958_, new_n9637_ );
or   ( new_n9960_, new_n9959_, new_n9955_ );
and  ( new_n9961_, new_n9960_, new_n9953_ );
or   ( new_n9962_, new_n9961_, new_n9952_ );
and  ( new_n9963_, new_n9962_, new_n9935_ );
or   ( new_n9964_, new_n9963_, new_n9934_ );
and  ( new_n9965_, new_n9964_, new_n9774_ );
or   ( new_n9966_, new_n9964_, new_n9774_ );
or   ( new_n9967_, new_n9287_, new_n9108_ );
and  ( new_n9968_, new_n9967_, new_n9140_ );
and  ( new_n9969_, new_n9285_, new_n9085_ );
and  ( new_n9970_, new_n9275_, new_n9107_ );
or   ( new_n9971_, new_n9970_, new_n9969_ );
and  ( new_n9972_, new_n9971_, new_n9300_ );
or   ( new_n9973_, new_n9972_, new_n9968_ );
and  ( new_n9974_, new_n9973_, new_n9966_ );
or   ( new_n9975_, new_n9974_, new_n9965_ );
and  ( new_n9976_, new_n9975_, new_n9749_ );
or   ( new_n9977_, new_n9975_, new_n9749_ );
or   ( new_n9978_, new_n9223_, new_n8971_ );
and  ( new_n9979_, new_n9978_, new_n8979_ );
and  ( new_n9980_, new_n9219_, new_n8970_ );
and  ( new_n9981_, new_n9222_, new_n8963_ );
or   ( new_n9982_, new_n9981_, new_n9980_ );
and  ( new_n9983_, new_n9982_, new_n9227_ );
or   ( new_n9984_, new_n9983_, new_n9979_ );
and  ( new_n9985_, new_n9984_, new_n9977_ );
or   ( new_n9986_, new_n9985_, new_n9976_ );
and  ( new_n9987_, new_n9986_, new_n9734_ );
or   ( new_n9988_, new_n9986_, new_n9734_ );
or   ( new_n9989_, new_n9702_, new_n9563_ );
and  ( new_n9990_, new_n9989_, new_n9571_ );
and  ( new_n9991_, new_n9701_, new_n9353_ );
and  ( new_n9992_, new_n9598_, new_n9562_ );
or   ( new_n9993_, new_n9992_, new_n9991_ );
and  ( new_n9994_, new_n9993_, new_n9706_ );
or   ( new_n9995_, new_n9994_, new_n9990_ );
and  ( new_n9996_, new_n9995_, new_n9988_ );
or   ( new_n9997_, new_n9996_, new_n9987_ );
and  ( new_n9998_, new_n9997_, new_n9719_ );
or   ( new_n9999_, new_n9997_, new_n9719_ );
and  ( new_n10000_, new_n9724_, new_n9169_ );
and  ( new_n10001_, new_n9720_, new_n9317_ );
or   ( new_n10002_, new_n10001_, new_n10000_ );
and  ( new_n10003_, new_n9731_, new_n9560_ );
and  ( new_n10004_, new_n9727_, new_n9699_ );
or   ( new_n10005_, new_n10004_, new_n10003_ );
and  ( new_n10006_, new_n10005_, new_n10002_ );
and  ( new_n10007_, new_n9739_, new_n9376_ );
and  ( new_n10008_, new_n9735_, new_n9692_ );
or   ( new_n10009_, new_n10008_, new_n10007_ );
and  ( new_n10010_, new_n9746_, new_n9549_ );
and  ( new_n10011_, new_n9742_, new_n9679_ );
or   ( new_n10012_, new_n10011_, new_n10010_ );
and  ( new_n10013_, new_n10012_, new_n10009_ );
and  ( new_n10014_, new_n9754_, new_n9105_ );
and  ( new_n10015_, new_n9750_, new_n9283_ );
or   ( new_n10016_, new_n10015_, new_n10014_ );
and  ( new_n10017_, new_n9761_, new_n9547_ );
and  ( new_n10018_, new_n9757_, new_n9677_ );
or   ( new_n10019_, new_n10018_, new_n10017_ );
and  ( new_n10020_, new_n10019_, new_n10016_ );
or   ( new_n10021_, new_n10019_, new_n10016_ );
and  ( new_n10022_, new_n9770_, new_n9423_ );
and  ( new_n10023_, new_n9766_, new_n9662_ );
or   ( new_n10024_, new_n10023_, new_n10022_ );
and  ( new_n10025_, new_n10024_, new_n10021_ );
or   ( new_n10026_, new_n10025_, new_n10020_ );
and  ( new_n10027_, new_n9781_, new_n1355_ );
and  ( new_n10028_, new_n9777_, new_n1267_ );
or   ( new_n10029_, new_n10028_, new_n10027_ );
and  ( new_n10030_, new_n9790_, new_n913_ );
and  ( new_n10031_, new_n9786_, new_n938_ );
or   ( new_n10032_, new_n10031_, new_n10030_ );
and  ( new_n10033_, new_n10032_, new_n10029_ );
or   ( new_n10034_, new_n10032_, new_n10029_ );
and  ( new_n10035_, new_n9801_, new_n428_ );
and  ( new_n10036_, new_n9797_, new_n457_ );
or   ( new_n10037_, new_n10036_, new_n10035_ );
and  ( new_n10038_, new_n10037_, new_n10034_ );
or   ( new_n10039_, new_n10038_, new_n10033_ );
and  ( new_n10040_, new_n9812_, new_n505_ );
and  ( new_n10041_, new_n9808_, new_n533_ );
or   ( new_n10042_, new_n10041_, new_n10040_ );
and  ( new_n10043_, new_n9821_, new_n590_ );
and  ( new_n10044_, new_n9817_, new_n619_ );
or   ( new_n10045_, new_n10044_, new_n10043_ );
and  ( new_n10046_, new_n10045_, new_n10042_ );
or   ( new_n10047_, new_n10045_, new_n10042_ );
and  ( new_n10048_, new_n9828_, new_n734_ );
and  ( new_n10049_, new_n9826_, new_n762_ );
or   ( new_n10050_, new_n10049_, new_n10048_ );
and  ( new_n10051_, new_n10050_, new_n10047_ );
or   ( new_n10052_, new_n10051_, new_n10046_ );
and  ( new_n10053_, new_n10052_, new_n10039_ );
or   ( new_n10054_, new_n10052_, new_n10039_ );
and  ( new_n10055_, new_n9841_, new_n590_ );
and  ( new_n10056_, new_n9837_, new_n619_ );
or   ( new_n10057_, new_n10056_, new_n10055_ );
and  ( new_n10058_, new_n10057_, new_n10054_ );
or   ( new_n10059_, new_n10058_, new_n10053_ );
and  ( new_n10060_, new_n9852_, new_n5182_ );
and  ( new_n10061_, new_n9848_, new_n5028_ );
or   ( new_n10062_, new_n10061_, new_n10060_ );
and  ( new_n10063_, new_n9861_, new_n4400_ );
and  ( new_n10064_, new_n9857_, new_n4215_ );
or   ( new_n10065_, new_n10064_, new_n10063_ );
and  ( new_n10066_, new_n10065_, new_n10062_ );
or   ( new_n10067_, new_n10065_, new_n10062_ );
and  ( new_n10068_, new_n9872_, new_n3695_ );
and  ( new_n10069_, new_n9868_, new_n3548_ );
or   ( new_n10070_, new_n10069_, new_n10068_ );
and  ( new_n10071_, new_n10070_, new_n10067_ );
or   ( new_n10072_, new_n10071_, new_n10066_ );
and  ( new_n10073_, new_n9883_, new_n5858_ );
and  ( new_n10074_, new_n9879_, new_n6037_ );
or   ( new_n10075_, new_n10074_, new_n10073_ );
or   ( new_n10076_, new_n10075_, new_n762_ );
and  ( new_n10077_, new_n10075_, new_n762_ );
and  ( new_n10078_, new_n9894_, new_n6039_ );
and  ( new_n10079_, new_n9890_, new_n5867_ );
or   ( new_n10080_, new_n10079_, new_n10078_ );
or   ( new_n10081_, new_n10080_, new_n10077_ );
and  ( new_n10082_, new_n10081_, new_n10076_ );
or   ( new_n10083_, new_n10082_, new_n10072_ );
and  ( new_n10084_, new_n10082_, new_n10072_ );
and  ( new_n10085_, new_n9907_, new_n3004_ );
and  ( new_n10086_, new_n9903_, new_n2868_ );
or   ( new_n10087_, new_n10086_, new_n10085_ );
and  ( new_n10088_, new_n9916_, new_n2334_ );
and  ( new_n10089_, new_n9912_, new_n2168_ );
or   ( new_n10090_, new_n10089_, new_n10088_ );
and  ( new_n10091_, new_n10090_, new_n10087_ );
or   ( new_n10092_, new_n10090_, new_n10087_ );
and  ( new_n10093_, new_n9927_, new_n1824_ );
and  ( new_n10094_, new_n9923_, new_n1717_ );
or   ( new_n10095_, new_n10094_, new_n10093_ );
and  ( new_n10096_, new_n10095_, new_n10092_ );
or   ( new_n10097_, new_n10096_, new_n10091_ );
or   ( new_n10098_, new_n10097_, new_n10084_ );
and  ( new_n10099_, new_n10098_, new_n10083_ );
or   ( new_n10100_, new_n10099_, new_n10059_ );
and  ( new_n10101_, new_n10099_, new_n10059_ );
and  ( new_n10102_, new_n9942_, new_n734_ );
and  ( new_n10103_, new_n9938_, new_n762_ );
or   ( new_n10104_, new_n10103_, new_n10102_ );
and  ( new_n10105_, new_n9949_, new_n9412_ );
and  ( new_n10106_, new_n9945_, new_n9655_ );
or   ( new_n10107_, new_n10106_, new_n10105_ );
and  ( new_n10108_, new_n10107_, new_n10104_ );
or   ( new_n10109_, new_n10107_, new_n10104_ );
and  ( new_n10110_, new_n9958_, new_n9518_ );
and  ( new_n10111_, new_n9954_, new_n9637_ );
or   ( new_n10112_, new_n10111_, new_n10110_ );
and  ( new_n10113_, new_n10112_, new_n10109_ );
or   ( new_n10114_, new_n10113_, new_n10108_ );
or   ( new_n10115_, new_n10114_, new_n10101_ );
and  ( new_n10116_, new_n10115_, new_n10100_ );
or   ( new_n10117_, new_n10116_, new_n10026_ );
and  ( new_n10118_, new_n10116_, new_n10026_ );
and  ( new_n10119_, new_n9971_, new_n9140_ );
and  ( new_n10120_, new_n9967_, new_n9300_ );
or   ( new_n10121_, new_n10120_, new_n10119_ );
or   ( new_n10122_, new_n10121_, new_n10118_ );
and  ( new_n10123_, new_n10122_, new_n10117_ );
or   ( new_n10124_, new_n10123_, new_n10013_ );
and  ( new_n10125_, new_n10123_, new_n10013_ );
and  ( new_n10126_, new_n9982_, new_n8979_ );
and  ( new_n10127_, new_n9978_, new_n9227_ );
or   ( new_n10128_, new_n10127_, new_n10126_ );
or   ( new_n10129_, new_n10128_, new_n10125_ );
and  ( new_n10130_, new_n10129_, new_n10124_ );
and  ( new_n10131_, new_n10130_, new_n10006_ );
or   ( new_n10132_, new_n10131_, new_n9987_ );
and  ( new_n10133_, new_n10132_, new_n9995_ );
and  ( new_n10134_, new_n10130_, new_n9734_ );
and  ( new_n10135_, new_n10006_, new_n9986_ );
or   ( new_n10136_, new_n10135_, new_n10134_ );
and  ( new_n10137_, new_n9993_, new_n9571_ );
and  ( new_n10138_, new_n9989_, new_n9706_ );
or   ( new_n10139_, new_n10138_, new_n10137_ );
and  ( new_n10140_, new_n10139_, new_n10136_ );
or   ( new_n10141_, new_n10140_, new_n10133_ );
and  ( new_n10142_, new_n9733_, new_n9726_ );
or   ( new_n10143_, new_n10142_, new_n10006_ );
and  ( new_n10144_, new_n9748_, new_n9741_ );
or   ( new_n10145_, new_n10144_, new_n10013_ );
or   ( new_n10146_, new_n7105_, new_n806_ );
or   ( new_n10147_, new_n7099_, new_n110_ );
and  ( new_n10148_, new_n10147_, new_n10146_ );
and  ( new_n10149_, new_n10148_, new_n5858_ );
and  ( new_n10150_, new_n7104_, RI2b1c4342d7b0_71 );
and  ( new_n10151_, new_n7110_, RI2b1c4342d828_72 );
or   ( new_n10152_, new_n10151_, new_n10150_ );
and  ( new_n10153_, new_n10152_, new_n6037_ );
or   ( new_n10154_, new_n10153_, new_n10149_ );
or   ( new_n10155_, new_n6156_, new_n859_ );
or   ( new_n10156_, new_n6160_, new_n105_ );
and  ( new_n10157_, new_n10156_, new_n10155_ );
and  ( new_n10158_, new_n10157_, new_n6039_ );
and  ( new_n10159_, new_n6164_, RI2b1c4342d918_74 );
and  ( new_n10160_, new_n6154_, RI2b1c4342d8a0_73 );
or   ( new_n10161_, new_n10160_, new_n10159_ );
and  ( new_n10162_, new_n10161_, new_n5867_ );
or   ( new_n10163_, new_n10162_, new_n10158_ );
and  ( new_n10164_, new_n10163_, new_n10154_ );
or   ( new_n10165_, new_n10163_, new_n10154_ );
or   ( new_n10166_, new_n5308_, new_n886_ );
or   ( new_n10167_, new_n5312_, new_n843_ );
and  ( new_n10168_, new_n10167_, new_n10166_ );
and  ( new_n10169_, new_n10168_, new_n5182_ );
and  ( new_n10170_, new_n5316_, RI2b1c4342da08_76 );
and  ( new_n10171_, new_n5306_, RI2b1c4342d990_75 );
or   ( new_n10172_, new_n10171_, new_n10170_ );
and  ( new_n10173_, new_n10172_, new_n5028_ );
or   ( new_n10174_, new_n10173_, new_n10169_ );
and  ( new_n10175_, new_n10174_, new_n10165_ );
or   ( new_n10176_, new_n10175_, new_n10164_ );
or   ( new_n10177_, new_n4535_, new_n1002_ );
or   ( new_n10178_, new_n4539_, new_n1004_ );
and  ( new_n10179_, new_n10178_, new_n10177_ );
and  ( new_n10180_, new_n10179_, new_n4400_ );
and  ( new_n10181_, new_n4543_, RI2b1c4342daf8_78 );
and  ( new_n10182_, new_n4533_, RI2b1c4342da80_77 );
or   ( new_n10183_, new_n10182_, new_n10181_ );
and  ( new_n10184_, new_n10183_, new_n4215_ );
or   ( new_n10185_, new_n10184_, new_n10180_ );
or   ( new_n10186_, new_n3802_, new_n1511_ );
or   ( new_n10187_, new_n3806_, new_n1310_ );
and  ( new_n10188_, new_n10187_, new_n10186_ );
and  ( new_n10189_, new_n10188_, new_n3695_ );
and  ( new_n10190_, new_n3810_, RI2b1c4342dbe8_80 );
and  ( new_n10191_, new_n3800_, RI2b1c4342db70_79 );
or   ( new_n10192_, new_n10191_, new_n10190_ );
and  ( new_n10193_, new_n10192_, new_n3548_ );
or   ( new_n10194_, new_n10193_, new_n10189_ );
and  ( new_n10195_, new_n10194_, new_n10185_ );
or   ( new_n10196_, new_n10194_, new_n10185_ );
or   ( new_n10197_, new_n3112_, new_n2119_ );
or   ( new_n10198_, new_n3116_, new_n126_ );
and  ( new_n10199_, new_n10198_, new_n10197_ );
and  ( new_n10200_, new_n10199_, new_n3004_ );
and  ( new_n10201_, new_n3120_, RI2b1c4342dcd8_82 );
and  ( new_n10202_, new_n3110_, RI2b1c4342dc60_81 );
or   ( new_n10203_, new_n10202_, new_n10201_ );
and  ( new_n10204_, new_n10203_, new_n2868_ );
or   ( new_n10205_, new_n10204_, new_n10200_ );
and  ( new_n10206_, new_n10205_, new_n10196_ );
or   ( new_n10207_, new_n10206_, new_n10195_ );
and  ( new_n10208_, new_n10207_, new_n10176_ );
or   ( new_n10209_, new_n10207_, new_n10176_ );
or   ( new_n10210_, new_n2450_, new_n2541_ );
or   ( new_n10211_, new_n2454_, new_n121_ );
and  ( new_n10212_, new_n10211_, new_n10210_ );
and  ( new_n10213_, new_n10212_, new_n2334_ );
and  ( new_n10214_, new_n2458_, RI2b1c4342ddc8_84 );
and  ( new_n10215_, new_n2448_, RI2b1c4342dd50_83 );
or   ( new_n10216_, new_n10215_, new_n10214_ );
and  ( new_n10217_, new_n10216_, new_n2168_ );
or   ( new_n10218_, new_n10217_, new_n10213_ );
or   ( new_n10219_, new_n1910_, new_n3239_ );
or   ( new_n10220_, new_n1914_, new_n2806_ );
and  ( new_n10221_, new_n10220_, new_n10219_ );
and  ( new_n10222_, new_n10221_, new_n1824_ );
and  ( new_n10223_, new_n1918_, RI2b1c4342deb8_86 );
and  ( new_n10224_, new_n1908_, RI2b1c4342de40_85 );
or   ( new_n10225_, new_n10224_, new_n10223_ );
and  ( new_n10226_, new_n10225_, new_n1717_ );
or   ( new_n10227_, new_n10226_, new_n10222_ );
and  ( new_n10228_, new_n10227_, new_n10218_ );
or   ( new_n10229_, new_n10227_, new_n10218_ );
or   ( new_n10230_, new_n1425_, new_n3902_ );
or   ( new_n10231_, new_n1429_, new_n3924_ );
and  ( new_n10232_, new_n10231_, new_n10230_ );
and  ( new_n10233_, new_n10232_, new_n1355_ );
and  ( new_n10234_, new_n1433_, RI2b1c4342dfa8_88 );
and  ( new_n10235_, new_n1423_, RI2b1c4342df30_87 );
or   ( new_n10236_, new_n10235_, new_n10234_ );
and  ( new_n10237_, new_n10236_, new_n1267_ );
or   ( new_n10238_, new_n10237_, new_n10233_ );
and  ( new_n10239_, new_n10238_, new_n10229_ );
or   ( new_n10240_, new_n10239_, new_n10228_ );
and  ( new_n10241_, new_n10240_, new_n10209_ );
or   ( new_n10242_, new_n10241_, new_n10208_ );
or   ( new_n10243_, new_n10046_, new_n9824_ );
and  ( new_n10244_, new_n10243_, new_n9830_ );
and  ( new_n10245_, new_n10042_, new_n9823_ );
and  ( new_n10246_, new_n10045_, new_n9814_ );
or   ( new_n10247_, new_n10246_, new_n10245_ );
and  ( new_n10248_, new_n10247_, new_n10050_ );
or   ( new_n10249_, new_n10248_, new_n10244_ );
or   ( new_n10250_, new_n934_, new_n4635_ );
or   ( new_n10251_, new_n940_, new_n132_ );
and  ( new_n10252_, new_n10251_, new_n10250_ );
and  ( new_n10253_, new_n10252_, new_n913_ );
and  ( new_n10254_, new_n944_, RI2b1c4342e098_90 );
and  ( new_n10255_, new_n932_, RI2b1c4342e020_89 );
or   ( new_n10256_, new_n10255_, new_n10254_ );
and  ( new_n10257_, new_n10256_, new_n938_ );
or   ( new_n10258_, new_n10257_, new_n10253_ );
or   ( new_n10259_, new_n453_, new_n5459_ );
or   ( new_n10260_, new_n459_, new_n117_ );
and  ( new_n10261_, new_n10260_, new_n10259_ );
and  ( new_n10262_, new_n10261_, new_n428_ );
and  ( new_n10263_, new_n463_, RI2b1c4342e188_92 );
and  ( new_n10264_, new_n451_, RI2b1c4342e110_91 );
or   ( new_n10265_, new_n10264_, new_n10263_ );
and  ( new_n10266_, new_n10265_, new_n457_ );
or   ( new_n10267_, new_n10266_, new_n10262_ );
and  ( new_n10268_, new_n10267_, new_n10258_ );
or   ( new_n10269_, new_n10267_, new_n10258_ );
or   ( new_n10270_, new_n524_, new_n6321_ );
or   ( new_n10271_, new_n528_, new_n6307_ );
and  ( new_n10272_, new_n10271_, new_n10270_ );
and  ( new_n10273_, new_n10272_, new_n505_ );
and  ( new_n10274_, new_n537_, RI2b1c4342e278_94 );
and  ( new_n10275_, new_n522_, RI2b1c4342e200_93 );
or   ( new_n10276_, new_n10275_, new_n10274_ );
and  ( new_n10277_, new_n10276_, new_n533_ );
or   ( new_n10278_, new_n10277_, new_n10273_ );
and  ( new_n10279_, new_n10278_, new_n10269_ );
or   ( new_n10280_, new_n10279_, new_n10268_ );
and  ( new_n10281_, new_n10280_, new_n10249_ );
or   ( new_n10282_, new_n10280_, new_n10249_ );
or   ( new_n10283_, new_n10033_, new_n9793_ );
and  ( new_n10284_, new_n10283_, new_n9803_ );
and  ( new_n10285_, new_n10029_, new_n9792_ );
and  ( new_n10286_, new_n10032_, new_n9783_ );
or   ( new_n10287_, new_n10286_, new_n10285_ );
and  ( new_n10288_, new_n10287_, new_n10037_ );
or   ( new_n10289_, new_n10288_, new_n10284_ );
and  ( new_n10290_, new_n10289_, new_n10282_ );
or   ( new_n10291_, new_n10290_, new_n10281_ );
and  ( new_n10292_, new_n10291_, new_n10242_ );
or   ( new_n10293_, new_n10291_, new_n10242_ );
or   ( new_n10294_, new_n10091_, new_n9919_ );
and  ( new_n10295_, new_n10294_, new_n9929_ );
and  ( new_n10296_, new_n10087_, new_n9918_ );
and  ( new_n10297_, new_n10090_, new_n9909_ );
or   ( new_n10298_, new_n10297_, new_n10296_ );
and  ( new_n10299_, new_n10298_, new_n10095_ );
or   ( new_n10300_, new_n10299_, new_n10295_ );
or   ( new_n10301_, new_n10066_, new_n9864_ );
and  ( new_n10302_, new_n10301_, new_n9874_ );
and  ( new_n10303_, new_n10062_, new_n9863_ );
and  ( new_n10304_, new_n10065_, new_n9854_ );
or   ( new_n10305_, new_n10304_, new_n10303_ );
and  ( new_n10306_, new_n10305_, new_n10070_ );
or   ( new_n10307_, new_n10306_, new_n10302_ );
and  ( new_n10308_, new_n10307_, new_n10300_ );
or   ( new_n10309_, new_n10307_, new_n10300_ );
or   ( new_n10310_, new_n10077_, new_n9886_ );
and  ( new_n10311_, new_n10310_, new_n9896_ );
and  ( new_n10312_, new_n9885_, new_n762_ );
and  ( new_n10313_, new_n10075_, new_n734_ );
or   ( new_n10314_, new_n10313_, new_n10312_ );
and  ( new_n10315_, new_n10314_, new_n10080_ );
or   ( new_n10316_, new_n10315_, new_n10311_ );
and  ( new_n10317_, new_n10316_, new_n10309_ );
or   ( new_n10318_, new_n10317_, new_n10308_ );
and  ( new_n10319_, new_n10318_, new_n10293_ );
or   ( new_n10320_, new_n10319_, new_n10292_ );
or   ( new_n10321_, new_n9618_, new_n9475_ );
and  ( new_n10322_, new_n10321_, new_n9485_ );
and  ( new_n10323_, new_n9614_, new_n9474_ );
and  ( new_n10324_, new_n9617_, new_n9465_ );
or   ( new_n10325_, new_n10324_, new_n10323_ );
and  ( new_n10326_, new_n10325_, new_n9622_ );
or   ( new_n10327_, new_n10326_, new_n10322_ );
or   ( new_n10328_, new_n9605_, new_n9444_ );
and  ( new_n10329_, new_n10328_, new_n9454_ );
and  ( new_n10330_, new_n9601_, new_n9443_ );
and  ( new_n10331_, new_n9604_, new_n9434_ );
or   ( new_n10332_, new_n10331_, new_n10330_ );
and  ( new_n10333_, new_n10332_, new_n9609_ );
or   ( new_n10334_, new_n10333_, new_n10329_ );
and  ( new_n10335_, new_n10334_, new_n10327_ );
or   ( new_n10336_, new_n10334_, new_n10327_ );
or   ( new_n10337_, new_n10108_, new_n9952_ );
and  ( new_n10338_, new_n10337_, new_n9960_ );
and  ( new_n10339_, new_n10104_, new_n9951_ );
and  ( new_n10340_, new_n10107_, new_n9944_ );
or   ( new_n10341_, new_n10340_, new_n10339_ );
and  ( new_n10342_, new_n10341_, new_n10112_ );
or   ( new_n10343_, new_n10342_, new_n10338_ );
and  ( new_n10344_, new_n10343_, new_n10336_ );
or   ( new_n10345_, new_n10344_, new_n10335_ );
and  ( new_n10346_, new_n10345_, new_n10320_ );
or   ( new_n10347_, new_n10345_, new_n10320_ );
or   ( new_n10348_, new_n9625_, new_n9488_ );
and  ( new_n10349_, new_n10348_, new_n9520_ );
and  ( new_n10350_, new_n9611_, new_n9487_ );
and  ( new_n10351_, new_n9624_, new_n9456_ );
or   ( new_n10352_, new_n10351_, new_n10350_ );
and  ( new_n10353_, new_n10352_, new_n9639_ );
or   ( new_n10354_, new_n10353_, new_n10349_ );
and  ( new_n10355_, new_n10354_, new_n10347_ );
or   ( new_n10356_, new_n10355_, new_n10346_ );
and  ( new_n10357_, new_n10356_, new_n10145_ );
or   ( new_n10358_, new_n10356_, new_n10145_ );
or   ( new_n10359_, new_n10118_, new_n9965_ );
and  ( new_n10360_, new_n10359_, new_n9973_ );
and  ( new_n10361_, new_n10116_, new_n9774_ );
and  ( new_n10362_, new_n10026_, new_n9964_ );
or   ( new_n10363_, new_n10362_, new_n10361_ );
and  ( new_n10364_, new_n10363_, new_n10121_ );
or   ( new_n10365_, new_n10364_, new_n10360_ );
and  ( new_n10366_, new_n10365_, new_n10358_ );
or   ( new_n10367_, new_n10366_, new_n10357_ );
and  ( new_n10368_, new_n10367_, new_n10143_ );
or   ( new_n10369_, new_n10367_, new_n10143_ );
or   ( new_n10370_, new_n10125_, new_n9976_ );
and  ( new_n10371_, new_n10370_, new_n9984_ );
and  ( new_n10372_, new_n10123_, new_n9749_ );
and  ( new_n10373_, new_n10013_, new_n9975_ );
or   ( new_n10374_, new_n10373_, new_n10372_ );
and  ( new_n10375_, new_n10374_, new_n10128_ );
or   ( new_n10376_, new_n10375_, new_n10371_ );
and  ( new_n10377_, new_n10376_, new_n10369_ );
or   ( new_n10378_, new_n10377_, new_n10368_ );
or   ( new_n10379_, new_n10378_, new_n10141_ );
and  ( new_n10380_, new_n10379_, new_n9999_ );
or   ( new_n10381_, new_n10380_, new_n9998_ );
and  ( new_n10382_, new_n10378_, new_n10141_ );
or   ( new_n10383_, new_n10382_, new_n9998_ );
and  ( new_n10384_, new_n10002_, new_n9733_ );
and  ( new_n10385_, new_n10005_, new_n9726_ );
or   ( new_n10386_, new_n10385_, new_n10384_ );
and  ( new_n10387_, new_n10009_, new_n9748_ );
and  ( new_n10388_, new_n10012_, new_n9741_ );
or   ( new_n10389_, new_n10388_, new_n10387_ );
and  ( new_n10390_, new_n10152_, new_n5858_ );
and  ( new_n10391_, new_n10148_, new_n6037_ );
or   ( new_n10392_, new_n10391_, new_n10390_ );
and  ( new_n10393_, new_n10161_, new_n6039_ );
and  ( new_n10394_, new_n10157_, new_n5867_ );
or   ( new_n10395_, new_n10394_, new_n10393_ );
and  ( new_n10396_, new_n10395_, new_n10392_ );
or   ( new_n10397_, new_n10395_, new_n10392_ );
and  ( new_n10398_, new_n10172_, new_n5182_ );
and  ( new_n10399_, new_n10168_, new_n5028_ );
or   ( new_n10400_, new_n10399_, new_n10398_ );
and  ( new_n10401_, new_n10400_, new_n10397_ );
or   ( new_n10402_, new_n10401_, new_n10396_ );
and  ( new_n10403_, new_n10183_, new_n4400_ );
and  ( new_n10404_, new_n10179_, new_n4215_ );
or   ( new_n10405_, new_n10404_, new_n10403_ );
and  ( new_n10406_, new_n10192_, new_n3695_ );
and  ( new_n10407_, new_n10188_, new_n3548_ );
or   ( new_n10408_, new_n10407_, new_n10406_ );
and  ( new_n10409_, new_n10408_, new_n10405_ );
or   ( new_n10410_, new_n10408_, new_n10405_ );
and  ( new_n10411_, new_n10203_, new_n3004_ );
and  ( new_n10412_, new_n10199_, new_n2868_ );
or   ( new_n10413_, new_n10412_, new_n10411_ );
and  ( new_n10414_, new_n10413_, new_n10410_ );
or   ( new_n10415_, new_n10414_, new_n10409_ );
and  ( new_n10416_, new_n10415_, new_n10402_ );
or   ( new_n10417_, new_n10415_, new_n10402_ );
and  ( new_n10418_, new_n10216_, new_n2334_ );
and  ( new_n10419_, new_n10212_, new_n2168_ );
or   ( new_n10420_, new_n10419_, new_n10418_ );
and  ( new_n10421_, new_n10225_, new_n1824_ );
and  ( new_n10422_, new_n10221_, new_n1717_ );
or   ( new_n10423_, new_n10422_, new_n10421_ );
and  ( new_n10424_, new_n10423_, new_n10420_ );
or   ( new_n10425_, new_n10423_, new_n10420_ );
and  ( new_n10426_, new_n10236_, new_n1355_ );
and  ( new_n10427_, new_n10232_, new_n1267_ );
or   ( new_n10428_, new_n10427_, new_n10426_ );
and  ( new_n10429_, new_n10428_, new_n10425_ );
or   ( new_n10430_, new_n10429_, new_n10424_ );
and  ( new_n10431_, new_n10430_, new_n10417_ );
or   ( new_n10432_, new_n10431_, new_n10416_ );
and  ( new_n10433_, new_n10247_, new_n9830_ );
and  ( new_n10434_, new_n10243_, new_n10050_ );
or   ( new_n10435_, new_n10434_, new_n10433_ );
and  ( new_n10436_, new_n10256_, new_n913_ );
and  ( new_n10437_, new_n10252_, new_n938_ );
or   ( new_n10438_, new_n10437_, new_n10436_ );
and  ( new_n10439_, new_n10265_, new_n428_ );
and  ( new_n10440_, new_n10261_, new_n457_ );
or   ( new_n10441_, new_n10440_, new_n10439_ );
and  ( new_n10442_, new_n10441_, new_n10438_ );
or   ( new_n10443_, new_n10441_, new_n10438_ );
and  ( new_n10444_, new_n10276_, new_n505_ );
and  ( new_n10445_, new_n10272_, new_n533_ );
or   ( new_n10446_, new_n10445_, new_n10444_ );
and  ( new_n10447_, new_n10446_, new_n10443_ );
or   ( new_n10448_, new_n10447_, new_n10442_ );
and  ( new_n10449_, new_n10448_, new_n10435_ );
or   ( new_n10450_, new_n10448_, new_n10435_ );
and  ( new_n10451_, new_n10287_, new_n9803_ );
and  ( new_n10452_, new_n10283_, new_n10037_ );
or   ( new_n10453_, new_n10452_, new_n10451_ );
and  ( new_n10454_, new_n10453_, new_n10450_ );
or   ( new_n10455_, new_n10454_, new_n10449_ );
and  ( new_n10456_, new_n10455_, new_n10432_ );
or   ( new_n10457_, new_n10455_, new_n10432_ );
and  ( new_n10458_, new_n10298_, new_n9929_ );
and  ( new_n10459_, new_n10294_, new_n10095_ );
or   ( new_n10460_, new_n10459_, new_n10458_ );
and  ( new_n10461_, new_n10305_, new_n9874_ );
and  ( new_n10462_, new_n10301_, new_n10070_ );
or   ( new_n10463_, new_n10462_, new_n10461_ );
and  ( new_n10464_, new_n10463_, new_n10460_ );
or   ( new_n10465_, new_n10463_, new_n10460_ );
and  ( new_n10466_, new_n10314_, new_n9896_ );
and  ( new_n10467_, new_n10310_, new_n10080_ );
or   ( new_n10468_, new_n10467_, new_n10466_ );
and  ( new_n10469_, new_n10468_, new_n10465_ );
or   ( new_n10470_, new_n10469_, new_n10464_ );
and  ( new_n10471_, new_n10470_, new_n10457_ );
or   ( new_n10472_, new_n10471_, new_n10456_ );
and  ( new_n10473_, new_n10325_, new_n9485_ );
and  ( new_n10474_, new_n10321_, new_n9622_ );
or   ( new_n10475_, new_n10474_, new_n10473_ );
and  ( new_n10476_, new_n10332_, new_n9454_ );
and  ( new_n10477_, new_n10328_, new_n9609_ );
or   ( new_n10478_, new_n10477_, new_n10476_ );
and  ( new_n10479_, new_n10478_, new_n10475_ );
or   ( new_n10480_, new_n10478_, new_n10475_ );
and  ( new_n10481_, new_n10341_, new_n9960_ );
and  ( new_n10482_, new_n10337_, new_n10112_ );
or   ( new_n10483_, new_n10482_, new_n10481_ );
and  ( new_n10484_, new_n10483_, new_n10480_ );
or   ( new_n10485_, new_n10484_, new_n10479_ );
and  ( new_n10486_, new_n10485_, new_n10472_ );
or   ( new_n10487_, new_n10485_, new_n10472_ );
and  ( new_n10488_, new_n10352_, new_n9520_ );
and  ( new_n10489_, new_n10348_, new_n9639_ );
or   ( new_n10490_, new_n10489_, new_n10488_ );
and  ( new_n10491_, new_n10490_, new_n10487_ );
or   ( new_n10492_, new_n10491_, new_n10486_ );
and  ( new_n10493_, new_n10492_, new_n10389_ );
or   ( new_n10494_, new_n10492_, new_n10389_ );
and  ( new_n10495_, new_n10363_, new_n9973_ );
and  ( new_n10496_, new_n10359_, new_n10121_ );
or   ( new_n10497_, new_n10496_, new_n10495_ );
and  ( new_n10498_, new_n10497_, new_n10494_ );
or   ( new_n10499_, new_n10498_, new_n10493_ );
and  ( new_n10500_, new_n10499_, new_n10386_ );
or   ( new_n10501_, new_n10500_, new_n10368_ );
and  ( new_n10502_, new_n10501_, new_n10376_ );
and  ( new_n10503_, new_n10499_, new_n10143_ );
and  ( new_n10504_, new_n10386_, new_n10367_ );
or   ( new_n10505_, new_n10504_, new_n10503_ );
and  ( new_n10506_, new_n10374_, new_n9984_ );
and  ( new_n10507_, new_n10370_, new_n10128_ );
or   ( new_n10508_, new_n10507_, new_n10506_ );
and  ( new_n10509_, new_n10508_, new_n10505_ );
or   ( new_n10510_, new_n10509_, new_n10502_ );
or   ( new_n10511_, new_n10101_, new_n9934_ );
and  ( new_n10512_, new_n10511_, new_n9962_ );
and  ( new_n10513_, new_n10099_, new_n9845_ );
and  ( new_n10514_, new_n10059_, new_n9933_ );
or   ( new_n10515_, new_n10514_, new_n10513_ );
and  ( new_n10516_, new_n10515_, new_n10114_ );
or   ( new_n10517_, new_n10516_, new_n10512_ );
or   ( new_n10518_, new_n10486_, new_n10346_ );
and  ( new_n10519_, new_n10518_, new_n10354_ );
and  ( new_n10520_, new_n10472_, new_n10345_ );
and  ( new_n10521_, new_n10485_, new_n10320_ );
or   ( new_n10522_, new_n10521_, new_n10520_ );
and  ( new_n10523_, new_n10522_, new_n10490_ );
or   ( new_n10524_, new_n10523_, new_n10519_ );
or   ( new_n10525_, new_n10524_, new_n10517_ );
or   ( new_n10526_, new_n10084_, new_n9899_ );
and  ( new_n10527_, new_n10526_, new_n9931_ );
and  ( new_n10528_, new_n10082_, new_n9876_ );
and  ( new_n10529_, new_n10072_, new_n9898_ );
or   ( new_n10530_, new_n10529_, new_n10528_ );
and  ( new_n10531_, new_n10530_, new_n10097_ );
or   ( new_n10532_, new_n10531_, new_n10527_ );
or   ( new_n10533_, new_n10479_, new_n10335_ );
and  ( new_n10534_, new_n10533_, new_n10343_ );
and  ( new_n10535_, new_n10475_, new_n10334_ );
and  ( new_n10536_, new_n10478_, new_n10327_ );
or   ( new_n10537_, new_n10536_, new_n10535_ );
and  ( new_n10538_, new_n10537_, new_n10483_ );
or   ( new_n10539_, new_n10538_, new_n10534_ );
and  ( new_n10540_, new_n10539_, new_n10532_ );
or   ( new_n10541_, new_n10539_, new_n10532_ );
or   ( new_n10542_, new_n10456_, new_n10292_ );
and  ( new_n10543_, new_n10542_, new_n10318_ );
and  ( new_n10544_, new_n10432_, new_n10291_ );
and  ( new_n10545_, new_n10455_, new_n10242_ );
or   ( new_n10546_, new_n10545_, new_n10544_ );
and  ( new_n10547_, new_n10546_, new_n10470_ );
or   ( new_n10548_, new_n10547_, new_n10543_ );
and  ( new_n10549_, new_n10548_, new_n10541_ );
or   ( new_n10550_, new_n10549_, new_n10540_ );
or   ( new_n10551_, new_n10464_, new_n10308_ );
and  ( new_n10552_, new_n10551_, new_n10316_ );
and  ( new_n10553_, new_n10460_, new_n10307_ );
and  ( new_n10554_, new_n10463_, new_n10300_ );
or   ( new_n10555_, new_n10554_, new_n10553_ );
and  ( new_n10556_, new_n10555_, new_n10468_ );
or   ( new_n10557_, new_n10556_, new_n10552_ );
or   ( new_n10558_, new_n10449_, new_n10281_ );
and  ( new_n10559_, new_n10558_, new_n10289_ );
and  ( new_n10560_, new_n10448_, new_n10249_ );
and  ( new_n10561_, new_n10435_, new_n10280_ );
or   ( new_n10562_, new_n10561_, new_n10560_ );
and  ( new_n10563_, new_n10562_, new_n10453_ );
or   ( new_n10564_, new_n10563_, new_n10559_ );
and  ( new_n10565_, new_n10564_, new_n10557_ );
or   ( new_n10566_, new_n10564_, new_n10557_ );
or   ( new_n10567_, new_n10416_, new_n10208_ );
and  ( new_n10568_, new_n10567_, new_n10240_ );
and  ( new_n10569_, new_n10402_, new_n10207_ );
and  ( new_n10570_, new_n10415_, new_n10176_ );
or   ( new_n10571_, new_n10570_, new_n10569_ );
and  ( new_n10572_, new_n10571_, new_n10430_ );
or   ( new_n10573_, new_n10572_, new_n10568_ );
and  ( new_n10574_, new_n10573_, new_n10566_ );
or   ( new_n10575_, new_n10574_, new_n10565_ );
or   ( new_n10576_, new_n524_, new_n124_ );
or   ( new_n10577_, new_n528_, new_n6321_ );
and  ( new_n10578_, new_n10577_, new_n10576_ );
and  ( new_n10579_, new_n10578_, new_n505_ );
and  ( new_n10580_, new_n537_, RI2b1c4342e2f0_95 );
and  ( new_n10581_, new_n522_, RI2b1c4342e278_94 );
or   ( new_n10582_, new_n10581_, new_n10580_ );
and  ( new_n10583_, new_n10582_, new_n533_ );
or   ( new_n10584_, new_n10583_, new_n10579_ );
or   ( new_n10585_, new_n614_, new_n7274_ );
and  ( new_n10586_, new_n10585_, new_n590_ );
and  ( new_n10587_, new_n608_, RI2b1c4342e368_96 );
and  ( new_n10588_, new_n10587_, new_n619_ );
or   ( new_n10589_, new_n10588_, new_n10586_ );
or   ( new_n10590_, new_n10589_, new_n10584_ );
or   ( new_n10591_, new_n1425_, new_n132_ );
or   ( new_n10592_, new_n1429_, new_n3902_ );
and  ( new_n10593_, new_n10592_, new_n10591_ );
and  ( new_n10594_, new_n10593_, new_n1355_ );
and  ( new_n10595_, new_n1433_, RI2b1c4342e020_89 );
and  ( new_n10596_, new_n1423_, RI2b1c4342dfa8_88 );
or   ( new_n10597_, new_n10596_, new_n10595_ );
and  ( new_n10598_, new_n10597_, new_n1267_ );
or   ( new_n10599_, new_n10598_, new_n10594_ );
or   ( new_n10600_, new_n934_, new_n117_ );
or   ( new_n10601_, new_n940_, new_n4635_ );
and  ( new_n10602_, new_n10601_, new_n10600_ );
and  ( new_n10603_, new_n10602_, new_n913_ );
and  ( new_n10604_, new_n944_, RI2b1c4342e110_91 );
and  ( new_n10605_, new_n932_, RI2b1c4342e098_90 );
or   ( new_n10606_, new_n10605_, new_n10604_ );
and  ( new_n10607_, new_n10606_, new_n938_ );
or   ( new_n10608_, new_n10607_, new_n10603_ );
and  ( new_n10609_, new_n10608_, new_n10599_ );
or   ( new_n10610_, new_n10608_, new_n10599_ );
or   ( new_n10611_, new_n453_, new_n6307_ );
or   ( new_n10612_, new_n459_, new_n5459_ );
and  ( new_n10613_, new_n10612_, new_n10611_ );
and  ( new_n10614_, new_n10613_, new_n428_ );
and  ( new_n10615_, new_n463_, RI2b1c4342e200_93 );
and  ( new_n10616_, new_n451_, RI2b1c4342e188_92 );
or   ( new_n10617_, new_n10616_, new_n10615_ );
and  ( new_n10618_, new_n10617_, new_n457_ );
or   ( new_n10619_, new_n10618_, new_n10614_ );
and  ( new_n10620_, new_n10619_, new_n10610_ );
or   ( new_n10621_, new_n10620_, new_n10609_ );
and  ( new_n10622_, new_n10621_, new_n10590_ );
or   ( new_n10623_, new_n10621_, new_n10590_ );
or   ( new_n10624_, new_n610_, new_n7274_ );
or   ( new_n10625_, new_n614_, new_n124_ );
and  ( new_n10626_, new_n10625_, new_n10624_ );
and  ( new_n10627_, new_n10626_, new_n590_ );
and  ( new_n10628_, new_n623_, RI2b1c4342e368_96 );
and  ( new_n10629_, new_n608_, RI2b1c4342e2f0_95 );
or   ( new_n10630_, new_n10629_, new_n10628_ );
and  ( new_n10631_, new_n10630_, new_n619_ );
or   ( new_n10632_, new_n10631_, new_n10627_ );
and  ( new_n10633_, new_n10632_, new_n10623_ );
or   ( new_n10634_, new_n10633_, new_n10622_ );
or   ( new_n10635_, new_n5308_, new_n1004_ );
or   ( new_n10636_, new_n5312_, new_n886_ );
and  ( new_n10637_, new_n10636_, new_n10635_ );
and  ( new_n10638_, new_n10637_, new_n5182_ );
and  ( new_n10639_, new_n5316_, RI2b1c4342da80_77 );
and  ( new_n10640_, new_n5306_, RI2b1c4342da08_76 );
or   ( new_n10641_, new_n10640_, new_n10639_ );
and  ( new_n10642_, new_n10641_, new_n5028_ );
or   ( new_n10643_, new_n10642_, new_n10638_ );
or   ( new_n10644_, new_n4535_, new_n1310_ );
or   ( new_n10645_, new_n4539_, new_n1002_ );
and  ( new_n10646_, new_n10645_, new_n10644_ );
and  ( new_n10647_, new_n10646_, new_n4400_ );
and  ( new_n10648_, new_n4543_, RI2b1c4342db70_79 );
and  ( new_n10649_, new_n4533_, RI2b1c4342daf8_78 );
or   ( new_n10650_, new_n10649_, new_n10648_ );
and  ( new_n10651_, new_n10650_, new_n4215_ );
or   ( new_n10652_, new_n10651_, new_n10647_ );
and  ( new_n10653_, new_n10652_, new_n10643_ );
or   ( new_n10654_, new_n10652_, new_n10643_ );
or   ( new_n10655_, new_n3802_, new_n126_ );
or   ( new_n10656_, new_n3806_, new_n1511_ );
and  ( new_n10657_, new_n10656_, new_n10655_ );
and  ( new_n10658_, new_n10657_, new_n3695_ );
and  ( new_n10659_, new_n3810_, RI2b1c4342dc60_81 );
and  ( new_n10660_, new_n3800_, RI2b1c4342dbe8_80 );
or   ( new_n10661_, new_n10660_, new_n10659_ );
and  ( new_n10662_, new_n10661_, new_n3548_ );
or   ( new_n10663_, new_n10662_, new_n10658_ );
and  ( new_n10664_, new_n10663_, new_n10654_ );
or   ( new_n10665_, new_n10664_, new_n10653_ );
or   ( new_n10666_, new_n7105_, new_n105_ );
or   ( new_n10667_, new_n7099_, new_n806_ );
and  ( new_n10668_, new_n10667_, new_n10666_ );
and  ( new_n10669_, new_n10668_, new_n5858_ );
and  ( new_n10670_, new_n7104_, RI2b1c4342d828_72 );
and  ( new_n10671_, new_n7110_, RI2b1c4342d8a0_73 );
or   ( new_n10672_, new_n10671_, new_n10670_ );
and  ( new_n10673_, new_n10672_, new_n6037_ );
or   ( new_n10674_, new_n10673_, new_n10669_ );
and  ( new_n10675_, new_n10674_, new_n590_ );
or   ( new_n10676_, new_n10674_, new_n590_ );
or   ( new_n10677_, new_n6156_, new_n843_ );
or   ( new_n10678_, new_n6160_, new_n859_ );
and  ( new_n10679_, new_n10678_, new_n10677_ );
and  ( new_n10680_, new_n10679_, new_n6039_ );
and  ( new_n10681_, new_n6164_, RI2b1c4342d990_75 );
and  ( new_n10682_, new_n6154_, RI2b1c4342d918_74 );
or   ( new_n10683_, new_n10682_, new_n10681_ );
and  ( new_n10684_, new_n10683_, new_n5867_ );
or   ( new_n10685_, new_n10684_, new_n10680_ );
and  ( new_n10686_, new_n10685_, new_n10676_ );
or   ( new_n10687_, new_n10686_, new_n10675_ );
and  ( new_n10688_, new_n10687_, new_n10665_ );
or   ( new_n10689_, new_n10687_, new_n10665_ );
or   ( new_n10690_, new_n3112_, new_n121_ );
or   ( new_n10691_, new_n3116_, new_n2119_ );
and  ( new_n10692_, new_n10691_, new_n10690_ );
and  ( new_n10693_, new_n10692_, new_n3004_ );
and  ( new_n10694_, new_n3120_, RI2b1c4342dd50_83 );
and  ( new_n10695_, new_n3110_, RI2b1c4342dcd8_82 );
or   ( new_n10696_, new_n10695_, new_n10694_ );
and  ( new_n10697_, new_n10696_, new_n2868_ );
or   ( new_n10698_, new_n10697_, new_n10693_ );
or   ( new_n10699_, new_n2450_, new_n2806_ );
or   ( new_n10700_, new_n2454_, new_n2541_ );
and  ( new_n10701_, new_n10700_, new_n10699_ );
and  ( new_n10702_, new_n10701_, new_n2334_ );
and  ( new_n10703_, new_n2458_, RI2b1c4342de40_85 );
and  ( new_n10704_, new_n2448_, RI2b1c4342ddc8_84 );
or   ( new_n10705_, new_n10704_, new_n10703_ );
and  ( new_n10706_, new_n10705_, new_n2168_ );
or   ( new_n10707_, new_n10706_, new_n10702_ );
and  ( new_n10708_, new_n10707_, new_n10698_ );
or   ( new_n10709_, new_n10707_, new_n10698_ );
or   ( new_n10710_, new_n1910_, new_n3924_ );
or   ( new_n10711_, new_n1914_, new_n3239_ );
and  ( new_n10712_, new_n10711_, new_n10710_ );
and  ( new_n10713_, new_n10712_, new_n1824_ );
and  ( new_n10714_, new_n1918_, RI2b1c4342df30_87 );
and  ( new_n10715_, new_n1908_, RI2b1c4342deb8_86 );
or   ( new_n10716_, new_n10715_, new_n10714_ );
and  ( new_n10717_, new_n10716_, new_n1717_ );
or   ( new_n10718_, new_n10717_, new_n10713_ );
and  ( new_n10719_, new_n10718_, new_n10709_ );
or   ( new_n10720_, new_n10719_, new_n10708_ );
and  ( new_n10721_, new_n10720_, new_n10689_ );
or   ( new_n10722_, new_n10721_, new_n10688_ );
and  ( new_n10723_, new_n10722_, new_n10634_ );
or   ( new_n10724_, new_n10722_, new_n10634_ );
or   ( new_n10725_, new_n10442_, new_n10268_ );
and  ( new_n10726_, new_n10725_, new_n10278_ );
and  ( new_n10727_, new_n10438_, new_n10267_ );
and  ( new_n10728_, new_n10441_, new_n10258_ );
or   ( new_n10729_, new_n10728_, new_n10727_ );
and  ( new_n10730_, new_n10729_, new_n10446_ );
or   ( new_n10731_, new_n10730_, new_n10726_ );
or   ( new_n10732_, new_n10424_, new_n10228_ );
and  ( new_n10733_, new_n10732_, new_n10238_ );
and  ( new_n10734_, new_n10420_, new_n10227_ );
and  ( new_n10735_, new_n10423_, new_n10218_ );
or   ( new_n10736_, new_n10735_, new_n10734_ );
and  ( new_n10737_, new_n10736_, new_n10428_ );
or   ( new_n10738_, new_n10737_, new_n10733_ );
and  ( new_n10739_, new_n10738_, new_n10731_ );
or   ( new_n10740_, new_n10738_, new_n10731_ );
or   ( new_n10741_, new_n10409_, new_n10195_ );
and  ( new_n10742_, new_n10741_, new_n10205_ );
and  ( new_n10743_, new_n10405_, new_n10194_ );
and  ( new_n10744_, new_n10408_, new_n10185_ );
or   ( new_n10745_, new_n10744_, new_n10743_ );
and  ( new_n10746_, new_n10745_, new_n10413_ );
or   ( new_n10747_, new_n10746_, new_n10742_ );
and  ( new_n10748_, new_n10747_, new_n10740_ );
or   ( new_n10749_, new_n10748_, new_n10739_ );
and  ( new_n10750_, new_n10749_, new_n10724_ );
or   ( new_n10751_, new_n10750_, new_n10723_ );
and  ( new_n10752_, new_n10751_, new_n10575_ );
or   ( new_n10753_, new_n10751_, new_n10575_ );
or   ( new_n10754_, new_n10053_, new_n9833_ );
and  ( new_n10755_, new_n10754_, new_n9843_ );
and  ( new_n10756_, new_n10039_, new_n9832_ );
and  ( new_n10757_, new_n10052_, new_n9805_ );
or   ( new_n10758_, new_n10757_, new_n10756_ );
and  ( new_n10759_, new_n10758_, new_n10057_ );
or   ( new_n10760_, new_n10759_, new_n10755_ );
and  ( new_n10761_, new_n10760_, new_n10753_ );
or   ( new_n10762_, new_n10761_, new_n10752_ );
and  ( new_n10763_, new_n10762_, new_n10550_ );
or   ( new_n10764_, new_n10762_, new_n10550_ );
or   ( new_n10765_, new_n10020_, new_n9764_ );
and  ( new_n10766_, new_n10765_, new_n9772_ );
and  ( new_n10767_, new_n10016_, new_n9763_ );
and  ( new_n10768_, new_n10019_, new_n9756_ );
or   ( new_n10769_, new_n10768_, new_n10767_ );
and  ( new_n10770_, new_n10769_, new_n10024_ );
or   ( new_n10771_, new_n10770_, new_n10766_ );
and  ( new_n10772_, new_n10771_, new_n10764_ );
or   ( new_n10773_, new_n10772_, new_n10763_ );
and  ( new_n10774_, new_n10773_, new_n10525_ );
or   ( new_n10775_, new_n10773_, new_n10525_ );
or   ( new_n10776_, new_n10493_, new_n10357_ );
and  ( new_n10777_, new_n10776_, new_n10365_ );
and  ( new_n10778_, new_n10492_, new_n10145_ );
and  ( new_n10779_, new_n10389_, new_n10356_ );
or   ( new_n10780_, new_n10779_, new_n10778_ );
and  ( new_n10781_, new_n10780_, new_n10497_ );
or   ( new_n10782_, new_n10781_, new_n10777_ );
and  ( new_n10783_, new_n10782_, new_n10775_ );
or   ( new_n10784_, new_n10783_, new_n10774_ );
and  ( new_n10785_, new_n10784_, new_n10510_ );
or   ( new_n10786_, new_n10784_, new_n10510_ );
and  ( new_n10787_, new_n10515_, new_n9962_ );
and  ( new_n10788_, new_n10511_, new_n10114_ );
or   ( new_n10789_, new_n10788_, new_n10787_ );
and  ( new_n10790_, new_n10522_, new_n10354_ );
and  ( new_n10791_, new_n10518_, new_n10490_ );
or   ( new_n10792_, new_n10791_, new_n10790_ );
and  ( new_n10793_, new_n10792_, new_n10789_ );
and  ( new_n10794_, new_n10530_, new_n9931_ );
and  ( new_n10795_, new_n10526_, new_n10097_ );
or   ( new_n10796_, new_n10795_, new_n10794_ );
and  ( new_n10797_, new_n10537_, new_n10343_ );
and  ( new_n10798_, new_n10533_, new_n10483_ );
or   ( new_n10799_, new_n10798_, new_n10797_ );
and  ( new_n10800_, new_n10799_, new_n10796_ );
or   ( new_n10801_, new_n10799_, new_n10796_ );
and  ( new_n10802_, new_n10546_, new_n10318_ );
and  ( new_n10803_, new_n10542_, new_n10470_ );
or   ( new_n10804_, new_n10803_, new_n10802_ );
and  ( new_n10805_, new_n10804_, new_n10801_ );
or   ( new_n10806_, new_n10805_, new_n10800_ );
and  ( new_n10807_, new_n10555_, new_n10316_ );
and  ( new_n10808_, new_n10551_, new_n10468_ );
or   ( new_n10809_, new_n10808_, new_n10807_ );
and  ( new_n10810_, new_n10562_, new_n10289_ );
and  ( new_n10811_, new_n10558_, new_n10453_ );
or   ( new_n10812_, new_n10811_, new_n10810_ );
and  ( new_n10813_, new_n10812_, new_n10809_ );
or   ( new_n10814_, new_n10812_, new_n10809_ );
and  ( new_n10815_, new_n10571_, new_n10240_ );
and  ( new_n10816_, new_n10567_, new_n10430_ );
or   ( new_n10817_, new_n10816_, new_n10815_ );
and  ( new_n10818_, new_n10817_, new_n10814_ );
or   ( new_n10819_, new_n10818_, new_n10813_ );
and  ( new_n10820_, new_n10582_, new_n505_ );
and  ( new_n10821_, new_n10578_, new_n533_ );
or   ( new_n10822_, new_n10821_, new_n10820_ );
and  ( new_n10823_, new_n10587_, new_n590_ );
and  ( new_n10824_, new_n10585_, new_n619_ );
or   ( new_n10825_, new_n10824_, new_n10823_ );
and  ( new_n10826_, new_n10825_, new_n10822_ );
and  ( new_n10827_, new_n10597_, new_n1355_ );
and  ( new_n10828_, new_n10593_, new_n1267_ );
or   ( new_n10829_, new_n10828_, new_n10827_ );
and  ( new_n10830_, new_n10606_, new_n913_ );
and  ( new_n10831_, new_n10602_, new_n938_ );
or   ( new_n10832_, new_n10831_, new_n10830_ );
and  ( new_n10833_, new_n10832_, new_n10829_ );
or   ( new_n10834_, new_n10832_, new_n10829_ );
and  ( new_n10835_, new_n10617_, new_n428_ );
and  ( new_n10836_, new_n10613_, new_n457_ );
or   ( new_n10837_, new_n10836_, new_n10835_ );
and  ( new_n10838_, new_n10837_, new_n10834_ );
or   ( new_n10839_, new_n10838_, new_n10833_ );
and  ( new_n10840_, new_n10839_, new_n10826_ );
or   ( new_n10841_, new_n10839_, new_n10826_ );
and  ( new_n10842_, new_n10630_, new_n590_ );
and  ( new_n10843_, new_n10626_, new_n619_ );
or   ( new_n10844_, new_n10843_, new_n10842_ );
and  ( new_n10845_, new_n10844_, new_n10841_ );
or   ( new_n10846_, new_n10845_, new_n10840_ );
and  ( new_n10847_, new_n10641_, new_n5182_ );
and  ( new_n10848_, new_n10637_, new_n5028_ );
or   ( new_n10849_, new_n10848_, new_n10847_ );
and  ( new_n10850_, new_n10650_, new_n4400_ );
and  ( new_n10851_, new_n10646_, new_n4215_ );
or   ( new_n10852_, new_n10851_, new_n10850_ );
and  ( new_n10853_, new_n10852_, new_n10849_ );
or   ( new_n10854_, new_n10852_, new_n10849_ );
and  ( new_n10855_, new_n10661_, new_n3695_ );
and  ( new_n10856_, new_n10657_, new_n3548_ );
or   ( new_n10857_, new_n10856_, new_n10855_ );
and  ( new_n10858_, new_n10857_, new_n10854_ );
or   ( new_n10859_, new_n10858_, new_n10853_ );
and  ( new_n10860_, new_n10672_, new_n5858_ );
and  ( new_n10861_, new_n10668_, new_n6037_ );
or   ( new_n10862_, new_n10861_, new_n10860_ );
or   ( new_n10863_, new_n10862_, new_n619_ );
and  ( new_n10864_, new_n10862_, new_n619_ );
and  ( new_n10865_, new_n10683_, new_n6039_ );
and  ( new_n10866_, new_n10679_, new_n5867_ );
or   ( new_n10867_, new_n10866_, new_n10865_ );
or   ( new_n10868_, new_n10867_, new_n10864_ );
and  ( new_n10869_, new_n10868_, new_n10863_ );
or   ( new_n10870_, new_n10869_, new_n10859_ );
and  ( new_n10871_, new_n10869_, new_n10859_ );
and  ( new_n10872_, new_n10696_, new_n3004_ );
and  ( new_n10873_, new_n10692_, new_n2868_ );
or   ( new_n10874_, new_n10873_, new_n10872_ );
and  ( new_n10875_, new_n10705_, new_n2334_ );
and  ( new_n10876_, new_n10701_, new_n2168_ );
or   ( new_n10877_, new_n10876_, new_n10875_ );
and  ( new_n10878_, new_n10877_, new_n10874_ );
or   ( new_n10879_, new_n10877_, new_n10874_ );
and  ( new_n10880_, new_n10716_, new_n1824_ );
and  ( new_n10881_, new_n10712_, new_n1717_ );
or   ( new_n10882_, new_n10881_, new_n10880_ );
and  ( new_n10883_, new_n10882_, new_n10879_ );
or   ( new_n10884_, new_n10883_, new_n10878_ );
or   ( new_n10885_, new_n10884_, new_n10871_ );
and  ( new_n10886_, new_n10885_, new_n10870_ );
or   ( new_n10887_, new_n10886_, new_n10846_ );
and  ( new_n10888_, new_n10886_, new_n10846_ );
and  ( new_n10889_, new_n10729_, new_n10278_ );
and  ( new_n10890_, new_n10725_, new_n10446_ );
or   ( new_n10891_, new_n10890_, new_n10889_ );
and  ( new_n10892_, new_n10736_, new_n10238_ );
and  ( new_n10893_, new_n10732_, new_n10428_ );
or   ( new_n10894_, new_n10893_, new_n10892_ );
and  ( new_n10895_, new_n10894_, new_n10891_ );
or   ( new_n10896_, new_n10894_, new_n10891_ );
and  ( new_n10897_, new_n10745_, new_n10205_ );
and  ( new_n10898_, new_n10741_, new_n10413_ );
or   ( new_n10899_, new_n10898_, new_n10897_ );
and  ( new_n10900_, new_n10899_, new_n10896_ );
or   ( new_n10901_, new_n10900_, new_n10895_ );
or   ( new_n10902_, new_n10901_, new_n10888_ );
and  ( new_n10903_, new_n10902_, new_n10887_ );
or   ( new_n10904_, new_n10903_, new_n10819_ );
and  ( new_n10905_, new_n10903_, new_n10819_ );
and  ( new_n10906_, new_n10758_, new_n9843_ );
and  ( new_n10907_, new_n10754_, new_n10057_ );
or   ( new_n10908_, new_n10907_, new_n10906_ );
or   ( new_n10909_, new_n10908_, new_n10905_ );
and  ( new_n10910_, new_n10909_, new_n10904_ );
or   ( new_n10911_, new_n10910_, new_n10806_ );
and  ( new_n10912_, new_n10910_, new_n10806_ );
and  ( new_n10913_, new_n10769_, new_n9772_ );
and  ( new_n10914_, new_n10765_, new_n10024_ );
or   ( new_n10915_, new_n10914_, new_n10913_ );
or   ( new_n10916_, new_n10915_, new_n10912_ );
and  ( new_n10917_, new_n10916_, new_n10911_ );
and  ( new_n10918_, new_n10917_, new_n10793_ );
or   ( new_n10919_, new_n10918_, new_n10774_ );
and  ( new_n10920_, new_n10919_, new_n10782_ );
and  ( new_n10921_, new_n10917_, new_n10525_ );
and  ( new_n10922_, new_n10793_, new_n10773_ );
or   ( new_n10923_, new_n10922_, new_n10921_ );
and  ( new_n10924_, new_n10780_, new_n10365_ );
and  ( new_n10925_, new_n10776_, new_n10497_ );
or   ( new_n10926_, new_n10925_, new_n10924_ );
and  ( new_n10927_, new_n10926_, new_n10923_ );
or   ( new_n10928_, new_n10927_, new_n10920_ );
and  ( new_n10929_, new_n10524_, new_n10517_ );
or   ( new_n10930_, new_n10929_, new_n10793_ );
or   ( new_n10931_, new_n10800_, new_n10540_ );
and  ( new_n10932_, new_n10931_, new_n10548_ );
and  ( new_n10933_, new_n10796_, new_n10539_ );
and  ( new_n10934_, new_n10799_, new_n10532_ );
or   ( new_n10935_, new_n10934_, new_n10933_ );
and  ( new_n10936_, new_n10935_, new_n10804_ );
or   ( new_n10937_, new_n10936_, new_n10932_ );
or   ( new_n10938_, new_n7105_, new_n859_ );
or   ( new_n10939_, new_n7099_, new_n105_ );
and  ( new_n10940_, new_n10939_, new_n10938_ );
and  ( new_n10941_, new_n10940_, new_n5858_ );
and  ( new_n10942_, new_n7104_, RI2b1c4342d8a0_73 );
and  ( new_n10943_, new_n7110_, RI2b1c4342d918_74 );
or   ( new_n10944_, new_n10943_, new_n10942_ );
and  ( new_n10945_, new_n10944_, new_n6037_ );
or   ( new_n10946_, new_n10945_, new_n10941_ );
or   ( new_n10947_, new_n6156_, new_n886_ );
or   ( new_n10948_, new_n6160_, new_n843_ );
and  ( new_n10949_, new_n10948_, new_n10947_ );
and  ( new_n10950_, new_n10949_, new_n6039_ );
and  ( new_n10951_, new_n6164_, RI2b1c4342da08_76 );
and  ( new_n10952_, new_n6154_, RI2b1c4342d990_75 );
or   ( new_n10953_, new_n10952_, new_n10951_ );
and  ( new_n10954_, new_n10953_, new_n5867_ );
or   ( new_n10955_, new_n10954_, new_n10950_ );
and  ( new_n10956_, new_n10955_, new_n10946_ );
or   ( new_n10957_, new_n10955_, new_n10946_ );
or   ( new_n10958_, new_n5308_, new_n1002_ );
or   ( new_n10959_, new_n5312_, new_n1004_ );
and  ( new_n10960_, new_n10959_, new_n10958_ );
and  ( new_n10961_, new_n10960_, new_n5182_ );
and  ( new_n10962_, new_n5316_, RI2b1c4342daf8_78 );
and  ( new_n10963_, new_n5306_, RI2b1c4342da80_77 );
or   ( new_n10964_, new_n10963_, new_n10962_ );
and  ( new_n10965_, new_n10964_, new_n5028_ );
or   ( new_n10966_, new_n10965_, new_n10961_ );
and  ( new_n10967_, new_n10966_, new_n10957_ );
or   ( new_n10968_, new_n10967_, new_n10956_ );
or   ( new_n10969_, new_n4535_, new_n1511_ );
or   ( new_n10970_, new_n4539_, new_n1310_ );
and  ( new_n10971_, new_n10970_, new_n10969_ );
and  ( new_n10972_, new_n10971_, new_n4400_ );
and  ( new_n10973_, new_n4543_, RI2b1c4342dbe8_80 );
and  ( new_n10974_, new_n4533_, RI2b1c4342db70_79 );
or   ( new_n10975_, new_n10974_, new_n10973_ );
and  ( new_n10976_, new_n10975_, new_n4215_ );
or   ( new_n10977_, new_n10976_, new_n10972_ );
or   ( new_n10978_, new_n3802_, new_n2119_ );
or   ( new_n10979_, new_n3806_, new_n126_ );
and  ( new_n10980_, new_n10979_, new_n10978_ );
and  ( new_n10981_, new_n10980_, new_n3695_ );
and  ( new_n10982_, new_n3810_, RI2b1c4342dcd8_82 );
and  ( new_n10983_, new_n3800_, RI2b1c4342dc60_81 );
or   ( new_n10984_, new_n10983_, new_n10982_ );
and  ( new_n10985_, new_n10984_, new_n3548_ );
or   ( new_n10986_, new_n10985_, new_n10981_ );
and  ( new_n10987_, new_n10986_, new_n10977_ );
or   ( new_n10988_, new_n10986_, new_n10977_ );
or   ( new_n10989_, new_n3112_, new_n2541_ );
or   ( new_n10990_, new_n3116_, new_n121_ );
and  ( new_n10991_, new_n10990_, new_n10989_ );
and  ( new_n10992_, new_n10991_, new_n3004_ );
and  ( new_n10993_, new_n3120_, RI2b1c4342ddc8_84 );
and  ( new_n10994_, new_n3110_, RI2b1c4342dd50_83 );
or   ( new_n10995_, new_n10994_, new_n10993_ );
and  ( new_n10996_, new_n10995_, new_n2868_ );
or   ( new_n10997_, new_n10996_, new_n10992_ );
and  ( new_n10998_, new_n10997_, new_n10988_ );
or   ( new_n10999_, new_n10998_, new_n10987_ );
and  ( new_n11000_, new_n10999_, new_n10968_ );
or   ( new_n11001_, new_n10999_, new_n10968_ );
or   ( new_n11002_, new_n2450_, new_n3239_ );
or   ( new_n11003_, new_n2454_, new_n2806_ );
and  ( new_n11004_, new_n11003_, new_n11002_ );
and  ( new_n11005_, new_n11004_, new_n2334_ );
and  ( new_n11006_, new_n2458_, RI2b1c4342deb8_86 );
and  ( new_n11007_, new_n2448_, RI2b1c4342de40_85 );
or   ( new_n11008_, new_n11007_, new_n11006_ );
and  ( new_n11009_, new_n11008_, new_n2168_ );
or   ( new_n11010_, new_n11009_, new_n11005_ );
or   ( new_n11011_, new_n1910_, new_n3902_ );
or   ( new_n11012_, new_n1914_, new_n3924_ );
and  ( new_n11013_, new_n11012_, new_n11011_ );
and  ( new_n11014_, new_n11013_, new_n1824_ );
and  ( new_n11015_, new_n1918_, RI2b1c4342dfa8_88 );
and  ( new_n11016_, new_n1908_, RI2b1c4342df30_87 );
or   ( new_n11017_, new_n11016_, new_n11015_ );
and  ( new_n11018_, new_n11017_, new_n1717_ );
or   ( new_n11019_, new_n11018_, new_n11014_ );
and  ( new_n11020_, new_n11019_, new_n11010_ );
or   ( new_n11021_, new_n11019_, new_n11010_ );
or   ( new_n11022_, new_n1425_, new_n4635_ );
or   ( new_n11023_, new_n1429_, new_n132_ );
and  ( new_n11024_, new_n11023_, new_n11022_ );
and  ( new_n11025_, new_n11024_, new_n1355_ );
and  ( new_n11026_, new_n1433_, RI2b1c4342e098_90 );
and  ( new_n11027_, new_n1423_, RI2b1c4342e020_89 );
or   ( new_n11028_, new_n11027_, new_n11026_ );
and  ( new_n11029_, new_n11028_, new_n1267_ );
or   ( new_n11030_, new_n11029_, new_n11025_ );
and  ( new_n11031_, new_n11030_, new_n11021_ );
or   ( new_n11032_, new_n11031_, new_n11020_ );
and  ( new_n11033_, new_n11032_, new_n11001_ );
or   ( new_n11034_, new_n11033_, new_n11000_ );
and  ( new_n11035_, new_n10589_, new_n10584_ );
or   ( new_n11036_, new_n11035_, new_n10826_ );
or   ( new_n11037_, new_n934_, new_n5459_ );
or   ( new_n11038_, new_n940_, new_n117_ );
and  ( new_n11039_, new_n11038_, new_n11037_ );
and  ( new_n11040_, new_n11039_, new_n913_ );
and  ( new_n11041_, new_n944_, RI2b1c4342e188_92 );
and  ( new_n11042_, new_n932_, RI2b1c4342e110_91 );
or   ( new_n11043_, new_n11042_, new_n11041_ );
and  ( new_n11044_, new_n11043_, new_n938_ );
or   ( new_n11045_, new_n11044_, new_n11040_ );
or   ( new_n11046_, new_n453_, new_n6321_ );
or   ( new_n11047_, new_n459_, new_n6307_ );
and  ( new_n11048_, new_n11047_, new_n11046_ );
and  ( new_n11049_, new_n11048_, new_n428_ );
and  ( new_n11050_, new_n463_, RI2b1c4342e278_94 );
and  ( new_n11051_, new_n451_, RI2b1c4342e200_93 );
or   ( new_n11052_, new_n11051_, new_n11050_ );
and  ( new_n11053_, new_n11052_, new_n457_ );
or   ( new_n11054_, new_n11053_, new_n11049_ );
and  ( new_n11055_, new_n11054_, new_n11045_ );
or   ( new_n11056_, new_n11054_, new_n11045_ );
or   ( new_n11057_, new_n524_, new_n7274_ );
or   ( new_n11058_, new_n528_, new_n124_ );
and  ( new_n11059_, new_n11058_, new_n11057_ );
and  ( new_n11060_, new_n11059_, new_n505_ );
and  ( new_n11061_, new_n537_, RI2b1c4342e368_96 );
and  ( new_n11062_, new_n522_, RI2b1c4342e2f0_95 );
or   ( new_n11063_, new_n11062_, new_n11061_ );
and  ( new_n11064_, new_n11063_, new_n533_ );
or   ( new_n11065_, new_n11064_, new_n11060_ );
and  ( new_n11066_, new_n11065_, new_n11056_ );
or   ( new_n11067_, new_n11066_, new_n11055_ );
and  ( new_n11068_, new_n11067_, new_n11036_ );
or   ( new_n11069_, new_n11067_, new_n11036_ );
or   ( new_n11070_, new_n10833_, new_n10609_ );
and  ( new_n11071_, new_n11070_, new_n10619_ );
and  ( new_n11072_, new_n10829_, new_n10608_ );
and  ( new_n11073_, new_n10832_, new_n10599_ );
or   ( new_n11074_, new_n11073_, new_n11072_ );
and  ( new_n11075_, new_n11074_, new_n10837_ );
or   ( new_n11076_, new_n11075_, new_n11071_ );
and  ( new_n11077_, new_n11076_, new_n11069_ );
or   ( new_n11078_, new_n11077_, new_n11068_ );
and  ( new_n11079_, new_n11078_, new_n11034_ );
or   ( new_n11080_, new_n11078_, new_n11034_ );
or   ( new_n11081_, new_n10878_, new_n10708_ );
and  ( new_n11082_, new_n11081_, new_n10718_ );
and  ( new_n11083_, new_n10874_, new_n10707_ );
and  ( new_n11084_, new_n10877_, new_n10698_ );
or   ( new_n11085_, new_n11084_, new_n11083_ );
and  ( new_n11086_, new_n11085_, new_n10882_ );
or   ( new_n11087_, new_n11086_, new_n11082_ );
or   ( new_n11088_, new_n10853_, new_n10653_ );
and  ( new_n11089_, new_n11088_, new_n10663_ );
and  ( new_n11090_, new_n10849_, new_n10652_ );
and  ( new_n11091_, new_n10852_, new_n10643_ );
or   ( new_n11092_, new_n11091_, new_n11090_ );
and  ( new_n11093_, new_n11092_, new_n10857_ );
or   ( new_n11094_, new_n11093_, new_n11089_ );
and  ( new_n11095_, new_n11094_, new_n11087_ );
or   ( new_n11096_, new_n11094_, new_n11087_ );
or   ( new_n11097_, new_n10864_, new_n10675_ );
and  ( new_n11098_, new_n11097_, new_n10685_ );
and  ( new_n11099_, new_n10674_, new_n619_ );
and  ( new_n11100_, new_n10862_, new_n590_ );
or   ( new_n11101_, new_n11100_, new_n11099_ );
and  ( new_n11102_, new_n11101_, new_n10867_ );
or   ( new_n11103_, new_n11102_, new_n11098_ );
and  ( new_n11104_, new_n11103_, new_n11096_ );
or   ( new_n11105_, new_n11104_, new_n11095_ );
and  ( new_n11106_, new_n11105_, new_n11080_ );
or   ( new_n11107_, new_n11106_, new_n11079_ );
or   ( new_n11108_, new_n10396_, new_n10164_ );
and  ( new_n11109_, new_n11108_, new_n10174_ );
and  ( new_n11110_, new_n10392_, new_n10163_ );
and  ( new_n11111_, new_n10395_, new_n10154_ );
or   ( new_n11112_, new_n11111_, new_n11110_ );
and  ( new_n11113_, new_n11112_, new_n10400_ );
or   ( new_n11114_, new_n11113_, new_n11109_ );
or   ( new_n11115_, new_n10895_, new_n10739_ );
and  ( new_n11116_, new_n11115_, new_n10747_ );
and  ( new_n11117_, new_n10891_, new_n10738_ );
and  ( new_n11118_, new_n10894_, new_n10731_ );
or   ( new_n11119_, new_n11118_, new_n11117_ );
and  ( new_n11120_, new_n11119_, new_n10899_ );
or   ( new_n11121_, new_n11120_, new_n11116_ );
and  ( new_n11122_, new_n11121_, new_n11114_ );
or   ( new_n11123_, new_n11121_, new_n11114_ );
or   ( new_n11124_, new_n10840_, new_n10622_ );
and  ( new_n11125_, new_n11124_, new_n10632_ );
and  ( new_n11126_, new_n10839_, new_n10590_ );
and  ( new_n11127_, new_n10826_, new_n10621_ );
or   ( new_n11128_, new_n11127_, new_n11126_ );
and  ( new_n11129_, new_n11128_, new_n10844_ );
or   ( new_n11130_, new_n11129_, new_n11125_ );
and  ( new_n11131_, new_n11130_, new_n11123_ );
or   ( new_n11132_, new_n11131_, new_n11122_ );
and  ( new_n11133_, new_n11132_, new_n11107_ );
or   ( new_n11134_, new_n11132_, new_n11107_ );
or   ( new_n11135_, new_n10813_, new_n10565_ );
and  ( new_n11136_, new_n11135_, new_n10573_ );
and  ( new_n11137_, new_n10809_, new_n10564_ );
and  ( new_n11138_, new_n10812_, new_n10557_ );
or   ( new_n11139_, new_n11138_, new_n11137_ );
and  ( new_n11140_, new_n11139_, new_n10817_ );
or   ( new_n11141_, new_n11140_, new_n11136_ );
and  ( new_n11142_, new_n11141_, new_n11134_ );
or   ( new_n11143_, new_n11142_, new_n11133_ );
and  ( new_n11144_, new_n11143_, new_n10937_ );
or   ( new_n11145_, new_n11143_, new_n10937_ );
or   ( new_n11146_, new_n10905_, new_n10752_ );
and  ( new_n11147_, new_n11146_, new_n10760_ );
and  ( new_n11148_, new_n10903_, new_n10575_ );
and  ( new_n11149_, new_n10819_, new_n10751_ );
or   ( new_n11150_, new_n11149_, new_n11148_ );
and  ( new_n11151_, new_n11150_, new_n10908_ );
or   ( new_n11152_, new_n11151_, new_n11147_ );
and  ( new_n11153_, new_n11152_, new_n11145_ );
or   ( new_n11154_, new_n11153_, new_n11144_ );
and  ( new_n11155_, new_n11154_, new_n10930_ );
or   ( new_n11156_, new_n11154_, new_n10930_ );
or   ( new_n11157_, new_n10912_, new_n10763_ );
and  ( new_n11158_, new_n11157_, new_n10771_ );
and  ( new_n11159_, new_n10910_, new_n10550_ );
and  ( new_n11160_, new_n10806_, new_n10762_ );
or   ( new_n11161_, new_n11160_, new_n11159_ );
and  ( new_n11162_, new_n11161_, new_n10915_ );
or   ( new_n11163_, new_n11162_, new_n11158_ );
and  ( new_n11164_, new_n11163_, new_n11156_ );
or   ( new_n11165_, new_n11164_, new_n11155_ );
or   ( new_n11166_, new_n11165_, new_n10928_ );
and  ( new_n11167_, new_n11166_, new_n10786_ );
or   ( new_n11168_, new_n11167_, new_n10785_ );
or   ( new_n11169_, new_n11168_, new_n10383_ );
and  ( new_n11170_, new_n11169_, new_n10381_ );
or   ( new_n11171_, new_n11170_, new_n9592_ );
and  ( new_n11172_, new_n11171_, new_n9589_ );
and  ( new_n11173_, new_n11165_, new_n10928_ );
or   ( new_n11174_, new_n11173_, new_n10785_ );
or   ( new_n11175_, new_n11174_, new_n10383_ );
and  ( new_n11176_, new_n10789_, new_n10524_ );
and  ( new_n11177_, new_n10792_, new_n10517_ );
or   ( new_n11178_, new_n11177_, new_n11176_ );
and  ( new_n11179_, new_n10935_, new_n10548_ );
and  ( new_n11180_, new_n10931_, new_n10804_ );
or   ( new_n11181_, new_n11180_, new_n11179_ );
and  ( new_n11182_, new_n10944_, new_n5858_ );
and  ( new_n11183_, new_n10940_, new_n6037_ );
or   ( new_n11184_, new_n11183_, new_n11182_ );
and  ( new_n11185_, new_n10953_, new_n6039_ );
and  ( new_n11186_, new_n10949_, new_n5867_ );
or   ( new_n11187_, new_n11186_, new_n11185_ );
and  ( new_n11188_, new_n11187_, new_n11184_ );
or   ( new_n11189_, new_n11187_, new_n11184_ );
and  ( new_n11190_, new_n10964_, new_n5182_ );
and  ( new_n11191_, new_n10960_, new_n5028_ );
or   ( new_n11192_, new_n11191_, new_n11190_ );
and  ( new_n11193_, new_n11192_, new_n11189_ );
or   ( new_n11194_, new_n11193_, new_n11188_ );
and  ( new_n11195_, new_n10975_, new_n4400_ );
and  ( new_n11196_, new_n10971_, new_n4215_ );
or   ( new_n11197_, new_n11196_, new_n11195_ );
and  ( new_n11198_, new_n10984_, new_n3695_ );
and  ( new_n11199_, new_n10980_, new_n3548_ );
or   ( new_n11200_, new_n11199_, new_n11198_ );
and  ( new_n11201_, new_n11200_, new_n11197_ );
or   ( new_n11202_, new_n11200_, new_n11197_ );
and  ( new_n11203_, new_n10995_, new_n3004_ );
and  ( new_n11204_, new_n10991_, new_n2868_ );
or   ( new_n11205_, new_n11204_, new_n11203_ );
and  ( new_n11206_, new_n11205_, new_n11202_ );
or   ( new_n11207_, new_n11206_, new_n11201_ );
and  ( new_n11208_, new_n11207_, new_n11194_ );
or   ( new_n11209_, new_n11207_, new_n11194_ );
and  ( new_n11210_, new_n11008_, new_n2334_ );
and  ( new_n11211_, new_n11004_, new_n2168_ );
or   ( new_n11212_, new_n11211_, new_n11210_ );
and  ( new_n11213_, new_n11017_, new_n1824_ );
and  ( new_n11214_, new_n11013_, new_n1717_ );
or   ( new_n11215_, new_n11214_, new_n11213_ );
and  ( new_n11216_, new_n11215_, new_n11212_ );
or   ( new_n11217_, new_n11215_, new_n11212_ );
and  ( new_n11218_, new_n11028_, new_n1355_ );
and  ( new_n11219_, new_n11024_, new_n1267_ );
or   ( new_n11220_, new_n11219_, new_n11218_ );
and  ( new_n11221_, new_n11220_, new_n11217_ );
or   ( new_n11222_, new_n11221_, new_n11216_ );
and  ( new_n11223_, new_n11222_, new_n11209_ );
or   ( new_n11224_, new_n11223_, new_n11208_ );
and  ( new_n11225_, new_n10822_, new_n10589_ );
and  ( new_n11226_, new_n10825_, new_n10584_ );
or   ( new_n11227_, new_n11226_, new_n11225_ );
and  ( new_n11228_, new_n11043_, new_n913_ );
and  ( new_n11229_, new_n11039_, new_n938_ );
or   ( new_n11230_, new_n11229_, new_n11228_ );
and  ( new_n11231_, new_n11052_, new_n428_ );
and  ( new_n11232_, new_n11048_, new_n457_ );
or   ( new_n11233_, new_n11232_, new_n11231_ );
and  ( new_n11234_, new_n11233_, new_n11230_ );
or   ( new_n11235_, new_n11233_, new_n11230_ );
and  ( new_n11236_, new_n11063_, new_n505_ );
and  ( new_n11237_, new_n11059_, new_n533_ );
or   ( new_n11238_, new_n11237_, new_n11236_ );
and  ( new_n11239_, new_n11238_, new_n11235_ );
or   ( new_n11240_, new_n11239_, new_n11234_ );
and  ( new_n11241_, new_n11240_, new_n11227_ );
or   ( new_n11242_, new_n11240_, new_n11227_ );
and  ( new_n11243_, new_n11074_, new_n10619_ );
and  ( new_n11244_, new_n11070_, new_n10837_ );
or   ( new_n11245_, new_n11244_, new_n11243_ );
and  ( new_n11246_, new_n11245_, new_n11242_ );
or   ( new_n11247_, new_n11246_, new_n11241_ );
and  ( new_n11248_, new_n11247_, new_n11224_ );
or   ( new_n11249_, new_n11247_, new_n11224_ );
and  ( new_n11250_, new_n11085_, new_n10718_ );
and  ( new_n11251_, new_n11081_, new_n10882_ );
or   ( new_n11252_, new_n11251_, new_n11250_ );
and  ( new_n11253_, new_n11092_, new_n10663_ );
and  ( new_n11254_, new_n11088_, new_n10857_ );
or   ( new_n11255_, new_n11254_, new_n11253_ );
and  ( new_n11256_, new_n11255_, new_n11252_ );
or   ( new_n11257_, new_n11255_, new_n11252_ );
and  ( new_n11258_, new_n11101_, new_n10685_ );
and  ( new_n11259_, new_n11097_, new_n10867_ );
or   ( new_n11260_, new_n11259_, new_n11258_ );
and  ( new_n11261_, new_n11260_, new_n11257_ );
or   ( new_n11262_, new_n11261_, new_n11256_ );
and  ( new_n11263_, new_n11262_, new_n11249_ );
or   ( new_n11264_, new_n11263_, new_n11248_ );
and  ( new_n11265_, new_n11112_, new_n10174_ );
and  ( new_n11266_, new_n11108_, new_n10400_ );
or   ( new_n11267_, new_n11266_, new_n11265_ );
and  ( new_n11268_, new_n11119_, new_n10747_ );
and  ( new_n11269_, new_n11115_, new_n10899_ );
or   ( new_n11270_, new_n11269_, new_n11268_ );
and  ( new_n11271_, new_n11270_, new_n11267_ );
or   ( new_n11272_, new_n11270_, new_n11267_ );
and  ( new_n11273_, new_n11128_, new_n10632_ );
and  ( new_n11274_, new_n11124_, new_n10844_ );
or   ( new_n11275_, new_n11274_, new_n11273_ );
and  ( new_n11276_, new_n11275_, new_n11272_ );
or   ( new_n11277_, new_n11276_, new_n11271_ );
and  ( new_n11278_, new_n11277_, new_n11264_ );
or   ( new_n11279_, new_n11277_, new_n11264_ );
and  ( new_n11280_, new_n11139_, new_n10573_ );
and  ( new_n11281_, new_n11135_, new_n10817_ );
or   ( new_n11282_, new_n11281_, new_n11280_ );
and  ( new_n11283_, new_n11282_, new_n11279_ );
or   ( new_n11284_, new_n11283_, new_n11278_ );
and  ( new_n11285_, new_n11284_, new_n11181_ );
or   ( new_n11286_, new_n11284_, new_n11181_ );
and  ( new_n11287_, new_n11150_, new_n10760_ );
and  ( new_n11288_, new_n11146_, new_n10908_ );
or   ( new_n11289_, new_n11288_, new_n11287_ );
and  ( new_n11290_, new_n11289_, new_n11286_ );
or   ( new_n11291_, new_n11290_, new_n11285_ );
and  ( new_n11292_, new_n11291_, new_n11178_ );
or   ( new_n11293_, new_n11292_, new_n11155_ );
and  ( new_n11294_, new_n11293_, new_n11163_ );
and  ( new_n11295_, new_n11291_, new_n10930_ );
and  ( new_n11296_, new_n11178_, new_n11154_ );
or   ( new_n11297_, new_n11296_, new_n11295_ );
and  ( new_n11298_, new_n11161_, new_n10771_ );
and  ( new_n11299_, new_n11157_, new_n10915_ );
or   ( new_n11300_, new_n11299_, new_n11298_ );
and  ( new_n11301_, new_n11300_, new_n11297_ );
or   ( new_n11302_, new_n11301_, new_n11294_ );
or   ( new_n11303_, new_n11285_, new_n11144_ );
and  ( new_n11304_, new_n11303_, new_n11152_ );
and  ( new_n11305_, new_n11284_, new_n10937_ );
and  ( new_n11306_, new_n11181_, new_n11143_ );
or   ( new_n11307_, new_n11306_, new_n11305_ );
and  ( new_n11308_, new_n11307_, new_n11289_ );
or   ( new_n11309_, new_n11308_, new_n11304_ );
or   ( new_n11310_, new_n11271_, new_n11122_ );
and  ( new_n11311_, new_n11310_, new_n11130_ );
and  ( new_n11312_, new_n11267_, new_n11121_ );
and  ( new_n11313_, new_n11270_, new_n11114_ );
or   ( new_n11314_, new_n11313_, new_n11312_ );
and  ( new_n11315_, new_n11314_, new_n11275_ );
or   ( new_n11316_, new_n11315_, new_n11311_ );
or   ( new_n11317_, new_n11248_, new_n11079_ );
and  ( new_n11318_, new_n11317_, new_n11105_ );
and  ( new_n11319_, new_n11224_, new_n11078_ );
and  ( new_n11320_, new_n11247_, new_n11034_ );
or   ( new_n11321_, new_n11320_, new_n11319_ );
and  ( new_n11322_, new_n11321_, new_n11262_ );
or   ( new_n11323_, new_n11322_, new_n11318_ );
or   ( new_n11324_, new_n11323_, new_n11316_ );
or   ( new_n11325_, new_n11256_, new_n11095_ );
and  ( new_n11326_, new_n11325_, new_n11103_ );
and  ( new_n11327_, new_n11252_, new_n11094_ );
and  ( new_n11328_, new_n11255_, new_n11087_ );
or   ( new_n11329_, new_n11328_, new_n11327_ );
and  ( new_n11330_, new_n11329_, new_n11260_ );
or   ( new_n11331_, new_n11330_, new_n11326_ );
or   ( new_n11332_, new_n11241_, new_n11068_ );
and  ( new_n11333_, new_n11332_, new_n11076_ );
and  ( new_n11334_, new_n11240_, new_n11036_ );
and  ( new_n11335_, new_n11227_, new_n11067_ );
or   ( new_n11336_, new_n11335_, new_n11334_ );
and  ( new_n11337_, new_n11336_, new_n11245_ );
or   ( new_n11338_, new_n11337_, new_n11333_ );
and  ( new_n11339_, new_n11338_, new_n11331_ );
or   ( new_n11340_, new_n11338_, new_n11331_ );
or   ( new_n11341_, new_n11208_, new_n11000_ );
and  ( new_n11342_, new_n11341_, new_n11032_ );
and  ( new_n11343_, new_n11194_, new_n10999_ );
and  ( new_n11344_, new_n11207_, new_n10968_ );
or   ( new_n11345_, new_n11344_, new_n11343_ );
and  ( new_n11346_, new_n11345_, new_n11222_ );
or   ( new_n11347_, new_n11346_, new_n11342_ );
and  ( new_n11348_, new_n11347_, new_n11340_ );
or   ( new_n11349_, new_n11348_, new_n11339_ );
or   ( new_n11350_, new_n11234_, new_n11055_ );
and  ( new_n11351_, new_n11350_, new_n11065_ );
and  ( new_n11352_, new_n11230_, new_n11054_ );
and  ( new_n11353_, new_n11233_, new_n11045_ );
or   ( new_n11354_, new_n11353_, new_n11352_ );
and  ( new_n11355_, new_n11354_, new_n11238_ );
or   ( new_n11356_, new_n11355_, new_n11351_ );
or   ( new_n11357_, new_n1425_, new_n117_ );
or   ( new_n11358_, new_n1429_, new_n4635_ );
and  ( new_n11359_, new_n11358_, new_n11357_ );
and  ( new_n11360_, new_n11359_, new_n1355_ );
and  ( new_n11361_, new_n1433_, RI2b1c4342e110_91 );
and  ( new_n11362_, new_n1423_, RI2b1c4342e098_90 );
or   ( new_n11363_, new_n11362_, new_n11361_ );
and  ( new_n11364_, new_n11363_, new_n1267_ );
or   ( new_n11365_, new_n11364_, new_n11360_ );
or   ( new_n11366_, new_n934_, new_n6307_ );
or   ( new_n11367_, new_n940_, new_n5459_ );
and  ( new_n11368_, new_n11367_, new_n11366_ );
and  ( new_n11369_, new_n11368_, new_n913_ );
and  ( new_n11370_, new_n944_, RI2b1c4342e200_93 );
and  ( new_n11371_, new_n932_, RI2b1c4342e188_92 );
or   ( new_n11372_, new_n11371_, new_n11370_ );
and  ( new_n11373_, new_n11372_, new_n938_ );
or   ( new_n11374_, new_n11373_, new_n11369_ );
and  ( new_n11375_, new_n11374_, new_n11365_ );
or   ( new_n11376_, new_n11374_, new_n11365_ );
or   ( new_n11377_, new_n453_, new_n124_ );
or   ( new_n11378_, new_n459_, new_n6321_ );
and  ( new_n11379_, new_n11378_, new_n11377_ );
and  ( new_n11380_, new_n11379_, new_n428_ );
and  ( new_n11381_, new_n463_, RI2b1c4342e2f0_95 );
and  ( new_n11382_, new_n451_, RI2b1c4342e278_94 );
or   ( new_n11383_, new_n11382_, new_n11381_ );
and  ( new_n11384_, new_n11383_, new_n457_ );
or   ( new_n11385_, new_n11384_, new_n11380_ );
and  ( new_n11386_, new_n11385_, new_n11376_ );
or   ( new_n11387_, new_n11386_, new_n11375_ );
and  ( new_n11388_, new_n11387_, new_n11356_ );
or   ( new_n11389_, new_n11387_, new_n11356_ );
or   ( new_n11390_, new_n11216_, new_n11020_ );
and  ( new_n11391_, new_n11390_, new_n11030_ );
and  ( new_n11392_, new_n11212_, new_n11019_ );
and  ( new_n11393_, new_n11215_, new_n11010_ );
or   ( new_n11394_, new_n11393_, new_n11392_ );
and  ( new_n11395_, new_n11394_, new_n11220_ );
or   ( new_n11396_, new_n11395_, new_n11391_ );
and  ( new_n11397_, new_n11396_, new_n11389_ );
or   ( new_n11398_, new_n11397_, new_n11388_ );
or   ( new_n11399_, new_n5308_, new_n1310_ );
or   ( new_n11400_, new_n5312_, new_n1002_ );
and  ( new_n11401_, new_n11400_, new_n11399_ );
and  ( new_n11402_, new_n11401_, new_n5182_ );
and  ( new_n11403_, new_n5316_, RI2b1c4342db70_79 );
and  ( new_n11404_, new_n5306_, RI2b1c4342daf8_78 );
or   ( new_n11405_, new_n11404_, new_n11403_ );
and  ( new_n11406_, new_n11405_, new_n5028_ );
or   ( new_n11407_, new_n11406_, new_n11402_ );
or   ( new_n11408_, new_n4535_, new_n126_ );
or   ( new_n11409_, new_n4539_, new_n1511_ );
and  ( new_n11410_, new_n11409_, new_n11408_ );
and  ( new_n11411_, new_n11410_, new_n4400_ );
and  ( new_n11412_, new_n4543_, RI2b1c4342dc60_81 );
and  ( new_n11413_, new_n4533_, RI2b1c4342dbe8_80 );
or   ( new_n11414_, new_n11413_, new_n11412_ );
and  ( new_n11415_, new_n11414_, new_n4215_ );
or   ( new_n11416_, new_n11415_, new_n11411_ );
and  ( new_n11417_, new_n11416_, new_n11407_ );
or   ( new_n11418_, new_n11416_, new_n11407_ );
or   ( new_n11419_, new_n3802_, new_n121_ );
or   ( new_n11420_, new_n3806_, new_n2119_ );
and  ( new_n11421_, new_n11420_, new_n11419_ );
and  ( new_n11422_, new_n11421_, new_n3695_ );
and  ( new_n11423_, new_n3810_, RI2b1c4342dd50_83 );
and  ( new_n11424_, new_n3800_, RI2b1c4342dcd8_82 );
or   ( new_n11425_, new_n11424_, new_n11423_ );
and  ( new_n11426_, new_n11425_, new_n3548_ );
or   ( new_n11427_, new_n11426_, new_n11422_ );
and  ( new_n11428_, new_n11427_, new_n11418_ );
or   ( new_n11429_, new_n11428_, new_n11417_ );
or   ( new_n11430_, new_n7105_, new_n843_ );
or   ( new_n11431_, new_n7099_, new_n859_ );
and  ( new_n11432_, new_n11431_, new_n11430_ );
and  ( new_n11433_, new_n11432_, new_n5858_ );
and  ( new_n11434_, new_n7104_, RI2b1c4342d918_74 );
and  ( new_n11435_, new_n7110_, RI2b1c4342d990_75 );
or   ( new_n11436_, new_n11435_, new_n11434_ );
and  ( new_n11437_, new_n11436_, new_n6037_ );
or   ( new_n11438_, new_n11437_, new_n11433_ );
and  ( new_n11439_, new_n11438_, new_n505_ );
or   ( new_n11440_, new_n11438_, new_n505_ );
or   ( new_n11441_, new_n6156_, new_n1004_ );
or   ( new_n11442_, new_n6160_, new_n886_ );
and  ( new_n11443_, new_n11442_, new_n11441_ );
and  ( new_n11444_, new_n11443_, new_n6039_ );
and  ( new_n11445_, new_n6164_, RI2b1c4342da80_77 );
and  ( new_n11446_, new_n6154_, RI2b1c4342da08_76 );
or   ( new_n11447_, new_n11446_, new_n11445_ );
and  ( new_n11448_, new_n11447_, new_n5867_ );
or   ( new_n11449_, new_n11448_, new_n11444_ );
and  ( new_n11450_, new_n11449_, new_n11440_ );
or   ( new_n11451_, new_n11450_, new_n11439_ );
and  ( new_n11452_, new_n11451_, new_n11429_ );
or   ( new_n11453_, new_n11451_, new_n11429_ );
or   ( new_n11454_, new_n3112_, new_n2806_ );
or   ( new_n11455_, new_n3116_, new_n2541_ );
and  ( new_n11456_, new_n11455_, new_n11454_ );
and  ( new_n11457_, new_n11456_, new_n3004_ );
and  ( new_n11458_, new_n3120_, RI2b1c4342de40_85 );
and  ( new_n11459_, new_n3110_, RI2b1c4342ddc8_84 );
or   ( new_n11460_, new_n11459_, new_n11458_ );
and  ( new_n11461_, new_n11460_, new_n2868_ );
or   ( new_n11462_, new_n11461_, new_n11457_ );
or   ( new_n11463_, new_n2450_, new_n3924_ );
or   ( new_n11464_, new_n2454_, new_n3239_ );
and  ( new_n11465_, new_n11464_, new_n11463_ );
and  ( new_n11466_, new_n11465_, new_n2334_ );
and  ( new_n11467_, new_n2458_, RI2b1c4342df30_87 );
and  ( new_n11468_, new_n2448_, RI2b1c4342deb8_86 );
or   ( new_n11469_, new_n11468_, new_n11467_ );
and  ( new_n11470_, new_n11469_, new_n2168_ );
or   ( new_n11471_, new_n11470_, new_n11466_ );
and  ( new_n11472_, new_n11471_, new_n11462_ );
or   ( new_n11473_, new_n11471_, new_n11462_ );
or   ( new_n11474_, new_n1910_, new_n132_ );
or   ( new_n11475_, new_n1914_, new_n3902_ );
and  ( new_n11476_, new_n11475_, new_n11474_ );
and  ( new_n11477_, new_n11476_, new_n1824_ );
and  ( new_n11478_, new_n1918_, RI2b1c4342e020_89 );
and  ( new_n11479_, new_n1908_, RI2b1c4342dfa8_88 );
or   ( new_n11480_, new_n11479_, new_n11478_ );
and  ( new_n11481_, new_n11480_, new_n1717_ );
or   ( new_n11482_, new_n11481_, new_n11477_ );
and  ( new_n11483_, new_n11482_, new_n11473_ );
or   ( new_n11484_, new_n11483_, new_n11472_ );
and  ( new_n11485_, new_n11484_, new_n11453_ );
or   ( new_n11486_, new_n11485_, new_n11452_ );
and  ( new_n11487_, new_n11486_, new_n11398_ );
or   ( new_n11488_, new_n11486_, new_n11398_ );
or   ( new_n11489_, new_n11201_, new_n10987_ );
and  ( new_n11490_, new_n11489_, new_n10997_ );
and  ( new_n11491_, new_n11197_, new_n10986_ );
and  ( new_n11492_, new_n11200_, new_n10977_ );
or   ( new_n11493_, new_n11492_, new_n11491_ );
and  ( new_n11494_, new_n11493_, new_n11205_ );
or   ( new_n11495_, new_n11494_, new_n11490_ );
or   ( new_n11496_, new_n11188_, new_n10956_ );
and  ( new_n11497_, new_n11496_, new_n10966_ );
and  ( new_n11498_, new_n11184_, new_n10955_ );
and  ( new_n11499_, new_n11187_, new_n10946_ );
or   ( new_n11500_, new_n11499_, new_n11498_ );
and  ( new_n11501_, new_n11500_, new_n11192_ );
or   ( new_n11502_, new_n11501_, new_n11497_ );
or   ( new_n11503_, new_n11502_, new_n11495_ );
and  ( new_n11504_, new_n11503_, new_n11488_ );
or   ( new_n11505_, new_n11504_, new_n11487_ );
and  ( new_n11506_, new_n11505_, new_n11349_ );
or   ( new_n11507_, new_n11505_, new_n11349_ );
or   ( new_n11508_, new_n10871_, new_n10688_ );
and  ( new_n11509_, new_n11508_, new_n10720_ );
and  ( new_n11510_, new_n10869_, new_n10665_ );
and  ( new_n11511_, new_n10859_, new_n10687_ );
or   ( new_n11512_, new_n11511_, new_n11510_ );
and  ( new_n11513_, new_n11512_, new_n10884_ );
or   ( new_n11514_, new_n11513_, new_n11509_ );
and  ( new_n11515_, new_n11514_, new_n11507_ );
or   ( new_n11516_, new_n11515_, new_n11506_ );
and  ( new_n11517_, new_n11516_, new_n11324_ );
or   ( new_n11518_, new_n11516_, new_n11324_ );
or   ( new_n11519_, new_n10888_, new_n10723_ );
and  ( new_n11520_, new_n11519_, new_n10749_ );
and  ( new_n11521_, new_n10886_, new_n10634_ );
and  ( new_n11522_, new_n10846_, new_n10722_ );
or   ( new_n11523_, new_n11522_, new_n11521_ );
and  ( new_n11524_, new_n11523_, new_n10901_ );
or   ( new_n11525_, new_n11524_, new_n11520_ );
and  ( new_n11526_, new_n11525_, new_n11518_ );
or   ( new_n11527_, new_n11526_, new_n11517_ );
or   ( new_n11528_, new_n11527_, new_n11309_ );
and  ( new_n11529_, new_n11528_, new_n11302_ );
or   ( new_n11530_, new_n11528_, new_n11302_ );
and  ( new_n11531_, new_n11527_, new_n11309_ );
and  ( new_n11532_, new_n11307_, new_n11152_ );
and  ( new_n11533_, new_n11303_, new_n11289_ );
or   ( new_n11534_, new_n11533_, new_n11532_ );
and  ( new_n11535_, new_n11314_, new_n11130_ );
and  ( new_n11536_, new_n11310_, new_n11275_ );
or   ( new_n11537_, new_n11536_, new_n11535_ );
and  ( new_n11538_, new_n11321_, new_n11105_ );
and  ( new_n11539_, new_n11317_, new_n11262_ );
or   ( new_n11540_, new_n11539_, new_n11538_ );
and  ( new_n11541_, new_n11540_, new_n11537_ );
and  ( new_n11542_, new_n11329_, new_n11103_ );
and  ( new_n11543_, new_n11325_, new_n11260_ );
or   ( new_n11544_, new_n11543_, new_n11542_ );
and  ( new_n11545_, new_n11336_, new_n11076_ );
and  ( new_n11546_, new_n11332_, new_n11245_ );
or   ( new_n11547_, new_n11546_, new_n11545_ );
and  ( new_n11548_, new_n11547_, new_n11544_ );
or   ( new_n11549_, new_n11547_, new_n11544_ );
and  ( new_n11550_, new_n11345_, new_n11032_ );
and  ( new_n11551_, new_n11341_, new_n11222_ );
or   ( new_n11552_, new_n11551_, new_n11550_ );
and  ( new_n11553_, new_n11552_, new_n11549_ );
or   ( new_n11554_, new_n11553_, new_n11548_ );
and  ( new_n11555_, new_n11354_, new_n11065_ );
and  ( new_n11556_, new_n11350_, new_n11238_ );
or   ( new_n11557_, new_n11556_, new_n11555_ );
and  ( new_n11558_, new_n11363_, new_n1355_ );
and  ( new_n11559_, new_n11359_, new_n1267_ );
or   ( new_n11560_, new_n11559_, new_n11558_ );
and  ( new_n11561_, new_n11372_, new_n913_ );
and  ( new_n11562_, new_n11368_, new_n938_ );
or   ( new_n11563_, new_n11562_, new_n11561_ );
and  ( new_n11564_, new_n11563_, new_n11560_ );
or   ( new_n11565_, new_n11563_, new_n11560_ );
and  ( new_n11566_, new_n11383_, new_n428_ );
and  ( new_n11567_, new_n11379_, new_n457_ );
or   ( new_n11568_, new_n11567_, new_n11566_ );
and  ( new_n11569_, new_n11568_, new_n11565_ );
or   ( new_n11570_, new_n11569_, new_n11564_ );
and  ( new_n11571_, new_n11570_, new_n11557_ );
or   ( new_n11572_, new_n11570_, new_n11557_ );
and  ( new_n11573_, new_n11394_, new_n11030_ );
and  ( new_n11574_, new_n11390_, new_n11220_ );
or   ( new_n11575_, new_n11574_, new_n11573_ );
and  ( new_n11576_, new_n11575_, new_n11572_ );
or   ( new_n11577_, new_n11576_, new_n11571_ );
and  ( new_n11578_, new_n11405_, new_n5182_ );
and  ( new_n11579_, new_n11401_, new_n5028_ );
or   ( new_n11580_, new_n11579_, new_n11578_ );
and  ( new_n11581_, new_n11414_, new_n4400_ );
and  ( new_n11582_, new_n11410_, new_n4215_ );
or   ( new_n11583_, new_n11582_, new_n11581_ );
and  ( new_n11584_, new_n11583_, new_n11580_ );
or   ( new_n11585_, new_n11583_, new_n11580_ );
and  ( new_n11586_, new_n11425_, new_n3695_ );
and  ( new_n11587_, new_n11421_, new_n3548_ );
or   ( new_n11588_, new_n11587_, new_n11586_ );
and  ( new_n11589_, new_n11588_, new_n11585_ );
or   ( new_n11590_, new_n11589_, new_n11584_ );
and  ( new_n11591_, new_n11436_, new_n5858_ );
and  ( new_n11592_, new_n11432_, new_n6037_ );
or   ( new_n11593_, new_n11592_, new_n11591_ );
or   ( new_n11594_, new_n11593_, new_n533_ );
and  ( new_n11595_, new_n11593_, new_n533_ );
and  ( new_n11596_, new_n11447_, new_n6039_ );
and  ( new_n11597_, new_n11443_, new_n5867_ );
or   ( new_n11598_, new_n11597_, new_n11596_ );
or   ( new_n11599_, new_n11598_, new_n11595_ );
and  ( new_n11600_, new_n11599_, new_n11594_ );
or   ( new_n11601_, new_n11600_, new_n11590_ );
and  ( new_n11602_, new_n11600_, new_n11590_ );
and  ( new_n11603_, new_n11460_, new_n3004_ );
and  ( new_n11604_, new_n11456_, new_n2868_ );
or   ( new_n11605_, new_n11604_, new_n11603_ );
and  ( new_n11606_, new_n11469_, new_n2334_ );
and  ( new_n11607_, new_n11465_, new_n2168_ );
or   ( new_n11608_, new_n11607_, new_n11606_ );
and  ( new_n11609_, new_n11608_, new_n11605_ );
or   ( new_n11610_, new_n11608_, new_n11605_ );
and  ( new_n11611_, new_n11480_, new_n1824_ );
and  ( new_n11612_, new_n11476_, new_n1717_ );
or   ( new_n11613_, new_n11612_, new_n11611_ );
and  ( new_n11614_, new_n11613_, new_n11610_ );
or   ( new_n11615_, new_n11614_, new_n11609_ );
or   ( new_n11616_, new_n11615_, new_n11602_ );
and  ( new_n11617_, new_n11616_, new_n11601_ );
or   ( new_n11618_, new_n11617_, new_n11577_ );
and  ( new_n11619_, new_n11617_, new_n11577_ );
and  ( new_n11620_, new_n11493_, new_n10997_ );
and  ( new_n11621_, new_n11489_, new_n11205_ );
or   ( new_n11622_, new_n11621_, new_n11620_ );
and  ( new_n11623_, new_n11500_, new_n10966_ );
and  ( new_n11624_, new_n11496_, new_n11192_ );
or   ( new_n11625_, new_n11624_, new_n11623_ );
and  ( new_n11626_, new_n11625_, new_n11622_ );
or   ( new_n11627_, new_n11626_, new_n11619_ );
and  ( new_n11628_, new_n11627_, new_n11618_ );
or   ( new_n11629_, new_n11628_, new_n11554_ );
and  ( new_n11630_, new_n11628_, new_n11554_ );
and  ( new_n11631_, new_n11512_, new_n10720_ );
and  ( new_n11632_, new_n11508_, new_n10884_ );
or   ( new_n11633_, new_n11632_, new_n11631_ );
or   ( new_n11634_, new_n11633_, new_n11630_ );
and  ( new_n11635_, new_n11634_, new_n11629_ );
or   ( new_n11636_, new_n11635_, new_n11541_ );
and  ( new_n11637_, new_n11635_, new_n11541_ );
and  ( new_n11638_, new_n11523_, new_n10749_ );
and  ( new_n11639_, new_n11519_, new_n10901_ );
or   ( new_n11640_, new_n11639_, new_n11638_ );
or   ( new_n11641_, new_n11640_, new_n11637_ );
and  ( new_n11642_, new_n11641_, new_n11636_ );
and  ( new_n11643_, new_n11642_, new_n11534_ );
or   ( new_n11644_, new_n11643_, new_n11531_ );
or   ( new_n11645_, new_n11278_, new_n11133_ );
and  ( new_n11646_, new_n11645_, new_n11141_ );
and  ( new_n11647_, new_n11264_, new_n11132_ );
and  ( new_n11648_, new_n11277_, new_n11107_ );
or   ( new_n11649_, new_n11648_, new_n11647_ );
and  ( new_n11650_, new_n11649_, new_n11282_ );
or   ( new_n11651_, new_n11650_, new_n11646_ );
or   ( new_n11652_, new_n11637_, new_n11517_ );
and  ( new_n11653_, new_n11652_, new_n11525_ );
and  ( new_n11654_, new_n11635_, new_n11324_ );
and  ( new_n11655_, new_n11541_, new_n11516_ );
or   ( new_n11656_, new_n11655_, new_n11654_ );
and  ( new_n11657_, new_n11656_, new_n11640_ );
or   ( new_n11658_, new_n11657_, new_n11653_ );
or   ( new_n11659_, new_n11658_, new_n11651_ );
or   ( new_n11660_, new_n11659_, new_n11644_ );
and  ( new_n11661_, new_n11660_, new_n11530_ );
or   ( new_n11662_, new_n11661_, new_n11529_ );
and  ( new_n11663_, new_n11659_, new_n11644_ );
or   ( new_n11664_, new_n11663_, new_n11529_ );
and  ( new_n11665_, new_n11658_, new_n11651_ );
and  ( new_n11666_, new_n11649_, new_n11141_ );
and  ( new_n11667_, new_n11645_, new_n11282_ );
or   ( new_n11668_, new_n11667_, new_n11666_ );
and  ( new_n11669_, new_n11656_, new_n11525_ );
and  ( new_n11670_, new_n11652_, new_n11640_ );
or   ( new_n11671_, new_n11670_, new_n11669_ );
and  ( new_n11672_, new_n11671_, new_n11668_ );
or   ( new_n11673_, new_n11672_, new_n11665_ );
and  ( new_n11674_, new_n11323_, new_n11316_ );
or   ( new_n11675_, new_n11674_, new_n11541_ );
or   ( new_n11676_, new_n7105_, new_n886_ );
or   ( new_n11677_, new_n7099_, new_n843_ );
and  ( new_n11678_, new_n11677_, new_n11676_ );
and  ( new_n11679_, new_n11678_, new_n5858_ );
and  ( new_n11680_, new_n7104_, RI2b1c4342d990_75 );
and  ( new_n11681_, new_n7110_, RI2b1c4342da08_76 );
or   ( new_n11682_, new_n11681_, new_n11680_ );
and  ( new_n11683_, new_n11682_, new_n6037_ );
or   ( new_n11684_, new_n11683_, new_n11679_ );
or   ( new_n11685_, new_n6156_, new_n1002_ );
or   ( new_n11686_, new_n6160_, new_n1004_ );
and  ( new_n11687_, new_n11686_, new_n11685_ );
and  ( new_n11688_, new_n11687_, new_n6039_ );
and  ( new_n11689_, new_n6164_, RI2b1c4342daf8_78 );
and  ( new_n11690_, new_n6154_, RI2b1c4342da80_77 );
or   ( new_n11691_, new_n11690_, new_n11689_ );
and  ( new_n11692_, new_n11691_, new_n5867_ );
or   ( new_n11693_, new_n11692_, new_n11688_ );
and  ( new_n11694_, new_n11693_, new_n11684_ );
or   ( new_n11695_, new_n11693_, new_n11684_ );
or   ( new_n11696_, new_n5308_, new_n1511_ );
or   ( new_n11697_, new_n5312_, new_n1310_ );
and  ( new_n11698_, new_n11697_, new_n11696_ );
and  ( new_n11699_, new_n11698_, new_n5182_ );
and  ( new_n11700_, new_n5316_, RI2b1c4342dbe8_80 );
and  ( new_n11701_, new_n5306_, RI2b1c4342db70_79 );
or   ( new_n11702_, new_n11701_, new_n11700_ );
and  ( new_n11703_, new_n11702_, new_n5028_ );
or   ( new_n11704_, new_n11703_, new_n11699_ );
and  ( new_n11705_, new_n11704_, new_n11695_ );
or   ( new_n11706_, new_n11705_, new_n11694_ );
or   ( new_n11707_, new_n4535_, new_n2119_ );
or   ( new_n11708_, new_n4539_, new_n126_ );
and  ( new_n11709_, new_n11708_, new_n11707_ );
and  ( new_n11710_, new_n11709_, new_n4400_ );
and  ( new_n11711_, new_n4543_, RI2b1c4342dcd8_82 );
and  ( new_n11712_, new_n4533_, RI2b1c4342dc60_81 );
or   ( new_n11713_, new_n11712_, new_n11711_ );
and  ( new_n11714_, new_n11713_, new_n4215_ );
or   ( new_n11715_, new_n11714_, new_n11710_ );
or   ( new_n11716_, new_n3802_, new_n2541_ );
or   ( new_n11717_, new_n3806_, new_n121_ );
and  ( new_n11718_, new_n11717_, new_n11716_ );
and  ( new_n11719_, new_n11718_, new_n3695_ );
and  ( new_n11720_, new_n3810_, RI2b1c4342ddc8_84 );
and  ( new_n11721_, new_n3800_, RI2b1c4342dd50_83 );
or   ( new_n11722_, new_n11721_, new_n11720_ );
and  ( new_n11723_, new_n11722_, new_n3548_ );
or   ( new_n11724_, new_n11723_, new_n11719_ );
and  ( new_n11725_, new_n11724_, new_n11715_ );
or   ( new_n11726_, new_n11724_, new_n11715_ );
or   ( new_n11727_, new_n3112_, new_n3239_ );
or   ( new_n11728_, new_n3116_, new_n2806_ );
and  ( new_n11729_, new_n11728_, new_n11727_ );
and  ( new_n11730_, new_n11729_, new_n3004_ );
and  ( new_n11731_, new_n3120_, RI2b1c4342deb8_86 );
and  ( new_n11732_, new_n3110_, RI2b1c4342de40_85 );
or   ( new_n11733_, new_n11732_, new_n11731_ );
and  ( new_n11734_, new_n11733_, new_n2868_ );
or   ( new_n11735_, new_n11734_, new_n11730_ );
and  ( new_n11736_, new_n11735_, new_n11726_ );
or   ( new_n11737_, new_n11736_, new_n11725_ );
and  ( new_n11738_, new_n11737_, new_n11706_ );
or   ( new_n11739_, new_n11737_, new_n11706_ );
or   ( new_n11740_, new_n2450_, new_n3902_ );
or   ( new_n11741_, new_n2454_, new_n3924_ );
and  ( new_n11742_, new_n11741_, new_n11740_ );
and  ( new_n11743_, new_n11742_, new_n2334_ );
and  ( new_n11744_, new_n2458_, RI2b1c4342dfa8_88 );
and  ( new_n11745_, new_n2448_, RI2b1c4342df30_87 );
or   ( new_n11746_, new_n11745_, new_n11744_ );
and  ( new_n11747_, new_n11746_, new_n2168_ );
or   ( new_n11748_, new_n11747_, new_n11743_ );
or   ( new_n11749_, new_n1910_, new_n4635_ );
or   ( new_n11750_, new_n1914_, new_n132_ );
and  ( new_n11751_, new_n11750_, new_n11749_ );
and  ( new_n11752_, new_n11751_, new_n1824_ );
and  ( new_n11753_, new_n1918_, RI2b1c4342e098_90 );
and  ( new_n11754_, new_n1908_, RI2b1c4342e020_89 );
or   ( new_n11755_, new_n11754_, new_n11753_ );
and  ( new_n11756_, new_n11755_, new_n1717_ );
or   ( new_n11757_, new_n11756_, new_n11752_ );
and  ( new_n11758_, new_n11757_, new_n11748_ );
or   ( new_n11759_, new_n11757_, new_n11748_ );
or   ( new_n11760_, new_n1425_, new_n5459_ );
or   ( new_n11761_, new_n1429_, new_n117_ );
and  ( new_n11762_, new_n11761_, new_n11760_ );
and  ( new_n11763_, new_n11762_, new_n1355_ );
and  ( new_n11764_, new_n1433_, RI2b1c4342e188_92 );
and  ( new_n11765_, new_n1423_, RI2b1c4342e110_91 );
or   ( new_n11766_, new_n11765_, new_n11764_ );
and  ( new_n11767_, new_n11766_, new_n1267_ );
or   ( new_n11768_, new_n11767_, new_n11763_ );
and  ( new_n11769_, new_n11768_, new_n11759_ );
or   ( new_n11770_, new_n11769_, new_n11758_ );
and  ( new_n11771_, new_n11770_, new_n11739_ );
or   ( new_n11772_, new_n11771_, new_n11738_ );
or   ( new_n11773_, new_n528_, new_n7274_ );
and  ( new_n11774_, new_n11773_, new_n505_ );
and  ( new_n11775_, new_n522_, RI2b1c4342e368_96 );
and  ( new_n11776_, new_n11775_, new_n533_ );
or   ( new_n11777_, new_n11776_, new_n11774_ );
or   ( new_n11778_, new_n11564_, new_n11375_ );
and  ( new_n11779_, new_n11778_, new_n11385_ );
and  ( new_n11780_, new_n11560_, new_n11374_ );
and  ( new_n11781_, new_n11563_, new_n11365_ );
or   ( new_n11782_, new_n11781_, new_n11780_ );
and  ( new_n11783_, new_n11782_, new_n11568_ );
or   ( new_n11784_, new_n11783_, new_n11779_ );
and  ( new_n11785_, new_n11784_, new_n11777_ );
or   ( new_n11786_, new_n11784_, new_n11777_ );
or   ( new_n11787_, new_n11609_, new_n11472_ );
and  ( new_n11788_, new_n11787_, new_n11482_ );
and  ( new_n11789_, new_n11605_, new_n11471_ );
and  ( new_n11790_, new_n11608_, new_n11462_ );
or   ( new_n11791_, new_n11790_, new_n11789_ );
and  ( new_n11792_, new_n11791_, new_n11613_ );
or   ( new_n11793_, new_n11792_, new_n11788_ );
and  ( new_n11794_, new_n11793_, new_n11786_ );
or   ( new_n11795_, new_n11794_, new_n11785_ );
and  ( new_n11796_, new_n11795_, new_n11772_ );
or   ( new_n11797_, new_n11795_, new_n11772_ );
or   ( new_n11798_, new_n11584_, new_n11417_ );
and  ( new_n11799_, new_n11798_, new_n11427_ );
and  ( new_n11800_, new_n11580_, new_n11416_ );
and  ( new_n11801_, new_n11583_, new_n11407_ );
or   ( new_n11802_, new_n11801_, new_n11800_ );
and  ( new_n11803_, new_n11802_, new_n11588_ );
or   ( new_n11804_, new_n11803_, new_n11799_ );
or   ( new_n11805_, new_n11595_, new_n11439_ );
and  ( new_n11806_, new_n11805_, new_n11449_ );
and  ( new_n11807_, new_n11438_, new_n533_ );
and  ( new_n11808_, new_n11593_, new_n505_ );
or   ( new_n11809_, new_n11808_, new_n11807_ );
and  ( new_n11810_, new_n11809_, new_n11598_ );
or   ( new_n11811_, new_n11810_, new_n11806_ );
or   ( new_n11812_, new_n11811_, new_n11804_ );
and  ( new_n11813_, new_n11812_, new_n11797_ );
or   ( new_n11814_, new_n11813_, new_n11796_ );
and  ( new_n11815_, new_n11502_, new_n11495_ );
or   ( new_n11816_, new_n11815_, new_n11626_ );
or   ( new_n11817_, new_n11571_, new_n11388_ );
and  ( new_n11818_, new_n11817_, new_n11396_ );
and  ( new_n11819_, new_n11570_, new_n11356_ );
and  ( new_n11820_, new_n11557_, new_n11387_ );
or   ( new_n11821_, new_n11820_, new_n11819_ );
and  ( new_n11822_, new_n11821_, new_n11575_ );
or   ( new_n11823_, new_n11822_, new_n11818_ );
and  ( new_n11824_, new_n11823_, new_n11816_ );
or   ( new_n11825_, new_n11823_, new_n11816_ );
or   ( new_n11826_, new_n11602_, new_n11452_ );
and  ( new_n11827_, new_n11826_, new_n11484_ );
and  ( new_n11828_, new_n11600_, new_n11429_ );
and  ( new_n11829_, new_n11590_, new_n11451_ );
or   ( new_n11830_, new_n11829_, new_n11828_ );
and  ( new_n11831_, new_n11830_, new_n11615_ );
or   ( new_n11832_, new_n11831_, new_n11827_ );
and  ( new_n11833_, new_n11832_, new_n11825_ );
or   ( new_n11834_, new_n11833_, new_n11824_ );
and  ( new_n11835_, new_n11834_, new_n11814_ );
or   ( new_n11836_, new_n11834_, new_n11814_ );
or   ( new_n11837_, new_n11548_, new_n11339_ );
and  ( new_n11838_, new_n11837_, new_n11347_ );
and  ( new_n11839_, new_n11544_, new_n11338_ );
and  ( new_n11840_, new_n11547_, new_n11331_ );
or   ( new_n11841_, new_n11840_, new_n11839_ );
and  ( new_n11842_, new_n11841_, new_n11552_ );
or   ( new_n11843_, new_n11842_, new_n11838_ );
and  ( new_n11844_, new_n11843_, new_n11836_ );
or   ( new_n11845_, new_n11844_, new_n11835_ );
and  ( new_n11846_, new_n11845_, new_n11675_ );
or   ( new_n11847_, new_n11845_, new_n11675_ );
or   ( new_n11848_, new_n11630_, new_n11506_ );
and  ( new_n11849_, new_n11848_, new_n11514_ );
and  ( new_n11850_, new_n11628_, new_n11349_ );
and  ( new_n11851_, new_n11554_, new_n11505_ );
or   ( new_n11852_, new_n11851_, new_n11850_ );
and  ( new_n11853_, new_n11852_, new_n11633_ );
or   ( new_n11854_, new_n11853_, new_n11849_ );
and  ( new_n11855_, new_n11854_, new_n11847_ );
or   ( new_n11856_, new_n11855_, new_n11846_ );
and  ( new_n11857_, new_n11856_, new_n11673_ );
or   ( new_n11858_, new_n11856_, new_n11673_ );
and  ( new_n11859_, new_n11537_, new_n11323_ );
and  ( new_n11860_, new_n11540_, new_n11316_ );
or   ( new_n11861_, new_n11860_, new_n11859_ );
and  ( new_n11862_, new_n11682_, new_n5858_ );
and  ( new_n11863_, new_n11678_, new_n6037_ );
or   ( new_n11864_, new_n11863_, new_n11862_ );
and  ( new_n11865_, new_n11691_, new_n6039_ );
and  ( new_n11866_, new_n11687_, new_n5867_ );
or   ( new_n11867_, new_n11866_, new_n11865_ );
and  ( new_n11868_, new_n11867_, new_n11864_ );
or   ( new_n11869_, new_n11867_, new_n11864_ );
and  ( new_n11870_, new_n11702_, new_n5182_ );
and  ( new_n11871_, new_n11698_, new_n5028_ );
or   ( new_n11872_, new_n11871_, new_n11870_ );
and  ( new_n11873_, new_n11872_, new_n11869_ );
or   ( new_n11874_, new_n11873_, new_n11868_ );
and  ( new_n11875_, new_n11713_, new_n4400_ );
and  ( new_n11876_, new_n11709_, new_n4215_ );
or   ( new_n11877_, new_n11876_, new_n11875_ );
and  ( new_n11878_, new_n11722_, new_n3695_ );
and  ( new_n11879_, new_n11718_, new_n3548_ );
or   ( new_n11880_, new_n11879_, new_n11878_ );
and  ( new_n11881_, new_n11880_, new_n11877_ );
or   ( new_n11882_, new_n11880_, new_n11877_ );
and  ( new_n11883_, new_n11733_, new_n3004_ );
and  ( new_n11884_, new_n11729_, new_n2868_ );
or   ( new_n11885_, new_n11884_, new_n11883_ );
and  ( new_n11886_, new_n11885_, new_n11882_ );
or   ( new_n11887_, new_n11886_, new_n11881_ );
and  ( new_n11888_, new_n11887_, new_n11874_ );
or   ( new_n11889_, new_n11887_, new_n11874_ );
and  ( new_n11890_, new_n11746_, new_n2334_ );
and  ( new_n11891_, new_n11742_, new_n2168_ );
or   ( new_n11892_, new_n11891_, new_n11890_ );
and  ( new_n11893_, new_n11755_, new_n1824_ );
and  ( new_n11894_, new_n11751_, new_n1717_ );
or   ( new_n11895_, new_n11894_, new_n11893_ );
and  ( new_n11896_, new_n11895_, new_n11892_ );
or   ( new_n11897_, new_n11895_, new_n11892_ );
and  ( new_n11898_, new_n11766_, new_n1355_ );
and  ( new_n11899_, new_n11762_, new_n1267_ );
or   ( new_n11900_, new_n11899_, new_n11898_ );
and  ( new_n11901_, new_n11900_, new_n11897_ );
or   ( new_n11902_, new_n11901_, new_n11896_ );
and  ( new_n11903_, new_n11902_, new_n11889_ );
or   ( new_n11904_, new_n11903_, new_n11888_ );
and  ( new_n11905_, new_n11775_, new_n505_ );
and  ( new_n11906_, new_n11773_, new_n533_ );
or   ( new_n11907_, new_n11906_, new_n11905_ );
and  ( new_n11908_, new_n11782_, new_n11385_ );
and  ( new_n11909_, new_n11778_, new_n11568_ );
or   ( new_n11910_, new_n11909_, new_n11908_ );
and  ( new_n11911_, new_n11910_, new_n11907_ );
or   ( new_n11912_, new_n11910_, new_n11907_ );
and  ( new_n11913_, new_n11791_, new_n11482_ );
and  ( new_n11914_, new_n11787_, new_n11613_ );
or   ( new_n11915_, new_n11914_, new_n11913_ );
and  ( new_n11916_, new_n11915_, new_n11912_ );
or   ( new_n11917_, new_n11916_, new_n11911_ );
and  ( new_n11918_, new_n11917_, new_n11904_ );
or   ( new_n11919_, new_n11917_, new_n11904_ );
and  ( new_n11920_, new_n11802_, new_n11427_ );
and  ( new_n11921_, new_n11798_, new_n11588_ );
or   ( new_n11922_, new_n11921_, new_n11920_ );
and  ( new_n11923_, new_n11809_, new_n11449_ );
and  ( new_n11924_, new_n11805_, new_n11598_ );
or   ( new_n11925_, new_n11924_, new_n11923_ );
and  ( new_n11926_, new_n11925_, new_n11922_ );
and  ( new_n11927_, new_n11926_, new_n11919_ );
or   ( new_n11928_, new_n11927_, new_n11918_ );
and  ( new_n11929_, new_n11622_, new_n11502_ );
and  ( new_n11930_, new_n11625_, new_n11495_ );
or   ( new_n11931_, new_n11930_, new_n11929_ );
and  ( new_n11932_, new_n11821_, new_n11396_ );
and  ( new_n11933_, new_n11817_, new_n11575_ );
or   ( new_n11934_, new_n11933_, new_n11932_ );
and  ( new_n11935_, new_n11934_, new_n11931_ );
or   ( new_n11936_, new_n11934_, new_n11931_ );
and  ( new_n11937_, new_n11830_, new_n11484_ );
and  ( new_n11938_, new_n11826_, new_n11615_ );
or   ( new_n11939_, new_n11938_, new_n11937_ );
and  ( new_n11940_, new_n11939_, new_n11936_ );
or   ( new_n11941_, new_n11940_, new_n11935_ );
and  ( new_n11942_, new_n11941_, new_n11928_ );
or   ( new_n11943_, new_n11941_, new_n11928_ );
and  ( new_n11944_, new_n11841_, new_n11347_ );
and  ( new_n11945_, new_n11837_, new_n11552_ );
or   ( new_n11946_, new_n11945_, new_n11944_ );
and  ( new_n11947_, new_n11946_, new_n11943_ );
or   ( new_n11948_, new_n11947_, new_n11942_ );
and  ( new_n11949_, new_n11948_, new_n11861_ );
or   ( new_n11950_, new_n11949_, new_n11846_ );
and  ( new_n11951_, new_n11950_, new_n11854_ );
and  ( new_n11952_, new_n11948_, new_n11675_ );
and  ( new_n11953_, new_n11861_, new_n11845_ );
or   ( new_n11954_, new_n11953_, new_n11952_ );
and  ( new_n11955_, new_n11852_, new_n11514_ );
and  ( new_n11956_, new_n11848_, new_n11633_ );
or   ( new_n11957_, new_n11956_, new_n11955_ );
and  ( new_n11958_, new_n11957_, new_n11954_ );
or   ( new_n11959_, new_n11958_, new_n11951_ );
or   ( new_n11960_, new_n11619_, new_n11487_ );
and  ( new_n11961_, new_n11960_, new_n11503_ );
and  ( new_n11962_, new_n11617_, new_n11398_ );
and  ( new_n11963_, new_n11577_, new_n11486_ );
or   ( new_n11964_, new_n11963_, new_n11962_ );
and  ( new_n11965_, new_n11964_, new_n11626_ );
or   ( new_n11966_, new_n11965_, new_n11961_ );
and  ( new_n11967_, new_n11811_, new_n11804_ );
or   ( new_n11968_, new_n11967_, new_n11926_ );
or   ( new_n11969_, new_n11911_, new_n11785_ );
and  ( new_n11970_, new_n11969_, new_n11793_ );
and  ( new_n11971_, new_n11907_, new_n11784_ );
and  ( new_n11972_, new_n11910_, new_n11777_ );
or   ( new_n11973_, new_n11972_, new_n11971_ );
and  ( new_n11974_, new_n11973_, new_n11915_ );
or   ( new_n11975_, new_n11974_, new_n11970_ );
and  ( new_n11976_, new_n11975_, new_n11968_ );
or   ( new_n11977_, new_n11975_, new_n11968_ );
or   ( new_n11978_, new_n11888_, new_n11738_ );
and  ( new_n11979_, new_n11978_, new_n11770_ );
and  ( new_n11980_, new_n11874_, new_n11737_ );
and  ( new_n11981_, new_n11887_, new_n11706_ );
or   ( new_n11982_, new_n11981_, new_n11980_ );
and  ( new_n11983_, new_n11982_, new_n11902_ );
or   ( new_n11984_, new_n11983_, new_n11979_ );
and  ( new_n11985_, new_n11984_, new_n11977_ );
or   ( new_n11986_, new_n11985_, new_n11976_ );
or   ( new_n11987_, new_n934_, new_n6321_ );
or   ( new_n11988_, new_n940_, new_n6307_ );
and  ( new_n11989_, new_n11988_, new_n11987_ );
and  ( new_n11990_, new_n11989_, new_n913_ );
and  ( new_n11991_, new_n944_, RI2b1c4342e278_94 );
and  ( new_n11992_, new_n932_, RI2b1c4342e200_93 );
or   ( new_n11993_, new_n11992_, new_n11991_ );
and  ( new_n11994_, new_n11993_, new_n938_ );
or   ( new_n11995_, new_n11994_, new_n11990_ );
or   ( new_n11996_, new_n1425_, new_n6307_ );
or   ( new_n11997_, new_n1429_, new_n5459_ );
and  ( new_n11998_, new_n11997_, new_n11996_ );
and  ( new_n11999_, new_n11998_, new_n1355_ );
and  ( new_n12000_, new_n1433_, RI2b1c4342e200_93 );
and  ( new_n12001_, new_n1423_, RI2b1c4342e188_92 );
or   ( new_n12002_, new_n12001_, new_n12000_ );
and  ( new_n12003_, new_n12002_, new_n1267_ );
or   ( new_n12004_, new_n12003_, new_n11999_ );
or   ( new_n12005_, new_n934_, new_n124_ );
or   ( new_n12006_, new_n940_, new_n6321_ );
and  ( new_n12007_, new_n12006_, new_n12005_ );
and  ( new_n12008_, new_n12007_, new_n913_ );
and  ( new_n12009_, new_n944_, RI2b1c4342e2f0_95 );
and  ( new_n12010_, new_n932_, RI2b1c4342e278_94 );
or   ( new_n12011_, new_n12010_, new_n12009_ );
and  ( new_n12012_, new_n12011_, new_n938_ );
or   ( new_n12013_, new_n12012_, new_n12008_ );
and  ( new_n12014_, new_n12013_, new_n12004_ );
or   ( new_n12015_, new_n12013_, new_n12004_ );
or   ( new_n12016_, new_n459_, new_n7274_ );
and  ( new_n12017_, new_n12016_, new_n428_ );
and  ( new_n12018_, new_n451_, RI2b1c4342e368_96 );
and  ( new_n12019_, new_n12018_, new_n457_ );
or   ( new_n12020_, new_n12019_, new_n12017_ );
and  ( new_n12021_, new_n12020_, new_n12015_ );
or   ( new_n12022_, new_n12021_, new_n12014_ );
and  ( new_n12023_, new_n12022_, new_n11995_ );
or   ( new_n12024_, new_n12022_, new_n11995_ );
or   ( new_n12025_, new_n453_, new_n7274_ );
or   ( new_n12026_, new_n459_, new_n124_ );
and  ( new_n12027_, new_n12026_, new_n12025_ );
and  ( new_n12028_, new_n12027_, new_n428_ );
and  ( new_n12029_, new_n463_, RI2b1c4342e368_96 );
and  ( new_n12030_, new_n451_, RI2b1c4342e2f0_95 );
or   ( new_n12031_, new_n12030_, new_n12029_ );
and  ( new_n12032_, new_n12031_, new_n457_ );
or   ( new_n12033_, new_n12032_, new_n12028_ );
and  ( new_n12034_, new_n12033_, new_n12024_ );
or   ( new_n12035_, new_n12034_, new_n12023_ );
or   ( new_n12036_, new_n5308_, new_n126_ );
or   ( new_n12037_, new_n5312_, new_n1511_ );
and  ( new_n12038_, new_n12037_, new_n12036_ );
and  ( new_n12039_, new_n12038_, new_n5182_ );
and  ( new_n12040_, new_n5316_, RI2b1c4342dc60_81 );
and  ( new_n12041_, new_n5306_, RI2b1c4342dbe8_80 );
or   ( new_n12042_, new_n12041_, new_n12040_ );
and  ( new_n12043_, new_n12042_, new_n5028_ );
or   ( new_n12044_, new_n12043_, new_n12039_ );
or   ( new_n12045_, new_n4535_, new_n121_ );
or   ( new_n12046_, new_n4539_, new_n2119_ );
and  ( new_n12047_, new_n12046_, new_n12045_ );
and  ( new_n12048_, new_n12047_, new_n4400_ );
and  ( new_n12049_, new_n4543_, RI2b1c4342dd50_83 );
and  ( new_n12050_, new_n4533_, RI2b1c4342dcd8_82 );
or   ( new_n12051_, new_n12050_, new_n12049_ );
and  ( new_n12052_, new_n12051_, new_n4215_ );
or   ( new_n12053_, new_n12052_, new_n12048_ );
and  ( new_n12054_, new_n12053_, new_n12044_ );
or   ( new_n12055_, new_n12053_, new_n12044_ );
or   ( new_n12056_, new_n3802_, new_n2806_ );
or   ( new_n12057_, new_n3806_, new_n2541_ );
and  ( new_n12058_, new_n12057_, new_n12056_ );
and  ( new_n12059_, new_n12058_, new_n3695_ );
and  ( new_n12060_, new_n3810_, RI2b1c4342de40_85 );
and  ( new_n12061_, new_n3800_, RI2b1c4342ddc8_84 );
or   ( new_n12062_, new_n12061_, new_n12060_ );
and  ( new_n12063_, new_n12062_, new_n3548_ );
or   ( new_n12064_, new_n12063_, new_n12059_ );
and  ( new_n12065_, new_n12064_, new_n12055_ );
or   ( new_n12066_, new_n12065_, new_n12054_ );
or   ( new_n12067_, new_n7105_, new_n1004_ );
or   ( new_n12068_, new_n7099_, new_n886_ );
and  ( new_n12069_, new_n12068_, new_n12067_ );
and  ( new_n12070_, new_n12069_, new_n5858_ );
and  ( new_n12071_, new_n7104_, RI2b1c4342da08_76 );
and  ( new_n12072_, new_n7110_, RI2b1c4342da80_77 );
or   ( new_n12073_, new_n12072_, new_n12071_ );
and  ( new_n12074_, new_n12073_, new_n6037_ );
or   ( new_n12075_, new_n12074_, new_n12070_ );
and  ( new_n12076_, new_n12075_, new_n428_ );
or   ( new_n12077_, new_n12075_, new_n428_ );
or   ( new_n12078_, new_n6156_, new_n1310_ );
or   ( new_n12079_, new_n6160_, new_n1002_ );
and  ( new_n12080_, new_n12079_, new_n12078_ );
and  ( new_n12081_, new_n12080_, new_n6039_ );
and  ( new_n12082_, new_n6164_, RI2b1c4342db70_79 );
and  ( new_n12083_, new_n6154_, RI2b1c4342daf8_78 );
or   ( new_n12084_, new_n12083_, new_n12082_ );
and  ( new_n12085_, new_n12084_, new_n5867_ );
or   ( new_n12086_, new_n12085_, new_n12081_ );
and  ( new_n12087_, new_n12086_, new_n12077_ );
or   ( new_n12088_, new_n12087_, new_n12076_ );
and  ( new_n12089_, new_n12088_, new_n12066_ );
or   ( new_n12090_, new_n12088_, new_n12066_ );
or   ( new_n12091_, new_n3112_, new_n3924_ );
or   ( new_n12092_, new_n3116_, new_n3239_ );
and  ( new_n12093_, new_n12092_, new_n12091_ );
and  ( new_n12094_, new_n12093_, new_n3004_ );
and  ( new_n12095_, new_n3120_, RI2b1c4342df30_87 );
and  ( new_n12096_, new_n3110_, RI2b1c4342deb8_86 );
or   ( new_n12097_, new_n12096_, new_n12095_ );
and  ( new_n12098_, new_n12097_, new_n2868_ );
or   ( new_n12099_, new_n12098_, new_n12094_ );
or   ( new_n12100_, new_n2450_, new_n132_ );
or   ( new_n12101_, new_n2454_, new_n3902_ );
and  ( new_n12102_, new_n12101_, new_n12100_ );
and  ( new_n12103_, new_n12102_, new_n2334_ );
and  ( new_n12104_, new_n2458_, RI2b1c4342e020_89 );
and  ( new_n12105_, new_n2448_, RI2b1c4342dfa8_88 );
or   ( new_n12106_, new_n12105_, new_n12104_ );
and  ( new_n12107_, new_n12106_, new_n2168_ );
or   ( new_n12108_, new_n12107_, new_n12103_ );
and  ( new_n12109_, new_n12108_, new_n12099_ );
or   ( new_n12110_, new_n12108_, new_n12099_ );
or   ( new_n12111_, new_n1910_, new_n117_ );
or   ( new_n12112_, new_n1914_, new_n4635_ );
and  ( new_n12113_, new_n12112_, new_n12111_ );
and  ( new_n12114_, new_n12113_, new_n1824_ );
and  ( new_n12115_, new_n1918_, RI2b1c4342e110_91 );
and  ( new_n12116_, new_n1908_, RI2b1c4342e098_90 );
or   ( new_n12117_, new_n12116_, new_n12115_ );
and  ( new_n12118_, new_n12117_, new_n1717_ );
or   ( new_n12119_, new_n12118_, new_n12114_ );
and  ( new_n12120_, new_n12119_, new_n12110_ );
or   ( new_n12121_, new_n12120_, new_n12109_ );
and  ( new_n12122_, new_n12121_, new_n12090_ );
or   ( new_n12123_, new_n12122_, new_n12089_ );
and  ( new_n12124_, new_n12123_, new_n12035_ );
or   ( new_n12125_, new_n12123_, new_n12035_ );
or   ( new_n12126_, new_n11896_, new_n11758_ );
and  ( new_n12127_, new_n12126_, new_n11768_ );
and  ( new_n12128_, new_n11892_, new_n11757_ );
and  ( new_n12129_, new_n11895_, new_n11748_ );
or   ( new_n12130_, new_n12129_, new_n12128_ );
and  ( new_n12131_, new_n12130_, new_n11900_ );
or   ( new_n12132_, new_n12131_, new_n12127_ );
or   ( new_n12133_, new_n11881_, new_n11725_ );
and  ( new_n12134_, new_n12133_, new_n11735_ );
and  ( new_n12135_, new_n11877_, new_n11724_ );
and  ( new_n12136_, new_n11880_, new_n11715_ );
or   ( new_n12137_, new_n12136_, new_n12135_ );
and  ( new_n12138_, new_n12137_, new_n11885_ );
or   ( new_n12139_, new_n12138_, new_n12134_ );
and  ( new_n12140_, new_n12139_, new_n12132_ );
or   ( new_n12141_, new_n12139_, new_n12132_ );
or   ( new_n12142_, new_n11868_, new_n11694_ );
and  ( new_n12143_, new_n12142_, new_n11704_ );
and  ( new_n12144_, new_n11864_, new_n11693_ );
and  ( new_n12145_, new_n11867_, new_n11684_ );
or   ( new_n12146_, new_n12145_, new_n12144_ );
and  ( new_n12147_, new_n12146_, new_n11872_ );
or   ( new_n12148_, new_n12147_, new_n12143_ );
and  ( new_n12149_, new_n12148_, new_n12141_ );
or   ( new_n12150_, new_n12149_, new_n12140_ );
and  ( new_n12151_, new_n12150_, new_n12125_ );
or   ( new_n12152_, new_n12151_, new_n12124_ );
and  ( new_n12153_, new_n12152_, new_n11986_ );
or   ( new_n12154_, new_n12152_, new_n11986_ );
or   ( new_n12155_, new_n11935_, new_n11824_ );
and  ( new_n12156_, new_n12155_, new_n11832_ );
and  ( new_n12157_, new_n11931_, new_n11823_ );
and  ( new_n12158_, new_n11934_, new_n11816_ );
or   ( new_n12159_, new_n12158_, new_n12157_ );
and  ( new_n12160_, new_n12159_, new_n11939_ );
or   ( new_n12161_, new_n12160_, new_n12156_ );
and  ( new_n12162_, new_n12161_, new_n12154_ );
or   ( new_n12163_, new_n12162_, new_n12153_ );
and  ( new_n12164_, new_n12163_, new_n11966_ );
or   ( new_n12165_, new_n12163_, new_n11966_ );
or   ( new_n12166_, new_n11942_, new_n11835_ );
and  ( new_n12167_, new_n12166_, new_n11843_ );
and  ( new_n12168_, new_n11928_, new_n11834_ );
and  ( new_n12169_, new_n11941_, new_n11814_ );
or   ( new_n12170_, new_n12169_, new_n12168_ );
and  ( new_n12171_, new_n12170_, new_n11946_ );
or   ( new_n12172_, new_n12171_, new_n12167_ );
and  ( new_n12173_, new_n12172_, new_n12165_ );
or   ( new_n12174_, new_n12173_, new_n12164_ );
or   ( new_n12175_, new_n12174_, new_n11959_ );
and  ( new_n12176_, new_n12175_, new_n11858_ );
or   ( new_n12177_, new_n12176_, new_n11857_ );
or   ( new_n12178_, new_n12177_, new_n11664_ );
and  ( new_n12179_, new_n12178_, new_n11662_ );
and  ( new_n12180_, new_n12174_, new_n11959_ );
or   ( new_n12181_, new_n12180_, new_n11857_ );
or   ( new_n12182_, new_n12181_, new_n11664_ );
and  ( new_n12183_, new_n11964_, new_n11503_ );
and  ( new_n12184_, new_n11960_, new_n11626_ );
or   ( new_n12185_, new_n12184_, new_n12183_ );
and  ( new_n12186_, new_n11922_, new_n11811_ );
and  ( new_n12187_, new_n11925_, new_n11804_ );
or   ( new_n12188_, new_n12187_, new_n12186_ );
and  ( new_n12189_, new_n11973_, new_n11793_ );
and  ( new_n12190_, new_n11969_, new_n11915_ );
or   ( new_n12191_, new_n12190_, new_n12189_ );
and  ( new_n12192_, new_n12191_, new_n12188_ );
or   ( new_n12193_, new_n12191_, new_n12188_ );
and  ( new_n12194_, new_n11982_, new_n11770_ );
and  ( new_n12195_, new_n11978_, new_n11902_ );
or   ( new_n12196_, new_n12195_, new_n12194_ );
and  ( new_n12197_, new_n12196_, new_n12193_ );
or   ( new_n12198_, new_n12197_, new_n12192_ );
and  ( new_n12199_, new_n11993_, new_n913_ );
and  ( new_n12200_, new_n11989_, new_n938_ );
or   ( new_n12201_, new_n12200_, new_n12199_ );
and  ( new_n12202_, new_n12002_, new_n1355_ );
and  ( new_n12203_, new_n11998_, new_n1267_ );
or   ( new_n12204_, new_n12203_, new_n12202_ );
and  ( new_n12205_, new_n12011_, new_n913_ );
and  ( new_n12206_, new_n12007_, new_n938_ );
or   ( new_n12207_, new_n12206_, new_n12205_ );
and  ( new_n12208_, new_n12207_, new_n12204_ );
or   ( new_n12209_, new_n12207_, new_n12204_ );
and  ( new_n12210_, new_n12018_, new_n428_ );
and  ( new_n12211_, new_n12016_, new_n457_ );
or   ( new_n12212_, new_n12211_, new_n12210_ );
and  ( new_n12213_, new_n12212_, new_n12209_ );
or   ( new_n12214_, new_n12213_, new_n12208_ );
and  ( new_n12215_, new_n12214_, new_n12201_ );
or   ( new_n12216_, new_n12214_, new_n12201_ );
and  ( new_n12217_, new_n12031_, new_n428_ );
and  ( new_n12218_, new_n12027_, new_n457_ );
or   ( new_n12219_, new_n12218_, new_n12217_ );
and  ( new_n12220_, new_n12219_, new_n12216_ );
or   ( new_n12221_, new_n12220_, new_n12215_ );
and  ( new_n12222_, new_n12042_, new_n5182_ );
and  ( new_n12223_, new_n12038_, new_n5028_ );
or   ( new_n12224_, new_n12223_, new_n12222_ );
and  ( new_n12225_, new_n12051_, new_n4400_ );
and  ( new_n12226_, new_n12047_, new_n4215_ );
or   ( new_n12227_, new_n12226_, new_n12225_ );
and  ( new_n12228_, new_n12227_, new_n12224_ );
or   ( new_n12229_, new_n12227_, new_n12224_ );
and  ( new_n12230_, new_n12062_, new_n3695_ );
and  ( new_n12231_, new_n12058_, new_n3548_ );
or   ( new_n12232_, new_n12231_, new_n12230_ );
and  ( new_n12233_, new_n12232_, new_n12229_ );
or   ( new_n12234_, new_n12233_, new_n12228_ );
and  ( new_n12235_, new_n12073_, new_n5858_ );
and  ( new_n12236_, new_n12069_, new_n6037_ );
or   ( new_n12237_, new_n12236_, new_n12235_ );
or   ( new_n12238_, new_n12237_, new_n457_ );
and  ( new_n12239_, new_n12237_, new_n457_ );
and  ( new_n12240_, new_n12084_, new_n6039_ );
and  ( new_n12241_, new_n12080_, new_n5867_ );
or   ( new_n12242_, new_n12241_, new_n12240_ );
or   ( new_n12243_, new_n12242_, new_n12239_ );
and  ( new_n12244_, new_n12243_, new_n12238_ );
or   ( new_n12245_, new_n12244_, new_n12234_ );
and  ( new_n12246_, new_n12244_, new_n12234_ );
and  ( new_n12247_, new_n12097_, new_n3004_ );
and  ( new_n12248_, new_n12093_, new_n2868_ );
or   ( new_n12249_, new_n12248_, new_n12247_ );
and  ( new_n12250_, new_n12106_, new_n2334_ );
and  ( new_n12251_, new_n12102_, new_n2168_ );
or   ( new_n12252_, new_n12251_, new_n12250_ );
and  ( new_n12253_, new_n12252_, new_n12249_ );
or   ( new_n12254_, new_n12252_, new_n12249_ );
and  ( new_n12255_, new_n12117_, new_n1824_ );
and  ( new_n12256_, new_n12113_, new_n1717_ );
or   ( new_n12257_, new_n12256_, new_n12255_ );
and  ( new_n12258_, new_n12257_, new_n12254_ );
or   ( new_n12259_, new_n12258_, new_n12253_ );
or   ( new_n12260_, new_n12259_, new_n12246_ );
and  ( new_n12261_, new_n12260_, new_n12245_ );
or   ( new_n12262_, new_n12261_, new_n12221_ );
and  ( new_n12263_, new_n12261_, new_n12221_ );
and  ( new_n12264_, new_n12130_, new_n11768_ );
and  ( new_n12265_, new_n12126_, new_n11900_ );
or   ( new_n12266_, new_n12265_, new_n12264_ );
and  ( new_n12267_, new_n12137_, new_n11735_ );
and  ( new_n12268_, new_n12133_, new_n11885_ );
or   ( new_n12269_, new_n12268_, new_n12267_ );
and  ( new_n12270_, new_n12269_, new_n12266_ );
or   ( new_n12271_, new_n12269_, new_n12266_ );
and  ( new_n12272_, new_n12146_, new_n11704_ );
and  ( new_n12273_, new_n12142_, new_n11872_ );
or   ( new_n12274_, new_n12273_, new_n12272_ );
and  ( new_n12275_, new_n12274_, new_n12271_ );
or   ( new_n12276_, new_n12275_, new_n12270_ );
or   ( new_n12277_, new_n12276_, new_n12263_ );
and  ( new_n12278_, new_n12277_, new_n12262_ );
or   ( new_n12279_, new_n12278_, new_n12198_ );
and  ( new_n12280_, new_n12278_, new_n12198_ );
and  ( new_n12281_, new_n12159_, new_n11832_ );
and  ( new_n12282_, new_n12155_, new_n11939_ );
or   ( new_n12283_, new_n12282_, new_n12281_ );
or   ( new_n12284_, new_n12283_, new_n12280_ );
and  ( new_n12285_, new_n12284_, new_n12279_ );
and  ( new_n12286_, new_n12285_, new_n12185_ );
or   ( new_n12287_, new_n12286_, new_n12164_ );
and  ( new_n12288_, new_n12287_, new_n12172_ );
and  ( new_n12289_, new_n12285_, new_n11966_ );
and  ( new_n12290_, new_n12185_, new_n12163_ );
or   ( new_n12291_, new_n12290_, new_n12289_ );
and  ( new_n12292_, new_n12170_, new_n11843_ );
and  ( new_n12293_, new_n12166_, new_n11946_ );
or   ( new_n12294_, new_n12293_, new_n12292_ );
and  ( new_n12295_, new_n12294_, new_n12291_ );
or   ( new_n12296_, new_n12295_, new_n12288_ );
or   ( new_n12297_, new_n11918_, new_n11796_ );
and  ( new_n12298_, new_n12297_, new_n11812_ );
and  ( new_n12299_, new_n11904_, new_n11795_ );
and  ( new_n12300_, new_n11917_, new_n11772_ );
or   ( new_n12301_, new_n12300_, new_n12299_ );
and  ( new_n12302_, new_n12301_, new_n11926_ );
or   ( new_n12303_, new_n12302_, new_n12298_ );
or   ( new_n12304_, new_n12192_, new_n11976_ );
and  ( new_n12305_, new_n12304_, new_n11984_ );
and  ( new_n12306_, new_n12188_, new_n11975_ );
and  ( new_n12307_, new_n12191_, new_n11968_ );
or   ( new_n12308_, new_n12307_, new_n12306_ );
and  ( new_n12309_, new_n12308_, new_n12196_ );
or   ( new_n12310_, new_n12309_, new_n12305_ );
or   ( new_n12311_, new_n7105_, new_n1002_ );
or   ( new_n12312_, new_n7099_, new_n1004_ );
and  ( new_n12313_, new_n12312_, new_n12311_ );
and  ( new_n12314_, new_n12313_, new_n5858_ );
and  ( new_n12315_, new_n7104_, RI2b1c4342da80_77 );
and  ( new_n12316_, new_n7110_, RI2b1c4342daf8_78 );
or   ( new_n12317_, new_n12316_, new_n12315_ );
and  ( new_n12318_, new_n12317_, new_n6037_ );
or   ( new_n12319_, new_n12318_, new_n12314_ );
or   ( new_n12320_, new_n6156_, new_n1511_ );
or   ( new_n12321_, new_n6160_, new_n1310_ );
and  ( new_n12322_, new_n12321_, new_n12320_ );
and  ( new_n12323_, new_n12322_, new_n6039_ );
and  ( new_n12324_, new_n6164_, RI2b1c4342dbe8_80 );
and  ( new_n12325_, new_n6154_, RI2b1c4342db70_79 );
or   ( new_n12326_, new_n12325_, new_n12324_ );
and  ( new_n12327_, new_n12326_, new_n5867_ );
or   ( new_n12328_, new_n12327_, new_n12323_ );
and  ( new_n12329_, new_n12328_, new_n12319_ );
or   ( new_n12330_, new_n12328_, new_n12319_ );
or   ( new_n12331_, new_n5308_, new_n2119_ );
or   ( new_n12332_, new_n5312_, new_n126_ );
and  ( new_n12333_, new_n12332_, new_n12331_ );
and  ( new_n12334_, new_n12333_, new_n5182_ );
and  ( new_n12335_, new_n5316_, RI2b1c4342dcd8_82 );
and  ( new_n12336_, new_n5306_, RI2b1c4342dc60_81 );
or   ( new_n12337_, new_n12336_, new_n12335_ );
and  ( new_n12338_, new_n12337_, new_n5028_ );
or   ( new_n12339_, new_n12338_, new_n12334_ );
and  ( new_n12340_, new_n12339_, new_n12330_ );
or   ( new_n12341_, new_n12340_, new_n12329_ );
or   ( new_n12342_, new_n4535_, new_n2541_ );
or   ( new_n12343_, new_n4539_, new_n121_ );
and  ( new_n12344_, new_n12343_, new_n12342_ );
and  ( new_n12345_, new_n12344_, new_n4400_ );
and  ( new_n12346_, new_n4543_, RI2b1c4342ddc8_84 );
and  ( new_n12347_, new_n4533_, RI2b1c4342dd50_83 );
or   ( new_n12348_, new_n12347_, new_n12346_ );
and  ( new_n12349_, new_n12348_, new_n4215_ );
or   ( new_n12350_, new_n12349_, new_n12345_ );
or   ( new_n12351_, new_n3802_, new_n3239_ );
or   ( new_n12352_, new_n3806_, new_n2806_ );
and  ( new_n12353_, new_n12352_, new_n12351_ );
and  ( new_n12354_, new_n12353_, new_n3695_ );
and  ( new_n12355_, new_n3810_, RI2b1c4342deb8_86 );
and  ( new_n12356_, new_n3800_, RI2b1c4342de40_85 );
or   ( new_n12357_, new_n12356_, new_n12355_ );
and  ( new_n12358_, new_n12357_, new_n3548_ );
or   ( new_n12359_, new_n12358_, new_n12354_ );
and  ( new_n12360_, new_n12359_, new_n12350_ );
or   ( new_n12361_, new_n12359_, new_n12350_ );
or   ( new_n12362_, new_n3112_, new_n3902_ );
or   ( new_n12363_, new_n3116_, new_n3924_ );
and  ( new_n12364_, new_n12363_, new_n12362_ );
and  ( new_n12365_, new_n12364_, new_n3004_ );
and  ( new_n12366_, new_n3120_, RI2b1c4342dfa8_88 );
and  ( new_n12367_, new_n3110_, RI2b1c4342df30_87 );
or   ( new_n12368_, new_n12367_, new_n12366_ );
and  ( new_n12369_, new_n12368_, new_n2868_ );
or   ( new_n12370_, new_n12369_, new_n12365_ );
and  ( new_n12371_, new_n12370_, new_n12361_ );
or   ( new_n12372_, new_n12371_, new_n12360_ );
and  ( new_n12373_, new_n12372_, new_n12341_ );
or   ( new_n12374_, new_n12372_, new_n12341_ );
or   ( new_n12375_, new_n2450_, new_n4635_ );
or   ( new_n12376_, new_n2454_, new_n132_ );
and  ( new_n12377_, new_n12376_, new_n12375_ );
and  ( new_n12378_, new_n12377_, new_n2334_ );
and  ( new_n12379_, new_n2458_, RI2b1c4342e098_90 );
and  ( new_n12380_, new_n2448_, RI2b1c4342e020_89 );
or   ( new_n12381_, new_n12380_, new_n12379_ );
and  ( new_n12382_, new_n12381_, new_n2168_ );
or   ( new_n12383_, new_n12382_, new_n12378_ );
or   ( new_n12384_, new_n1910_, new_n5459_ );
or   ( new_n12385_, new_n1914_, new_n117_ );
and  ( new_n12386_, new_n12385_, new_n12384_ );
and  ( new_n12387_, new_n12386_, new_n1824_ );
and  ( new_n12388_, new_n1918_, RI2b1c4342e188_92 );
and  ( new_n12389_, new_n1908_, RI2b1c4342e110_91 );
or   ( new_n12390_, new_n12389_, new_n12388_ );
and  ( new_n12391_, new_n12390_, new_n1717_ );
or   ( new_n12392_, new_n12391_, new_n12387_ );
and  ( new_n12393_, new_n12392_, new_n12383_ );
or   ( new_n12394_, new_n12392_, new_n12383_ );
or   ( new_n12395_, new_n1425_, new_n6321_ );
or   ( new_n12396_, new_n1429_, new_n6307_ );
and  ( new_n12397_, new_n12396_, new_n12395_ );
and  ( new_n12398_, new_n12397_, new_n1355_ );
and  ( new_n12399_, new_n1433_, RI2b1c4342e278_94 );
and  ( new_n12400_, new_n1423_, RI2b1c4342e200_93 );
or   ( new_n12401_, new_n12400_, new_n12399_ );
and  ( new_n12402_, new_n12401_, new_n1267_ );
or   ( new_n12403_, new_n12402_, new_n12398_ );
and  ( new_n12404_, new_n12403_, new_n12394_ );
or   ( new_n12405_, new_n12404_, new_n12393_ );
and  ( new_n12406_, new_n12405_, new_n12374_ );
or   ( new_n12407_, new_n12406_, new_n12373_ );
or   ( new_n12408_, new_n12208_, new_n12014_ );
and  ( new_n12409_, new_n12408_, new_n12020_ );
and  ( new_n12410_, new_n12204_, new_n12013_ );
and  ( new_n12411_, new_n12207_, new_n12004_ );
or   ( new_n12412_, new_n12411_, new_n12410_ );
and  ( new_n12413_, new_n12412_, new_n12212_ );
or   ( new_n12414_, new_n12413_, new_n12409_ );
or   ( new_n12415_, new_n12253_, new_n12109_ );
and  ( new_n12416_, new_n12415_, new_n12119_ );
and  ( new_n12417_, new_n12249_, new_n12108_ );
and  ( new_n12418_, new_n12252_, new_n12099_ );
or   ( new_n12419_, new_n12418_, new_n12417_ );
and  ( new_n12420_, new_n12419_, new_n12257_ );
or   ( new_n12421_, new_n12420_, new_n12416_ );
and  ( new_n12422_, new_n12421_, new_n12414_ );
or   ( new_n12423_, new_n12421_, new_n12414_ );
or   ( new_n12424_, new_n12228_, new_n12054_ );
and  ( new_n12425_, new_n12424_, new_n12064_ );
and  ( new_n12426_, new_n12224_, new_n12053_ );
and  ( new_n12427_, new_n12227_, new_n12044_ );
or   ( new_n12428_, new_n12427_, new_n12426_ );
and  ( new_n12429_, new_n12428_, new_n12232_ );
or   ( new_n12430_, new_n12429_, new_n12425_ );
and  ( new_n12431_, new_n12430_, new_n12423_ );
or   ( new_n12432_, new_n12431_, new_n12422_ );
and  ( new_n12433_, new_n12432_, new_n12407_ );
or   ( new_n12434_, new_n12432_, new_n12407_ );
or   ( new_n12435_, new_n12270_, new_n12140_ );
and  ( new_n12436_, new_n12435_, new_n12148_ );
and  ( new_n12437_, new_n12266_, new_n12139_ );
and  ( new_n12438_, new_n12269_, new_n12132_ );
or   ( new_n12439_, new_n12438_, new_n12437_ );
and  ( new_n12440_, new_n12439_, new_n12274_ );
or   ( new_n12441_, new_n12440_, new_n12436_ );
and  ( new_n12442_, new_n12441_, new_n12434_ );
or   ( new_n12443_, new_n12442_, new_n12433_ );
and  ( new_n12444_, new_n12443_, new_n12310_ );
or   ( new_n12445_, new_n12443_, new_n12310_ );
or   ( new_n12446_, new_n12263_, new_n12124_ );
and  ( new_n12447_, new_n12446_, new_n12150_ );
and  ( new_n12448_, new_n12261_, new_n12035_ );
and  ( new_n12449_, new_n12221_, new_n12123_ );
or   ( new_n12450_, new_n12449_, new_n12448_ );
and  ( new_n12451_, new_n12450_, new_n12276_ );
or   ( new_n12452_, new_n12451_, new_n12447_ );
and  ( new_n12453_, new_n12452_, new_n12445_ );
or   ( new_n12454_, new_n12453_, new_n12444_ );
and  ( new_n12455_, new_n12454_, new_n12303_ );
or   ( new_n12456_, new_n12454_, new_n12303_ );
or   ( new_n12457_, new_n12280_, new_n12153_ );
and  ( new_n12458_, new_n12457_, new_n12161_ );
and  ( new_n12459_, new_n12278_, new_n11986_ );
and  ( new_n12460_, new_n12198_, new_n12152_ );
or   ( new_n12461_, new_n12460_, new_n12459_ );
and  ( new_n12462_, new_n12461_, new_n12283_ );
or   ( new_n12463_, new_n12462_, new_n12458_ );
and  ( new_n12464_, new_n12463_, new_n12456_ );
or   ( new_n12465_, new_n12464_, new_n12455_ );
and  ( new_n12466_, new_n12465_, new_n12296_ );
and  ( new_n12467_, new_n12301_, new_n11812_ );
and  ( new_n12468_, new_n12297_, new_n11926_ );
or   ( new_n12469_, new_n12468_, new_n12467_ );
and  ( new_n12470_, new_n12308_, new_n11984_ );
and  ( new_n12471_, new_n12304_, new_n12196_ );
or   ( new_n12472_, new_n12471_, new_n12470_ );
and  ( new_n12473_, new_n12317_, new_n5858_ );
and  ( new_n12474_, new_n12313_, new_n6037_ );
or   ( new_n12475_, new_n12474_, new_n12473_ );
and  ( new_n12476_, new_n12326_, new_n6039_ );
and  ( new_n12477_, new_n12322_, new_n5867_ );
or   ( new_n12478_, new_n12477_, new_n12476_ );
and  ( new_n12479_, new_n12478_, new_n12475_ );
or   ( new_n12480_, new_n12478_, new_n12475_ );
and  ( new_n12481_, new_n12337_, new_n5182_ );
and  ( new_n12482_, new_n12333_, new_n5028_ );
or   ( new_n12483_, new_n12482_, new_n12481_ );
and  ( new_n12484_, new_n12483_, new_n12480_ );
or   ( new_n12485_, new_n12484_, new_n12479_ );
and  ( new_n12486_, new_n12348_, new_n4400_ );
and  ( new_n12487_, new_n12344_, new_n4215_ );
or   ( new_n12488_, new_n12487_, new_n12486_ );
and  ( new_n12489_, new_n12357_, new_n3695_ );
and  ( new_n12490_, new_n12353_, new_n3548_ );
or   ( new_n12491_, new_n12490_, new_n12489_ );
and  ( new_n12492_, new_n12491_, new_n12488_ );
or   ( new_n12493_, new_n12491_, new_n12488_ );
and  ( new_n12494_, new_n12368_, new_n3004_ );
and  ( new_n12495_, new_n12364_, new_n2868_ );
or   ( new_n12496_, new_n12495_, new_n12494_ );
and  ( new_n12497_, new_n12496_, new_n12493_ );
or   ( new_n12498_, new_n12497_, new_n12492_ );
and  ( new_n12499_, new_n12498_, new_n12485_ );
or   ( new_n12500_, new_n12498_, new_n12485_ );
and  ( new_n12501_, new_n12381_, new_n2334_ );
and  ( new_n12502_, new_n12377_, new_n2168_ );
or   ( new_n12503_, new_n12502_, new_n12501_ );
and  ( new_n12504_, new_n12390_, new_n1824_ );
and  ( new_n12505_, new_n12386_, new_n1717_ );
or   ( new_n12506_, new_n12505_, new_n12504_ );
and  ( new_n12507_, new_n12506_, new_n12503_ );
or   ( new_n12508_, new_n12506_, new_n12503_ );
and  ( new_n12509_, new_n12401_, new_n1355_ );
and  ( new_n12510_, new_n12397_, new_n1267_ );
or   ( new_n12511_, new_n12510_, new_n12509_ );
and  ( new_n12512_, new_n12511_, new_n12508_ );
or   ( new_n12513_, new_n12512_, new_n12507_ );
and  ( new_n12514_, new_n12513_, new_n12500_ );
or   ( new_n12515_, new_n12514_, new_n12499_ );
and  ( new_n12516_, new_n12412_, new_n12020_ );
and  ( new_n12517_, new_n12408_, new_n12212_ );
or   ( new_n12518_, new_n12517_, new_n12516_ );
and  ( new_n12519_, new_n12419_, new_n12119_ );
and  ( new_n12520_, new_n12415_, new_n12257_ );
or   ( new_n12521_, new_n12520_, new_n12519_ );
and  ( new_n12522_, new_n12521_, new_n12518_ );
or   ( new_n12523_, new_n12521_, new_n12518_ );
and  ( new_n12524_, new_n12428_, new_n12064_ );
and  ( new_n12525_, new_n12424_, new_n12232_ );
or   ( new_n12526_, new_n12525_, new_n12524_ );
and  ( new_n12527_, new_n12526_, new_n12523_ );
or   ( new_n12528_, new_n12527_, new_n12522_ );
and  ( new_n12529_, new_n12528_, new_n12515_ );
or   ( new_n12530_, new_n12528_, new_n12515_ );
and  ( new_n12531_, new_n12439_, new_n12148_ );
and  ( new_n12532_, new_n12435_, new_n12274_ );
or   ( new_n12533_, new_n12532_, new_n12531_ );
and  ( new_n12534_, new_n12533_, new_n12530_ );
or   ( new_n12535_, new_n12534_, new_n12529_ );
and  ( new_n12536_, new_n12535_, new_n12472_ );
or   ( new_n12537_, new_n12535_, new_n12472_ );
and  ( new_n12538_, new_n12450_, new_n12150_ );
and  ( new_n12539_, new_n12446_, new_n12276_ );
or   ( new_n12540_, new_n12539_, new_n12538_ );
and  ( new_n12541_, new_n12540_, new_n12537_ );
or   ( new_n12542_, new_n12541_, new_n12536_ );
and  ( new_n12543_, new_n12542_, new_n12469_ );
or   ( new_n12544_, new_n12543_, new_n12455_ );
and  ( new_n12545_, new_n12544_, new_n12463_ );
and  ( new_n12546_, new_n12542_, new_n12303_ );
and  ( new_n12547_, new_n12469_, new_n12454_ );
or   ( new_n12548_, new_n12547_, new_n12546_ );
and  ( new_n12549_, new_n12461_, new_n12161_ );
and  ( new_n12550_, new_n12457_, new_n12283_ );
or   ( new_n12551_, new_n12550_, new_n12549_ );
and  ( new_n12552_, new_n12551_, new_n12548_ );
or   ( new_n12553_, new_n12552_, new_n12545_ );
or   ( new_n12554_, new_n12246_, new_n12089_ );
and  ( new_n12555_, new_n12554_, new_n12121_ );
and  ( new_n12556_, new_n12244_, new_n12066_ );
and  ( new_n12557_, new_n12234_, new_n12088_ );
or   ( new_n12558_, new_n12557_, new_n12556_ );
and  ( new_n12559_, new_n12558_, new_n12259_ );
or   ( new_n12560_, new_n12559_, new_n12555_ );
or   ( new_n12561_, new_n12529_, new_n12433_ );
and  ( new_n12562_, new_n12561_, new_n12441_ );
and  ( new_n12563_, new_n12515_, new_n12432_ );
and  ( new_n12564_, new_n12528_, new_n12407_ );
or   ( new_n12565_, new_n12564_, new_n12563_ );
and  ( new_n12566_, new_n12565_, new_n12533_ );
or   ( new_n12567_, new_n12566_, new_n12562_ );
or   ( new_n12568_, new_n12567_, new_n12560_ );
or   ( new_n12569_, new_n12522_, new_n12422_ );
and  ( new_n12570_, new_n12569_, new_n12430_ );
and  ( new_n12571_, new_n12518_, new_n12421_ );
and  ( new_n12572_, new_n12521_, new_n12414_ );
or   ( new_n12573_, new_n12572_, new_n12571_ );
and  ( new_n12574_, new_n12573_, new_n12526_ );
or   ( new_n12575_, new_n12574_, new_n12570_ );
or   ( new_n12576_, new_n12499_, new_n12373_ );
and  ( new_n12577_, new_n12576_, new_n12405_ );
and  ( new_n12578_, new_n12485_, new_n12372_ );
and  ( new_n12579_, new_n12498_, new_n12341_ );
or   ( new_n12580_, new_n12579_, new_n12578_ );
and  ( new_n12581_, new_n12580_, new_n12513_ );
or   ( new_n12582_, new_n12581_, new_n12577_ );
or   ( new_n12583_, new_n12582_, new_n12575_ );
or   ( new_n12584_, new_n5308_, new_n121_ );
or   ( new_n12585_, new_n5312_, new_n2119_ );
and  ( new_n12586_, new_n12585_, new_n12584_ );
and  ( new_n12587_, new_n12586_, new_n5182_ );
and  ( new_n12588_, new_n5316_, RI2b1c4342dd50_83 );
and  ( new_n12589_, new_n5306_, RI2b1c4342dcd8_82 );
or   ( new_n12590_, new_n12589_, new_n12588_ );
and  ( new_n12591_, new_n12590_, new_n5028_ );
or   ( new_n12592_, new_n12591_, new_n12587_ );
or   ( new_n12593_, new_n4535_, new_n2806_ );
or   ( new_n12594_, new_n4539_, new_n2541_ );
and  ( new_n12595_, new_n12594_, new_n12593_ );
and  ( new_n12596_, new_n12595_, new_n4400_ );
and  ( new_n12597_, new_n4543_, RI2b1c4342de40_85 );
and  ( new_n12598_, new_n4533_, RI2b1c4342ddc8_84 );
or   ( new_n12599_, new_n12598_, new_n12597_ );
and  ( new_n12600_, new_n12599_, new_n4215_ );
or   ( new_n12601_, new_n12600_, new_n12596_ );
and  ( new_n12602_, new_n12601_, new_n12592_ );
or   ( new_n12603_, new_n12601_, new_n12592_ );
or   ( new_n12604_, new_n3802_, new_n3924_ );
or   ( new_n12605_, new_n3806_, new_n3239_ );
and  ( new_n12606_, new_n12605_, new_n12604_ );
and  ( new_n12607_, new_n12606_, new_n3695_ );
and  ( new_n12608_, new_n3810_, RI2b1c4342df30_87 );
and  ( new_n12609_, new_n3800_, RI2b1c4342deb8_86 );
or   ( new_n12610_, new_n12609_, new_n12608_ );
and  ( new_n12611_, new_n12610_, new_n3548_ );
or   ( new_n12612_, new_n12611_, new_n12607_ );
and  ( new_n12613_, new_n12612_, new_n12603_ );
or   ( new_n12614_, new_n12613_, new_n12602_ );
or   ( new_n12615_, new_n7105_, new_n1310_ );
or   ( new_n12616_, new_n7099_, new_n1002_ );
and  ( new_n12617_, new_n12616_, new_n12615_ );
and  ( new_n12618_, new_n12617_, new_n5858_ );
and  ( new_n12619_, new_n7104_, RI2b1c4342daf8_78 );
and  ( new_n12620_, new_n7110_, RI2b1c4342db70_79 );
or   ( new_n12621_, new_n12620_, new_n12619_ );
and  ( new_n12622_, new_n12621_, new_n6037_ );
or   ( new_n12623_, new_n12622_, new_n12618_ );
and  ( new_n12624_, new_n12623_, new_n913_ );
or   ( new_n12625_, new_n12623_, new_n913_ );
or   ( new_n12626_, new_n6156_, new_n126_ );
or   ( new_n12627_, new_n6160_, new_n1511_ );
and  ( new_n12628_, new_n12627_, new_n12626_ );
and  ( new_n12629_, new_n12628_, new_n6039_ );
and  ( new_n12630_, new_n6164_, RI2b1c4342dc60_81 );
and  ( new_n12631_, new_n6154_, RI2b1c4342dbe8_80 );
or   ( new_n12632_, new_n12631_, new_n12630_ );
and  ( new_n12633_, new_n12632_, new_n5867_ );
or   ( new_n12634_, new_n12633_, new_n12629_ );
and  ( new_n12635_, new_n12634_, new_n12625_ );
or   ( new_n12636_, new_n12635_, new_n12624_ );
and  ( new_n12637_, new_n12636_, new_n12614_ );
or   ( new_n12638_, new_n12636_, new_n12614_ );
or   ( new_n12639_, new_n3112_, new_n132_ );
or   ( new_n12640_, new_n3116_, new_n3902_ );
and  ( new_n12641_, new_n12640_, new_n12639_ );
and  ( new_n12642_, new_n12641_, new_n3004_ );
and  ( new_n12643_, new_n3120_, RI2b1c4342e020_89 );
and  ( new_n12644_, new_n3110_, RI2b1c4342dfa8_88 );
or   ( new_n12645_, new_n12644_, new_n12643_ );
and  ( new_n12646_, new_n12645_, new_n2868_ );
or   ( new_n12647_, new_n12646_, new_n12642_ );
or   ( new_n12648_, new_n2450_, new_n117_ );
or   ( new_n12649_, new_n2454_, new_n4635_ );
and  ( new_n12650_, new_n12649_, new_n12648_ );
and  ( new_n12651_, new_n12650_, new_n2334_ );
and  ( new_n12652_, new_n2458_, RI2b1c4342e110_91 );
and  ( new_n12653_, new_n2448_, RI2b1c4342e098_90 );
or   ( new_n12654_, new_n12653_, new_n12652_ );
and  ( new_n12655_, new_n12654_, new_n2168_ );
or   ( new_n12656_, new_n12655_, new_n12651_ );
and  ( new_n12657_, new_n12656_, new_n12647_ );
or   ( new_n12658_, new_n12656_, new_n12647_ );
or   ( new_n12659_, new_n1910_, new_n6307_ );
or   ( new_n12660_, new_n1914_, new_n5459_ );
and  ( new_n12661_, new_n12660_, new_n12659_ );
and  ( new_n12662_, new_n12661_, new_n1824_ );
and  ( new_n12663_, new_n1918_, RI2b1c4342e200_93 );
and  ( new_n12664_, new_n1908_, RI2b1c4342e188_92 );
or   ( new_n12665_, new_n12664_, new_n12663_ );
and  ( new_n12666_, new_n12665_, new_n1717_ );
or   ( new_n12667_, new_n12666_, new_n12662_ );
and  ( new_n12668_, new_n12667_, new_n12658_ );
or   ( new_n12669_, new_n12668_, new_n12657_ );
and  ( new_n12670_, new_n12669_, new_n12638_ );
or   ( new_n12671_, new_n12670_, new_n12637_ );
or   ( new_n12672_, new_n934_, new_n7274_ );
or   ( new_n12673_, new_n940_, new_n124_ );
and  ( new_n12674_, new_n12673_, new_n12672_ );
and  ( new_n12675_, new_n12674_, new_n913_ );
and  ( new_n12676_, new_n944_, RI2b1c4342e368_96 );
and  ( new_n12677_, new_n932_, RI2b1c4342e2f0_95 );
or   ( new_n12678_, new_n12677_, new_n12676_ );
and  ( new_n12679_, new_n12678_, new_n938_ );
or   ( new_n12680_, new_n12679_, new_n12675_ );
or   ( new_n12681_, new_n12507_, new_n12393_ );
and  ( new_n12682_, new_n12681_, new_n12403_ );
and  ( new_n12683_, new_n12503_, new_n12392_ );
and  ( new_n12684_, new_n12506_, new_n12383_ );
or   ( new_n12685_, new_n12684_, new_n12683_ );
and  ( new_n12686_, new_n12685_, new_n12511_ );
or   ( new_n12687_, new_n12686_, new_n12682_ );
and  ( new_n12688_, new_n12687_, new_n12680_ );
or   ( new_n12689_, new_n12687_, new_n12680_ );
or   ( new_n12690_, new_n12492_, new_n12360_ );
and  ( new_n12691_, new_n12690_, new_n12370_ );
and  ( new_n12692_, new_n12488_, new_n12359_ );
and  ( new_n12693_, new_n12491_, new_n12350_ );
or   ( new_n12694_, new_n12693_, new_n12692_ );
and  ( new_n12695_, new_n12694_, new_n12496_ );
or   ( new_n12696_, new_n12695_, new_n12691_ );
and  ( new_n12697_, new_n12696_, new_n12689_ );
or   ( new_n12698_, new_n12697_, new_n12688_ );
and  ( new_n12699_, new_n12698_, new_n12671_ );
or   ( new_n12700_, new_n12698_, new_n12671_ );
or   ( new_n12701_, new_n12239_, new_n12076_ );
and  ( new_n12702_, new_n12701_, new_n12086_ );
and  ( new_n12703_, new_n12075_, new_n457_ );
and  ( new_n12704_, new_n12237_, new_n428_ );
or   ( new_n12705_, new_n12704_, new_n12703_ );
and  ( new_n12706_, new_n12705_, new_n12242_ );
or   ( new_n12707_, new_n12706_, new_n12702_ );
and  ( new_n12708_, new_n12707_, new_n12700_ );
or   ( new_n12709_, new_n12708_, new_n12699_ );
and  ( new_n12710_, new_n12709_, new_n12583_ );
or   ( new_n12711_, new_n12709_, new_n12583_ );
or   ( new_n12712_, new_n12215_, new_n12023_ );
and  ( new_n12713_, new_n12712_, new_n12033_ );
and  ( new_n12714_, new_n12214_, new_n11995_ );
and  ( new_n12715_, new_n12201_, new_n12022_ );
or   ( new_n12716_, new_n12715_, new_n12714_ );
and  ( new_n12717_, new_n12716_, new_n12219_ );
or   ( new_n12718_, new_n12717_, new_n12713_ );
and  ( new_n12719_, new_n12718_, new_n12711_ );
or   ( new_n12720_, new_n12719_, new_n12710_ );
and  ( new_n12721_, new_n12720_, new_n12568_ );
or   ( new_n12722_, new_n12720_, new_n12568_ );
or   ( new_n12723_, new_n12536_, new_n12444_ );
and  ( new_n12724_, new_n12723_, new_n12452_ );
and  ( new_n12725_, new_n12535_, new_n12310_ );
and  ( new_n12726_, new_n12472_, new_n12443_ );
or   ( new_n12727_, new_n12726_, new_n12725_ );
and  ( new_n12728_, new_n12727_, new_n12540_ );
or   ( new_n12729_, new_n12728_, new_n12724_ );
and  ( new_n12730_, new_n12729_, new_n12722_ );
or   ( new_n12731_, new_n12730_, new_n12721_ );
and  ( new_n12732_, new_n12731_, new_n12553_ );
or   ( new_n12733_, new_n12732_, new_n12466_ );
and  ( new_n12734_, new_n12558_, new_n12121_ );
and  ( new_n12735_, new_n12554_, new_n12259_ );
or   ( new_n12736_, new_n12735_, new_n12734_ );
and  ( new_n12737_, new_n12565_, new_n12441_ );
and  ( new_n12738_, new_n12561_, new_n12533_ );
or   ( new_n12739_, new_n12738_, new_n12737_ );
and  ( new_n12740_, new_n12739_, new_n12736_ );
and  ( new_n12741_, new_n12573_, new_n12430_ );
and  ( new_n12742_, new_n12569_, new_n12526_ );
or   ( new_n12743_, new_n12742_, new_n12741_ );
and  ( new_n12744_, new_n12580_, new_n12405_ );
and  ( new_n12745_, new_n12576_, new_n12513_ );
or   ( new_n12746_, new_n12745_, new_n12744_ );
and  ( new_n12747_, new_n12746_, new_n12743_ );
and  ( new_n12748_, new_n12678_, new_n913_ );
and  ( new_n12749_, new_n12674_, new_n938_ );
or   ( new_n12750_, new_n12749_, new_n12748_ );
and  ( new_n12751_, new_n12685_, new_n12403_ );
and  ( new_n12752_, new_n12681_, new_n12511_ );
or   ( new_n12753_, new_n12752_, new_n12751_ );
and  ( new_n12754_, new_n12753_, new_n12750_ );
or   ( new_n12755_, new_n12753_, new_n12750_ );
and  ( new_n12756_, new_n12694_, new_n12370_ );
and  ( new_n12757_, new_n12690_, new_n12496_ );
or   ( new_n12758_, new_n12757_, new_n12756_ );
and  ( new_n12759_, new_n12758_, new_n12755_ );
or   ( new_n12760_, new_n12759_, new_n12754_ );
and  ( new_n12761_, new_n12590_, new_n5182_ );
and  ( new_n12762_, new_n12586_, new_n5028_ );
or   ( new_n12763_, new_n12762_, new_n12761_ );
and  ( new_n12764_, new_n12599_, new_n4400_ );
and  ( new_n12765_, new_n12595_, new_n4215_ );
or   ( new_n12766_, new_n12765_, new_n12764_ );
and  ( new_n12767_, new_n12766_, new_n12763_ );
or   ( new_n12768_, new_n12766_, new_n12763_ );
and  ( new_n12769_, new_n12610_, new_n3695_ );
and  ( new_n12770_, new_n12606_, new_n3548_ );
or   ( new_n12771_, new_n12770_, new_n12769_ );
and  ( new_n12772_, new_n12771_, new_n12768_ );
or   ( new_n12773_, new_n12772_, new_n12767_ );
and  ( new_n12774_, new_n12621_, new_n5858_ );
and  ( new_n12775_, new_n12617_, new_n6037_ );
or   ( new_n12776_, new_n12775_, new_n12774_ );
or   ( new_n12777_, new_n12776_, new_n938_ );
and  ( new_n12778_, new_n12776_, new_n938_ );
and  ( new_n12779_, new_n12632_, new_n6039_ );
and  ( new_n12780_, new_n12628_, new_n5867_ );
or   ( new_n12781_, new_n12780_, new_n12779_ );
or   ( new_n12782_, new_n12781_, new_n12778_ );
and  ( new_n12783_, new_n12782_, new_n12777_ );
or   ( new_n12784_, new_n12783_, new_n12773_ );
and  ( new_n12785_, new_n12783_, new_n12773_ );
and  ( new_n12786_, new_n12645_, new_n3004_ );
and  ( new_n12787_, new_n12641_, new_n2868_ );
or   ( new_n12788_, new_n12787_, new_n12786_ );
and  ( new_n12789_, new_n12654_, new_n2334_ );
and  ( new_n12790_, new_n12650_, new_n2168_ );
or   ( new_n12791_, new_n12790_, new_n12789_ );
and  ( new_n12792_, new_n12791_, new_n12788_ );
or   ( new_n12793_, new_n12791_, new_n12788_ );
and  ( new_n12794_, new_n12665_, new_n1824_ );
and  ( new_n12795_, new_n12661_, new_n1717_ );
or   ( new_n12796_, new_n12795_, new_n12794_ );
and  ( new_n12797_, new_n12796_, new_n12793_ );
or   ( new_n12798_, new_n12797_, new_n12792_ );
or   ( new_n12799_, new_n12798_, new_n12785_ );
and  ( new_n12800_, new_n12799_, new_n12784_ );
or   ( new_n12801_, new_n12800_, new_n12760_ );
and  ( new_n12802_, new_n12800_, new_n12760_ );
and  ( new_n12803_, new_n12705_, new_n12086_ );
and  ( new_n12804_, new_n12701_, new_n12242_ );
or   ( new_n12805_, new_n12804_, new_n12803_ );
or   ( new_n12806_, new_n12805_, new_n12802_ );
and  ( new_n12807_, new_n12806_, new_n12801_ );
or   ( new_n12808_, new_n12807_, new_n12747_ );
and  ( new_n12809_, new_n12807_, new_n12747_ );
and  ( new_n12810_, new_n12716_, new_n12033_ );
and  ( new_n12811_, new_n12712_, new_n12219_ );
or   ( new_n12812_, new_n12811_, new_n12810_ );
or   ( new_n12813_, new_n12812_, new_n12809_ );
and  ( new_n12814_, new_n12813_, new_n12808_ );
and  ( new_n12815_, new_n12814_, new_n12740_ );
or   ( new_n12816_, new_n12815_, new_n12721_ );
and  ( new_n12817_, new_n12816_, new_n12729_ );
and  ( new_n12818_, new_n12814_, new_n12568_ );
and  ( new_n12819_, new_n12740_, new_n12720_ );
or   ( new_n12820_, new_n12819_, new_n12818_ );
and  ( new_n12821_, new_n12727_, new_n12452_ );
and  ( new_n12822_, new_n12723_, new_n12540_ );
or   ( new_n12823_, new_n12822_, new_n12821_ );
and  ( new_n12824_, new_n12823_, new_n12820_ );
or   ( new_n12825_, new_n12824_, new_n12817_ );
and  ( new_n12826_, new_n12567_, new_n12560_ );
or   ( new_n12827_, new_n12826_, new_n12740_ );
and  ( new_n12828_, new_n12582_, new_n12575_ );
or   ( new_n12829_, new_n12828_, new_n12747_ );
or   ( new_n12830_, new_n7105_, new_n1511_ );
or   ( new_n12831_, new_n7099_, new_n1310_ );
and  ( new_n12832_, new_n12831_, new_n12830_ );
and  ( new_n12833_, new_n12832_, new_n5858_ );
and  ( new_n12834_, new_n7104_, RI2b1c4342db70_79 );
and  ( new_n12835_, new_n7110_, RI2b1c4342dbe8_80 );
or   ( new_n12836_, new_n12835_, new_n12834_ );
and  ( new_n12837_, new_n12836_, new_n6037_ );
or   ( new_n12838_, new_n12837_, new_n12833_ );
or   ( new_n12839_, new_n6156_, new_n2119_ );
or   ( new_n12840_, new_n6160_, new_n126_ );
and  ( new_n12841_, new_n12840_, new_n12839_ );
and  ( new_n12842_, new_n12841_, new_n6039_ );
and  ( new_n12843_, new_n6164_, RI2b1c4342dcd8_82 );
and  ( new_n12844_, new_n6154_, RI2b1c4342dc60_81 );
or   ( new_n12845_, new_n12844_, new_n12843_ );
and  ( new_n12846_, new_n12845_, new_n5867_ );
or   ( new_n12847_, new_n12846_, new_n12842_ );
and  ( new_n12848_, new_n12847_, new_n12838_ );
or   ( new_n12849_, new_n12847_, new_n12838_ );
or   ( new_n12850_, new_n5308_, new_n2541_ );
or   ( new_n12851_, new_n5312_, new_n121_ );
and  ( new_n12852_, new_n12851_, new_n12850_ );
and  ( new_n12853_, new_n12852_, new_n5182_ );
and  ( new_n12854_, new_n5316_, RI2b1c4342ddc8_84 );
and  ( new_n12855_, new_n5306_, RI2b1c4342dd50_83 );
or   ( new_n12856_, new_n12855_, new_n12854_ );
and  ( new_n12857_, new_n12856_, new_n5028_ );
or   ( new_n12858_, new_n12857_, new_n12853_ );
and  ( new_n12859_, new_n12858_, new_n12849_ );
or   ( new_n12860_, new_n12859_, new_n12848_ );
or   ( new_n12861_, new_n4535_, new_n3239_ );
or   ( new_n12862_, new_n4539_, new_n2806_ );
and  ( new_n12863_, new_n12862_, new_n12861_ );
and  ( new_n12864_, new_n12863_, new_n4400_ );
and  ( new_n12865_, new_n4543_, RI2b1c4342deb8_86 );
and  ( new_n12866_, new_n4533_, RI2b1c4342de40_85 );
or   ( new_n12867_, new_n12866_, new_n12865_ );
and  ( new_n12868_, new_n12867_, new_n4215_ );
or   ( new_n12869_, new_n12868_, new_n12864_ );
or   ( new_n12870_, new_n3802_, new_n3902_ );
or   ( new_n12871_, new_n3806_, new_n3924_ );
and  ( new_n12872_, new_n12871_, new_n12870_ );
and  ( new_n12873_, new_n12872_, new_n3695_ );
and  ( new_n12874_, new_n3810_, RI2b1c4342dfa8_88 );
and  ( new_n12875_, new_n3800_, RI2b1c4342df30_87 );
or   ( new_n12876_, new_n12875_, new_n12874_ );
and  ( new_n12877_, new_n12876_, new_n3548_ );
or   ( new_n12878_, new_n12877_, new_n12873_ );
and  ( new_n12879_, new_n12878_, new_n12869_ );
or   ( new_n12880_, new_n12878_, new_n12869_ );
or   ( new_n12881_, new_n3112_, new_n4635_ );
or   ( new_n12882_, new_n3116_, new_n132_ );
and  ( new_n12883_, new_n12882_, new_n12881_ );
and  ( new_n12884_, new_n12883_, new_n3004_ );
and  ( new_n12885_, new_n3120_, RI2b1c4342e098_90 );
and  ( new_n12886_, new_n3110_, RI2b1c4342e020_89 );
or   ( new_n12887_, new_n12886_, new_n12885_ );
and  ( new_n12888_, new_n12887_, new_n2868_ );
or   ( new_n12889_, new_n12888_, new_n12884_ );
and  ( new_n12890_, new_n12889_, new_n12880_ );
or   ( new_n12891_, new_n12890_, new_n12879_ );
and  ( new_n12892_, new_n12891_, new_n12860_ );
or   ( new_n12893_, new_n12891_, new_n12860_ );
or   ( new_n12894_, new_n2450_, new_n5459_ );
or   ( new_n12895_, new_n2454_, new_n117_ );
and  ( new_n12896_, new_n12895_, new_n12894_ );
and  ( new_n12897_, new_n12896_, new_n2334_ );
and  ( new_n12898_, new_n2458_, RI2b1c4342e188_92 );
and  ( new_n12899_, new_n2448_, RI2b1c4342e110_91 );
or   ( new_n12900_, new_n12899_, new_n12898_ );
and  ( new_n12901_, new_n12900_, new_n2168_ );
or   ( new_n12902_, new_n12901_, new_n12897_ );
or   ( new_n12903_, new_n1910_, new_n6321_ );
or   ( new_n12904_, new_n1914_, new_n6307_ );
and  ( new_n12905_, new_n12904_, new_n12903_ );
and  ( new_n12906_, new_n12905_, new_n1824_ );
and  ( new_n12907_, new_n1918_, RI2b1c4342e278_94 );
and  ( new_n12908_, new_n1908_, RI2b1c4342e200_93 );
or   ( new_n12909_, new_n12908_, new_n12907_ );
and  ( new_n12910_, new_n12909_, new_n1717_ );
or   ( new_n12911_, new_n12910_, new_n12906_ );
and  ( new_n12912_, new_n12911_, new_n12902_ );
or   ( new_n12913_, new_n12911_, new_n12902_ );
or   ( new_n12914_, new_n1425_, new_n7274_ );
or   ( new_n12915_, new_n1429_, new_n124_ );
and  ( new_n12916_, new_n12915_, new_n12914_ );
and  ( new_n12917_, new_n12916_, new_n1355_ );
and  ( new_n12918_, new_n1433_, RI2b1c4342e368_96 );
and  ( new_n12919_, new_n1423_, RI2b1c4342e2f0_95 );
or   ( new_n12920_, new_n12919_, new_n12918_ );
and  ( new_n12921_, new_n12920_, new_n1267_ );
or   ( new_n12922_, new_n12921_, new_n12917_ );
and  ( new_n12923_, new_n12922_, new_n12913_ );
or   ( new_n12924_, new_n12923_, new_n12912_ );
and  ( new_n12925_, new_n12924_, new_n12893_ );
or   ( new_n12926_, new_n12925_, new_n12892_ );
or   ( new_n12927_, new_n1425_, new_n124_ );
or   ( new_n12928_, new_n1429_, new_n6321_ );
and  ( new_n12929_, new_n12928_, new_n12927_ );
and  ( new_n12930_, new_n12929_, new_n1355_ );
and  ( new_n12931_, new_n1433_, RI2b1c4342e2f0_95 );
and  ( new_n12932_, new_n1423_, RI2b1c4342e278_94 );
or   ( new_n12933_, new_n12932_, new_n12931_ );
and  ( new_n12934_, new_n12933_, new_n1267_ );
or   ( new_n12935_, new_n12934_, new_n12930_ );
or   ( new_n12936_, new_n940_, new_n7274_ );
and  ( new_n12937_, new_n12936_, new_n913_ );
and  ( new_n12938_, new_n932_, RI2b1c4342e368_96 );
and  ( new_n12939_, new_n12938_, new_n938_ );
or   ( new_n12940_, new_n12939_, new_n12937_ );
and  ( new_n12941_, new_n12940_, new_n12935_ );
or   ( new_n12942_, new_n12940_, new_n12935_ );
or   ( new_n12943_, new_n12792_, new_n12657_ );
and  ( new_n12944_, new_n12943_, new_n12667_ );
and  ( new_n12945_, new_n12788_, new_n12656_ );
and  ( new_n12946_, new_n12791_, new_n12647_ );
or   ( new_n12947_, new_n12946_, new_n12945_ );
and  ( new_n12948_, new_n12947_, new_n12796_ );
or   ( new_n12949_, new_n12948_, new_n12944_ );
and  ( new_n12950_, new_n12949_, new_n12942_ );
or   ( new_n12951_, new_n12950_, new_n12941_ );
and  ( new_n12952_, new_n12951_, new_n12926_ );
or   ( new_n12953_, new_n12951_, new_n12926_ );
or   ( new_n12954_, new_n12479_, new_n12329_ );
and  ( new_n12955_, new_n12954_, new_n12339_ );
and  ( new_n12956_, new_n12475_, new_n12328_ );
and  ( new_n12957_, new_n12478_, new_n12319_ );
or   ( new_n12958_, new_n12957_, new_n12956_ );
and  ( new_n12959_, new_n12958_, new_n12483_ );
or   ( new_n12960_, new_n12959_, new_n12955_ );
and  ( new_n12961_, new_n12960_, new_n12953_ );
or   ( new_n12962_, new_n12961_, new_n12952_ );
and  ( new_n12963_, new_n12962_, new_n12829_ );
or   ( new_n12964_, new_n12962_, new_n12829_ );
or   ( new_n12965_, new_n12802_, new_n12699_ );
and  ( new_n12966_, new_n12965_, new_n12707_ );
and  ( new_n12967_, new_n12800_, new_n12698_ );
and  ( new_n12968_, new_n12760_, new_n12671_ );
or   ( new_n12969_, new_n12968_, new_n12967_ );
and  ( new_n12970_, new_n12969_, new_n12805_ );
or   ( new_n12971_, new_n12970_, new_n12966_ );
and  ( new_n12972_, new_n12971_, new_n12964_ );
or   ( new_n12973_, new_n12972_, new_n12963_ );
and  ( new_n12974_, new_n12973_, new_n12827_ );
or   ( new_n12975_, new_n12973_, new_n12827_ );
or   ( new_n12976_, new_n12809_, new_n12710_ );
and  ( new_n12977_, new_n12976_, new_n12718_ );
and  ( new_n12978_, new_n12807_, new_n12583_ );
and  ( new_n12979_, new_n12747_, new_n12709_ );
or   ( new_n12980_, new_n12979_, new_n12978_ );
and  ( new_n12981_, new_n12980_, new_n12812_ );
or   ( new_n12982_, new_n12981_, new_n12977_ );
and  ( new_n12983_, new_n12982_, new_n12975_ );
or   ( new_n12984_, new_n12983_, new_n12974_ );
and  ( new_n12985_, new_n12984_, new_n12825_ );
and  ( new_n12986_, new_n12736_, new_n12567_ );
and  ( new_n12987_, new_n12739_, new_n12560_ );
or   ( new_n12988_, new_n12987_, new_n12986_ );
and  ( new_n12989_, new_n12743_, new_n12582_ );
and  ( new_n12990_, new_n12746_, new_n12575_ );
or   ( new_n12991_, new_n12990_, new_n12989_ );
and  ( new_n12992_, new_n12836_, new_n5858_ );
and  ( new_n12993_, new_n12832_, new_n6037_ );
or   ( new_n12994_, new_n12993_, new_n12992_ );
and  ( new_n12995_, new_n12845_, new_n6039_ );
and  ( new_n12996_, new_n12841_, new_n5867_ );
or   ( new_n12997_, new_n12996_, new_n12995_ );
and  ( new_n12998_, new_n12997_, new_n12994_ );
or   ( new_n12999_, new_n12997_, new_n12994_ );
and  ( new_n13000_, new_n12856_, new_n5182_ );
and  ( new_n13001_, new_n12852_, new_n5028_ );
or   ( new_n13002_, new_n13001_, new_n13000_ );
and  ( new_n13003_, new_n13002_, new_n12999_ );
or   ( new_n13004_, new_n13003_, new_n12998_ );
and  ( new_n13005_, new_n12867_, new_n4400_ );
and  ( new_n13006_, new_n12863_, new_n4215_ );
or   ( new_n13007_, new_n13006_, new_n13005_ );
and  ( new_n13008_, new_n12876_, new_n3695_ );
and  ( new_n13009_, new_n12872_, new_n3548_ );
or   ( new_n13010_, new_n13009_, new_n13008_ );
and  ( new_n13011_, new_n13010_, new_n13007_ );
or   ( new_n13012_, new_n13010_, new_n13007_ );
and  ( new_n13013_, new_n12887_, new_n3004_ );
and  ( new_n13014_, new_n12883_, new_n2868_ );
or   ( new_n13015_, new_n13014_, new_n13013_ );
and  ( new_n13016_, new_n13015_, new_n13012_ );
or   ( new_n13017_, new_n13016_, new_n13011_ );
and  ( new_n13018_, new_n13017_, new_n13004_ );
or   ( new_n13019_, new_n13017_, new_n13004_ );
and  ( new_n13020_, new_n12900_, new_n2334_ );
and  ( new_n13021_, new_n12896_, new_n2168_ );
or   ( new_n13022_, new_n13021_, new_n13020_ );
and  ( new_n13023_, new_n12909_, new_n1824_ );
and  ( new_n13024_, new_n12905_, new_n1717_ );
or   ( new_n13025_, new_n13024_, new_n13023_ );
and  ( new_n13026_, new_n13025_, new_n13022_ );
or   ( new_n13027_, new_n13025_, new_n13022_ );
and  ( new_n13028_, new_n12920_, new_n1355_ );
and  ( new_n13029_, new_n12916_, new_n1267_ );
or   ( new_n13030_, new_n13029_, new_n13028_ );
and  ( new_n13031_, new_n13030_, new_n13027_ );
or   ( new_n13032_, new_n13031_, new_n13026_ );
and  ( new_n13033_, new_n13032_, new_n13019_ );
or   ( new_n13034_, new_n13033_, new_n13018_ );
and  ( new_n13035_, new_n12933_, new_n1355_ );
and  ( new_n13036_, new_n12929_, new_n1267_ );
or   ( new_n13037_, new_n13036_, new_n13035_ );
and  ( new_n13038_, new_n12938_, new_n913_ );
and  ( new_n13039_, new_n12936_, new_n938_ );
or   ( new_n13040_, new_n13039_, new_n13038_ );
and  ( new_n13041_, new_n13040_, new_n13037_ );
or   ( new_n13042_, new_n13040_, new_n13037_ );
and  ( new_n13043_, new_n12947_, new_n12667_ );
and  ( new_n13044_, new_n12943_, new_n12796_ );
or   ( new_n13045_, new_n13044_, new_n13043_ );
and  ( new_n13046_, new_n13045_, new_n13042_ );
or   ( new_n13047_, new_n13046_, new_n13041_ );
and  ( new_n13048_, new_n13047_, new_n13034_ );
or   ( new_n13049_, new_n13047_, new_n13034_ );
and  ( new_n13050_, new_n12958_, new_n12339_ );
and  ( new_n13051_, new_n12954_, new_n12483_ );
or   ( new_n13052_, new_n13051_, new_n13050_ );
and  ( new_n13053_, new_n13052_, new_n13049_ );
or   ( new_n13054_, new_n13053_, new_n13048_ );
and  ( new_n13055_, new_n13054_, new_n12991_ );
or   ( new_n13056_, new_n13054_, new_n12991_ );
and  ( new_n13057_, new_n12969_, new_n12707_ );
and  ( new_n13058_, new_n12965_, new_n12805_ );
or   ( new_n13059_, new_n13058_, new_n13057_ );
and  ( new_n13060_, new_n13059_, new_n13056_ );
or   ( new_n13061_, new_n13060_, new_n13055_ );
and  ( new_n13062_, new_n13061_, new_n12988_ );
or   ( new_n13063_, new_n13062_, new_n12974_ );
and  ( new_n13064_, new_n13063_, new_n12982_ );
and  ( new_n13065_, new_n13061_, new_n12827_ );
and  ( new_n13066_, new_n12988_, new_n12973_ );
or   ( new_n13067_, new_n13066_, new_n13065_ );
and  ( new_n13068_, new_n12980_, new_n12718_ );
and  ( new_n13069_, new_n12976_, new_n12812_ );
or   ( new_n13070_, new_n13069_, new_n13068_ );
and  ( new_n13071_, new_n13070_, new_n13067_ );
or   ( new_n13072_, new_n13071_, new_n13064_ );
or   ( new_n13073_, new_n12785_, new_n12637_ );
and  ( new_n13074_, new_n13073_, new_n12669_ );
and  ( new_n13075_, new_n12783_, new_n12614_ );
and  ( new_n13076_, new_n12773_, new_n12636_ );
or   ( new_n13077_, new_n13076_, new_n13075_ );
and  ( new_n13078_, new_n13077_, new_n12798_ );
or   ( new_n13079_, new_n13078_, new_n13074_ );
or   ( new_n13080_, new_n13048_, new_n12952_ );
and  ( new_n13081_, new_n13080_, new_n12960_ );
and  ( new_n13082_, new_n13034_, new_n12951_ );
and  ( new_n13083_, new_n13047_, new_n12926_ );
or   ( new_n13084_, new_n13083_, new_n13082_ );
and  ( new_n13085_, new_n13084_, new_n13052_ );
or   ( new_n13086_, new_n13085_, new_n13081_ );
or   ( new_n13087_, new_n13086_, new_n13079_ );
or   ( new_n13088_, new_n12778_, new_n12624_ );
and  ( new_n13089_, new_n13088_, new_n12634_ );
and  ( new_n13090_, new_n12623_, new_n938_ );
and  ( new_n13091_, new_n12776_, new_n913_ );
or   ( new_n13092_, new_n13091_, new_n13090_ );
and  ( new_n13093_, new_n13092_, new_n12781_ );
or   ( new_n13094_, new_n13093_, new_n13089_ );
or   ( new_n13095_, new_n13041_, new_n12941_ );
and  ( new_n13096_, new_n13095_, new_n12949_ );
and  ( new_n13097_, new_n13037_, new_n12940_ );
and  ( new_n13098_, new_n13040_, new_n12935_ );
or   ( new_n13099_, new_n13098_, new_n13097_ );
and  ( new_n13100_, new_n13099_, new_n13045_ );
or   ( new_n13101_, new_n13100_, new_n13096_ );
and  ( new_n13102_, new_n13101_, new_n13094_ );
or   ( new_n13103_, new_n13101_, new_n13094_ );
or   ( new_n13104_, new_n13018_, new_n12892_ );
and  ( new_n13105_, new_n13104_, new_n12924_ );
and  ( new_n13106_, new_n13004_, new_n12891_ );
and  ( new_n13107_, new_n13017_, new_n12860_ );
or   ( new_n13108_, new_n13107_, new_n13106_ );
and  ( new_n13109_, new_n13108_, new_n13032_ );
or   ( new_n13110_, new_n13109_, new_n13105_ );
and  ( new_n13111_, new_n13110_, new_n13103_ );
or   ( new_n13112_, new_n13111_, new_n13102_ );
or   ( new_n13113_, new_n13026_, new_n12912_ );
and  ( new_n13114_, new_n13113_, new_n12922_ );
and  ( new_n13115_, new_n13022_, new_n12911_ );
and  ( new_n13116_, new_n13025_, new_n12902_ );
or   ( new_n13117_, new_n13116_, new_n13115_ );
and  ( new_n13118_, new_n13117_, new_n13030_ );
or   ( new_n13119_, new_n13118_, new_n13114_ );
or   ( new_n13120_, new_n13011_, new_n12879_ );
and  ( new_n13121_, new_n13120_, new_n12889_ );
and  ( new_n13122_, new_n13007_, new_n12878_ );
and  ( new_n13123_, new_n13010_, new_n12869_ );
or   ( new_n13124_, new_n13123_, new_n13122_ );
and  ( new_n13125_, new_n13124_, new_n13015_ );
or   ( new_n13126_, new_n13125_, new_n13121_ );
and  ( new_n13127_, new_n13126_, new_n13119_ );
or   ( new_n13128_, new_n13126_, new_n13119_ );
or   ( new_n13129_, new_n12998_, new_n12848_ );
and  ( new_n13130_, new_n13129_, new_n12858_ );
and  ( new_n13131_, new_n12994_, new_n12847_ );
and  ( new_n13132_, new_n12997_, new_n12838_ );
or   ( new_n13133_, new_n13132_, new_n13131_ );
and  ( new_n13134_, new_n13133_, new_n13002_ );
or   ( new_n13135_, new_n13134_, new_n13130_ );
and  ( new_n13136_, new_n13135_, new_n13128_ );
or   ( new_n13137_, new_n13136_, new_n13127_ );
or   ( new_n13138_, new_n5308_, new_n2806_ );
or   ( new_n13139_, new_n5312_, new_n2541_ );
and  ( new_n13140_, new_n13139_, new_n13138_ );
and  ( new_n13141_, new_n13140_, new_n5182_ );
and  ( new_n13142_, new_n5316_, RI2b1c4342de40_85 );
and  ( new_n13143_, new_n5306_, RI2b1c4342ddc8_84 );
or   ( new_n13144_, new_n13143_, new_n13142_ );
and  ( new_n13145_, new_n13144_, new_n5028_ );
or   ( new_n13146_, new_n13145_, new_n13141_ );
or   ( new_n13147_, new_n4535_, new_n3924_ );
or   ( new_n13148_, new_n4539_, new_n3239_ );
and  ( new_n13149_, new_n13148_, new_n13147_ );
and  ( new_n13150_, new_n13149_, new_n4400_ );
and  ( new_n13151_, new_n4543_, RI2b1c4342df30_87 );
and  ( new_n13152_, new_n4533_, RI2b1c4342deb8_86 );
or   ( new_n13153_, new_n13152_, new_n13151_ );
and  ( new_n13154_, new_n13153_, new_n4215_ );
or   ( new_n13155_, new_n13154_, new_n13150_ );
and  ( new_n13156_, new_n13155_, new_n13146_ );
or   ( new_n13157_, new_n13155_, new_n13146_ );
or   ( new_n13158_, new_n3802_, new_n132_ );
or   ( new_n13159_, new_n3806_, new_n3902_ );
and  ( new_n13160_, new_n13159_, new_n13158_ );
and  ( new_n13161_, new_n13160_, new_n3695_ );
and  ( new_n13162_, new_n3810_, RI2b1c4342e020_89 );
and  ( new_n13163_, new_n3800_, RI2b1c4342dfa8_88 );
or   ( new_n13164_, new_n13163_, new_n13162_ );
and  ( new_n13165_, new_n13164_, new_n3548_ );
or   ( new_n13166_, new_n13165_, new_n13161_ );
and  ( new_n13167_, new_n13166_, new_n13157_ );
or   ( new_n13168_, new_n13167_, new_n13156_ );
or   ( new_n13169_, new_n7105_, new_n126_ );
or   ( new_n13170_, new_n7099_, new_n1511_ );
and  ( new_n13171_, new_n13170_, new_n13169_ );
and  ( new_n13172_, new_n13171_, new_n5858_ );
and  ( new_n13173_, new_n7104_, RI2b1c4342dbe8_80 );
and  ( new_n13174_, new_n7110_, RI2b1c4342dc60_81 );
or   ( new_n13175_, new_n13174_, new_n13173_ );
and  ( new_n13176_, new_n13175_, new_n6037_ );
or   ( new_n13177_, new_n13176_, new_n13172_ );
and  ( new_n13178_, new_n13177_, new_n1355_ );
or   ( new_n13179_, new_n13177_, new_n1355_ );
or   ( new_n13180_, new_n6156_, new_n121_ );
or   ( new_n13181_, new_n6160_, new_n2119_ );
and  ( new_n13182_, new_n13181_, new_n13180_ );
and  ( new_n13183_, new_n13182_, new_n6039_ );
and  ( new_n13184_, new_n6164_, RI2b1c4342dd50_83 );
and  ( new_n13185_, new_n6154_, RI2b1c4342dcd8_82 );
or   ( new_n13186_, new_n13185_, new_n13184_ );
and  ( new_n13187_, new_n13186_, new_n5867_ );
or   ( new_n13188_, new_n13187_, new_n13183_ );
and  ( new_n13189_, new_n13188_, new_n13179_ );
or   ( new_n13190_, new_n13189_, new_n13178_ );
and  ( new_n13191_, new_n13190_, new_n13168_ );
or   ( new_n13192_, new_n13190_, new_n13168_ );
or   ( new_n13193_, new_n3112_, new_n117_ );
or   ( new_n13194_, new_n3116_, new_n4635_ );
and  ( new_n13195_, new_n13194_, new_n13193_ );
and  ( new_n13196_, new_n13195_, new_n3004_ );
and  ( new_n13197_, new_n3120_, RI2b1c4342e110_91 );
and  ( new_n13198_, new_n3110_, RI2b1c4342e098_90 );
or   ( new_n13199_, new_n13198_, new_n13197_ );
and  ( new_n13200_, new_n13199_, new_n2868_ );
or   ( new_n13201_, new_n13200_, new_n13196_ );
or   ( new_n13202_, new_n2450_, new_n6307_ );
or   ( new_n13203_, new_n2454_, new_n5459_ );
and  ( new_n13204_, new_n13203_, new_n13202_ );
and  ( new_n13205_, new_n13204_, new_n2334_ );
and  ( new_n13206_, new_n2458_, RI2b1c4342e200_93 );
and  ( new_n13207_, new_n2448_, RI2b1c4342e188_92 );
or   ( new_n13208_, new_n13207_, new_n13206_ );
and  ( new_n13209_, new_n13208_, new_n2168_ );
or   ( new_n13210_, new_n13209_, new_n13205_ );
and  ( new_n13211_, new_n13210_, new_n13201_ );
or   ( new_n13212_, new_n13210_, new_n13201_ );
or   ( new_n13213_, new_n1910_, new_n124_ );
or   ( new_n13214_, new_n1914_, new_n6321_ );
and  ( new_n13215_, new_n13214_, new_n13213_ );
and  ( new_n13216_, new_n13215_, new_n1824_ );
and  ( new_n13217_, new_n1918_, RI2b1c4342e2f0_95 );
and  ( new_n13218_, new_n1908_, RI2b1c4342e278_94 );
or   ( new_n13219_, new_n13218_, new_n13217_ );
and  ( new_n13220_, new_n13219_, new_n1717_ );
or   ( new_n13221_, new_n13220_, new_n13216_ );
and  ( new_n13222_, new_n13221_, new_n13212_ );
or   ( new_n13223_, new_n13222_, new_n13211_ );
and  ( new_n13224_, new_n13223_, new_n13192_ );
or   ( new_n13225_, new_n13224_, new_n13191_ );
and  ( new_n13226_, new_n13225_, new_n13137_ );
or   ( new_n13227_, new_n13225_, new_n13137_ );
or   ( new_n13228_, new_n12767_, new_n12602_ );
and  ( new_n13229_, new_n13228_, new_n12612_ );
and  ( new_n13230_, new_n12763_, new_n12601_ );
and  ( new_n13231_, new_n12766_, new_n12592_ );
or   ( new_n13232_, new_n13231_, new_n13230_ );
and  ( new_n13233_, new_n13232_, new_n12771_ );
or   ( new_n13234_, new_n13233_, new_n13229_ );
and  ( new_n13235_, new_n13234_, new_n13227_ );
or   ( new_n13236_, new_n13235_, new_n13226_ );
and  ( new_n13237_, new_n13236_, new_n13112_ );
or   ( new_n13238_, new_n13236_, new_n13112_ );
or   ( new_n13239_, new_n12754_, new_n12688_ );
and  ( new_n13240_, new_n13239_, new_n12696_ );
and  ( new_n13241_, new_n12750_, new_n12687_ );
and  ( new_n13242_, new_n12753_, new_n12680_ );
or   ( new_n13243_, new_n13242_, new_n13241_ );
and  ( new_n13244_, new_n13243_, new_n12758_ );
or   ( new_n13245_, new_n13244_, new_n13240_ );
and  ( new_n13246_, new_n13245_, new_n13238_ );
or   ( new_n13247_, new_n13246_, new_n13237_ );
and  ( new_n13248_, new_n13247_, new_n13087_ );
or   ( new_n13249_, new_n13247_, new_n13087_ );
or   ( new_n13250_, new_n13055_, new_n12963_ );
and  ( new_n13251_, new_n13250_, new_n12971_ );
and  ( new_n13252_, new_n13054_, new_n12829_ );
and  ( new_n13253_, new_n12991_, new_n12962_ );
or   ( new_n13254_, new_n13253_, new_n13252_ );
and  ( new_n13255_, new_n13254_, new_n13059_ );
or   ( new_n13256_, new_n13255_, new_n13251_ );
and  ( new_n13257_, new_n13256_, new_n13249_ );
or   ( new_n13258_, new_n13257_, new_n13248_ );
and  ( new_n13259_, new_n13258_, new_n13072_ );
or   ( new_n13260_, new_n13259_, new_n12985_ );
and  ( new_n13261_, new_n13077_, new_n12669_ );
and  ( new_n13262_, new_n13073_, new_n12798_ );
or   ( new_n13263_, new_n13262_, new_n13261_ );
and  ( new_n13264_, new_n13084_, new_n12960_ );
and  ( new_n13265_, new_n13080_, new_n13052_ );
or   ( new_n13266_, new_n13265_, new_n13264_ );
and  ( new_n13267_, new_n13266_, new_n13263_ );
and  ( new_n13268_, new_n13092_, new_n12634_ );
and  ( new_n13269_, new_n13088_, new_n12781_ );
or   ( new_n13270_, new_n13269_, new_n13268_ );
and  ( new_n13271_, new_n13099_, new_n12949_ );
and  ( new_n13272_, new_n13095_, new_n13045_ );
or   ( new_n13273_, new_n13272_, new_n13271_ );
and  ( new_n13274_, new_n13273_, new_n13270_ );
or   ( new_n13275_, new_n13273_, new_n13270_ );
and  ( new_n13276_, new_n13108_, new_n12924_ );
and  ( new_n13277_, new_n13104_, new_n13032_ );
or   ( new_n13278_, new_n13277_, new_n13276_ );
and  ( new_n13279_, new_n13278_, new_n13275_ );
or   ( new_n13280_, new_n13279_, new_n13274_ );
and  ( new_n13281_, new_n13117_, new_n12922_ );
and  ( new_n13282_, new_n13113_, new_n13030_ );
or   ( new_n13283_, new_n13282_, new_n13281_ );
and  ( new_n13284_, new_n13124_, new_n12889_ );
and  ( new_n13285_, new_n13120_, new_n13015_ );
or   ( new_n13286_, new_n13285_, new_n13284_ );
and  ( new_n13287_, new_n13286_, new_n13283_ );
or   ( new_n13288_, new_n13286_, new_n13283_ );
and  ( new_n13289_, new_n13133_, new_n12858_ );
and  ( new_n13290_, new_n13129_, new_n13002_ );
or   ( new_n13291_, new_n13290_, new_n13289_ );
and  ( new_n13292_, new_n13291_, new_n13288_ );
or   ( new_n13293_, new_n13292_, new_n13287_ );
and  ( new_n13294_, new_n13144_, new_n5182_ );
and  ( new_n13295_, new_n13140_, new_n5028_ );
or   ( new_n13296_, new_n13295_, new_n13294_ );
and  ( new_n13297_, new_n13153_, new_n4400_ );
and  ( new_n13298_, new_n13149_, new_n4215_ );
or   ( new_n13299_, new_n13298_, new_n13297_ );
and  ( new_n13300_, new_n13299_, new_n13296_ );
or   ( new_n13301_, new_n13299_, new_n13296_ );
and  ( new_n13302_, new_n13164_, new_n3695_ );
and  ( new_n13303_, new_n13160_, new_n3548_ );
or   ( new_n13304_, new_n13303_, new_n13302_ );
and  ( new_n13305_, new_n13304_, new_n13301_ );
or   ( new_n13306_, new_n13305_, new_n13300_ );
and  ( new_n13307_, new_n13175_, new_n5858_ );
and  ( new_n13308_, new_n13171_, new_n6037_ );
or   ( new_n13309_, new_n13308_, new_n13307_ );
or   ( new_n13310_, new_n13309_, new_n1267_ );
and  ( new_n13311_, new_n13309_, new_n1267_ );
and  ( new_n13312_, new_n13186_, new_n6039_ );
and  ( new_n13313_, new_n13182_, new_n5867_ );
or   ( new_n13314_, new_n13313_, new_n13312_ );
or   ( new_n13315_, new_n13314_, new_n13311_ );
and  ( new_n13316_, new_n13315_, new_n13310_ );
or   ( new_n13317_, new_n13316_, new_n13306_ );
and  ( new_n13318_, new_n13316_, new_n13306_ );
and  ( new_n13319_, new_n13199_, new_n3004_ );
and  ( new_n13320_, new_n13195_, new_n2868_ );
or   ( new_n13321_, new_n13320_, new_n13319_ );
and  ( new_n13322_, new_n13208_, new_n2334_ );
and  ( new_n13323_, new_n13204_, new_n2168_ );
or   ( new_n13324_, new_n13323_, new_n13322_ );
and  ( new_n13325_, new_n13324_, new_n13321_ );
or   ( new_n13326_, new_n13324_, new_n13321_ );
and  ( new_n13327_, new_n13219_, new_n1824_ );
and  ( new_n13328_, new_n13215_, new_n1717_ );
or   ( new_n13329_, new_n13328_, new_n13327_ );
and  ( new_n13330_, new_n13329_, new_n13326_ );
or   ( new_n13331_, new_n13330_, new_n13325_ );
or   ( new_n13332_, new_n13331_, new_n13318_ );
and  ( new_n13333_, new_n13332_, new_n13317_ );
or   ( new_n13334_, new_n13333_, new_n13293_ );
and  ( new_n13335_, new_n13333_, new_n13293_ );
and  ( new_n13336_, new_n13232_, new_n12612_ );
and  ( new_n13337_, new_n13228_, new_n12771_ );
or   ( new_n13338_, new_n13337_, new_n13336_ );
or   ( new_n13339_, new_n13338_, new_n13335_ );
and  ( new_n13340_, new_n13339_, new_n13334_ );
or   ( new_n13341_, new_n13340_, new_n13280_ );
and  ( new_n13342_, new_n13340_, new_n13280_ );
and  ( new_n13343_, new_n13243_, new_n12696_ );
and  ( new_n13344_, new_n13239_, new_n12758_ );
or   ( new_n13345_, new_n13344_, new_n13343_ );
or   ( new_n13346_, new_n13345_, new_n13342_ );
and  ( new_n13347_, new_n13346_, new_n13341_ );
and  ( new_n13348_, new_n13347_, new_n13267_ );
or   ( new_n13349_, new_n13348_, new_n13248_ );
and  ( new_n13350_, new_n13349_, new_n13256_ );
and  ( new_n13351_, new_n13347_, new_n13087_ );
and  ( new_n13352_, new_n13267_, new_n13247_ );
or   ( new_n13353_, new_n13352_, new_n13351_ );
and  ( new_n13354_, new_n13254_, new_n12971_ );
and  ( new_n13355_, new_n13250_, new_n13059_ );
or   ( new_n13356_, new_n13355_, new_n13354_ );
and  ( new_n13357_, new_n13356_, new_n13353_ );
or   ( new_n13358_, new_n13357_, new_n13350_ );
and  ( new_n13359_, new_n13086_, new_n13079_ );
or   ( new_n13360_, new_n13359_, new_n13267_ );
or   ( new_n13361_, new_n13274_, new_n13102_ );
and  ( new_n13362_, new_n13361_, new_n13110_ );
and  ( new_n13363_, new_n13270_, new_n13101_ );
and  ( new_n13364_, new_n13273_, new_n13094_ );
or   ( new_n13365_, new_n13364_, new_n13363_ );
and  ( new_n13366_, new_n13365_, new_n13278_ );
or   ( new_n13367_, new_n13366_, new_n13362_ );
or   ( new_n13368_, new_n7105_, new_n2119_ );
or   ( new_n13369_, new_n7099_, new_n126_ );
and  ( new_n13370_, new_n13369_, new_n13368_ );
and  ( new_n13371_, new_n13370_, new_n5858_ );
and  ( new_n13372_, new_n7104_, RI2b1c4342dc60_81 );
and  ( new_n13373_, new_n7110_, RI2b1c4342dcd8_82 );
or   ( new_n13374_, new_n13373_, new_n13372_ );
and  ( new_n13375_, new_n13374_, new_n6037_ );
or   ( new_n13376_, new_n13375_, new_n13371_ );
or   ( new_n13377_, new_n6156_, new_n2541_ );
or   ( new_n13378_, new_n6160_, new_n121_ );
and  ( new_n13379_, new_n13378_, new_n13377_ );
and  ( new_n13380_, new_n13379_, new_n6039_ );
and  ( new_n13381_, new_n6164_, RI2b1c4342ddc8_84 );
and  ( new_n13382_, new_n6154_, RI2b1c4342dd50_83 );
or   ( new_n13383_, new_n13382_, new_n13381_ );
and  ( new_n13384_, new_n13383_, new_n5867_ );
or   ( new_n13385_, new_n13384_, new_n13380_ );
and  ( new_n13386_, new_n13385_, new_n13376_ );
or   ( new_n13387_, new_n13385_, new_n13376_ );
or   ( new_n13388_, new_n5308_, new_n3239_ );
or   ( new_n13389_, new_n5312_, new_n2806_ );
and  ( new_n13390_, new_n13389_, new_n13388_ );
and  ( new_n13391_, new_n13390_, new_n5182_ );
and  ( new_n13392_, new_n5316_, RI2b1c4342deb8_86 );
and  ( new_n13393_, new_n5306_, RI2b1c4342de40_85 );
or   ( new_n13394_, new_n13393_, new_n13392_ );
and  ( new_n13395_, new_n13394_, new_n5028_ );
or   ( new_n13396_, new_n13395_, new_n13391_ );
and  ( new_n13397_, new_n13396_, new_n13387_ );
or   ( new_n13398_, new_n13397_, new_n13386_ );
or   ( new_n13399_, new_n4535_, new_n3902_ );
or   ( new_n13400_, new_n4539_, new_n3924_ );
and  ( new_n13401_, new_n13400_, new_n13399_ );
and  ( new_n13402_, new_n13401_, new_n4400_ );
and  ( new_n13403_, new_n4543_, RI2b1c4342dfa8_88 );
and  ( new_n13404_, new_n4533_, RI2b1c4342df30_87 );
or   ( new_n13405_, new_n13404_, new_n13403_ );
and  ( new_n13406_, new_n13405_, new_n4215_ );
or   ( new_n13407_, new_n13406_, new_n13402_ );
or   ( new_n13408_, new_n3802_, new_n4635_ );
or   ( new_n13409_, new_n3806_, new_n132_ );
and  ( new_n13410_, new_n13409_, new_n13408_ );
and  ( new_n13411_, new_n13410_, new_n3695_ );
and  ( new_n13412_, new_n3810_, RI2b1c4342e098_90 );
and  ( new_n13413_, new_n3800_, RI2b1c4342e020_89 );
or   ( new_n13414_, new_n13413_, new_n13412_ );
and  ( new_n13415_, new_n13414_, new_n3548_ );
or   ( new_n13416_, new_n13415_, new_n13411_ );
and  ( new_n13417_, new_n13416_, new_n13407_ );
or   ( new_n13418_, new_n13416_, new_n13407_ );
or   ( new_n13419_, new_n3112_, new_n5459_ );
or   ( new_n13420_, new_n3116_, new_n117_ );
and  ( new_n13421_, new_n13420_, new_n13419_ );
and  ( new_n13422_, new_n13421_, new_n3004_ );
and  ( new_n13423_, new_n3120_, RI2b1c4342e188_92 );
and  ( new_n13424_, new_n3110_, RI2b1c4342e110_91 );
or   ( new_n13425_, new_n13424_, new_n13423_ );
and  ( new_n13426_, new_n13425_, new_n2868_ );
or   ( new_n13427_, new_n13426_, new_n13422_ );
and  ( new_n13428_, new_n13427_, new_n13418_ );
or   ( new_n13429_, new_n13428_, new_n13417_ );
and  ( new_n13430_, new_n13429_, new_n13398_ );
or   ( new_n13431_, new_n13429_, new_n13398_ );
or   ( new_n13432_, new_n2450_, new_n6321_ );
or   ( new_n13433_, new_n2454_, new_n6307_ );
and  ( new_n13434_, new_n13433_, new_n13432_ );
and  ( new_n13435_, new_n13434_, new_n2334_ );
and  ( new_n13436_, new_n2458_, RI2b1c4342e278_94 );
and  ( new_n13437_, new_n2448_, RI2b1c4342e200_93 );
or   ( new_n13438_, new_n13437_, new_n13436_ );
and  ( new_n13439_, new_n13438_, new_n2168_ );
or   ( new_n13440_, new_n13439_, new_n13435_ );
or   ( new_n13441_, new_n1910_, new_n7274_ );
or   ( new_n13442_, new_n1914_, new_n124_ );
and  ( new_n13443_, new_n13442_, new_n13441_ );
and  ( new_n13444_, new_n13443_, new_n1824_ );
and  ( new_n13445_, new_n1918_, RI2b1c4342e368_96 );
and  ( new_n13446_, new_n1908_, RI2b1c4342e2f0_95 );
or   ( new_n13447_, new_n13446_, new_n13445_ );
and  ( new_n13448_, new_n13447_, new_n1717_ );
or   ( new_n13449_, new_n13448_, new_n13444_ );
or   ( new_n13450_, new_n13449_, new_n13440_ );
and  ( new_n13451_, new_n13450_, new_n13431_ );
or   ( new_n13452_, new_n13451_, new_n13430_ );
or   ( new_n13453_, new_n1429_, new_n7274_ );
and  ( new_n13454_, new_n13453_, new_n1355_ );
and  ( new_n13455_, new_n1423_, RI2b1c4342e368_96 );
and  ( new_n13456_, new_n13455_, new_n1267_ );
or   ( new_n13457_, new_n13456_, new_n13454_ );
or   ( new_n13458_, new_n13325_, new_n13211_ );
and  ( new_n13459_, new_n13458_, new_n13221_ );
and  ( new_n13460_, new_n13321_, new_n13210_ );
and  ( new_n13461_, new_n13324_, new_n13201_ );
or   ( new_n13462_, new_n13461_, new_n13460_ );
and  ( new_n13463_, new_n13462_, new_n13329_ );
or   ( new_n13464_, new_n13463_, new_n13459_ );
and  ( new_n13465_, new_n13464_, new_n13457_ );
or   ( new_n13466_, new_n13464_, new_n13457_ );
or   ( new_n13467_, new_n13300_, new_n13156_ );
and  ( new_n13468_, new_n13467_, new_n13166_ );
and  ( new_n13469_, new_n13296_, new_n13155_ );
and  ( new_n13470_, new_n13299_, new_n13146_ );
or   ( new_n13471_, new_n13470_, new_n13469_ );
and  ( new_n13472_, new_n13471_, new_n13304_ );
or   ( new_n13473_, new_n13472_, new_n13468_ );
and  ( new_n13474_, new_n13473_, new_n13466_ );
or   ( new_n13475_, new_n13474_, new_n13465_ );
and  ( new_n13476_, new_n13475_, new_n13452_ );
or   ( new_n13477_, new_n13475_, new_n13452_ );
or   ( new_n13478_, new_n13287_, new_n13127_ );
and  ( new_n13479_, new_n13478_, new_n13135_ );
and  ( new_n13480_, new_n13283_, new_n13126_ );
and  ( new_n13481_, new_n13286_, new_n13119_ );
or   ( new_n13482_, new_n13481_, new_n13480_ );
and  ( new_n13483_, new_n13482_, new_n13291_ );
or   ( new_n13484_, new_n13483_, new_n13479_ );
and  ( new_n13485_, new_n13484_, new_n13477_ );
or   ( new_n13486_, new_n13485_, new_n13476_ );
and  ( new_n13487_, new_n13486_, new_n13367_ );
or   ( new_n13488_, new_n13486_, new_n13367_ );
or   ( new_n13489_, new_n13335_, new_n13226_ );
and  ( new_n13490_, new_n13489_, new_n13234_ );
and  ( new_n13491_, new_n13333_, new_n13137_ );
and  ( new_n13492_, new_n13293_, new_n13225_ );
or   ( new_n13493_, new_n13492_, new_n13491_ );
and  ( new_n13494_, new_n13493_, new_n13338_ );
or   ( new_n13495_, new_n13494_, new_n13490_ );
and  ( new_n13496_, new_n13495_, new_n13488_ );
or   ( new_n13497_, new_n13496_, new_n13487_ );
and  ( new_n13498_, new_n13497_, new_n13360_ );
or   ( new_n13499_, new_n13497_, new_n13360_ );
or   ( new_n13500_, new_n13342_, new_n13237_ );
and  ( new_n13501_, new_n13500_, new_n13245_ );
and  ( new_n13502_, new_n13340_, new_n13112_ );
and  ( new_n13503_, new_n13280_, new_n13236_ );
or   ( new_n13504_, new_n13503_, new_n13502_ );
and  ( new_n13505_, new_n13504_, new_n13345_ );
or   ( new_n13506_, new_n13505_, new_n13501_ );
and  ( new_n13507_, new_n13506_, new_n13499_ );
or   ( new_n13508_, new_n13507_, new_n13498_ );
and  ( new_n13509_, new_n13508_, new_n13358_ );
and  ( new_n13510_, new_n13263_, new_n13086_ );
and  ( new_n13511_, new_n13266_, new_n13079_ );
or   ( new_n13512_, new_n13511_, new_n13510_ );
and  ( new_n13513_, new_n13365_, new_n13110_ );
and  ( new_n13514_, new_n13361_, new_n13278_ );
or   ( new_n13515_, new_n13514_, new_n13513_ );
and  ( new_n13516_, new_n13374_, new_n5858_ );
and  ( new_n13517_, new_n13370_, new_n6037_ );
or   ( new_n13518_, new_n13517_, new_n13516_ );
and  ( new_n13519_, new_n13383_, new_n6039_ );
and  ( new_n13520_, new_n13379_, new_n5867_ );
or   ( new_n13521_, new_n13520_, new_n13519_ );
and  ( new_n13522_, new_n13521_, new_n13518_ );
or   ( new_n13523_, new_n13521_, new_n13518_ );
and  ( new_n13524_, new_n13394_, new_n5182_ );
and  ( new_n13525_, new_n13390_, new_n5028_ );
or   ( new_n13526_, new_n13525_, new_n13524_ );
and  ( new_n13527_, new_n13526_, new_n13523_ );
or   ( new_n13528_, new_n13527_, new_n13522_ );
and  ( new_n13529_, new_n13405_, new_n4400_ );
and  ( new_n13530_, new_n13401_, new_n4215_ );
or   ( new_n13531_, new_n13530_, new_n13529_ );
and  ( new_n13532_, new_n13414_, new_n3695_ );
and  ( new_n13533_, new_n13410_, new_n3548_ );
or   ( new_n13534_, new_n13533_, new_n13532_ );
and  ( new_n13535_, new_n13534_, new_n13531_ );
or   ( new_n13536_, new_n13534_, new_n13531_ );
and  ( new_n13537_, new_n13425_, new_n3004_ );
and  ( new_n13538_, new_n13421_, new_n2868_ );
or   ( new_n13539_, new_n13538_, new_n13537_ );
and  ( new_n13540_, new_n13539_, new_n13536_ );
or   ( new_n13541_, new_n13540_, new_n13535_ );
and  ( new_n13542_, new_n13541_, new_n13528_ );
or   ( new_n13543_, new_n13541_, new_n13528_ );
and  ( new_n13544_, new_n13438_, new_n2334_ );
and  ( new_n13545_, new_n13434_, new_n2168_ );
or   ( new_n13546_, new_n13545_, new_n13544_ );
and  ( new_n13547_, new_n13447_, new_n1824_ );
and  ( new_n13548_, new_n13443_, new_n1717_ );
or   ( new_n13549_, new_n13548_, new_n13547_ );
and  ( new_n13550_, new_n13549_, new_n13546_ );
and  ( new_n13551_, new_n13550_, new_n13543_ );
or   ( new_n13552_, new_n13551_, new_n13542_ );
and  ( new_n13553_, new_n13455_, new_n1355_ );
and  ( new_n13554_, new_n13453_, new_n1267_ );
or   ( new_n13555_, new_n13554_, new_n13553_ );
and  ( new_n13556_, new_n13462_, new_n13221_ );
and  ( new_n13557_, new_n13458_, new_n13329_ );
or   ( new_n13558_, new_n13557_, new_n13556_ );
and  ( new_n13559_, new_n13558_, new_n13555_ );
or   ( new_n13560_, new_n13558_, new_n13555_ );
and  ( new_n13561_, new_n13471_, new_n13166_ );
and  ( new_n13562_, new_n13467_, new_n13304_ );
or   ( new_n13563_, new_n13562_, new_n13561_ );
and  ( new_n13564_, new_n13563_, new_n13560_ );
or   ( new_n13565_, new_n13564_, new_n13559_ );
and  ( new_n13566_, new_n13565_, new_n13552_ );
or   ( new_n13567_, new_n13565_, new_n13552_ );
and  ( new_n13568_, new_n13482_, new_n13135_ );
and  ( new_n13569_, new_n13478_, new_n13291_ );
or   ( new_n13570_, new_n13569_, new_n13568_ );
and  ( new_n13571_, new_n13570_, new_n13567_ );
or   ( new_n13572_, new_n13571_, new_n13566_ );
and  ( new_n13573_, new_n13572_, new_n13515_ );
or   ( new_n13574_, new_n13572_, new_n13515_ );
and  ( new_n13575_, new_n13493_, new_n13234_ );
and  ( new_n13576_, new_n13489_, new_n13338_ );
or   ( new_n13577_, new_n13576_, new_n13575_ );
and  ( new_n13578_, new_n13577_, new_n13574_ );
or   ( new_n13579_, new_n13578_, new_n13573_ );
and  ( new_n13580_, new_n13579_, new_n13512_ );
or   ( new_n13581_, new_n13580_, new_n13498_ );
and  ( new_n13582_, new_n13581_, new_n13506_ );
and  ( new_n13583_, new_n13579_, new_n13360_ );
and  ( new_n13584_, new_n13512_, new_n13497_ );
or   ( new_n13585_, new_n13584_, new_n13583_ );
and  ( new_n13586_, new_n13504_, new_n13245_ );
and  ( new_n13587_, new_n13500_, new_n13345_ );
or   ( new_n13588_, new_n13587_, new_n13586_ );
and  ( new_n13589_, new_n13588_, new_n13585_ );
or   ( new_n13590_, new_n13589_, new_n13582_ );
or   ( new_n13591_, new_n13573_, new_n13487_ );
and  ( new_n13592_, new_n13591_, new_n13495_ );
and  ( new_n13593_, new_n13572_, new_n13367_ );
and  ( new_n13594_, new_n13515_, new_n13486_ );
or   ( new_n13595_, new_n13594_, new_n13593_ );
and  ( new_n13596_, new_n13595_, new_n13577_ );
or   ( new_n13597_, new_n13596_, new_n13592_ );
or   ( new_n13598_, new_n13559_, new_n13465_ );
and  ( new_n13599_, new_n13598_, new_n13473_ );
and  ( new_n13600_, new_n13555_, new_n13464_ );
and  ( new_n13601_, new_n13558_, new_n13457_ );
or   ( new_n13602_, new_n13601_, new_n13600_ );
and  ( new_n13603_, new_n13602_, new_n13563_ );
or   ( new_n13604_, new_n13603_, new_n13599_ );
or   ( new_n13605_, new_n13542_, new_n13430_ );
and  ( new_n13606_, new_n13605_, new_n13450_ );
and  ( new_n13607_, new_n13528_, new_n13429_ );
and  ( new_n13608_, new_n13541_, new_n13398_ );
or   ( new_n13609_, new_n13608_, new_n13607_ );
and  ( new_n13610_, new_n13609_, new_n13550_ );
or   ( new_n13611_, new_n13610_, new_n13606_ );
or   ( new_n13612_, new_n13611_, new_n13604_ );
and  ( new_n13613_, new_n13449_, new_n13440_ );
or   ( new_n13614_, new_n13613_, new_n13550_ );
or   ( new_n13615_, new_n13535_, new_n13417_ );
and  ( new_n13616_, new_n13615_, new_n13427_ );
and  ( new_n13617_, new_n13531_, new_n13416_ );
and  ( new_n13618_, new_n13534_, new_n13407_ );
or   ( new_n13619_, new_n13618_, new_n13617_ );
and  ( new_n13620_, new_n13619_, new_n13539_ );
or   ( new_n13621_, new_n13620_, new_n13616_ );
and  ( new_n13622_, new_n13621_, new_n13614_ );
or   ( new_n13623_, new_n13621_, new_n13614_ );
or   ( new_n13624_, new_n13522_, new_n13386_ );
and  ( new_n13625_, new_n13624_, new_n13396_ );
and  ( new_n13626_, new_n13518_, new_n13385_ );
and  ( new_n13627_, new_n13521_, new_n13376_ );
or   ( new_n13628_, new_n13627_, new_n13626_ );
and  ( new_n13629_, new_n13628_, new_n13526_ );
or   ( new_n13630_, new_n13629_, new_n13625_ );
and  ( new_n13631_, new_n13630_, new_n13623_ );
or   ( new_n13632_, new_n13631_, new_n13622_ );
or   ( new_n13633_, new_n4535_, new_n132_ );
or   ( new_n13634_, new_n4539_, new_n3902_ );
and  ( new_n13635_, new_n13634_, new_n13633_ );
and  ( new_n13636_, new_n13635_, new_n4400_ );
and  ( new_n13637_, new_n4543_, RI2b1c4342e020_89 );
and  ( new_n13638_, new_n4533_, RI2b1c4342dfa8_88 );
or   ( new_n13639_, new_n13638_, new_n13637_ );
and  ( new_n13640_, new_n13639_, new_n4215_ );
or   ( new_n13641_, new_n13640_, new_n13636_ );
or   ( new_n13642_, new_n5308_, new_n3924_ );
or   ( new_n13643_, new_n5312_, new_n3239_ );
and  ( new_n13644_, new_n13643_, new_n13642_ );
and  ( new_n13645_, new_n13644_, new_n5182_ );
and  ( new_n13646_, new_n5316_, RI2b1c4342df30_87 );
and  ( new_n13647_, new_n5306_, RI2b1c4342deb8_86 );
or   ( new_n13648_, new_n13647_, new_n13646_ );
and  ( new_n13649_, new_n13648_, new_n5028_ );
or   ( new_n13650_, new_n13649_, new_n13645_ );
and  ( new_n13651_, new_n13650_, new_n13641_ );
or   ( new_n13652_, new_n13650_, new_n13641_ );
or   ( new_n13653_, new_n3802_, new_n117_ );
or   ( new_n13654_, new_n3806_, new_n4635_ );
and  ( new_n13655_, new_n13654_, new_n13653_ );
and  ( new_n13656_, new_n13655_, new_n3695_ );
and  ( new_n13657_, new_n3810_, RI2b1c4342e110_91 );
and  ( new_n13658_, new_n3800_, RI2b1c4342e098_90 );
or   ( new_n13659_, new_n13658_, new_n13657_ );
and  ( new_n13660_, new_n13659_, new_n3548_ );
or   ( new_n13661_, new_n13660_, new_n13656_ );
and  ( new_n13662_, new_n13661_, new_n13652_ );
or   ( new_n13663_, new_n13662_, new_n13651_ );
or   ( new_n13664_, new_n7105_, new_n121_ );
or   ( new_n13665_, new_n7099_, new_n2119_ );
and  ( new_n13666_, new_n13665_, new_n13664_ );
and  ( new_n13667_, new_n13666_, new_n5858_ );
and  ( new_n13668_, new_n7104_, RI2b1c4342dcd8_82 );
and  ( new_n13669_, new_n7110_, RI2b1c4342dd50_83 );
or   ( new_n13670_, new_n13669_, new_n13668_ );
and  ( new_n13671_, new_n13670_, new_n6037_ );
or   ( new_n13672_, new_n13671_, new_n13667_ );
and  ( new_n13673_, new_n13672_, new_n1824_ );
or   ( new_n13674_, new_n13672_, new_n1824_ );
or   ( new_n13675_, new_n6156_, new_n2806_ );
or   ( new_n13676_, new_n6160_, new_n2541_ );
and  ( new_n13677_, new_n13676_, new_n13675_ );
and  ( new_n13678_, new_n13677_, new_n6039_ );
and  ( new_n13679_, new_n6164_, RI2b1c4342de40_85 );
and  ( new_n13680_, new_n6154_, RI2b1c4342ddc8_84 );
or   ( new_n13681_, new_n13680_, new_n13679_ );
and  ( new_n13682_, new_n13681_, new_n5867_ );
or   ( new_n13683_, new_n13682_, new_n13678_ );
and  ( new_n13684_, new_n13683_, new_n13674_ );
or   ( new_n13685_, new_n13684_, new_n13673_ );
and  ( new_n13686_, new_n13685_, new_n13663_ );
or   ( new_n13687_, new_n13685_, new_n13663_ );
or   ( new_n13688_, new_n3112_, new_n6307_ );
or   ( new_n13689_, new_n3116_, new_n5459_ );
and  ( new_n13690_, new_n13689_, new_n13688_ );
and  ( new_n13691_, new_n13690_, new_n3004_ );
and  ( new_n13692_, new_n3120_, RI2b1c4342e200_93 );
and  ( new_n13693_, new_n3110_, RI2b1c4342e188_92 );
or   ( new_n13694_, new_n13693_, new_n13692_ );
and  ( new_n13695_, new_n13694_, new_n2868_ );
or   ( new_n13696_, new_n13695_, new_n13691_ );
or   ( new_n13697_, new_n2450_, new_n124_ );
or   ( new_n13698_, new_n2454_, new_n6321_ );
and  ( new_n13699_, new_n13698_, new_n13697_ );
and  ( new_n13700_, new_n13699_, new_n2334_ );
and  ( new_n13701_, new_n2458_, RI2b1c4342e2f0_95 );
and  ( new_n13702_, new_n2448_, RI2b1c4342e278_94 );
or   ( new_n13703_, new_n13702_, new_n13701_ );
and  ( new_n13704_, new_n13703_, new_n2168_ );
or   ( new_n13705_, new_n13704_, new_n13700_ );
and  ( new_n13706_, new_n13705_, new_n13696_ );
or   ( new_n13707_, new_n13705_, new_n13696_ );
or   ( new_n13708_, new_n1914_, new_n7274_ );
and  ( new_n13709_, new_n13708_, new_n1824_ );
and  ( new_n13710_, new_n1908_, RI2b1c4342e368_96 );
and  ( new_n13711_, new_n13710_, new_n1717_ );
or   ( new_n13712_, new_n13711_, new_n13709_ );
and  ( new_n13713_, new_n13712_, new_n13707_ );
or   ( new_n13714_, new_n13713_, new_n13706_ );
and  ( new_n13715_, new_n13714_, new_n13687_ );
or   ( new_n13716_, new_n13715_, new_n13686_ );
and  ( new_n13717_, new_n13716_, new_n13632_ );
or   ( new_n13718_, new_n13716_, new_n13632_ );
or   ( new_n13719_, new_n13311_, new_n13178_ );
and  ( new_n13720_, new_n13719_, new_n13188_ );
and  ( new_n13721_, new_n13177_, new_n1267_ );
and  ( new_n13722_, new_n13309_, new_n1355_ );
or   ( new_n13723_, new_n13722_, new_n13721_ );
and  ( new_n13724_, new_n13723_, new_n13314_ );
or   ( new_n13725_, new_n13724_, new_n13720_ );
and  ( new_n13726_, new_n13725_, new_n13718_ );
or   ( new_n13727_, new_n13726_, new_n13717_ );
and  ( new_n13728_, new_n13727_, new_n13612_ );
or   ( new_n13729_, new_n13727_, new_n13612_ );
or   ( new_n13730_, new_n13318_, new_n13191_ );
and  ( new_n13731_, new_n13730_, new_n13223_ );
and  ( new_n13732_, new_n13316_, new_n13168_ );
and  ( new_n13733_, new_n13306_, new_n13190_ );
or   ( new_n13734_, new_n13733_, new_n13732_ );
and  ( new_n13735_, new_n13734_, new_n13331_ );
or   ( new_n13736_, new_n13735_, new_n13731_ );
and  ( new_n13737_, new_n13736_, new_n13729_ );
or   ( new_n13738_, new_n13737_, new_n13728_ );
or   ( new_n13739_, new_n13738_, new_n13597_ );
and  ( new_n13740_, new_n13739_, new_n13590_ );
or   ( new_n13741_, new_n13740_, new_n13509_ );
or   ( new_n13742_, new_n13566_, new_n13476_ );
and  ( new_n13743_, new_n13742_, new_n13484_ );
and  ( new_n13744_, new_n13552_, new_n13475_ );
and  ( new_n13745_, new_n13565_, new_n13452_ );
or   ( new_n13746_, new_n13745_, new_n13744_ );
and  ( new_n13747_, new_n13746_, new_n13570_ );
or   ( new_n13748_, new_n13747_, new_n13743_ );
and  ( new_n13749_, new_n13602_, new_n13473_ );
and  ( new_n13750_, new_n13598_, new_n13563_ );
or   ( new_n13751_, new_n13750_, new_n13749_ );
and  ( new_n13752_, new_n13609_, new_n13450_ );
and  ( new_n13753_, new_n13605_, new_n13550_ );
or   ( new_n13754_, new_n13753_, new_n13752_ );
and  ( new_n13755_, new_n13754_, new_n13751_ );
and  ( new_n13756_, new_n13546_, new_n13449_ );
and  ( new_n13757_, new_n13549_, new_n13440_ );
or   ( new_n13758_, new_n13757_, new_n13756_ );
and  ( new_n13759_, new_n13619_, new_n13427_ );
and  ( new_n13760_, new_n13615_, new_n13539_ );
or   ( new_n13761_, new_n13760_, new_n13759_ );
and  ( new_n13762_, new_n13761_, new_n13758_ );
or   ( new_n13763_, new_n13761_, new_n13758_ );
and  ( new_n13764_, new_n13628_, new_n13396_ );
and  ( new_n13765_, new_n13624_, new_n13526_ );
or   ( new_n13766_, new_n13765_, new_n13764_ );
and  ( new_n13767_, new_n13766_, new_n13763_ );
or   ( new_n13768_, new_n13767_, new_n13762_ );
and  ( new_n13769_, new_n13648_, new_n5182_ );
and  ( new_n13770_, new_n13644_, new_n5028_ );
or   ( new_n13771_, new_n13770_, new_n13769_ );
and  ( new_n13772_, new_n13639_, new_n4400_ );
and  ( new_n13773_, new_n13635_, new_n4215_ );
or   ( new_n13774_, new_n13773_, new_n13772_ );
and  ( new_n13775_, new_n13774_, new_n13771_ );
or   ( new_n13776_, new_n13774_, new_n13771_ );
and  ( new_n13777_, new_n13659_, new_n3695_ );
and  ( new_n13778_, new_n13655_, new_n3548_ );
or   ( new_n13779_, new_n13778_, new_n13777_ );
and  ( new_n13780_, new_n13779_, new_n13776_ );
or   ( new_n13781_, new_n13780_, new_n13775_ );
and  ( new_n13782_, new_n13670_, new_n5858_ );
and  ( new_n13783_, new_n13666_, new_n6037_ );
or   ( new_n13784_, new_n13783_, new_n13782_ );
or   ( new_n13785_, new_n13784_, new_n1717_ );
and  ( new_n13786_, new_n13784_, new_n1717_ );
and  ( new_n13787_, new_n13681_, new_n6039_ );
and  ( new_n13788_, new_n13677_, new_n5867_ );
or   ( new_n13789_, new_n13788_, new_n13787_ );
or   ( new_n13790_, new_n13789_, new_n13786_ );
and  ( new_n13791_, new_n13790_, new_n13785_ );
or   ( new_n13792_, new_n13791_, new_n13781_ );
and  ( new_n13793_, new_n13791_, new_n13781_ );
and  ( new_n13794_, new_n13694_, new_n3004_ );
and  ( new_n13795_, new_n13690_, new_n2868_ );
or   ( new_n13796_, new_n13795_, new_n13794_ );
and  ( new_n13797_, new_n13703_, new_n2334_ );
and  ( new_n13798_, new_n13699_, new_n2168_ );
or   ( new_n13799_, new_n13798_, new_n13797_ );
and  ( new_n13800_, new_n13799_, new_n13796_ );
or   ( new_n13801_, new_n13799_, new_n13796_ );
and  ( new_n13802_, new_n13710_, new_n1824_ );
and  ( new_n13803_, new_n13708_, new_n1717_ );
or   ( new_n13804_, new_n13803_, new_n13802_ );
and  ( new_n13805_, new_n13804_, new_n13801_ );
or   ( new_n13806_, new_n13805_, new_n13800_ );
or   ( new_n13807_, new_n13806_, new_n13793_ );
and  ( new_n13808_, new_n13807_, new_n13792_ );
or   ( new_n13809_, new_n13808_, new_n13768_ );
and  ( new_n13810_, new_n13808_, new_n13768_ );
and  ( new_n13811_, new_n13723_, new_n13188_ );
and  ( new_n13812_, new_n13719_, new_n13314_ );
or   ( new_n13813_, new_n13812_, new_n13811_ );
or   ( new_n13814_, new_n13813_, new_n13810_ );
and  ( new_n13815_, new_n13814_, new_n13809_ );
and  ( new_n13816_, new_n13815_, new_n13755_ );
or   ( new_n13817_, new_n13816_, new_n13728_ );
and  ( new_n13818_, new_n13817_, new_n13736_ );
and  ( new_n13819_, new_n13815_, new_n13612_ );
and  ( new_n13820_, new_n13755_, new_n13727_ );
or   ( new_n13821_, new_n13820_, new_n13819_ );
and  ( new_n13822_, new_n13734_, new_n13223_ );
and  ( new_n13823_, new_n13730_, new_n13331_ );
or   ( new_n13824_, new_n13823_, new_n13822_ );
and  ( new_n13825_, new_n13824_, new_n13821_ );
or   ( new_n13826_, new_n13825_, new_n13818_ );
and  ( new_n13827_, new_n13826_, new_n13748_ );
and  ( new_n13828_, new_n13746_, new_n13484_ );
and  ( new_n13829_, new_n13742_, new_n13570_ );
or   ( new_n13830_, new_n13829_, new_n13828_ );
and  ( new_n13831_, new_n13821_, new_n13736_ );
and  ( new_n13832_, new_n13824_, new_n13817_ );
or   ( new_n13833_, new_n13832_, new_n13831_ );
and  ( new_n13834_, new_n13833_, new_n13830_ );
or   ( new_n13835_, new_n13834_, new_n13827_ );
and  ( new_n13836_, new_n13611_, new_n13604_ );
or   ( new_n13837_, new_n13836_, new_n13755_ );
or   ( new_n13838_, new_n13786_, new_n13673_ );
and  ( new_n13839_, new_n13838_, new_n13683_ );
and  ( new_n13840_, new_n13672_, new_n1717_ );
and  ( new_n13841_, new_n13784_, new_n1824_ );
or   ( new_n13842_, new_n13841_, new_n13840_ );
and  ( new_n13843_, new_n13842_, new_n13789_ );
or   ( new_n13844_, new_n13843_, new_n13839_ );
or   ( new_n13845_, new_n13775_, new_n13651_ );
and  ( new_n13846_, new_n13845_, new_n13661_ );
and  ( new_n13847_, new_n13771_, new_n13641_ );
and  ( new_n13848_, new_n13774_, new_n13650_ );
or   ( new_n13849_, new_n13848_, new_n13847_ );
and  ( new_n13850_, new_n13849_, new_n13779_ );
or   ( new_n13851_, new_n13850_, new_n13846_ );
or   ( new_n13852_, new_n13851_, new_n13844_ );
or   ( new_n13853_, new_n7105_, new_n2541_ );
or   ( new_n13854_, new_n7099_, new_n121_ );
and  ( new_n13855_, new_n13854_, new_n13853_ );
and  ( new_n13856_, new_n13855_, new_n5858_ );
and  ( new_n13857_, new_n7104_, RI2b1c4342dd50_83 );
and  ( new_n13858_, new_n7110_, RI2b1c4342ddc8_84 );
or   ( new_n13859_, new_n13858_, new_n13857_ );
and  ( new_n13860_, new_n13859_, new_n6037_ );
or   ( new_n13861_, new_n13860_, new_n13856_ );
or   ( new_n13862_, new_n6156_, new_n3239_ );
or   ( new_n13863_, new_n6160_, new_n2806_ );
and  ( new_n13864_, new_n13863_, new_n13862_ );
and  ( new_n13865_, new_n13864_, new_n6039_ );
and  ( new_n13866_, new_n6164_, RI2b1c4342deb8_86 );
and  ( new_n13867_, new_n6154_, RI2b1c4342de40_85 );
or   ( new_n13868_, new_n13867_, new_n13866_ );
and  ( new_n13869_, new_n13868_, new_n5867_ );
or   ( new_n13870_, new_n13869_, new_n13865_ );
and  ( new_n13871_, new_n13870_, new_n13861_ );
or   ( new_n13872_, new_n13870_, new_n13861_ );
or   ( new_n13873_, new_n5308_, new_n3902_ );
or   ( new_n13874_, new_n5312_, new_n3924_ );
and  ( new_n13875_, new_n13874_, new_n13873_ );
and  ( new_n13876_, new_n13875_, new_n5182_ );
and  ( new_n13877_, new_n5316_, RI2b1c4342dfa8_88 );
and  ( new_n13878_, new_n5306_, RI2b1c4342df30_87 );
or   ( new_n13879_, new_n13878_, new_n13877_ );
and  ( new_n13880_, new_n13879_, new_n5028_ );
or   ( new_n13881_, new_n13880_, new_n13876_ );
and  ( new_n13882_, new_n13881_, new_n13872_ );
or   ( new_n13883_, new_n13882_, new_n13871_ );
or   ( new_n13884_, new_n4535_, new_n4635_ );
or   ( new_n13885_, new_n4539_, new_n132_ );
and  ( new_n13886_, new_n13885_, new_n13884_ );
and  ( new_n13887_, new_n13886_, new_n4400_ );
and  ( new_n13888_, new_n4543_, RI2b1c4342e098_90 );
and  ( new_n13889_, new_n4533_, RI2b1c4342e020_89 );
or   ( new_n13890_, new_n13889_, new_n13888_ );
and  ( new_n13891_, new_n13890_, new_n4215_ );
or   ( new_n13892_, new_n13891_, new_n13887_ );
or   ( new_n13893_, new_n3802_, new_n5459_ );
or   ( new_n13894_, new_n3806_, new_n117_ );
and  ( new_n13895_, new_n13894_, new_n13893_ );
and  ( new_n13896_, new_n13895_, new_n3695_ );
and  ( new_n13897_, new_n3810_, RI2b1c4342e188_92 );
and  ( new_n13898_, new_n3800_, RI2b1c4342e110_91 );
or   ( new_n13899_, new_n13898_, new_n13897_ );
and  ( new_n13900_, new_n13899_, new_n3548_ );
or   ( new_n13901_, new_n13900_, new_n13896_ );
and  ( new_n13902_, new_n13901_, new_n13892_ );
or   ( new_n13903_, new_n13901_, new_n13892_ );
or   ( new_n13904_, new_n3112_, new_n6321_ );
or   ( new_n13905_, new_n3116_, new_n6307_ );
and  ( new_n13906_, new_n13905_, new_n13904_ );
and  ( new_n13907_, new_n13906_, new_n3004_ );
and  ( new_n13908_, new_n3120_, RI2b1c4342e278_94 );
and  ( new_n13909_, new_n3110_, RI2b1c4342e200_93 );
or   ( new_n13910_, new_n13909_, new_n13908_ );
and  ( new_n13911_, new_n13910_, new_n2868_ );
or   ( new_n13912_, new_n13911_, new_n13907_ );
and  ( new_n13913_, new_n13912_, new_n13903_ );
or   ( new_n13914_, new_n13913_, new_n13902_ );
and  ( new_n13915_, new_n13914_, new_n13883_ );
or   ( new_n13916_, new_n13914_, new_n13883_ );
or   ( new_n13917_, new_n13800_, new_n13706_ );
and  ( new_n13918_, new_n13917_, new_n13712_ );
and  ( new_n13919_, new_n13796_, new_n13705_ );
and  ( new_n13920_, new_n13799_, new_n13696_ );
or   ( new_n13921_, new_n13920_, new_n13919_ );
and  ( new_n13922_, new_n13921_, new_n13804_ );
or   ( new_n13923_, new_n13922_, new_n13918_ );
and  ( new_n13924_, new_n13923_, new_n13916_ );
or   ( new_n13925_, new_n13924_, new_n13915_ );
and  ( new_n13926_, new_n13925_, new_n13852_ );
or   ( new_n13927_, new_n13925_, new_n13852_ );
or   ( new_n13928_, new_n13762_, new_n13622_ );
and  ( new_n13929_, new_n13928_, new_n13630_ );
and  ( new_n13930_, new_n13758_, new_n13621_ );
and  ( new_n13931_, new_n13761_, new_n13614_ );
or   ( new_n13932_, new_n13931_, new_n13930_ );
and  ( new_n13933_, new_n13932_, new_n13766_ );
or   ( new_n13934_, new_n13933_, new_n13929_ );
and  ( new_n13935_, new_n13934_, new_n13927_ );
or   ( new_n13936_, new_n13935_, new_n13926_ );
and  ( new_n13937_, new_n13936_, new_n13837_ );
or   ( new_n13938_, new_n13936_, new_n13837_ );
or   ( new_n13939_, new_n13810_, new_n13717_ );
and  ( new_n13940_, new_n13939_, new_n13725_ );
and  ( new_n13941_, new_n13808_, new_n13632_ );
and  ( new_n13942_, new_n13768_, new_n13716_ );
or   ( new_n13943_, new_n13942_, new_n13941_ );
and  ( new_n13944_, new_n13943_, new_n13813_ );
or   ( new_n13945_, new_n13944_, new_n13940_ );
and  ( new_n13946_, new_n13945_, new_n13938_ );
or   ( new_n13947_, new_n13946_, new_n13937_ );
and  ( new_n13948_, new_n13947_, new_n13835_ );
and  ( new_n13949_, new_n13738_, new_n13597_ );
and  ( new_n13950_, new_n13595_, new_n13495_ );
and  ( new_n13951_, new_n13591_, new_n13577_ );
or   ( new_n13952_, new_n13951_, new_n13950_ );
or   ( new_n13953_, new_n13815_, new_n13755_ );
or   ( new_n13954_, new_n13824_, new_n13816_ );
and  ( new_n13955_, new_n13954_, new_n13953_ );
and  ( new_n13956_, new_n13955_, new_n13952_ );
or   ( new_n13957_, new_n13956_, new_n13949_ );
or   ( new_n13958_, new_n13826_, new_n13748_ );
and  ( new_n13959_, new_n13958_, new_n13957_ );
or   ( new_n13960_, new_n13959_, new_n13948_ );
and  ( new_n13961_, new_n13751_, new_n13611_ );
and  ( new_n13962_, new_n13754_, new_n13604_ );
or   ( new_n13963_, new_n13962_, new_n13961_ );
and  ( new_n13964_, new_n13849_, new_n13661_ );
and  ( new_n13965_, new_n13845_, new_n13779_ );
or   ( new_n13966_, new_n13965_, new_n13964_ );
and  ( new_n13967_, new_n13842_, new_n13683_ );
and  ( new_n13968_, new_n13838_, new_n13789_ );
or   ( new_n13969_, new_n13968_, new_n13967_ );
and  ( new_n13970_, new_n13969_, new_n13966_ );
and  ( new_n13971_, new_n13859_, new_n5858_ );
and  ( new_n13972_, new_n13855_, new_n6037_ );
or   ( new_n13973_, new_n13972_, new_n13971_ );
and  ( new_n13974_, new_n13868_, new_n6039_ );
and  ( new_n13975_, new_n13864_, new_n5867_ );
or   ( new_n13976_, new_n13975_, new_n13974_ );
and  ( new_n13977_, new_n13976_, new_n13973_ );
or   ( new_n13978_, new_n13976_, new_n13973_ );
and  ( new_n13979_, new_n13879_, new_n5182_ );
and  ( new_n13980_, new_n13875_, new_n5028_ );
or   ( new_n13981_, new_n13980_, new_n13979_ );
and  ( new_n13982_, new_n13981_, new_n13978_ );
or   ( new_n13983_, new_n13982_, new_n13977_ );
and  ( new_n13984_, new_n13890_, new_n4400_ );
and  ( new_n13985_, new_n13886_, new_n4215_ );
or   ( new_n13986_, new_n13985_, new_n13984_ );
and  ( new_n13987_, new_n13899_, new_n3695_ );
and  ( new_n13988_, new_n13895_, new_n3548_ );
or   ( new_n13989_, new_n13988_, new_n13987_ );
and  ( new_n13990_, new_n13989_, new_n13986_ );
or   ( new_n13991_, new_n13989_, new_n13986_ );
and  ( new_n13992_, new_n13910_, new_n3004_ );
and  ( new_n13993_, new_n13906_, new_n2868_ );
or   ( new_n13994_, new_n13993_, new_n13992_ );
and  ( new_n13995_, new_n13994_, new_n13991_ );
or   ( new_n13996_, new_n13995_, new_n13990_ );
and  ( new_n13997_, new_n13996_, new_n13983_ );
or   ( new_n13998_, new_n13996_, new_n13983_ );
and  ( new_n13999_, new_n13921_, new_n13712_ );
and  ( new_n14000_, new_n13917_, new_n13804_ );
or   ( new_n14001_, new_n14000_, new_n13999_ );
and  ( new_n14002_, new_n14001_, new_n13998_ );
or   ( new_n14003_, new_n14002_, new_n13997_ );
and  ( new_n14004_, new_n14003_, new_n13970_ );
or   ( new_n14005_, new_n14003_, new_n13970_ );
and  ( new_n14006_, new_n13932_, new_n13630_ );
and  ( new_n14007_, new_n13928_, new_n13766_ );
or   ( new_n14008_, new_n14007_, new_n14006_ );
and  ( new_n14009_, new_n14008_, new_n14005_ );
or   ( new_n14010_, new_n14009_, new_n14004_ );
and  ( new_n14011_, new_n14010_, new_n13963_ );
or   ( new_n14012_, new_n14011_, new_n13937_ );
and  ( new_n14013_, new_n14012_, new_n13945_ );
and  ( new_n14014_, new_n14010_, new_n13837_ );
and  ( new_n14015_, new_n13963_, new_n13936_ );
or   ( new_n14016_, new_n14015_, new_n14014_ );
and  ( new_n14017_, new_n13943_, new_n13725_ );
and  ( new_n14018_, new_n13939_, new_n13813_ );
or   ( new_n14019_, new_n14018_, new_n14017_ );
and  ( new_n14020_, new_n14019_, new_n14016_ );
or   ( new_n14021_, new_n14020_, new_n14013_ );
or   ( new_n14022_, new_n13793_, new_n13686_ );
and  ( new_n14023_, new_n14022_, new_n13714_ );
and  ( new_n14024_, new_n13791_, new_n13663_ );
and  ( new_n14025_, new_n13781_, new_n13685_ );
or   ( new_n14026_, new_n14025_, new_n14024_ );
and  ( new_n14027_, new_n14026_, new_n13806_ );
or   ( new_n14028_, new_n14027_, new_n14023_ );
and  ( new_n14029_, new_n13851_, new_n13844_ );
or   ( new_n14030_, new_n14029_, new_n13970_ );
or   ( new_n14031_, new_n5308_, new_n132_ );
or   ( new_n14032_, new_n5312_, new_n3902_ );
and  ( new_n14033_, new_n14032_, new_n14031_ );
and  ( new_n14034_, new_n14033_, new_n5182_ );
and  ( new_n14035_, new_n5316_, RI2b1c4342e020_89 );
and  ( new_n14036_, new_n5306_, RI2b1c4342dfa8_88 );
or   ( new_n14037_, new_n14036_, new_n14035_ );
and  ( new_n14038_, new_n14037_, new_n5028_ );
or   ( new_n14039_, new_n14038_, new_n14034_ );
or   ( new_n14040_, new_n4535_, new_n117_ );
or   ( new_n14041_, new_n4539_, new_n4635_ );
and  ( new_n14042_, new_n14041_, new_n14040_ );
and  ( new_n14043_, new_n14042_, new_n4400_ );
and  ( new_n14044_, new_n4543_, RI2b1c4342e110_91 );
and  ( new_n14045_, new_n4533_, RI2b1c4342e098_90 );
or   ( new_n14046_, new_n14045_, new_n14044_ );
and  ( new_n14047_, new_n14046_, new_n4215_ );
or   ( new_n14048_, new_n14047_, new_n14043_ );
and  ( new_n14049_, new_n14048_, new_n14039_ );
or   ( new_n14050_, new_n14048_, new_n14039_ );
or   ( new_n14051_, new_n3802_, new_n6307_ );
or   ( new_n14052_, new_n3806_, new_n5459_ );
and  ( new_n14053_, new_n14052_, new_n14051_ );
and  ( new_n14054_, new_n14053_, new_n3695_ );
and  ( new_n14055_, new_n3810_, RI2b1c4342e200_93 );
and  ( new_n14056_, new_n3800_, RI2b1c4342e188_92 );
or   ( new_n14057_, new_n14056_, new_n14055_ );
and  ( new_n14058_, new_n14057_, new_n3548_ );
or   ( new_n14059_, new_n14058_, new_n14054_ );
and  ( new_n14060_, new_n14059_, new_n14050_ );
or   ( new_n14061_, new_n14060_, new_n14049_ );
or   ( new_n14062_, new_n7105_, new_n2806_ );
or   ( new_n14063_, new_n7099_, new_n2541_ );
and  ( new_n14064_, new_n14063_, new_n14062_ );
and  ( new_n14065_, new_n14064_, new_n5858_ );
and  ( new_n14066_, new_n7104_, RI2b1c4342ddc8_84 );
and  ( new_n14067_, new_n7110_, RI2b1c4342de40_85 );
or   ( new_n14068_, new_n14067_, new_n14066_ );
and  ( new_n14069_, new_n14068_, new_n6037_ );
or   ( new_n14070_, new_n14069_, new_n14065_ );
and  ( new_n14071_, new_n14070_, new_n2334_ );
or   ( new_n14072_, new_n14070_, new_n2334_ );
or   ( new_n14073_, new_n6156_, new_n3924_ );
or   ( new_n14074_, new_n6160_, new_n3239_ );
and  ( new_n14075_, new_n14074_, new_n14073_ );
and  ( new_n14076_, new_n14075_, new_n6039_ );
and  ( new_n14077_, new_n6164_, RI2b1c4342df30_87 );
and  ( new_n14078_, new_n6154_, RI2b1c4342deb8_86 );
or   ( new_n14079_, new_n14078_, new_n14077_ );
and  ( new_n14080_, new_n14079_, new_n5867_ );
or   ( new_n14081_, new_n14080_, new_n14076_ );
and  ( new_n14082_, new_n14081_, new_n14072_ );
or   ( new_n14083_, new_n14082_, new_n14071_ );
and  ( new_n14084_, new_n14083_, new_n14061_ );
or   ( new_n14085_, new_n14083_, new_n14061_ );
or   ( new_n14086_, new_n2450_, new_n7274_ );
or   ( new_n14087_, new_n2454_, new_n124_ );
and  ( new_n14088_, new_n14087_, new_n14086_ );
and  ( new_n14089_, new_n14088_, new_n2334_ );
and  ( new_n14090_, new_n2458_, RI2b1c4342e368_96 );
and  ( new_n14091_, new_n2448_, RI2b1c4342e2f0_95 );
or   ( new_n14092_, new_n14091_, new_n14090_ );
and  ( new_n14093_, new_n14092_, new_n2168_ );
or   ( new_n14094_, new_n14093_, new_n14089_ );
and  ( new_n14095_, new_n14094_, new_n14085_ );
or   ( new_n14096_, new_n14095_, new_n14084_ );
and  ( new_n14097_, new_n14096_, new_n14030_ );
or   ( new_n14098_, new_n14096_, new_n14030_ );
or   ( new_n14099_, new_n13997_, new_n13915_ );
and  ( new_n14100_, new_n14099_, new_n13923_ );
and  ( new_n14101_, new_n13983_, new_n13914_ );
and  ( new_n14102_, new_n13996_, new_n13883_ );
or   ( new_n14103_, new_n14102_, new_n14101_ );
and  ( new_n14104_, new_n14103_, new_n14001_ );
or   ( new_n14105_, new_n14104_, new_n14100_ );
and  ( new_n14106_, new_n14105_, new_n14098_ );
or   ( new_n14107_, new_n14106_, new_n14097_ );
and  ( new_n14108_, new_n14107_, new_n14028_ );
or   ( new_n14109_, new_n14107_, new_n14028_ );
or   ( new_n14110_, new_n14004_, new_n13926_ );
and  ( new_n14111_, new_n14110_, new_n13934_ );
and  ( new_n14112_, new_n14003_, new_n13852_ );
and  ( new_n14113_, new_n13970_, new_n13925_ );
or   ( new_n14114_, new_n14113_, new_n14112_ );
and  ( new_n14115_, new_n14114_, new_n14008_ );
or   ( new_n14116_, new_n14115_, new_n14111_ );
and  ( new_n14117_, new_n14116_, new_n14109_ );
or   ( new_n14118_, new_n14117_, new_n14108_ );
and  ( new_n14119_, new_n14118_, new_n14021_ );
and  ( new_n14120_, new_n14026_, new_n13714_ );
and  ( new_n14121_, new_n14022_, new_n13806_ );
or   ( new_n14122_, new_n14121_, new_n14120_ );
and  ( new_n14123_, new_n13966_, new_n13844_ );
and  ( new_n14124_, new_n13969_, new_n13851_ );
or   ( new_n14125_, new_n14124_, new_n14123_ );
and  ( new_n14126_, new_n14037_, new_n5182_ );
and  ( new_n14127_, new_n14033_, new_n5028_ );
or   ( new_n14128_, new_n14127_, new_n14126_ );
and  ( new_n14129_, new_n14046_, new_n4400_ );
and  ( new_n14130_, new_n14042_, new_n4215_ );
or   ( new_n14131_, new_n14130_, new_n14129_ );
and  ( new_n14132_, new_n14131_, new_n14128_ );
or   ( new_n14133_, new_n14131_, new_n14128_ );
and  ( new_n14134_, new_n14057_, new_n3695_ );
and  ( new_n14135_, new_n14053_, new_n3548_ );
or   ( new_n14136_, new_n14135_, new_n14134_ );
and  ( new_n14137_, new_n14136_, new_n14133_ );
or   ( new_n14138_, new_n14137_, new_n14132_ );
and  ( new_n14139_, new_n14068_, new_n5858_ );
and  ( new_n14140_, new_n14064_, new_n6037_ );
or   ( new_n14141_, new_n14140_, new_n14139_ );
or   ( new_n14142_, new_n14141_, new_n2168_ );
and  ( new_n14143_, new_n14141_, new_n2168_ );
and  ( new_n14144_, new_n14079_, new_n6039_ );
and  ( new_n14145_, new_n14075_, new_n5867_ );
or   ( new_n14146_, new_n14145_, new_n14144_ );
or   ( new_n14147_, new_n14146_, new_n14143_ );
and  ( new_n14148_, new_n14147_, new_n14142_ );
or   ( new_n14149_, new_n14148_, new_n14138_ );
and  ( new_n14150_, new_n14148_, new_n14138_ );
and  ( new_n14151_, new_n14092_, new_n2334_ );
and  ( new_n14152_, new_n14088_, new_n2168_ );
or   ( new_n14153_, new_n14152_, new_n14151_ );
or   ( new_n14154_, new_n14153_, new_n14150_ );
and  ( new_n14155_, new_n14154_, new_n14149_ );
or   ( new_n14156_, new_n14155_, new_n14125_ );
and  ( new_n14157_, new_n14155_, new_n14125_ );
and  ( new_n14158_, new_n14103_, new_n13923_ );
and  ( new_n14159_, new_n14099_, new_n14001_ );
or   ( new_n14160_, new_n14159_, new_n14158_ );
or   ( new_n14161_, new_n14160_, new_n14157_ );
and  ( new_n14162_, new_n14161_, new_n14156_ );
and  ( new_n14163_, new_n14162_, new_n14122_ );
or   ( new_n14164_, new_n14163_, new_n14108_ );
and  ( new_n14165_, new_n14164_, new_n14116_ );
and  ( new_n14166_, new_n14162_, new_n14028_ );
and  ( new_n14167_, new_n14122_, new_n14107_ );
or   ( new_n14168_, new_n14167_, new_n14166_ );
and  ( new_n14169_, new_n14114_, new_n13934_ );
and  ( new_n14170_, new_n14110_, new_n14008_ );
or   ( new_n14171_, new_n14170_, new_n14169_ );
and  ( new_n14172_, new_n14171_, new_n14168_ );
or   ( new_n14173_, new_n14172_, new_n14165_ );
or   ( new_n14174_, new_n13977_, new_n13871_ );
and  ( new_n14175_, new_n14174_, new_n13881_ );
and  ( new_n14176_, new_n13973_, new_n13870_ );
and  ( new_n14177_, new_n13976_, new_n13861_ );
or   ( new_n14178_, new_n14177_, new_n14176_ );
and  ( new_n14179_, new_n14178_, new_n13981_ );
or   ( new_n14180_, new_n14179_, new_n14175_ );
or   ( new_n14181_, new_n14150_, new_n14084_ );
and  ( new_n14182_, new_n14181_, new_n14094_ );
and  ( new_n14183_, new_n14148_, new_n14061_ );
and  ( new_n14184_, new_n14138_, new_n14083_ );
or   ( new_n14185_, new_n14184_, new_n14183_ );
and  ( new_n14186_, new_n14185_, new_n14153_ );
or   ( new_n14187_, new_n14186_, new_n14182_ );
or   ( new_n14188_, new_n14187_, new_n14180_ );
or   ( new_n14189_, new_n7105_, new_n3239_ );
or   ( new_n14190_, new_n7099_, new_n2806_ );
and  ( new_n14191_, new_n14190_, new_n14189_ );
and  ( new_n14192_, new_n14191_, new_n5858_ );
and  ( new_n14193_, new_n7104_, RI2b1c4342de40_85 );
and  ( new_n14194_, new_n7110_, RI2b1c4342deb8_86 );
or   ( new_n14195_, new_n14194_, new_n14193_ );
and  ( new_n14196_, new_n14195_, new_n6037_ );
or   ( new_n14197_, new_n14196_, new_n14192_ );
or   ( new_n14198_, new_n6156_, new_n3902_ );
or   ( new_n14199_, new_n6160_, new_n3924_ );
and  ( new_n14200_, new_n14199_, new_n14198_ );
and  ( new_n14201_, new_n14200_, new_n6039_ );
and  ( new_n14202_, new_n6164_, RI2b1c4342dfa8_88 );
and  ( new_n14203_, new_n6154_, RI2b1c4342df30_87 );
or   ( new_n14204_, new_n14203_, new_n14202_ );
and  ( new_n14205_, new_n14204_, new_n5867_ );
or   ( new_n14206_, new_n14205_, new_n14201_ );
and  ( new_n14207_, new_n14206_, new_n14197_ );
or   ( new_n14208_, new_n14206_, new_n14197_ );
or   ( new_n14209_, new_n5308_, new_n4635_ );
or   ( new_n14210_, new_n5312_, new_n132_ );
and  ( new_n14211_, new_n14210_, new_n14209_ );
and  ( new_n14212_, new_n14211_, new_n5182_ );
and  ( new_n14213_, new_n5316_, RI2b1c4342e098_90 );
and  ( new_n14214_, new_n5306_, RI2b1c4342e020_89 );
or   ( new_n14215_, new_n14214_, new_n14213_ );
and  ( new_n14216_, new_n14215_, new_n5028_ );
or   ( new_n14217_, new_n14216_, new_n14212_ );
and  ( new_n14218_, new_n14217_, new_n14208_ );
or   ( new_n14219_, new_n14218_, new_n14207_ );
or   ( new_n14220_, new_n4535_, new_n5459_ );
or   ( new_n14221_, new_n4539_, new_n117_ );
and  ( new_n14222_, new_n14221_, new_n14220_ );
and  ( new_n14223_, new_n14222_, new_n4400_ );
and  ( new_n14224_, new_n4543_, RI2b1c4342e188_92 );
and  ( new_n14225_, new_n4533_, RI2b1c4342e110_91 );
or   ( new_n14226_, new_n14225_, new_n14224_ );
and  ( new_n14227_, new_n14226_, new_n4215_ );
or   ( new_n14228_, new_n14227_, new_n14223_ );
or   ( new_n14229_, new_n3802_, new_n6321_ );
or   ( new_n14230_, new_n3806_, new_n6307_ );
and  ( new_n14231_, new_n14230_, new_n14229_ );
and  ( new_n14232_, new_n14231_, new_n3695_ );
and  ( new_n14233_, new_n3810_, RI2b1c4342e278_94 );
and  ( new_n14234_, new_n3800_, RI2b1c4342e200_93 );
or   ( new_n14235_, new_n14234_, new_n14233_ );
and  ( new_n14236_, new_n14235_, new_n3548_ );
or   ( new_n14237_, new_n14236_, new_n14232_ );
and  ( new_n14238_, new_n14237_, new_n14228_ );
or   ( new_n14239_, new_n14237_, new_n14228_ );
or   ( new_n14240_, new_n3112_, new_n7274_ );
or   ( new_n14241_, new_n3116_, new_n124_ );
and  ( new_n14242_, new_n14241_, new_n14240_ );
and  ( new_n14243_, new_n14242_, new_n3004_ );
and  ( new_n14244_, new_n3120_, RI2b1c4342e368_96 );
and  ( new_n14245_, new_n3110_, RI2b1c4342e2f0_95 );
or   ( new_n14246_, new_n14245_, new_n14244_ );
and  ( new_n14247_, new_n14246_, new_n2868_ );
or   ( new_n14248_, new_n14247_, new_n14243_ );
and  ( new_n14249_, new_n14248_, new_n14239_ );
or   ( new_n14250_, new_n14249_, new_n14238_ );
and  ( new_n14251_, new_n14250_, new_n14219_ );
or   ( new_n14252_, new_n14250_, new_n14219_ );
or   ( new_n14253_, new_n3112_, new_n124_ );
or   ( new_n14254_, new_n3116_, new_n6321_ );
and  ( new_n14255_, new_n14254_, new_n14253_ );
and  ( new_n14256_, new_n14255_, new_n3004_ );
and  ( new_n14257_, new_n3120_, RI2b1c4342e2f0_95 );
and  ( new_n14258_, new_n3110_, RI2b1c4342e278_94 );
or   ( new_n14259_, new_n14258_, new_n14257_ );
and  ( new_n14260_, new_n14259_, new_n2868_ );
or   ( new_n14261_, new_n14260_, new_n14256_ );
and  ( new_n14262_, new_n14261_, new_n14252_ );
or   ( new_n14263_, new_n14262_, new_n14251_ );
or   ( new_n14264_, new_n2454_, new_n7274_ );
and  ( new_n14265_, new_n14264_, new_n2334_ );
and  ( new_n14266_, new_n2448_, RI2b1c4342e368_96 );
and  ( new_n14267_, new_n14266_, new_n2168_ );
or   ( new_n14268_, new_n14267_, new_n14265_ );
or   ( new_n14269_, new_n14132_, new_n14049_ );
and  ( new_n14270_, new_n14269_, new_n14059_ );
and  ( new_n14271_, new_n14128_, new_n14048_ );
and  ( new_n14272_, new_n14131_, new_n14039_ );
or   ( new_n14273_, new_n14272_, new_n14271_ );
and  ( new_n14274_, new_n14273_, new_n14136_ );
or   ( new_n14275_, new_n14274_, new_n14270_ );
and  ( new_n14276_, new_n14275_, new_n14268_ );
or   ( new_n14277_, new_n14275_, new_n14268_ );
or   ( new_n14278_, new_n14143_, new_n14071_ );
and  ( new_n14279_, new_n14278_, new_n14081_ );
and  ( new_n14280_, new_n14070_, new_n2168_ );
and  ( new_n14281_, new_n14141_, new_n2334_ );
or   ( new_n14282_, new_n14281_, new_n14280_ );
and  ( new_n14283_, new_n14282_, new_n14146_ );
or   ( new_n14284_, new_n14283_, new_n14279_ );
and  ( new_n14285_, new_n14284_, new_n14277_ );
or   ( new_n14286_, new_n14285_, new_n14276_ );
and  ( new_n14287_, new_n14286_, new_n14263_ );
or   ( new_n14288_, new_n14286_, new_n14263_ );
or   ( new_n14289_, new_n13990_, new_n13902_ );
and  ( new_n14290_, new_n14289_, new_n13912_ );
and  ( new_n14291_, new_n13986_, new_n13901_ );
and  ( new_n14292_, new_n13989_, new_n13892_ );
or   ( new_n14293_, new_n14292_, new_n14291_ );
and  ( new_n14294_, new_n14293_, new_n13994_ );
or   ( new_n14295_, new_n14294_, new_n14290_ );
and  ( new_n14296_, new_n14295_, new_n14288_ );
or   ( new_n14297_, new_n14296_, new_n14287_ );
and  ( new_n14298_, new_n14297_, new_n14188_ );
or   ( new_n14299_, new_n14297_, new_n14188_ );
or   ( new_n14300_, new_n14157_, new_n14097_ );
and  ( new_n14301_, new_n14300_, new_n14105_ );
and  ( new_n14302_, new_n14155_, new_n14030_ );
and  ( new_n14303_, new_n14125_, new_n14096_ );
or   ( new_n14304_, new_n14303_, new_n14302_ );
and  ( new_n14305_, new_n14304_, new_n14160_ );
or   ( new_n14306_, new_n14305_, new_n14301_ );
and  ( new_n14307_, new_n14306_, new_n14299_ );
or   ( new_n14308_, new_n14307_, new_n14298_ );
and  ( new_n14309_, new_n14308_, new_n14173_ );
or   ( new_n14310_, new_n14309_, new_n14119_ );
and  ( new_n14311_, new_n14187_, new_n14180_ );
and  ( new_n14312_, new_n14178_, new_n13881_ );
and  ( new_n14313_, new_n14174_, new_n13981_ );
or   ( new_n14314_, new_n14313_, new_n14312_ );
and  ( new_n14315_, new_n14185_, new_n14094_ );
and  ( new_n14316_, new_n14181_, new_n14153_ );
or   ( new_n14317_, new_n14316_, new_n14315_ );
and  ( new_n14318_, new_n14317_, new_n14314_ );
or   ( new_n14319_, new_n14318_, new_n14311_ );
and  ( new_n14320_, new_n14266_, new_n2334_ );
and  ( new_n14321_, new_n14264_, new_n2168_ );
or   ( new_n14322_, new_n14321_, new_n14320_ );
and  ( new_n14323_, new_n14273_, new_n14059_ );
and  ( new_n14324_, new_n14269_, new_n14136_ );
or   ( new_n14325_, new_n14324_, new_n14323_ );
and  ( new_n14326_, new_n14325_, new_n14322_ );
or   ( new_n14327_, new_n14326_, new_n14276_ );
and  ( new_n14328_, new_n14327_, new_n14284_ );
and  ( new_n14329_, new_n14322_, new_n14275_ );
and  ( new_n14330_, new_n14325_, new_n14268_ );
or   ( new_n14331_, new_n14330_, new_n14329_ );
and  ( new_n14332_, new_n14282_, new_n14081_ );
and  ( new_n14333_, new_n14278_, new_n14146_ );
or   ( new_n14334_, new_n14333_, new_n14332_ );
and  ( new_n14335_, new_n14334_, new_n14331_ );
or   ( new_n14336_, new_n14335_, new_n14328_ );
or   ( new_n14337_, new_n5308_, new_n117_ );
or   ( new_n14338_, new_n5312_, new_n4635_ );
and  ( new_n14339_, new_n14338_, new_n14337_ );
and  ( new_n14340_, new_n14339_, new_n5182_ );
and  ( new_n14341_, new_n5316_, RI2b1c4342e110_91 );
and  ( new_n14342_, new_n5306_, RI2b1c4342e098_90 );
or   ( new_n14343_, new_n14342_, new_n14341_ );
and  ( new_n14344_, new_n14343_, new_n5028_ );
or   ( new_n14345_, new_n14344_, new_n14340_ );
or   ( new_n14346_, new_n4535_, new_n6307_ );
or   ( new_n14347_, new_n4539_, new_n5459_ );
and  ( new_n14348_, new_n14347_, new_n14346_ );
and  ( new_n14349_, new_n14348_, new_n4400_ );
and  ( new_n14350_, new_n4543_, RI2b1c4342e200_93 );
and  ( new_n14351_, new_n4533_, RI2b1c4342e188_92 );
or   ( new_n14352_, new_n14351_, new_n14350_ );
and  ( new_n14353_, new_n14352_, new_n4215_ );
or   ( new_n14354_, new_n14353_, new_n14349_ );
and  ( new_n14355_, new_n14354_, new_n14345_ );
or   ( new_n14356_, new_n14354_, new_n14345_ );
or   ( new_n14357_, new_n3802_, new_n124_ );
or   ( new_n14358_, new_n3806_, new_n6321_ );
and  ( new_n14359_, new_n14358_, new_n14357_ );
and  ( new_n14360_, new_n14359_, new_n3695_ );
and  ( new_n14361_, new_n3810_, RI2b1c4342e2f0_95 );
and  ( new_n14362_, new_n3800_, RI2b1c4342e278_94 );
or   ( new_n14363_, new_n14362_, new_n14361_ );
and  ( new_n14364_, new_n14363_, new_n3548_ );
or   ( new_n14365_, new_n14364_, new_n14360_ );
and  ( new_n14366_, new_n14365_, new_n14356_ );
or   ( new_n14367_, new_n14366_, new_n14355_ );
or   ( new_n14368_, new_n7105_, new_n3924_ );
or   ( new_n14369_, new_n7099_, new_n3239_ );
and  ( new_n14370_, new_n14369_, new_n14368_ );
and  ( new_n14371_, new_n14370_, new_n5858_ );
and  ( new_n14372_, new_n7104_, RI2b1c4342deb8_86 );
and  ( new_n14373_, new_n7110_, RI2b1c4342df30_87 );
or   ( new_n14374_, new_n14373_, new_n14372_ );
and  ( new_n14375_, new_n14374_, new_n6037_ );
or   ( new_n14376_, new_n14375_, new_n14371_ );
and  ( new_n14377_, new_n14376_, new_n3004_ );
or   ( new_n14378_, new_n14376_, new_n3004_ );
or   ( new_n14379_, new_n6156_, new_n132_ );
or   ( new_n14380_, new_n6160_, new_n3902_ );
and  ( new_n14381_, new_n14380_, new_n14379_ );
and  ( new_n14382_, new_n14381_, new_n6039_ );
and  ( new_n14383_, new_n6164_, RI2b1c4342e020_89 );
and  ( new_n14384_, new_n6154_, RI2b1c4342dfa8_88 );
or   ( new_n14385_, new_n14384_, new_n14383_ );
and  ( new_n14386_, new_n14385_, new_n5867_ );
or   ( new_n14387_, new_n14386_, new_n14382_ );
and  ( new_n14388_, new_n14387_, new_n14378_ );
or   ( new_n14389_, new_n14388_, new_n14377_ );
and  ( new_n14390_, new_n14389_, new_n14367_ );
or   ( new_n14391_, new_n14389_, new_n14367_ );
and  ( new_n14392_, new_n14226_, new_n4400_ );
and  ( new_n14393_, new_n14222_, new_n4215_ );
or   ( new_n14394_, new_n14393_, new_n14392_ );
and  ( new_n14395_, new_n14235_, new_n3695_ );
and  ( new_n14396_, new_n14231_, new_n3548_ );
or   ( new_n14397_, new_n14396_, new_n14395_ );
and  ( new_n14398_, new_n14397_, new_n14394_ );
or   ( new_n14399_, new_n14398_, new_n14238_ );
and  ( new_n14400_, new_n14399_, new_n14248_ );
and  ( new_n14401_, new_n14394_, new_n14237_ );
and  ( new_n14402_, new_n14397_, new_n14228_ );
or   ( new_n14403_, new_n14402_, new_n14401_ );
and  ( new_n14404_, new_n14246_, new_n3004_ );
and  ( new_n14405_, new_n14242_, new_n2868_ );
or   ( new_n14406_, new_n14405_, new_n14404_ );
and  ( new_n14407_, new_n14406_, new_n14403_ );
or   ( new_n14408_, new_n14407_, new_n14400_ );
and  ( new_n14409_, new_n14408_, new_n14391_ );
or   ( new_n14410_, new_n14409_, new_n14390_ );
and  ( new_n14411_, new_n14410_, new_n14336_ );
or   ( new_n14412_, new_n14410_, new_n14336_ );
and  ( new_n14413_, new_n14195_, new_n5858_ );
and  ( new_n14414_, new_n14191_, new_n6037_ );
or   ( new_n14415_, new_n14414_, new_n14413_ );
and  ( new_n14416_, new_n14204_, new_n6039_ );
and  ( new_n14417_, new_n14200_, new_n5867_ );
or   ( new_n14418_, new_n14417_, new_n14416_ );
and  ( new_n14419_, new_n14418_, new_n14415_ );
or   ( new_n14420_, new_n14418_, new_n14415_ );
and  ( new_n14421_, new_n14215_, new_n5182_ );
and  ( new_n14422_, new_n14211_, new_n5028_ );
or   ( new_n14423_, new_n14422_, new_n14421_ );
and  ( new_n14424_, new_n14423_, new_n14420_ );
or   ( new_n14425_, new_n14424_, new_n14419_ );
or   ( new_n14426_, new_n14397_, new_n14394_ );
and  ( new_n14427_, new_n14426_, new_n14406_ );
or   ( new_n14428_, new_n14427_, new_n14398_ );
and  ( new_n14429_, new_n14428_, new_n14425_ );
or   ( new_n14430_, new_n14429_, new_n14251_ );
and  ( new_n14431_, new_n14430_, new_n14261_ );
and  ( new_n14432_, new_n14425_, new_n14250_ );
and  ( new_n14433_, new_n14428_, new_n14219_ );
or   ( new_n14434_, new_n14433_, new_n14432_ );
and  ( new_n14435_, new_n14259_, new_n3004_ );
and  ( new_n14436_, new_n14255_, new_n2868_ );
or   ( new_n14437_, new_n14436_, new_n14435_ );
and  ( new_n14438_, new_n14437_, new_n14434_ );
or   ( new_n14439_, new_n14438_, new_n14431_ );
and  ( new_n14440_, new_n14439_, new_n14412_ );
or   ( new_n14441_, new_n14440_, new_n14411_ );
and  ( new_n14442_, new_n14441_, new_n14319_ );
and  ( new_n14443_, new_n14314_, new_n14187_ );
and  ( new_n14444_, new_n14317_, new_n14180_ );
or   ( new_n14445_, new_n14444_, new_n14443_ );
and  ( new_n14446_, new_n14331_, new_n14284_ );
and  ( new_n14447_, new_n14334_, new_n14327_ );
or   ( new_n14448_, new_n14447_, new_n14446_ );
and  ( new_n14449_, new_n14343_, new_n5182_ );
and  ( new_n14450_, new_n14339_, new_n5028_ );
or   ( new_n14451_, new_n14450_, new_n14449_ );
and  ( new_n14452_, new_n14352_, new_n4400_ );
and  ( new_n14453_, new_n14348_, new_n4215_ );
or   ( new_n14454_, new_n14453_, new_n14452_ );
and  ( new_n14455_, new_n14454_, new_n14451_ );
or   ( new_n14456_, new_n14454_, new_n14451_ );
and  ( new_n14457_, new_n14363_, new_n3695_ );
and  ( new_n14458_, new_n14359_, new_n3548_ );
or   ( new_n14459_, new_n14458_, new_n14457_ );
and  ( new_n14460_, new_n14459_, new_n14456_ );
or   ( new_n14461_, new_n14460_, new_n14455_ );
and  ( new_n14462_, new_n14374_, new_n5858_ );
and  ( new_n14463_, new_n14370_, new_n6037_ );
or   ( new_n14464_, new_n14463_, new_n14462_ );
or   ( new_n14465_, new_n14464_, new_n2868_ );
and  ( new_n14466_, new_n14464_, new_n2868_ );
and  ( new_n14467_, new_n14385_, new_n6039_ );
and  ( new_n14468_, new_n14381_, new_n5867_ );
or   ( new_n14469_, new_n14468_, new_n14467_ );
or   ( new_n14470_, new_n14469_, new_n14466_ );
and  ( new_n14471_, new_n14470_, new_n14465_ );
or   ( new_n14472_, new_n14471_, new_n14461_ );
and  ( new_n14473_, new_n14471_, new_n14461_ );
and  ( new_n14474_, new_n14403_, new_n14248_ );
and  ( new_n14475_, new_n14406_, new_n14399_ );
or   ( new_n14476_, new_n14475_, new_n14474_ );
or   ( new_n14477_, new_n14476_, new_n14473_ );
and  ( new_n14478_, new_n14477_, new_n14472_ );
or   ( new_n14479_, new_n14478_, new_n14448_ );
and  ( new_n14480_, new_n14478_, new_n14448_ );
and  ( new_n14481_, new_n14434_, new_n14261_ );
and  ( new_n14482_, new_n14437_, new_n14430_ );
or   ( new_n14483_, new_n14482_, new_n14481_ );
or   ( new_n14484_, new_n14483_, new_n14480_ );
and  ( new_n14485_, new_n14484_, new_n14479_ );
and  ( new_n14486_, new_n14485_, new_n14445_ );
or   ( new_n14487_, new_n14486_, new_n14442_ );
or   ( new_n14488_, new_n14428_, new_n14425_ );
and  ( new_n14489_, new_n14488_, new_n14437_ );
or   ( new_n14490_, new_n14489_, new_n14429_ );
or   ( new_n14491_, new_n14325_, new_n14322_ );
and  ( new_n14492_, new_n14491_, new_n14334_ );
or   ( new_n14493_, new_n14492_, new_n14326_ );
and  ( new_n14494_, new_n14493_, new_n14490_ );
or   ( new_n14495_, new_n14494_, new_n14287_ );
and  ( new_n14496_, new_n14495_, new_n14295_ );
and  ( new_n14497_, new_n14490_, new_n14286_ );
and  ( new_n14498_, new_n14493_, new_n14263_ );
or   ( new_n14499_, new_n14498_, new_n14497_ );
and  ( new_n14500_, new_n14293_, new_n13912_ );
and  ( new_n14501_, new_n14289_, new_n13994_ );
or   ( new_n14502_, new_n14501_, new_n14500_ );
and  ( new_n14503_, new_n14502_, new_n14499_ );
or   ( new_n14504_, new_n14503_, new_n14496_ );
and  ( new_n14505_, new_n14504_, new_n14487_ );
and  ( new_n14506_, new_n14485_, new_n14319_ );
and  ( new_n14507_, new_n14445_, new_n14441_ );
or   ( new_n14508_, new_n14507_, new_n14506_ );
and  ( new_n14509_, new_n14499_, new_n14295_ );
and  ( new_n14510_, new_n14502_, new_n14495_ );
or   ( new_n14511_, new_n14510_, new_n14509_ );
and  ( new_n14512_, new_n14511_, new_n14508_ );
or   ( new_n14513_, new_n14512_, new_n14505_ );
or   ( new_n14514_, new_n14480_, new_n14411_ );
and  ( new_n14515_, new_n14514_, new_n14439_ );
and  ( new_n14516_, new_n14478_, new_n14336_ );
and  ( new_n14517_, new_n14448_, new_n14410_ );
or   ( new_n14518_, new_n14517_, new_n14516_ );
and  ( new_n14519_, new_n14518_, new_n14483_ );
or   ( new_n14520_, new_n14519_, new_n14515_ );
or   ( new_n14521_, new_n14419_, new_n14207_ );
and  ( new_n14522_, new_n14521_, new_n14217_ );
and  ( new_n14523_, new_n14415_, new_n14206_ );
and  ( new_n14524_, new_n14418_, new_n14197_ );
or   ( new_n14525_, new_n14524_, new_n14523_ );
and  ( new_n14526_, new_n14525_, new_n14423_ );
or   ( new_n14527_, new_n14526_, new_n14522_ );
or   ( new_n14528_, new_n3116_, new_n7274_ );
and  ( new_n14529_, new_n14528_, new_n3004_ );
and  ( new_n14530_, new_n3110_, RI2b1c4342e368_96 );
and  ( new_n14531_, new_n14530_, new_n2868_ );
or   ( new_n14532_, new_n14531_, new_n14529_ );
or   ( new_n14533_, new_n7105_, new_n3902_ );
or   ( new_n14534_, new_n7099_, new_n3924_ );
and  ( new_n14535_, new_n14534_, new_n14533_ );
and  ( new_n14536_, new_n14535_, new_n5858_ );
and  ( new_n14537_, new_n7104_, RI2b1c4342df30_87 );
and  ( new_n14538_, new_n7110_, RI2b1c4342dfa8_88 );
or   ( new_n14539_, new_n14538_, new_n14537_ );
and  ( new_n14540_, new_n14539_, new_n6037_ );
or   ( new_n14541_, new_n14540_, new_n14536_ );
or   ( new_n14542_, new_n6156_, new_n4635_ );
or   ( new_n14543_, new_n6160_, new_n132_ );
and  ( new_n14544_, new_n14543_, new_n14542_ );
and  ( new_n14545_, new_n14544_, new_n6039_ );
and  ( new_n14546_, new_n6164_, RI2b1c4342e098_90 );
and  ( new_n14547_, new_n6154_, RI2b1c4342e020_89 );
or   ( new_n14548_, new_n14547_, new_n14546_ );
and  ( new_n14549_, new_n14548_, new_n5867_ );
or   ( new_n14550_, new_n14549_, new_n14545_ );
and  ( new_n14551_, new_n14550_, new_n14541_ );
or   ( new_n14552_, new_n14550_, new_n14541_ );
or   ( new_n14553_, new_n5308_, new_n5459_ );
or   ( new_n14554_, new_n5312_, new_n117_ );
and  ( new_n14555_, new_n14554_, new_n14553_ );
and  ( new_n14556_, new_n14555_, new_n5182_ );
and  ( new_n14557_, new_n5316_, RI2b1c4342e188_92 );
and  ( new_n14558_, new_n5306_, RI2b1c4342e110_91 );
or   ( new_n14559_, new_n14558_, new_n14557_ );
and  ( new_n14560_, new_n14559_, new_n5028_ );
or   ( new_n14561_, new_n14560_, new_n14556_ );
and  ( new_n14562_, new_n14561_, new_n14552_ );
or   ( new_n14563_, new_n14562_, new_n14551_ );
and  ( new_n14564_, new_n14563_, new_n14532_ );
or   ( new_n14565_, new_n14563_, new_n14532_ );
or   ( new_n14566_, new_n14455_, new_n14355_ );
and  ( new_n14567_, new_n14566_, new_n14365_ );
and  ( new_n14568_, new_n14451_, new_n14354_ );
and  ( new_n14569_, new_n14454_, new_n14345_ );
or   ( new_n14570_, new_n14569_, new_n14568_ );
and  ( new_n14571_, new_n14570_, new_n14459_ );
or   ( new_n14572_, new_n14571_, new_n14567_ );
and  ( new_n14573_, new_n14572_, new_n14565_ );
or   ( new_n14574_, new_n14573_, new_n14564_ );
and  ( new_n14575_, new_n14574_, new_n14527_ );
or   ( new_n14576_, new_n14574_, new_n14527_ );
or   ( new_n14577_, new_n14473_, new_n14390_ );
and  ( new_n14578_, new_n14577_, new_n14408_ );
and  ( new_n14579_, new_n14471_, new_n14367_ );
and  ( new_n14580_, new_n14461_, new_n14389_ );
or   ( new_n14581_, new_n14580_, new_n14579_ );
and  ( new_n14582_, new_n14581_, new_n14476_ );
or   ( new_n14583_, new_n14582_, new_n14578_ );
and  ( new_n14584_, new_n14583_, new_n14576_ );
or   ( new_n14585_, new_n14584_, new_n14575_ );
or   ( new_n14586_, new_n14585_, new_n14520_ );
and  ( new_n14587_, new_n14586_, new_n14513_ );
or   ( new_n14588_, new_n14493_, new_n14490_ );
and  ( new_n14589_, new_n14588_, new_n14502_ );
or   ( new_n14590_, new_n14589_, new_n14494_ );
and  ( new_n14591_, new_n14590_, new_n14318_ );
or   ( new_n14592_, new_n14591_, new_n14298_ );
and  ( new_n14593_, new_n14592_, new_n14306_ );
and  ( new_n14594_, new_n14590_, new_n14188_ );
and  ( new_n14595_, new_n14318_, new_n14297_ );
or   ( new_n14596_, new_n14595_, new_n14594_ );
and  ( new_n14597_, new_n14304_, new_n14105_ );
and  ( new_n14598_, new_n14300_, new_n14160_ );
or   ( new_n14599_, new_n14598_, new_n14597_ );
and  ( new_n14600_, new_n14599_, new_n14596_ );
or   ( new_n14601_, new_n14600_, new_n14593_ );
or   ( new_n14602_, new_n14441_, new_n14319_ );
and  ( new_n14603_, new_n14602_, new_n14504_ );
or   ( new_n14604_, new_n14603_, new_n14442_ );
and  ( new_n14605_, new_n14604_, new_n14601_ );
or   ( new_n14606_, new_n14605_, new_n14587_ );
and  ( new_n14607_, new_n14585_, new_n14520_ );
and  ( new_n14608_, new_n14518_, new_n14439_ );
and  ( new_n14609_, new_n14514_, new_n14483_ );
or   ( new_n14610_, new_n14609_, new_n14608_ );
and  ( new_n14611_, new_n14525_, new_n14217_ );
and  ( new_n14612_, new_n14521_, new_n14423_ );
or   ( new_n14613_, new_n14612_, new_n14611_ );
and  ( new_n14614_, new_n14530_, new_n3004_ );
and  ( new_n14615_, new_n14528_, new_n2868_ );
or   ( new_n14616_, new_n14615_, new_n14614_ );
and  ( new_n14617_, new_n14539_, new_n5858_ );
and  ( new_n14618_, new_n14535_, new_n6037_ );
or   ( new_n14619_, new_n14618_, new_n14617_ );
and  ( new_n14620_, new_n14548_, new_n6039_ );
and  ( new_n14621_, new_n14544_, new_n5867_ );
or   ( new_n14622_, new_n14621_, new_n14620_ );
and  ( new_n14623_, new_n14622_, new_n14619_ );
or   ( new_n14624_, new_n14622_, new_n14619_ );
and  ( new_n14625_, new_n14559_, new_n5182_ );
and  ( new_n14626_, new_n14555_, new_n5028_ );
or   ( new_n14627_, new_n14626_, new_n14625_ );
and  ( new_n14628_, new_n14627_, new_n14624_ );
or   ( new_n14629_, new_n14628_, new_n14623_ );
and  ( new_n14630_, new_n14629_, new_n14616_ );
or   ( new_n14631_, new_n14629_, new_n14616_ );
and  ( new_n14632_, new_n14570_, new_n14365_ );
and  ( new_n14633_, new_n14566_, new_n14459_ );
or   ( new_n14634_, new_n14633_, new_n14632_ );
and  ( new_n14635_, new_n14634_, new_n14631_ );
or   ( new_n14636_, new_n14635_, new_n14630_ );
and  ( new_n14637_, new_n14636_, new_n14613_ );
or   ( new_n14638_, new_n14636_, new_n14613_ );
and  ( new_n14639_, new_n14581_, new_n14408_ );
and  ( new_n14640_, new_n14577_, new_n14476_ );
or   ( new_n14641_, new_n14640_, new_n14639_ );
and  ( new_n14642_, new_n14641_, new_n14638_ );
or   ( new_n14643_, new_n14642_, new_n14637_ );
and  ( new_n14644_, new_n14643_, new_n14610_ );
or   ( new_n14645_, new_n14644_, new_n14607_ );
or   ( new_n14646_, new_n14637_, new_n14575_ );
and  ( new_n14647_, new_n14646_, new_n14583_ );
and  ( new_n14648_, new_n14636_, new_n14527_ );
and  ( new_n14649_, new_n14613_, new_n14574_ );
or   ( new_n14650_, new_n14649_, new_n14648_ );
and  ( new_n14651_, new_n14650_, new_n14641_ );
or   ( new_n14652_, new_n14651_, new_n14647_ );
or   ( new_n14653_, new_n3802_, new_n7274_ );
or   ( new_n14654_, new_n3806_, new_n124_ );
and  ( new_n14655_, new_n14654_, new_n14653_ );
and  ( new_n14656_, new_n14655_, new_n3695_ );
and  ( new_n14657_, new_n3810_, RI2b1c4342e368_96 );
and  ( new_n14658_, new_n3800_, RI2b1c4342e2f0_95 );
or   ( new_n14659_, new_n14658_, new_n14657_ );
and  ( new_n14660_, new_n14659_, new_n3548_ );
or   ( new_n14661_, new_n14660_, new_n14656_ );
or   ( new_n14662_, new_n14623_, new_n14551_ );
and  ( new_n14663_, new_n14662_, new_n14561_ );
and  ( new_n14664_, new_n14619_, new_n14550_ );
and  ( new_n14665_, new_n14622_, new_n14541_ );
or   ( new_n14666_, new_n14665_, new_n14664_ );
and  ( new_n14667_, new_n14666_, new_n14627_ );
or   ( new_n14668_, new_n14667_, new_n14663_ );
or   ( new_n14669_, new_n14668_, new_n14661_ );
or   ( new_n14670_, new_n5308_, new_n6307_ );
or   ( new_n14671_, new_n5312_, new_n5459_ );
and  ( new_n14672_, new_n14671_, new_n14670_ );
and  ( new_n14673_, new_n14672_, new_n5182_ );
and  ( new_n14674_, new_n5316_, RI2b1c4342e200_93 );
and  ( new_n14675_, new_n5306_, RI2b1c4342e188_92 );
or   ( new_n14676_, new_n14675_, new_n14674_ );
and  ( new_n14677_, new_n14676_, new_n5028_ );
or   ( new_n14678_, new_n14677_, new_n14673_ );
or   ( new_n14679_, new_n4535_, new_n124_ );
or   ( new_n14680_, new_n4539_, new_n6321_ );
and  ( new_n14681_, new_n14680_, new_n14679_ );
and  ( new_n14682_, new_n14681_, new_n4400_ );
and  ( new_n14683_, new_n4543_, RI2b1c4342e2f0_95 );
and  ( new_n14684_, new_n4533_, RI2b1c4342e278_94 );
or   ( new_n14685_, new_n14684_, new_n14683_ );
and  ( new_n14686_, new_n14685_, new_n4215_ );
or   ( new_n14687_, new_n14686_, new_n14682_ );
and  ( new_n14688_, new_n14687_, new_n14678_ );
or   ( new_n14689_, new_n14687_, new_n14678_ );
or   ( new_n14690_, new_n3806_, new_n7274_ );
and  ( new_n14691_, new_n14690_, new_n3695_ );
and  ( new_n14692_, new_n3800_, RI2b1c4342e368_96 );
and  ( new_n14693_, new_n14692_, new_n3548_ );
or   ( new_n14694_, new_n14693_, new_n14691_ );
and  ( new_n14695_, new_n14694_, new_n14689_ );
or   ( new_n14696_, new_n14695_, new_n14688_ );
or   ( new_n14697_, new_n7105_, new_n132_ );
or   ( new_n14698_, new_n7099_, new_n3902_ );
and  ( new_n14699_, new_n14698_, new_n14697_ );
and  ( new_n14700_, new_n14699_, new_n5858_ );
and  ( new_n14701_, new_n7104_, RI2b1c4342dfa8_88 );
and  ( new_n14702_, new_n7110_, RI2b1c4342e020_89 );
or   ( new_n14703_, new_n14702_, new_n14701_ );
and  ( new_n14704_, new_n14703_, new_n6037_ );
or   ( new_n14705_, new_n14704_, new_n14700_ );
and  ( new_n14706_, new_n14705_, new_n3695_ );
or   ( new_n14707_, new_n14705_, new_n3695_ );
or   ( new_n14708_, new_n6156_, new_n117_ );
or   ( new_n14709_, new_n6160_, new_n4635_ );
and  ( new_n14710_, new_n14709_, new_n14708_ );
and  ( new_n14711_, new_n14710_, new_n6039_ );
and  ( new_n14712_, new_n6164_, RI2b1c4342e110_91 );
and  ( new_n14713_, new_n6154_, RI2b1c4342e098_90 );
or   ( new_n14714_, new_n14713_, new_n14712_ );
and  ( new_n14715_, new_n14714_, new_n5867_ );
or   ( new_n14716_, new_n14715_, new_n14711_ );
and  ( new_n14717_, new_n14716_, new_n14707_ );
or   ( new_n14718_, new_n14717_, new_n14706_ );
and  ( new_n14719_, new_n14718_, new_n14696_ );
or   ( new_n14720_, new_n14718_, new_n14696_ );
or   ( new_n14721_, new_n4535_, new_n6321_ );
or   ( new_n14722_, new_n4539_, new_n6307_ );
and  ( new_n14723_, new_n14722_, new_n14721_ );
and  ( new_n14724_, new_n14723_, new_n4400_ );
and  ( new_n14725_, new_n4543_, RI2b1c4342e278_94 );
and  ( new_n14726_, new_n4533_, RI2b1c4342e200_93 );
or   ( new_n14727_, new_n14726_, new_n14725_ );
and  ( new_n14728_, new_n14727_, new_n4215_ );
or   ( new_n14729_, new_n14728_, new_n14724_ );
and  ( new_n14730_, new_n14729_, new_n14720_ );
or   ( new_n14731_, new_n14730_, new_n14719_ );
and  ( new_n14732_, new_n14731_, new_n14669_ );
or   ( new_n14733_, new_n14731_, new_n14669_ );
or   ( new_n14734_, new_n14466_, new_n14377_ );
and  ( new_n14735_, new_n14734_, new_n14387_ );
and  ( new_n14736_, new_n14376_, new_n2868_ );
and  ( new_n14737_, new_n14464_, new_n3004_ );
or   ( new_n14738_, new_n14737_, new_n14736_ );
and  ( new_n14739_, new_n14738_, new_n14469_ );
or   ( new_n14740_, new_n14739_, new_n14735_ );
and  ( new_n14741_, new_n14740_, new_n14733_ );
or   ( new_n14742_, new_n14741_, new_n14732_ );
or   ( new_n14743_, new_n14742_, new_n14652_ );
and  ( new_n14744_, new_n14743_, new_n14645_ );
and  ( new_n14745_, new_n14742_, new_n14652_ );
and  ( new_n14746_, new_n14650_, new_n14583_ );
and  ( new_n14747_, new_n14646_, new_n14641_ );
or   ( new_n14748_, new_n14747_, new_n14746_ );
and  ( new_n14749_, new_n14659_, new_n3695_ );
and  ( new_n14750_, new_n14655_, new_n3548_ );
or   ( new_n14751_, new_n14750_, new_n14749_ );
and  ( new_n14752_, new_n14666_, new_n14561_ );
and  ( new_n14753_, new_n14662_, new_n14627_ );
or   ( new_n14754_, new_n14753_, new_n14752_ );
and  ( new_n14755_, new_n14754_, new_n14751_ );
and  ( new_n14756_, new_n14676_, new_n5182_ );
and  ( new_n14757_, new_n14672_, new_n5028_ );
or   ( new_n14758_, new_n14757_, new_n14756_ );
and  ( new_n14759_, new_n14685_, new_n4400_ );
and  ( new_n14760_, new_n14681_, new_n4215_ );
or   ( new_n14761_, new_n14760_, new_n14759_ );
and  ( new_n14762_, new_n14761_, new_n14758_ );
or   ( new_n14763_, new_n14761_, new_n14758_ );
and  ( new_n14764_, new_n14692_, new_n3695_ );
and  ( new_n14765_, new_n14690_, new_n3548_ );
or   ( new_n14766_, new_n14765_, new_n14764_ );
and  ( new_n14767_, new_n14766_, new_n14763_ );
or   ( new_n14768_, new_n14767_, new_n14762_ );
and  ( new_n14769_, new_n14703_, new_n5858_ );
and  ( new_n14770_, new_n14699_, new_n6037_ );
or   ( new_n14771_, new_n14770_, new_n14769_ );
or   ( new_n14772_, new_n14771_, new_n3548_ );
and  ( new_n14773_, new_n14771_, new_n3548_ );
and  ( new_n14774_, new_n14714_, new_n6039_ );
and  ( new_n14775_, new_n14710_, new_n5867_ );
or   ( new_n14776_, new_n14775_, new_n14774_ );
or   ( new_n14777_, new_n14776_, new_n14773_ );
and  ( new_n14778_, new_n14777_, new_n14772_ );
or   ( new_n14779_, new_n14778_, new_n14768_ );
and  ( new_n14780_, new_n14778_, new_n14768_ );
and  ( new_n14781_, new_n14727_, new_n4400_ );
and  ( new_n14782_, new_n14723_, new_n4215_ );
or   ( new_n14783_, new_n14782_, new_n14781_ );
or   ( new_n14784_, new_n14783_, new_n14780_ );
and  ( new_n14785_, new_n14784_, new_n14779_ );
or   ( new_n14786_, new_n14785_, new_n14755_ );
and  ( new_n14787_, new_n14785_, new_n14755_ );
and  ( new_n14788_, new_n14738_, new_n14387_ );
and  ( new_n14789_, new_n14734_, new_n14469_ );
or   ( new_n14790_, new_n14789_, new_n14788_ );
or   ( new_n14791_, new_n14790_, new_n14787_ );
and  ( new_n14792_, new_n14791_, new_n14786_ );
and  ( new_n14793_, new_n14792_, new_n14748_ );
or   ( new_n14794_, new_n14793_, new_n14745_ );
or   ( new_n14795_, new_n14630_, new_n14564_ );
and  ( new_n14796_, new_n14795_, new_n14572_ );
and  ( new_n14797_, new_n14629_, new_n14532_ );
and  ( new_n14798_, new_n14616_, new_n14563_ );
or   ( new_n14799_, new_n14798_, new_n14797_ );
and  ( new_n14800_, new_n14799_, new_n14634_ );
or   ( new_n14801_, new_n14800_, new_n14796_ );
or   ( new_n14802_, new_n14787_, new_n14732_ );
and  ( new_n14803_, new_n14802_, new_n14740_ );
and  ( new_n14804_, new_n14785_, new_n14669_ );
and  ( new_n14805_, new_n14755_, new_n14731_ );
or   ( new_n14806_, new_n14805_, new_n14804_ );
and  ( new_n14807_, new_n14806_, new_n14790_ );
or   ( new_n14808_, new_n14807_, new_n14803_ );
or   ( new_n14809_, new_n14808_, new_n14801_ );
and  ( new_n14810_, new_n14809_, new_n14794_ );
or   ( new_n14811_, new_n14810_, new_n14744_ );
and  ( new_n14812_, new_n14668_, new_n14661_ );
or   ( new_n14813_, new_n14812_, new_n14755_ );
or   ( new_n14814_, new_n14762_, new_n14688_ );
and  ( new_n14815_, new_n14814_, new_n14694_ );
and  ( new_n14816_, new_n14758_, new_n14687_ );
and  ( new_n14817_, new_n14761_, new_n14678_ );
or   ( new_n14818_, new_n14817_, new_n14816_ );
and  ( new_n14819_, new_n14818_, new_n14766_ );
or   ( new_n14820_, new_n14819_, new_n14815_ );
or   ( new_n14821_, new_n7105_, new_n4635_ );
or   ( new_n14822_, new_n7099_, new_n132_ );
and  ( new_n14823_, new_n14822_, new_n14821_ );
and  ( new_n14824_, new_n14823_, new_n5858_ );
and  ( new_n14825_, new_n7104_, RI2b1c4342e020_89 );
and  ( new_n14826_, new_n7110_, RI2b1c4342e098_90 );
or   ( new_n14827_, new_n14826_, new_n14825_ );
and  ( new_n14828_, new_n14827_, new_n6037_ );
or   ( new_n14829_, new_n14828_, new_n14824_ );
or   ( new_n14830_, new_n6156_, new_n5459_ );
or   ( new_n14831_, new_n6160_, new_n117_ );
and  ( new_n14832_, new_n14831_, new_n14830_ );
and  ( new_n14833_, new_n14832_, new_n6039_ );
and  ( new_n14834_, new_n6164_, RI2b1c4342e188_92 );
and  ( new_n14835_, new_n6154_, RI2b1c4342e110_91 );
or   ( new_n14836_, new_n14835_, new_n14834_ );
and  ( new_n14837_, new_n14836_, new_n5867_ );
or   ( new_n14838_, new_n14837_, new_n14833_ );
and  ( new_n14839_, new_n14838_, new_n14829_ );
or   ( new_n14840_, new_n14838_, new_n14829_ );
or   ( new_n14841_, new_n5308_, new_n6321_ );
or   ( new_n14842_, new_n5312_, new_n6307_ );
and  ( new_n14843_, new_n14842_, new_n14841_ );
and  ( new_n14844_, new_n14843_, new_n5182_ );
and  ( new_n14845_, new_n5316_, RI2b1c4342e278_94 );
and  ( new_n14846_, new_n5306_, RI2b1c4342e200_93 );
or   ( new_n14847_, new_n14846_, new_n14845_ );
and  ( new_n14848_, new_n14847_, new_n5028_ );
or   ( new_n14849_, new_n14848_, new_n14844_ );
and  ( new_n14850_, new_n14849_, new_n14840_ );
or   ( new_n14851_, new_n14850_, new_n14839_ );
and  ( new_n14852_, new_n14851_, new_n14820_ );
or   ( new_n14853_, new_n14851_, new_n14820_ );
or   ( new_n14854_, new_n14773_, new_n14706_ );
and  ( new_n14855_, new_n14854_, new_n14716_ );
and  ( new_n14856_, new_n14705_, new_n3548_ );
and  ( new_n14857_, new_n14771_, new_n3695_ );
or   ( new_n14858_, new_n14857_, new_n14856_ );
and  ( new_n14859_, new_n14858_, new_n14776_ );
or   ( new_n14860_, new_n14859_, new_n14855_ );
and  ( new_n14861_, new_n14860_, new_n14853_ );
or   ( new_n14862_, new_n14861_, new_n14852_ );
and  ( new_n14863_, new_n14862_, new_n14813_ );
and  ( new_n14864_, new_n14751_, new_n14668_ );
and  ( new_n14865_, new_n14754_, new_n14661_ );
or   ( new_n14866_, new_n14865_, new_n14864_ );
and  ( new_n14867_, new_n14818_, new_n14694_ );
and  ( new_n14868_, new_n14814_, new_n14766_ );
or   ( new_n14869_, new_n14868_, new_n14867_ );
and  ( new_n14870_, new_n14827_, new_n5858_ );
and  ( new_n14871_, new_n14823_, new_n6037_ );
or   ( new_n14872_, new_n14871_, new_n14870_ );
and  ( new_n14873_, new_n14836_, new_n6039_ );
and  ( new_n14874_, new_n14832_, new_n5867_ );
or   ( new_n14875_, new_n14874_, new_n14873_ );
and  ( new_n14876_, new_n14875_, new_n14872_ );
or   ( new_n14877_, new_n14875_, new_n14872_ );
and  ( new_n14878_, new_n14847_, new_n5182_ );
and  ( new_n14879_, new_n14843_, new_n5028_ );
or   ( new_n14880_, new_n14879_, new_n14878_ );
and  ( new_n14881_, new_n14880_, new_n14877_ );
or   ( new_n14882_, new_n14881_, new_n14876_ );
and  ( new_n14883_, new_n14882_, new_n14869_ );
or   ( new_n14884_, new_n14882_, new_n14869_ );
and  ( new_n14885_, new_n14858_, new_n14716_ );
and  ( new_n14886_, new_n14854_, new_n14776_ );
or   ( new_n14887_, new_n14886_, new_n14885_ );
and  ( new_n14888_, new_n14887_, new_n14884_ );
or   ( new_n14889_, new_n14888_, new_n14883_ );
and  ( new_n14890_, new_n14889_, new_n14866_ );
or   ( new_n14891_, new_n14890_, new_n14863_ );
or   ( new_n14892_, new_n14780_, new_n14719_ );
and  ( new_n14893_, new_n14892_, new_n14729_ );
and  ( new_n14894_, new_n14778_, new_n14696_ );
and  ( new_n14895_, new_n14768_, new_n14718_ );
or   ( new_n14896_, new_n14895_, new_n14894_ );
and  ( new_n14897_, new_n14896_, new_n14783_ );
or   ( new_n14898_, new_n14897_, new_n14893_ );
and  ( new_n14899_, new_n14898_, new_n14891_ );
and  ( new_n14900_, new_n14889_, new_n14813_ );
and  ( new_n14901_, new_n14866_, new_n14862_ );
or   ( new_n14902_, new_n14901_, new_n14900_ );
and  ( new_n14903_, new_n14896_, new_n14729_ );
and  ( new_n14904_, new_n14892_, new_n14783_ );
or   ( new_n14905_, new_n14904_, new_n14903_ );
and  ( new_n14906_, new_n14905_, new_n14902_ );
or   ( new_n14907_, new_n14906_, new_n14899_ );
or   ( new_n14908_, new_n14883_, new_n14852_ );
and  ( new_n14909_, new_n14908_, new_n14860_ );
and  ( new_n14910_, new_n14882_, new_n14820_ );
and  ( new_n14911_, new_n14869_, new_n14851_ );
or   ( new_n14912_, new_n14911_, new_n14910_ );
and  ( new_n14913_, new_n14912_, new_n14887_ );
or   ( new_n14914_, new_n14913_, new_n14909_ );
or   ( new_n14915_, new_n5308_, new_n124_ );
or   ( new_n14916_, new_n5312_, new_n6321_ );
and  ( new_n14917_, new_n14916_, new_n14915_ );
and  ( new_n14918_, new_n14917_, new_n5182_ );
and  ( new_n14919_, new_n5316_, RI2b1c4342e2f0_95 );
and  ( new_n14920_, new_n5306_, RI2b1c4342e278_94 );
or   ( new_n14921_, new_n14920_, new_n14919_ );
and  ( new_n14922_, new_n14921_, new_n5028_ );
or   ( new_n14923_, new_n14922_, new_n14918_ );
or   ( new_n14924_, new_n4539_, new_n7274_ );
and  ( new_n14925_, new_n14924_, new_n4400_ );
and  ( new_n14926_, new_n4533_, RI2b1c4342e368_96 );
and  ( new_n14927_, new_n14926_, new_n4215_ );
or   ( new_n14928_, new_n14927_, new_n14925_ );
or   ( new_n14929_, new_n14928_, new_n14923_ );
or   ( new_n14930_, new_n7105_, new_n117_ );
or   ( new_n14931_, new_n7099_, new_n4635_ );
and  ( new_n14932_, new_n14931_, new_n14930_ );
and  ( new_n14933_, new_n14932_, new_n5858_ );
and  ( new_n14934_, new_n7104_, RI2b1c4342e098_90 );
and  ( new_n14935_, new_n7110_, RI2b1c4342e110_91 );
or   ( new_n14936_, new_n14935_, new_n14934_ );
and  ( new_n14937_, new_n14936_, new_n6037_ );
or   ( new_n14938_, new_n14937_, new_n14933_ );
and  ( new_n14939_, new_n14938_, new_n4400_ );
or   ( new_n14940_, new_n14938_, new_n4400_ );
or   ( new_n14941_, new_n6156_, new_n6307_ );
or   ( new_n14942_, new_n6160_, new_n5459_ );
and  ( new_n14943_, new_n14942_, new_n14941_ );
and  ( new_n14944_, new_n14943_, new_n6039_ );
and  ( new_n14945_, new_n6164_, RI2b1c4342e200_93 );
and  ( new_n14946_, new_n6154_, RI2b1c4342e188_92 );
or   ( new_n14947_, new_n14946_, new_n14945_ );
and  ( new_n14948_, new_n14947_, new_n5867_ );
or   ( new_n14949_, new_n14948_, new_n14944_ );
and  ( new_n14950_, new_n14949_, new_n14940_ );
or   ( new_n14951_, new_n14950_, new_n14939_ );
and  ( new_n14952_, new_n14951_, new_n14929_ );
or   ( new_n14953_, new_n14951_, new_n14929_ );
or   ( new_n14954_, new_n4535_, new_n7274_ );
or   ( new_n14955_, new_n4539_, new_n124_ );
and  ( new_n14956_, new_n14955_, new_n14954_ );
and  ( new_n14957_, new_n14956_, new_n4400_ );
and  ( new_n14958_, new_n4543_, RI2b1c4342e368_96 );
and  ( new_n14959_, new_n4533_, RI2b1c4342e2f0_95 );
or   ( new_n14960_, new_n14959_, new_n14958_ );
and  ( new_n14961_, new_n14960_, new_n4215_ );
or   ( new_n14962_, new_n14961_, new_n14957_ );
and  ( new_n14963_, new_n14962_, new_n14953_ );
or   ( new_n14964_, new_n14963_, new_n14952_ );
or   ( new_n14965_, new_n14964_, new_n14914_ );
and  ( new_n14966_, new_n14965_, new_n14907_ );
and  ( new_n14967_, new_n14808_, new_n14801_ );
and  ( new_n14968_, new_n14799_, new_n14572_ );
and  ( new_n14969_, new_n14795_, new_n14634_ );
or   ( new_n14970_, new_n14969_, new_n14968_ );
and  ( new_n14971_, new_n14806_, new_n14740_ );
and  ( new_n14972_, new_n14802_, new_n14790_ );
or   ( new_n14973_, new_n14972_, new_n14971_ );
and  ( new_n14974_, new_n14973_, new_n14970_ );
or   ( new_n14975_, new_n14974_, new_n14967_ );
or   ( new_n14976_, new_n14862_, new_n14813_ );
and  ( new_n14977_, new_n14976_, new_n14898_ );
or   ( new_n14978_, new_n14977_, new_n14863_ );
and  ( new_n14979_, new_n14978_, new_n14975_ );
or   ( new_n14980_, new_n14979_, new_n14966_ );
and  ( new_n14981_, new_n14964_, new_n14914_ );
and  ( new_n14982_, new_n14912_, new_n14860_ );
and  ( new_n14983_, new_n14908_, new_n14887_ );
or   ( new_n14984_, new_n14983_, new_n14982_ );
and  ( new_n14985_, new_n14921_, new_n5182_ );
and  ( new_n14986_, new_n14917_, new_n5028_ );
or   ( new_n14987_, new_n14986_, new_n14985_ );
and  ( new_n14988_, new_n14926_, new_n4400_ );
and  ( new_n14989_, new_n14924_, new_n4215_ );
or   ( new_n14990_, new_n14989_, new_n14988_ );
and  ( new_n14991_, new_n14990_, new_n14987_ );
and  ( new_n14992_, new_n14936_, new_n5858_ );
and  ( new_n14993_, new_n14932_, new_n6037_ );
or   ( new_n14994_, new_n14993_, new_n14992_ );
or   ( new_n14995_, new_n14994_, new_n4215_ );
and  ( new_n14996_, new_n14994_, new_n4215_ );
and  ( new_n14997_, new_n14947_, new_n6039_ );
and  ( new_n14998_, new_n14943_, new_n5867_ );
or   ( new_n14999_, new_n14998_, new_n14997_ );
or   ( new_n15000_, new_n14999_, new_n14996_ );
and  ( new_n15001_, new_n15000_, new_n14995_ );
or   ( new_n15002_, new_n15001_, new_n14991_ );
and  ( new_n15003_, new_n15001_, new_n14991_ );
and  ( new_n15004_, new_n14960_, new_n4400_ );
and  ( new_n15005_, new_n14956_, new_n4215_ );
or   ( new_n15006_, new_n15005_, new_n15004_ );
or   ( new_n15007_, new_n15006_, new_n15003_ );
and  ( new_n15008_, new_n15007_, new_n15002_ );
and  ( new_n15009_, new_n15008_, new_n14984_ );
or   ( new_n15010_, new_n15009_, new_n14981_ );
or   ( new_n15011_, new_n14876_, new_n14839_ );
and  ( new_n15012_, new_n15011_, new_n14849_ );
and  ( new_n15013_, new_n14872_, new_n14838_ );
and  ( new_n15014_, new_n14875_, new_n14829_ );
or   ( new_n15015_, new_n15014_, new_n15013_ );
and  ( new_n15016_, new_n15015_, new_n14880_ );
or   ( new_n15017_, new_n15016_, new_n15012_ );
or   ( new_n15018_, new_n15003_, new_n14952_ );
and  ( new_n15019_, new_n15018_, new_n14962_ );
and  ( new_n15020_, new_n15001_, new_n14929_ );
and  ( new_n15021_, new_n14991_, new_n14951_ );
or   ( new_n15022_, new_n15021_, new_n15020_ );
and  ( new_n15023_, new_n15022_, new_n15006_ );
or   ( new_n15024_, new_n15023_, new_n15019_ );
or   ( new_n15025_, new_n15024_, new_n15017_ );
and  ( new_n15026_, new_n15025_, new_n15010_ );
or   ( new_n15027_, new_n15025_, new_n15010_ );
and  ( new_n15028_, new_n15024_, new_n15017_ );
and  ( new_n15029_, new_n15015_, new_n14849_ );
and  ( new_n15030_, new_n15011_, new_n14880_ );
or   ( new_n15031_, new_n15030_, new_n15029_ );
and  ( new_n15032_, new_n15022_, new_n14962_ );
and  ( new_n15033_, new_n15018_, new_n15006_ );
or   ( new_n15034_, new_n15033_, new_n15032_ );
and  ( new_n15035_, new_n15034_, new_n15031_ );
or   ( new_n15036_, new_n15035_, new_n15028_ );
and  ( new_n15037_, new_n14928_, new_n14923_ );
or   ( new_n15038_, new_n15037_, new_n14991_ );
or   ( new_n15039_, new_n7105_, new_n5459_ );
or   ( new_n15040_, new_n7099_, new_n117_ );
and  ( new_n15041_, new_n15040_, new_n15039_ );
and  ( new_n15042_, new_n15041_, new_n5858_ );
and  ( new_n15043_, new_n7104_, RI2b1c4342e110_91 );
and  ( new_n15044_, new_n7110_, RI2b1c4342e188_92 );
or   ( new_n15045_, new_n15044_, new_n15043_ );
and  ( new_n15046_, new_n15045_, new_n6037_ );
or   ( new_n15047_, new_n15046_, new_n15042_ );
or   ( new_n15048_, new_n6156_, new_n6321_ );
or   ( new_n15049_, new_n6160_, new_n6307_ );
and  ( new_n15050_, new_n15049_, new_n15048_ );
and  ( new_n15051_, new_n15050_, new_n6039_ );
and  ( new_n15052_, new_n6164_, RI2b1c4342e278_94 );
and  ( new_n15053_, new_n6154_, RI2b1c4342e200_93 );
or   ( new_n15054_, new_n15053_, new_n15052_ );
and  ( new_n15055_, new_n15054_, new_n5867_ );
or   ( new_n15056_, new_n15055_, new_n15051_ );
and  ( new_n15057_, new_n15056_, new_n15047_ );
or   ( new_n15058_, new_n15056_, new_n15047_ );
or   ( new_n15059_, new_n5308_, new_n7274_ );
or   ( new_n15060_, new_n5312_, new_n124_ );
and  ( new_n15061_, new_n15060_, new_n15059_ );
and  ( new_n15062_, new_n15061_, new_n5182_ );
and  ( new_n15063_, new_n5316_, RI2b1c4342e368_96 );
and  ( new_n15064_, new_n5306_, RI2b1c4342e2f0_95 );
or   ( new_n15065_, new_n15064_, new_n15063_ );
and  ( new_n15066_, new_n15065_, new_n5028_ );
or   ( new_n15067_, new_n15066_, new_n15062_ );
and  ( new_n15068_, new_n15067_, new_n15058_ );
or   ( new_n15069_, new_n15068_, new_n15057_ );
and  ( new_n15070_, new_n15069_, new_n15038_ );
or   ( new_n15071_, new_n15069_, new_n15038_ );
or   ( new_n15072_, new_n14996_, new_n14939_ );
and  ( new_n15073_, new_n15072_, new_n14949_ );
and  ( new_n15074_, new_n14938_, new_n4215_ );
and  ( new_n15075_, new_n14994_, new_n4400_ );
or   ( new_n15076_, new_n15075_, new_n15074_ );
and  ( new_n15077_, new_n15076_, new_n14999_ );
or   ( new_n15078_, new_n15077_, new_n15073_ );
and  ( new_n15079_, new_n15078_, new_n15071_ );
or   ( new_n15080_, new_n15079_, new_n15070_ );
or   ( new_n15081_, new_n15080_, new_n15036_ );
and  ( new_n15082_, new_n15081_, new_n15027_ );
or   ( new_n15083_, new_n15082_, new_n15026_ );
and  ( new_n15084_, new_n15080_, new_n15036_ );
or   ( new_n15085_, new_n15084_, new_n15026_ );
and  ( new_n15086_, new_n14987_, new_n14928_ );
and  ( new_n15087_, new_n14990_, new_n14923_ );
or   ( new_n15088_, new_n15087_, new_n15086_ );
and  ( new_n15089_, new_n15045_, new_n5858_ );
and  ( new_n15090_, new_n15041_, new_n6037_ );
or   ( new_n15091_, new_n15090_, new_n15089_ );
and  ( new_n15092_, new_n15054_, new_n6039_ );
and  ( new_n15093_, new_n15050_, new_n5867_ );
or   ( new_n15094_, new_n15093_, new_n15092_ );
and  ( new_n15095_, new_n15094_, new_n15091_ );
or   ( new_n15096_, new_n15094_, new_n15091_ );
and  ( new_n15097_, new_n15065_, new_n5182_ );
and  ( new_n15098_, new_n15061_, new_n5028_ );
or   ( new_n15099_, new_n15098_, new_n15097_ );
and  ( new_n15100_, new_n15099_, new_n15096_ );
or   ( new_n15101_, new_n15100_, new_n15095_ );
and  ( new_n15102_, new_n15101_, new_n15088_ );
or   ( new_n15103_, new_n15102_, new_n15070_ );
and  ( new_n15104_, new_n15103_, new_n15078_ );
and  ( new_n15105_, new_n15101_, new_n15038_ );
and  ( new_n15106_, new_n15088_, new_n15069_ );
or   ( new_n15107_, new_n15106_, new_n15105_ );
and  ( new_n15108_, new_n15076_, new_n14949_ );
and  ( new_n15109_, new_n15072_, new_n14999_ );
or   ( new_n15110_, new_n15109_, new_n15108_ );
and  ( new_n15111_, new_n15110_, new_n15107_ );
or   ( new_n15112_, new_n15111_, new_n15104_ );
or   ( new_n15113_, new_n15095_, new_n15057_ );
and  ( new_n15114_, new_n15113_, new_n15067_ );
and  ( new_n15115_, new_n15091_, new_n15056_ );
and  ( new_n15116_, new_n15094_, new_n15047_ );
or   ( new_n15117_, new_n15116_, new_n15115_ );
and  ( new_n15118_, new_n15117_, new_n15099_ );
or   ( new_n15119_, new_n15118_, new_n15114_ );
or   ( new_n15120_, new_n7105_, new_n6307_ );
or   ( new_n15121_, new_n7099_, new_n5459_ );
and  ( new_n15122_, new_n15121_, new_n15120_ );
and  ( new_n15123_, new_n15122_, new_n5858_ );
and  ( new_n15124_, new_n7104_, RI2b1c4342e188_92 );
and  ( new_n15125_, new_n7110_, RI2b1c4342e200_93 );
or   ( new_n15126_, new_n15125_, new_n15124_ );
and  ( new_n15127_, new_n15126_, new_n6037_ );
or   ( new_n15128_, new_n15127_, new_n15123_ );
and  ( new_n15129_, new_n15128_, new_n5182_ );
or   ( new_n15130_, new_n15128_, new_n5182_ );
or   ( new_n15131_, new_n6156_, new_n124_ );
or   ( new_n15132_, new_n6160_, new_n6321_ );
and  ( new_n15133_, new_n15132_, new_n15131_ );
and  ( new_n15134_, new_n15133_, new_n6039_ );
and  ( new_n15135_, new_n6164_, RI2b1c4342e2f0_95 );
and  ( new_n15136_, new_n6154_, RI2b1c4342e278_94 );
or   ( new_n15137_, new_n15136_, new_n15135_ );
and  ( new_n15138_, new_n15137_, new_n5867_ );
or   ( new_n15139_, new_n15138_, new_n15134_ );
and  ( new_n15140_, new_n15139_, new_n15130_ );
or   ( new_n15141_, new_n15140_, new_n15129_ );
or   ( new_n15142_, new_n15141_, new_n15119_ );
and  ( new_n15143_, new_n15142_, new_n15112_ );
or   ( new_n15144_, new_n15142_, new_n15112_ );
and  ( new_n15145_, new_n15141_, new_n15119_ );
and  ( new_n15146_, new_n15117_, new_n15067_ );
and  ( new_n15147_, new_n15113_, new_n15099_ );
or   ( new_n15148_, new_n15147_, new_n15146_ );
and  ( new_n15149_, new_n15126_, new_n5858_ );
and  ( new_n15150_, new_n15122_, new_n6037_ );
or   ( new_n15151_, new_n15150_, new_n15149_ );
and  ( new_n15152_, new_n15151_, new_n5028_ );
or   ( new_n15153_, new_n15151_, new_n5028_ );
and  ( new_n15154_, new_n15137_, new_n6039_ );
and  ( new_n15155_, new_n15133_, new_n5867_ );
or   ( new_n15156_, new_n15155_, new_n15154_ );
and  ( new_n15157_, new_n15156_, new_n15153_ );
or   ( new_n15158_, new_n15157_, new_n15152_ );
and  ( new_n15159_, new_n15158_, new_n15148_ );
or   ( new_n15160_, new_n15159_, new_n15145_ );
or   ( new_n15161_, new_n5312_, new_n7274_ );
and  ( new_n15162_, new_n15161_, new_n5182_ );
and  ( new_n15163_, new_n5306_, RI2b1c4342e368_96 );
and  ( new_n15164_, new_n15163_, new_n5028_ );
or   ( new_n15165_, new_n15164_, new_n15162_ );
or   ( new_n15166_, new_n15152_, new_n15129_ );
and  ( new_n15167_, new_n15166_, new_n15139_ );
and  ( new_n15168_, new_n15128_, new_n5028_ );
and  ( new_n15169_, new_n15151_, new_n5182_ );
or   ( new_n15170_, new_n15169_, new_n15168_ );
and  ( new_n15171_, new_n15170_, new_n15156_ );
or   ( new_n15172_, new_n15171_, new_n15167_ );
or   ( new_n15173_, new_n15172_, new_n15165_ );
or   ( new_n15174_, new_n15173_, new_n15160_ );
and  ( new_n15175_, new_n15174_, new_n15144_ );
or   ( new_n15176_, new_n15175_, new_n15143_ );
and  ( new_n15177_, new_n15173_, new_n15160_ );
and  ( new_n15178_, new_n15172_, new_n15165_ );
and  ( new_n15179_, new_n15163_, new_n5182_ );
and  ( new_n15180_, new_n15161_, new_n5028_ );
or   ( new_n15181_, new_n15180_, new_n15179_ );
and  ( new_n15182_, new_n15170_, new_n15139_ );
and  ( new_n15183_, new_n15166_, new_n15156_ );
or   ( new_n15184_, new_n15183_, new_n15182_ );
and  ( new_n15185_, new_n15184_, new_n15181_ );
or   ( new_n15186_, new_n15185_, new_n15178_ );
or   ( new_n15187_, new_n7105_, new_n6321_ );
or   ( new_n15188_, new_n7099_, new_n6307_ );
and  ( new_n15189_, new_n15188_, new_n15187_ );
and  ( new_n15190_, new_n15189_, new_n5858_ );
and  ( new_n15191_, new_n7104_, RI2b1c4342e200_93 );
and  ( new_n15192_, new_n7110_, RI2b1c4342e278_94 );
or   ( new_n15193_, new_n15192_, new_n15191_ );
and  ( new_n15194_, new_n15193_, new_n6037_ );
or   ( new_n15195_, new_n15194_, new_n15190_ );
or   ( new_n15196_, new_n6156_, new_n7274_ );
or   ( new_n15197_, new_n6160_, new_n124_ );
and  ( new_n15198_, new_n15197_, new_n15196_ );
and  ( new_n15199_, new_n15198_, new_n6039_ );
and  ( new_n15200_, new_n6164_, RI2b1c4342e368_96 );
and  ( new_n15201_, new_n6154_, RI2b1c4342e2f0_95 );
or   ( new_n15202_, new_n15201_, new_n15200_ );
and  ( new_n15203_, new_n15202_, new_n5867_ );
or   ( new_n15204_, new_n15203_, new_n15199_ );
or   ( new_n15205_, new_n15204_, new_n15195_ );
and  ( new_n15206_, new_n15205_, new_n15186_ );
or   ( new_n15207_, new_n15206_, new_n15177_ );
or   ( new_n15208_, new_n15205_, new_n15186_ );
and  ( new_n15209_, new_n15204_, new_n15195_ );
and  ( new_n15210_, new_n15193_, new_n5858_ );
and  ( new_n15211_, new_n15189_, new_n6037_ );
or   ( new_n15212_, new_n15211_, new_n15210_ );
and  ( new_n15213_, new_n15202_, new_n6039_ );
and  ( new_n15214_, new_n15198_, new_n5867_ );
or   ( new_n15215_, new_n15214_, new_n15213_ );
and  ( new_n15216_, new_n15215_, new_n15212_ );
or   ( new_n15217_, new_n15216_, new_n15209_ );
or   ( new_n15218_, new_n7105_, new_n124_ );
or   ( new_n15219_, new_n7099_, new_n6321_ );
and  ( new_n15220_, new_n15219_, new_n15218_ );
and  ( new_n15221_, new_n15220_, new_n5858_ );
and  ( new_n15222_, new_n7104_, RI2b1c4342e278_94 );
and  ( new_n15223_, new_n7110_, RI2b1c4342e2f0_95 );
or   ( new_n15224_, new_n15223_, new_n15222_ );
and  ( new_n15225_, new_n15224_, new_n6037_ );
or   ( new_n15226_, new_n15225_, new_n15221_ );
or   ( new_n15227_, new_n15226_, new_n6039_ );
and  ( new_n15228_, new_n15227_, new_n15217_ );
and  ( new_n15229_, new_n15226_, new_n6039_ );
and  ( new_n15230_, new_n15224_, new_n5858_ );
and  ( new_n15231_, new_n15220_, new_n6037_ );
or   ( new_n15232_, new_n15231_, new_n15230_ );
and  ( new_n15233_, new_n15232_, new_n5867_ );
or   ( new_n15234_, new_n15233_, new_n15229_ );
or   ( new_n15235_, new_n6160_, new_n7274_ );
and  ( new_n15236_, new_n15235_, new_n6039_ );
and  ( new_n15237_, new_n6154_, RI2b1c4342e368_96 );
and  ( new_n15238_, new_n15237_, new_n5867_ );
or   ( new_n15239_, new_n15238_, new_n15236_ );
or   ( new_n15240_, new_n15239_, new_n15234_ );
or   ( new_n15241_, new_n15227_, new_n15217_ );
and  ( new_n15242_, new_n15241_, new_n15240_ );
or   ( new_n15243_, new_n15242_, new_n15228_ );
and  ( new_n15244_, new_n15239_, new_n15234_ );
and  ( new_n15245_, new_n7274_, new_n124_ );
not  ( new_n15246_, new_n7104_ );
nor  ( new_n15247_, new_n15246_, new_n15245_ );
and  ( new_n15248_, new_n7110_, RI2b1c4342e368_96 );
or   ( new_n15249_, new_n15248_, new_n15247_ );
and  ( new_n15250_, new_n15249_, new_n6037_ );
or   ( new_n15251_, new_n15250_, new_n5858_ );
or   ( new_n15252_, new_n15251_, new_n15244_ );
or   ( new_n15253_, new_n15252_, new_n15228_ );
and  ( new_n15254_, new_n15253_, new_n15243_ );
and  ( new_n15255_, new_n15254_, new_n15208_ );
or   ( new_n15256_, new_n15255_, new_n15207_ );
or   ( new_n15257_, new_n15256_, new_n15143_ );
and  ( new_n15258_, new_n15257_, new_n15176_ );
or   ( new_n15259_, new_n15258_, new_n15085_ );
and  ( new_n15260_, new_n15259_, new_n15083_ );
or   ( new_n15261_, new_n15260_, new_n14980_ );
or   ( new_n15262_, new_n15261_, new_n14811_ );
or   ( new_n15263_, new_n14743_, new_n14645_ );
or   ( new_n15264_, new_n14809_, new_n14794_ );
and  ( new_n15265_, new_n15264_, new_n15263_ );
or   ( new_n15266_, new_n15265_, new_n14744_ );
or   ( new_n15267_, new_n14978_, new_n14975_ );
or   ( new_n15268_, new_n14965_, new_n14907_ );
and  ( new_n15269_, new_n15268_, new_n15267_ );
or   ( new_n15270_, new_n15269_, new_n14979_ );
or   ( new_n15271_, new_n15270_, new_n14811_ );
and  ( new_n15272_, new_n15271_, new_n15266_ );
and  ( new_n15273_, new_n15272_, new_n15262_ );
or   ( new_n15274_, new_n15273_, new_n14606_ );
or   ( new_n15275_, new_n15274_, new_n14310_ );
or   ( new_n15276_, new_n14118_, new_n14021_ );
or   ( new_n15277_, new_n14308_, new_n14173_ );
and  ( new_n15278_, new_n15277_, new_n15276_ );
or   ( new_n15279_, new_n15278_, new_n14119_ );
or   ( new_n15280_, new_n14604_, new_n14601_ );
or   ( new_n15281_, new_n14586_, new_n14513_ );
and  ( new_n15282_, new_n15281_, new_n15280_ );
or   ( new_n15283_, new_n15282_, new_n14605_ );
or   ( new_n15284_, new_n15283_, new_n14310_ );
and  ( new_n15285_, new_n15284_, new_n15279_ );
and  ( new_n15286_, new_n15285_, new_n15275_ );
or   ( new_n15287_, new_n15286_, new_n13960_ );
or   ( new_n15288_, new_n15287_, new_n13741_ );
or   ( new_n15289_, new_n13508_, new_n13358_ );
or   ( new_n15290_, new_n13739_, new_n13590_ );
and  ( new_n15291_, new_n15290_, new_n15289_ );
or   ( new_n15292_, new_n15291_, new_n13509_ );
or   ( new_n15293_, new_n13958_, new_n13957_ );
or   ( new_n15294_, new_n13947_, new_n13835_ );
and  ( new_n15295_, new_n15294_, new_n15293_ );
or   ( new_n15296_, new_n15295_, new_n13959_ );
or   ( new_n15297_, new_n15296_, new_n13741_ );
and  ( new_n15298_, new_n15297_, new_n15292_ );
and  ( new_n15299_, new_n15298_, new_n15288_ );
or   ( new_n15300_, new_n15299_, new_n13260_ );
or   ( new_n15301_, new_n15300_, new_n12733_ );
or   ( new_n15302_, new_n12465_, new_n12296_ );
or   ( new_n15303_, new_n12731_, new_n12553_ );
and  ( new_n15304_, new_n15303_, new_n15302_ );
or   ( new_n15305_, new_n15304_, new_n12466_ );
or   ( new_n15306_, new_n12984_, new_n12825_ );
or   ( new_n15307_, new_n13258_, new_n13072_ );
and  ( new_n15308_, new_n15307_, new_n15306_ );
or   ( new_n15309_, new_n15308_, new_n12985_ );
or   ( new_n15310_, new_n15309_, new_n12733_ );
and  ( new_n15311_, new_n15310_, new_n15305_ );
and  ( new_n15312_, new_n15311_, new_n15301_ );
or   ( new_n15313_, new_n15312_, new_n12182_ );
and  ( new_n15314_, new_n15313_, new_n12179_ );
or   ( new_n15315_, new_n15314_, new_n11175_ );
or   ( new_n15316_, new_n15315_, new_n9592_ );
and  ( new_n15317_, new_n15316_, new_n11172_ );
and  ( new_n15318_, new_n7853_, new_n7569_ );
or   ( new_n15319_, new_n15318_, new_n7406_ );
or   ( new_n15320_, new_n15319_, new_n6907_ );
or   ( new_n15321_, new_n15320_, new_n5994_ );
or   ( new_n15322_, new_n15321_, new_n15317_ );
and  ( new_n15323_, new_n15322_, new_n7860_ );
or   ( new_n15324_, new_n15323_, new_n4382_ );
and  ( new_n15325_, new_n15324_, new_n4378_ );
or   ( new_n15326_, new_n841_, new_n843_ );
or   ( new_n15327_, new_n857_, new_n859_ );
or   ( new_n15328_, new_n861_, new_n105_ );
and  ( new_n15329_, new_n15328_, new_n15327_ );
and  ( new_n15330_, new_n15329_, new_n842_ );
and  ( new_n15331_, new_n870_, RI2b1c4342d918_74 );
and  ( new_n15332_, new_n855_, RI2b1c4342d8a0_73 );
or   ( new_n15333_, new_n15332_, new_n15331_ );
and  ( new_n15334_, new_n15333_, new_n866_ );
or   ( new_n15335_, new_n15334_, new_n15330_ );
or   ( new_n15336_, new_n753_, new_n755_ );
or   ( new_n15337_, new_n757_, new_n591_ );
and  ( new_n15338_, new_n15337_, new_n15336_ );
and  ( new_n15339_, new_n15338_, new_n734_ );
and  ( new_n15340_, new_n766_, RI2b1c4342d738_70 );
and  ( new_n15341_, new_n751_, RI2b1c4342d6c0_69 );
or   ( new_n15342_, new_n15341_, new_n15340_ );
and  ( new_n15343_, new_n15342_, new_n762_ );
or   ( new_n15344_, new_n15343_, new_n15339_ );
or   ( new_n15345_, new_n804_, new_n806_ );
or   ( new_n15346_, new_n808_, new_n110_ );
and  ( new_n15347_, new_n15346_, new_n15345_ );
and  ( new_n15348_, new_n15347_, new_n785_ );
and  ( new_n15349_, new_n817_, RI2b1c4342d828_72 );
and  ( new_n15350_, new_n802_, RI2b1c4342d7b0_71 );
or   ( new_n15351_, new_n15350_, new_n15349_ );
and  ( new_n15352_, new_n15351_, new_n813_ );
or   ( new_n15353_, new_n15352_, new_n15348_ );
and  ( new_n15354_, new_n15353_, new_n15344_ );
and  ( new_n15355_, new_n15342_, new_n734_ );
and  ( new_n15356_, new_n15338_, new_n762_ );
or   ( new_n15357_, new_n15356_, new_n15355_ );
and  ( new_n15358_, new_n15351_, new_n785_ );
and  ( new_n15359_, new_n15347_, new_n813_ );
or   ( new_n15360_, new_n15359_, new_n15358_ );
and  ( new_n15361_, new_n15360_, new_n15357_ );
or   ( new_n15362_, new_n15361_, new_n15354_ );
and  ( new_n15363_, new_n15362_, new_n15335_ );
and  ( new_n15364_, new_n15333_, new_n842_ );
and  ( new_n15365_, new_n15329_, new_n866_ );
or   ( new_n15366_, new_n15365_, new_n15364_ );
and  ( new_n15367_, new_n15357_, new_n15353_ );
and  ( new_n15368_, new_n15360_, new_n15344_ );
or   ( new_n15369_, new_n15368_, new_n15367_ );
and  ( new_n15370_, new_n15369_, new_n15366_ );
or   ( new_n15371_, new_n15370_, new_n15363_ );
and  ( new_n15372_, new_n15371_, new_n15326_ );
and  ( new_n15373_, new_n720_, RI2b1c4342d990_75 );
and  ( new_n15374_, new_n15369_, new_n15335_ );
and  ( new_n15375_, new_n15366_, new_n15362_ );
or   ( new_n15376_, new_n15375_, new_n15374_ );
and  ( new_n15377_, new_n15376_, new_n15373_ );
or   ( new_n15378_, new_n15377_, new_n15372_ );
or   ( new_n15379_, new_n610_, new_n612_ );
or   ( new_n15380_, new_n614_, new_n112_ );
and  ( new_n15381_, new_n15380_, new_n15379_ );
and  ( new_n15382_, new_n15381_, new_n590_ );
and  ( new_n15383_, new_n623_, RI2b1c4342d648_68 );
and  ( new_n15384_, new_n608_, RI2b1c4342d5d0_67 );
or   ( new_n15385_, new_n15384_, new_n15383_ );
and  ( new_n15386_, new_n15385_, new_n619_ );
or   ( new_n15387_, new_n15386_, new_n15382_ );
and  ( new_n15388_, new_n537_, RI2b1c4342d558_66 );
and  ( new_n15389_, new_n522_, RI2b1c4342d4e0_65 );
or   ( new_n15390_, new_n15389_, new_n15388_ );
and  ( new_n15391_, new_n15390_, new_n505_ );
or   ( new_n15392_, new_n524_, new_n526_ );
or   ( new_n15393_, new_n528_, new_n99_ );
and  ( new_n15394_, new_n15393_, new_n15392_ );
and  ( new_n15395_, new_n15394_, new_n533_ );
or   ( new_n15396_, new_n15395_, new_n15391_ );
and  ( new_n15397_, new_n15396_, new_n428_ );
and  ( new_n15398_, new_n15394_, new_n505_ );
and  ( new_n15399_, new_n15390_, new_n533_ );
or   ( new_n15400_, new_n15399_, new_n15398_ );
and  ( new_n15401_, new_n15400_, new_n457_ );
or   ( new_n15402_, new_n15401_, new_n15397_ );
and  ( new_n15403_, new_n15402_, new_n15387_ );
and  ( new_n15404_, new_n15385_, new_n590_ );
and  ( new_n15405_, new_n15381_, new_n619_ );
or   ( new_n15406_, new_n15405_, new_n15404_ );
and  ( new_n15407_, new_n15400_, new_n428_ );
and  ( new_n15408_, new_n15396_, new_n457_ );
or   ( new_n15409_, new_n15408_, new_n15407_ );
and  ( new_n15410_, new_n15409_, new_n15406_ );
or   ( new_n15411_, new_n15410_, new_n15403_ );
and  ( new_n15412_, new_n15411_, new_n15378_ );
and  ( new_n15413_, new_n15373_, new_n15371_ );
and  ( new_n15414_, new_n15376_, new_n15326_ );
or   ( new_n15415_, new_n15414_, new_n15413_ );
and  ( new_n15416_, new_n15409_, new_n15387_ );
and  ( new_n15417_, new_n15406_, new_n15402_ );
or   ( new_n15418_, new_n15417_, new_n15416_ );
and  ( new_n15419_, new_n15418_, new_n15415_ );
or   ( new_n15420_, new_n15419_, new_n15412_ );
or   ( new_n15421_, new_n1183_, new_n1180_ );
and  ( new_n15422_, new_n15421_, new_n1177_ );
or   ( new_n15423_, new_n15422_, new_n1184_ );
or   ( new_n15424_, new_n884_, new_n721_ );
and  ( new_n15425_, new_n15424_, new_n637_ );
or   ( new_n15426_, new_n15425_, new_n885_ );
and  ( new_n15427_, new_n15426_, new_n15423_ );
or   ( new_n15428_, new_n890_, new_n887_ );
and  ( new_n15429_, new_n15428_, new_n896_ );
or   ( new_n15430_, new_n15429_, new_n891_ );
or   ( new_n15431_, new_n1190_, new_n1187_ );
or   ( new_n15432_, new_n1191_, new_n1028_ );
and  ( new_n15433_, new_n15432_, new_n15431_ );
and  ( new_n15434_, new_n15433_, new_n15430_ );
or   ( new_n15435_, new_n15434_, new_n15427_ );
and  ( new_n15436_, new_n15435_, new_n15420_ );
and  ( new_n15437_, new_n15415_, new_n15411_ );
and  ( new_n15438_, new_n15418_, new_n15378_ );
or   ( new_n15439_, new_n15438_, new_n15437_ );
and  ( new_n15440_, new_n15433_, new_n15426_ );
and  ( new_n15441_, new_n15430_, new_n15423_ );
or   ( new_n15442_, new_n15441_, new_n15440_ );
and  ( new_n15443_, new_n15442_, new_n15439_ );
or   ( new_n15444_, new_n15443_, new_n15436_ );
or   ( new_n15445_, new_n542_, new_n466_ );
and  ( new_n15446_, new_n15445_, new_n628_ );
or   ( new_n15447_, new_n15446_, new_n543_ );
or   ( new_n15448_, new_n822_, new_n771_ );
and  ( new_n15449_, new_n15448_, new_n875_ );
or   ( new_n15450_, new_n15449_, new_n823_ );
and  ( new_n15451_, new_n15450_, new_n15447_ );
or   ( new_n15452_, new_n549_, new_n546_ );
and  ( new_n15453_, new_n15452_, new_n635_ );
or   ( new_n15454_, new_n15453_, new_n550_ );
or   ( new_n15455_, new_n829_, new_n826_ );
and  ( new_n15456_, new_n15455_, new_n882_ );
or   ( new_n15457_, new_n15456_, new_n830_ );
and  ( new_n15458_, new_n15457_, new_n15454_ );
or   ( new_n15459_, new_n15458_, new_n15451_ );
and  ( new_n15460_, new_n15459_, new_n887_ );
and  ( new_n15461_, new_n15454_, new_n15450_ );
and  ( new_n15462_, new_n15457_, new_n15447_ );
or   ( new_n15463_, new_n15462_, new_n15461_ );
and  ( new_n15464_, new_n15463_, new_n721_ );
or   ( new_n15465_, new_n15464_, new_n15460_ );
or   ( new_n15466_, new_n1165_, new_n1152_ );
and  ( new_n15467_, new_n15466_, new_n1171_ );
or   ( new_n15468_, new_n15467_, new_n1166_ );
and  ( new_n15469_, new_n15468_, new_n15465_ );
or   ( new_n15470_, new_n1116_, new_n1017_ );
and  ( new_n15471_, new_n15470_, new_n901_ );
or   ( new_n15472_, new_n15471_, new_n1117_ );
and  ( new_n15473_, new_n15463_, new_n887_ );
and  ( new_n15474_, new_n15459_, new_n721_ );
or   ( new_n15475_, new_n15474_, new_n15473_ );
and  ( new_n15476_, new_n15475_, new_n15472_ );
or   ( new_n15477_, new_n15476_, new_n15469_ );
and  ( new_n15478_, new_n15477_, new_n15444_ );
and  ( new_n15479_, new_n15442_, new_n15420_ );
and  ( new_n15480_, new_n15439_, new_n15435_ );
or   ( new_n15481_, new_n15480_, new_n15479_ );
and  ( new_n15482_, new_n15472_, new_n15465_ );
and  ( new_n15483_, new_n15475_, new_n15468_ );
or   ( new_n15484_, new_n15483_, new_n15482_ );
and  ( new_n15485_, new_n15484_, new_n15481_ );
or   ( new_n15486_, new_n15485_, new_n15478_ );
or   ( new_n15487_, new_n1400_, new_n1332_ );
or   ( new_n15488_, new_n1406_, new_n1401_ );
and  ( new_n15489_, new_n15488_, new_n15487_ );
and  ( new_n15490_, new_n15489_, new_n15486_ );
and  ( new_n15491_, new_n15484_, new_n15444_ );
and  ( new_n15492_, new_n15481_, new_n15477_ );
or   ( new_n15493_, new_n15492_, new_n15491_ );
or   ( new_n15494_, new_n1328_, new_n1198_ );
and  ( new_n15495_, new_n15494_, new_n1176_ );
or   ( new_n15496_, new_n15495_, new_n1329_ );
and  ( new_n15497_, new_n15496_, new_n15493_ );
or   ( new_n15498_, new_n15497_, new_n15490_ );
or   ( new_n15499_, new_n1564_, new_n1411_ );
or   ( new_n15500_, new_n15499_, new_n15498_ );
and  ( new_n15501_, new_n15493_, new_n15489_ );
and  ( new_n15502_, new_n15496_, new_n15486_ );
or   ( new_n15503_, new_n15502_, new_n15501_ );
or   ( new_n15504_, new_n15503_, new_n1640_ );
and  ( new_n15505_, new_n15504_, new_n15500_ );
and  ( new_n15506_, new_n15505_, new_n15325_ );
and  ( new_n15507_, new_n15499_, new_n15498_ );
and  ( new_n15508_, new_n15503_, new_n1640_ );
or   ( new_n15509_, new_n15508_, new_n15507_ );
and  ( new_n15510_, new_n1639_, new_n1411_ );
and  ( new_n15511_, new_n1568_, new_n1564_ );
or   ( new_n15512_, new_n15511_, new_n15510_ );
and  ( new_n15513_, new_n15512_, new_n1879_ );
or   ( new_n15514_, new_n15512_, new_n1879_ );
and  ( new_n15515_, new_n1878_, new_n1648_ );
and  ( new_n15516_, new_n1802_, new_n1796_ );
or   ( new_n15517_, new_n15516_, new_n15515_ );
or   ( new_n15518_, new_n2414_, new_n2411_ );
and  ( new_n15519_, new_n15518_, new_n2420_ );
or   ( new_n15520_, new_n15519_, new_n2415_ );
and  ( new_n15521_, new_n15520_, new_n15517_ );
and  ( new_n15522_, new_n15521_, new_n15514_ );
or   ( new_n15523_, new_n15522_, new_n15513_ );
or   ( new_n15524_, new_n15520_, new_n15517_ );
and  ( new_n15525_, new_n15524_, new_n15514_ );
and  ( new_n15526_, new_n2423_, new_n2301_ );
and  ( new_n15527_, new_n2420_, new_n2416_ );
or   ( new_n15528_, new_n15527_, new_n15526_ );
and  ( new_n15529_, new_n15528_, new_n2743_ );
or   ( new_n15530_, new_n15528_, new_n2743_ );
and  ( new_n15531_, new_n2742_, new_n2432_ );
and  ( new_n15532_, new_n2640_, new_n2633_ );
or   ( new_n15533_, new_n15532_, new_n15531_ );
and  ( new_n15534_, new_n15533_, new_n3090_ );
and  ( new_n15535_, new_n15534_, new_n15530_ );
or   ( new_n15536_, new_n15535_, new_n15529_ );
and  ( new_n15537_, new_n15536_, new_n15525_ );
or   ( new_n15538_, new_n15537_, new_n15523_ );
and  ( new_n15539_, new_n3089_, new_n2751_ );
and  ( new_n15540_, new_n2976_, new_n2966_ );
or   ( new_n15541_, new_n15540_, new_n15539_ );
and  ( new_n15542_, new_n15541_, new_n3427_ );
or   ( new_n15543_, new_n15541_, new_n3427_ );
and  ( new_n15544_, new_n3426_, new_n3098_ );
and  ( new_n15545_, new_n3321_, new_n3314_ );
or   ( new_n15546_, new_n15545_, new_n15544_ );
and  ( new_n15547_, new_n15546_, new_n3780_ );
and  ( new_n15548_, new_n15547_, new_n15543_ );
or   ( new_n15549_, new_n15548_, new_n15542_ );
and  ( new_n15550_, new_n3779_, new_n3435_ );
and  ( new_n15551_, new_n3664_, new_n3656_ );
or   ( new_n15552_, new_n15551_, new_n15550_ );
and  ( new_n15553_, new_n15552_, new_n4128_ );
or   ( new_n15554_, new_n15552_, new_n4128_ );
and  ( new_n15555_, new_n4127_, new_n3788_ );
and  ( new_n15556_, new_n4019_, new_n4012_ );
or   ( new_n15557_, new_n15556_, new_n15555_ );
and  ( new_n15558_, new_n15557_, new_n4505_ );
and  ( new_n15559_, new_n15558_, new_n15554_ );
or   ( new_n15560_, new_n15559_, new_n15553_ );
or   ( new_n15561_, new_n15546_, new_n3780_ );
and  ( new_n15562_, new_n15561_, new_n15543_ );
and  ( new_n15563_, new_n15562_, new_n15560_ );
or   ( new_n15564_, new_n15563_, new_n15549_ );
or   ( new_n15565_, new_n15533_, new_n3090_ );
and  ( new_n15566_, new_n15565_, new_n15530_ );
and  ( new_n15567_, new_n15566_, new_n15525_ );
and  ( new_n15568_, new_n15567_, new_n15564_ );
or   ( new_n15569_, new_n15568_, new_n15538_ );
or   ( new_n15570_, new_n15557_, new_n4505_ );
and  ( new_n15571_, new_n15570_, new_n15554_ );
and  ( new_n15572_, new_n15571_, new_n15562_ );
and  ( new_n15573_, new_n15572_, new_n15567_ );
and  ( new_n15574_, new_n4504_, new_n4136_ );
and  ( new_n15575_, new_n4386_, new_n4365_ );
or   ( new_n15576_, new_n15575_, new_n15574_ );
and  ( new_n15577_, new_n15576_, new_n4885_ );
or   ( new_n15578_, new_n15576_, new_n4885_ );
and  ( new_n15579_, new_n4884_, new_n4513_ );
and  ( new_n15580_, new_n4767_, new_n4760_ );
or   ( new_n15581_, new_n15580_, new_n15579_ );
or   ( new_n15582_, new_n5283_, new_n5155_ );
or   ( new_n15583_, new_n5292_, new_n5284_ );
and  ( new_n15584_, new_n15583_, new_n15582_ );
and  ( new_n15585_, new_n15584_, new_n15581_ );
and  ( new_n15586_, new_n15585_, new_n15578_ );
or   ( new_n15587_, new_n15586_, new_n15577_ );
or   ( new_n15588_, new_n15584_, new_n15581_ );
and  ( new_n15589_, new_n15588_, new_n15578_ );
and  ( new_n15590_, new_n5289_, new_n5145_ );
and  ( new_n15591_, new_n5292_, new_n5285_ );
or   ( new_n15592_, new_n15591_, new_n15590_ );
and  ( new_n15593_, new_n15592_, new_n5713_ );
or   ( new_n15594_, new_n15592_, new_n5713_ );
and  ( new_n15595_, new_n5712_, new_n5301_ );
and  ( new_n15596_, new_n5581_, new_n5574_ );
or   ( new_n15597_, new_n15596_, new_n15595_ );
or   ( new_n15598_, new_n6123_, new_n5997_ );
and  ( new_n15599_, new_n15598_, new_n6132_ );
or   ( new_n15600_, new_n15599_, new_n6124_ );
and  ( new_n15601_, new_n15600_, new_n15597_ );
and  ( new_n15602_, new_n15601_, new_n15594_ );
or   ( new_n15603_, new_n15602_, new_n15593_ );
and  ( new_n15604_, new_n15603_, new_n15589_ );
or   ( new_n15605_, new_n15604_, new_n15587_ );
or   ( new_n15606_, new_n15600_, new_n15597_ );
and  ( new_n15607_, new_n15606_, new_n15594_ );
and  ( new_n15608_, new_n15607_, new_n15589_ );
and  ( new_n15609_, new_n6129_, new_n5984_ );
and  ( new_n15610_, new_n6132_, new_n6125_ );
or   ( new_n15611_, new_n15610_, new_n15609_ );
or   ( new_n15612_, new_n6619_, new_n6471_ );
or   ( new_n15613_, new_n6628_, new_n6620_ );
and  ( new_n15614_, new_n15613_, new_n15612_ );
or   ( new_n15615_, new_n15614_, new_n15611_ );
and  ( new_n15616_, new_n15614_, new_n15611_ );
and  ( new_n15617_, new_n6625_, new_n6460_ );
and  ( new_n15618_, new_n6628_, new_n6621_ );
or   ( new_n15619_, new_n15618_, new_n15617_ );
or   ( new_n15620_, new_n7039_, new_n6910_ );
and  ( new_n15621_, new_n15620_, new_n7048_ );
or   ( new_n15622_, new_n15621_, new_n7040_ );
and  ( new_n15623_, new_n15622_, new_n15619_ );
or   ( new_n15624_, new_n15623_, new_n15616_ );
and  ( new_n15625_, new_n15624_, new_n15615_ );
or   ( new_n15626_, new_n15622_, new_n15619_ );
and  ( new_n15627_, new_n15626_, new_n15615_ );
and  ( new_n15628_, new_n7045_, new_n6900_ );
and  ( new_n15629_, new_n7048_, new_n7041_ );
or   ( new_n15630_, new_n15629_, new_n15628_ );
or   ( new_n15631_, new_n7558_, new_n7414_ );
or   ( new_n15632_, new_n7567_, new_n7559_ );
and  ( new_n15633_, new_n15632_, new_n15631_ );
or   ( new_n15634_, new_n15633_, new_n15630_ );
and  ( new_n15635_, new_n15633_, new_n15630_ );
and  ( new_n15636_, new_n7564_, new_n7402_ );
and  ( new_n15637_, new_n7567_, new_n7560_ );
or   ( new_n15638_, new_n15637_, new_n15636_ );
or   ( new_n15639_, new_n7996_, new_n7863_ );
and  ( new_n15640_, new_n15639_, new_n8005_ );
or   ( new_n15641_, new_n15640_, new_n7997_ );
and  ( new_n15642_, new_n15641_, new_n15638_ );
or   ( new_n15643_, new_n15642_, new_n15635_ );
and  ( new_n15644_, new_n15643_, new_n15634_ );
and  ( new_n15645_, new_n15644_, new_n15627_ );
or   ( new_n15646_, new_n15645_, new_n15625_ );
and  ( new_n15647_, new_n15646_, new_n15608_ );
or   ( new_n15648_, new_n15647_, new_n15605_ );
and  ( new_n15649_, new_n8002_, new_n7851_ );
and  ( new_n15650_, new_n8005_, new_n7998_ );
or   ( new_n15651_, new_n15650_, new_n15649_ );
or   ( new_n15652_, new_n8431_, new_n8297_ );
or   ( new_n15653_, new_n8440_, new_n8432_ );
and  ( new_n15654_, new_n15653_, new_n15652_ );
or   ( new_n15655_, new_n15654_, new_n15651_ );
and  ( new_n15656_, new_n15654_, new_n15651_ );
and  ( new_n15657_, new_n8437_, new_n8290_ );
and  ( new_n15658_, new_n8440_, new_n8433_ );
or   ( new_n15659_, new_n15658_, new_n15657_ );
or   ( new_n15660_, new_n8923_, new_n8770_ );
and  ( new_n15661_, new_n15660_, new_n8932_ );
or   ( new_n15662_, new_n15661_, new_n8924_ );
and  ( new_n15663_, new_n15662_, new_n15659_ );
or   ( new_n15664_, new_n15663_, new_n15656_ );
and  ( new_n15665_, new_n15664_, new_n15655_ );
or   ( new_n15666_, new_n15662_, new_n15659_ );
and  ( new_n15667_, new_n15666_, new_n15655_ );
and  ( new_n15668_, new_n8929_, new_n8760_ );
and  ( new_n15669_, new_n8932_, new_n8925_ );
or   ( new_n15670_, new_n15669_, new_n15668_ );
or   ( new_n15671_, new_n9333_, new_n9209_ );
or   ( new_n15672_, new_n9342_, new_n9334_ );
and  ( new_n15673_, new_n15672_, new_n15671_ );
or   ( new_n15674_, new_n15673_, new_n15670_ );
and  ( new_n15675_, new_n15673_, new_n15670_ );
and  ( new_n15676_, new_n9339_, new_n9202_ );
and  ( new_n15677_, new_n9342_, new_n9335_ );
or   ( new_n15678_, new_n15677_, new_n15676_ );
or   ( new_n15679_, new_n9708_, new_n9595_ );
and  ( new_n15680_, new_n15679_, new_n9717_ );
or   ( new_n15681_, new_n15680_, new_n9709_ );
and  ( new_n15682_, new_n15681_, new_n15678_ );
or   ( new_n15683_, new_n15682_, new_n15675_ );
and  ( new_n15684_, new_n15683_, new_n15674_ );
and  ( new_n15685_, new_n15684_, new_n15667_ );
or   ( new_n15686_, new_n15685_, new_n15665_ );
or   ( new_n15687_, new_n15681_, new_n15678_ );
and  ( new_n15688_, new_n15687_, new_n15674_ );
and  ( new_n15689_, new_n15688_, new_n15667_ );
and  ( new_n15690_, new_n9714_, new_n9582_ );
and  ( new_n15691_, new_n9717_, new_n9710_ );
or   ( new_n15692_, new_n15691_, new_n15690_ );
or   ( new_n15693_, new_n10130_, new_n10006_ );
or   ( new_n15694_, new_n10139_, new_n10131_ );
and  ( new_n15695_, new_n15694_, new_n15693_ );
or   ( new_n15696_, new_n15695_, new_n15692_ );
and  ( new_n15697_, new_n15695_, new_n15692_ );
and  ( new_n15698_, new_n10136_, new_n9995_ );
and  ( new_n15699_, new_n10139_, new_n10132_ );
or   ( new_n15700_, new_n15699_, new_n15698_ );
or   ( new_n15701_, new_n10499_, new_n10386_ );
and  ( new_n15702_, new_n15701_, new_n10508_ );
or   ( new_n15703_, new_n15702_, new_n10500_ );
and  ( new_n15704_, new_n15703_, new_n15700_ );
or   ( new_n15705_, new_n15704_, new_n15697_ );
and  ( new_n15706_, new_n15705_, new_n15696_ );
or   ( new_n15707_, new_n15703_, new_n15700_ );
and  ( new_n15708_, new_n15707_, new_n15696_ );
and  ( new_n15709_, new_n10505_, new_n10376_ );
and  ( new_n15710_, new_n10508_, new_n10501_ );
or   ( new_n15711_, new_n15710_, new_n15709_ );
or   ( new_n15712_, new_n10917_, new_n10793_ );
or   ( new_n15713_, new_n10926_, new_n10918_ );
and  ( new_n15714_, new_n15713_, new_n15712_ );
or   ( new_n15715_, new_n15714_, new_n15711_ );
and  ( new_n15716_, new_n15714_, new_n15711_ );
and  ( new_n15717_, new_n10923_, new_n10782_ );
and  ( new_n15718_, new_n10926_, new_n10919_ );
or   ( new_n15719_, new_n15718_, new_n15717_ );
or   ( new_n15720_, new_n11291_, new_n11178_ );
and  ( new_n15721_, new_n15720_, new_n11300_ );
or   ( new_n15722_, new_n15721_, new_n11292_ );
and  ( new_n15723_, new_n15722_, new_n15719_ );
or   ( new_n15724_, new_n15723_, new_n15716_ );
and  ( new_n15725_, new_n15724_, new_n15715_ );
and  ( new_n15726_, new_n15725_, new_n15708_ );
or   ( new_n15727_, new_n15726_, new_n15706_ );
and  ( new_n15728_, new_n15727_, new_n15689_ );
or   ( new_n15729_, new_n15728_, new_n15686_ );
or   ( new_n15730_, new_n15722_, new_n15719_ );
and  ( new_n15731_, new_n15730_, new_n15715_ );
and  ( new_n15732_, new_n15731_, new_n15708_ );
and  ( new_n15733_, new_n11297_, new_n11163_ );
and  ( new_n15734_, new_n11300_, new_n11293_ );
or   ( new_n15735_, new_n15734_, new_n15733_ );
and  ( new_n15736_, new_n15735_, new_n11643_ );
or   ( new_n15737_, new_n15735_, new_n11643_ );
and  ( new_n15738_, new_n11642_, new_n11309_ );
and  ( new_n15739_, new_n11534_, new_n11527_ );
or   ( new_n15740_, new_n15739_, new_n15738_ );
and  ( new_n15741_, new_n15740_, new_n11672_ );
and  ( new_n15742_, new_n15741_, new_n15737_ );
or   ( new_n15743_, new_n15742_, new_n15736_ );
or   ( new_n15744_, new_n15740_, new_n11672_ );
and  ( new_n15745_, new_n15744_, new_n15737_ );
and  ( new_n15746_, new_n11668_, new_n11658_ );
and  ( new_n15747_, new_n11671_, new_n11651_ );
or   ( new_n15748_, new_n15747_, new_n15746_ );
or   ( new_n15749_, new_n11948_, new_n11861_ );
and  ( new_n15750_, new_n15749_, new_n11957_ );
or   ( new_n15751_, new_n15750_, new_n11949_ );
and  ( new_n15752_, new_n15751_, new_n15748_ );
or   ( new_n15753_, new_n15751_, new_n15748_ );
and  ( new_n15754_, new_n11954_, new_n11854_ );
and  ( new_n15755_, new_n11957_, new_n11950_ );
or   ( new_n15756_, new_n15755_, new_n15754_ );
or   ( new_n15757_, new_n12285_, new_n12185_ );
or   ( new_n15758_, new_n12294_, new_n12286_ );
and  ( new_n15759_, new_n15758_, new_n15757_ );
and  ( new_n15760_, new_n15759_, new_n15756_ );
and  ( new_n15761_, new_n15760_, new_n15753_ );
or   ( new_n15762_, new_n15761_, new_n15752_ );
and  ( new_n15763_, new_n15762_, new_n15745_ );
or   ( new_n15764_, new_n15763_, new_n15743_ );
or   ( new_n15765_, new_n15759_, new_n15756_ );
and  ( new_n15766_, new_n15765_, new_n15753_ );
and  ( new_n15767_, new_n15766_, new_n15745_ );
and  ( new_n15768_, new_n12291_, new_n12172_ );
and  ( new_n15769_, new_n12294_, new_n12287_ );
or   ( new_n15770_, new_n15769_, new_n15768_ );
or   ( new_n15771_, new_n12542_, new_n12469_ );
and  ( new_n15772_, new_n15771_, new_n12551_ );
or   ( new_n15773_, new_n15772_, new_n12543_ );
or   ( new_n15774_, new_n15773_, new_n15770_ );
and  ( new_n15775_, new_n12548_, new_n12463_ );
and  ( new_n15776_, new_n12551_, new_n12544_ );
or   ( new_n15777_, new_n15776_, new_n15775_ );
or   ( new_n15778_, new_n12814_, new_n12740_ );
or   ( new_n15779_, new_n12823_, new_n12815_ );
and  ( new_n15780_, new_n15779_, new_n15778_ );
or   ( new_n15781_, new_n15780_, new_n15777_ );
and  ( new_n15782_, new_n15781_, new_n15774_ );
and  ( new_n15783_, new_n12820_, new_n12729_ );
and  ( new_n15784_, new_n12823_, new_n12816_ );
or   ( new_n15785_, new_n15784_, new_n15783_ );
or   ( new_n15786_, new_n13061_, new_n12988_ );
and  ( new_n15787_, new_n15786_, new_n13070_ );
or   ( new_n15788_, new_n15787_, new_n13062_ );
or   ( new_n15789_, new_n15788_, new_n15785_ );
and  ( new_n15790_, new_n13067_, new_n12982_ );
and  ( new_n15791_, new_n13070_, new_n13063_ );
or   ( new_n15792_, new_n15791_, new_n15790_ );
or   ( new_n15793_, new_n13347_, new_n13267_ );
or   ( new_n15794_, new_n13356_, new_n13348_ );
and  ( new_n15795_, new_n15794_, new_n15793_ );
or   ( new_n15796_, new_n15795_, new_n15792_ );
and  ( new_n15797_, new_n15796_, new_n15789_ );
and  ( new_n15798_, new_n13353_, new_n13256_ );
and  ( new_n15799_, new_n13356_, new_n13349_ );
or   ( new_n15800_, new_n15799_, new_n15798_ );
or   ( new_n15801_, new_n13579_, new_n13512_ );
and  ( new_n15802_, new_n15801_, new_n13588_ );
or   ( new_n15803_, new_n15802_, new_n13580_ );
or   ( new_n15804_, new_n15803_, new_n15800_ );
and  ( new_n15805_, new_n13585_, new_n13506_ );
and  ( new_n15806_, new_n13588_, new_n13581_ );
or   ( new_n15807_, new_n15806_, new_n15805_ );
or   ( new_n15808_, new_n15807_, new_n13956_ );
and  ( new_n15809_, new_n15808_, new_n15804_ );
and  ( new_n15810_, new_n13830_, new_n13826_ );
and  ( new_n15811_, new_n13833_, new_n13748_ );
or   ( new_n15812_, new_n15811_, new_n15810_ );
or   ( new_n15813_, new_n14010_, new_n13963_ );
and  ( new_n15814_, new_n15813_, new_n14019_ );
or   ( new_n15815_, new_n15814_, new_n14011_ );
or   ( new_n15816_, new_n15815_, new_n15812_ );
and  ( new_n15817_, new_n13955_, new_n13597_ );
and  ( new_n15818_, new_n13952_, new_n13738_ );
or   ( new_n15819_, new_n15818_, new_n15817_ );
or   ( new_n15820_, new_n15819_, new_n13834_ );
and  ( new_n15821_, new_n15820_, new_n15816_ );
and  ( new_n15822_, new_n14016_, new_n13945_ );
and  ( new_n15823_, new_n14019_, new_n14012_ );
or   ( new_n15824_, new_n15823_, new_n15822_ );
or   ( new_n15825_, new_n14162_, new_n14122_ );
or   ( new_n15826_, new_n14171_, new_n14163_ );
and  ( new_n15827_, new_n15826_, new_n15825_ );
or   ( new_n15828_, new_n15827_, new_n15824_ );
and  ( new_n15829_, new_n14168_, new_n14116_ );
and  ( new_n15830_, new_n14171_, new_n14164_ );
or   ( new_n15831_, new_n15830_, new_n15829_ );
or   ( new_n15832_, new_n14590_, new_n14318_ );
and  ( new_n15833_, new_n15832_, new_n14599_ );
or   ( new_n15834_, new_n15833_, new_n14591_ );
or   ( new_n15835_, new_n15834_, new_n15831_ );
and  ( new_n15836_, new_n15835_, new_n15828_ );
and  ( new_n15837_, new_n14508_, new_n14504_ );
and  ( new_n15838_, new_n14511_, new_n14487_ );
or   ( new_n15839_, new_n15838_, new_n15837_ );
or   ( new_n15840_, new_n15839_, new_n14644_ );
and  ( new_n15841_, new_n14596_, new_n14306_ );
and  ( new_n15842_, new_n14599_, new_n14592_ );
or   ( new_n15843_, new_n15842_, new_n15841_ );
or   ( new_n15844_, new_n14485_, new_n14445_ );
or   ( new_n15845_, new_n14511_, new_n14486_ );
and  ( new_n15846_, new_n15845_, new_n15844_ );
or   ( new_n15847_, new_n15846_, new_n15843_ );
and  ( new_n15848_, new_n15847_, new_n15840_ );
and  ( new_n15849_, new_n14643_, new_n14520_ );
and  ( new_n15850_, new_n14610_, new_n14585_ );
or   ( new_n15851_, new_n15850_, new_n15849_ );
or   ( new_n15852_, new_n15851_, new_n14793_ );
and  ( new_n15853_, new_n14792_, new_n14652_ );
and  ( new_n15854_, new_n14748_, new_n14742_ );
or   ( new_n15855_, new_n15854_, new_n15853_ );
or   ( new_n15856_, new_n15855_, new_n14974_ );
and  ( new_n15857_, new_n15856_, new_n15852_ );
and  ( new_n15858_, new_n14902_, new_n14898_ );
and  ( new_n15859_, new_n14905_, new_n14891_ );
or   ( new_n15860_, new_n15859_, new_n15858_ );
or   ( new_n15861_, new_n15860_, new_n15009_ );
and  ( new_n15862_, new_n14970_, new_n14808_ );
and  ( new_n15863_, new_n14973_, new_n14801_ );
or   ( new_n15864_, new_n15863_, new_n15862_ );
or   ( new_n15865_, new_n14889_, new_n14866_ );
and  ( new_n15866_, new_n15865_, new_n14905_ );
or   ( new_n15867_, new_n15866_, new_n14890_ );
or   ( new_n15868_, new_n15867_, new_n15864_ );
and  ( new_n15869_, new_n15868_, new_n15861_ );
and  ( new_n15870_, new_n15008_, new_n14914_ );
and  ( new_n15871_, new_n14984_, new_n14964_ );
or   ( new_n15872_, new_n15871_, new_n15870_ );
and  ( new_n15873_, new_n15872_, new_n15035_ );
or   ( new_n15874_, new_n15872_, new_n15035_ );
and  ( new_n15875_, new_n15031_, new_n15024_ );
and  ( new_n15876_, new_n15034_, new_n15017_ );
or   ( new_n15877_, new_n15876_, new_n15875_ );
or   ( new_n15878_, new_n15101_, new_n15088_ );
and  ( new_n15879_, new_n15878_, new_n15110_ );
or   ( new_n15880_, new_n15879_, new_n15102_ );
and  ( new_n15881_, new_n15880_, new_n15877_ );
and  ( new_n15882_, new_n15881_, new_n15874_ );
or   ( new_n15883_, new_n15882_, new_n15873_ );
or   ( new_n15884_, new_n15880_, new_n15877_ );
and  ( new_n15885_, new_n15884_, new_n15874_ );
and  ( new_n15886_, new_n15107_, new_n15078_ );
and  ( new_n15887_, new_n15110_, new_n15103_ );
or   ( new_n15888_, new_n15887_, new_n15886_ );
or   ( new_n15889_, new_n15888_, new_n15159_ );
and  ( new_n15890_, new_n15158_, new_n15119_ );
and  ( new_n15891_, new_n15148_, new_n15141_ );
or   ( new_n15892_, new_n15891_, new_n15890_ );
or   ( new_n15893_, new_n15892_, new_n15185_ );
and  ( new_n15894_, new_n15181_, new_n15172_ );
and  ( new_n15895_, new_n15184_, new_n15165_ );
or   ( new_n15896_, new_n15895_, new_n15894_ );
and  ( new_n15897_, new_n15896_, new_n15216_ );
or   ( new_n15898_, new_n15896_, new_n15216_ );
and  ( new_n15899_, new_n15212_, new_n15204_ );
and  ( new_n15900_, new_n15215_, new_n15195_ );
or   ( new_n15901_, new_n15900_, new_n15899_ );
or   ( new_n15902_, new_n15901_, new_n15233_ );
and  ( new_n15903_, new_n15232_, new_n6039_ );
and  ( new_n15904_, new_n15226_, new_n5867_ );
or   ( new_n15905_, new_n15904_, new_n15903_ );
and  ( new_n15906_, new_n15237_, new_n6039_ );
and  ( new_n15907_, new_n15235_, new_n5867_ );
or   ( new_n15908_, new_n15907_, new_n15906_ );
or   ( new_n15909_, new_n15908_, new_n15905_ );
or   ( new_n15910_, new_n7099_, new_n124_ );
and  ( new_n15911_, new_n15910_, new_n7274_ );
or   ( new_n15912_, new_n7099_, new_n5854_ );
and  ( new_n15913_, new_n15912_, new_n7105_ );
or   ( new_n15914_, new_n15913_, new_n15911_ );
and  ( new_n15915_, new_n15914_, new_n6037_ );
and  ( new_n15916_, new_n15915_, new_n15909_ );
and  ( new_n15917_, new_n15916_, new_n15902_ );
and  ( new_n15918_, new_n15901_, new_n15233_ );
and  ( new_n15919_, new_n15908_, new_n15905_ );
and  ( new_n15920_, new_n15919_, new_n15902_ );
or   ( new_n15921_, new_n15920_, new_n15918_ );
or   ( new_n15922_, new_n15921_, new_n15917_ );
and  ( new_n15923_, new_n15922_, new_n15898_ );
or   ( new_n15924_, new_n15923_, new_n15897_ );
and  ( new_n15925_, new_n15924_, new_n15893_ );
and  ( new_n15926_, new_n15925_, new_n15889_ );
and  ( new_n15927_, new_n15888_, new_n15159_ );
and  ( new_n15928_, new_n15892_, new_n15185_ );
and  ( new_n15929_, new_n15928_, new_n15889_ );
or   ( new_n15930_, new_n15929_, new_n15927_ );
or   ( new_n15931_, new_n15930_, new_n15926_ );
and  ( new_n15932_, new_n15931_, new_n15885_ );
or   ( new_n15933_, new_n15932_, new_n15883_ );
and  ( new_n15934_, new_n15933_, new_n15869_ );
and  ( new_n15935_, new_n15934_, new_n15857_ );
and  ( new_n15936_, new_n15851_, new_n14793_ );
and  ( new_n15937_, new_n15855_, new_n14974_ );
and  ( new_n15938_, new_n15937_, new_n15852_ );
or   ( new_n15939_, new_n15938_, new_n15936_ );
and  ( new_n15940_, new_n15867_, new_n15864_ );
and  ( new_n15941_, new_n15860_, new_n15009_ );
and  ( new_n15942_, new_n15941_, new_n15868_ );
or   ( new_n15943_, new_n15942_, new_n15940_ );
and  ( new_n15944_, new_n15943_, new_n15857_ );
or   ( new_n15945_, new_n15944_, new_n15939_ );
or   ( new_n15946_, new_n15945_, new_n15935_ );
and  ( new_n15947_, new_n15946_, new_n15848_ );
and  ( new_n15948_, new_n15947_, new_n15836_ );
and  ( new_n15949_, new_n15827_, new_n15824_ );
and  ( new_n15950_, new_n15834_, new_n15831_ );
or   ( new_n15951_, new_n15950_, new_n15949_ );
and  ( new_n15952_, new_n15951_, new_n15828_ );
and  ( new_n15953_, new_n15846_, new_n15843_ );
and  ( new_n15954_, new_n15839_, new_n14644_ );
or   ( new_n15955_, new_n15954_, new_n15953_ );
and  ( new_n15956_, new_n15955_, new_n15847_ );
and  ( new_n15957_, new_n15956_, new_n15836_ );
or   ( new_n15958_, new_n15957_, new_n15952_ );
or   ( new_n15959_, new_n15958_, new_n15948_ );
and  ( new_n15960_, new_n15959_, new_n15821_ );
and  ( new_n15961_, new_n15960_, new_n15809_ );
and  ( new_n15962_, new_n15803_, new_n15800_ );
and  ( new_n15963_, new_n15807_, new_n13956_ );
and  ( new_n15964_, new_n15963_, new_n15804_ );
or   ( new_n15965_, new_n15964_, new_n15962_ );
and  ( new_n15966_, new_n15819_, new_n13834_ );
and  ( new_n15967_, new_n15815_, new_n15812_ );
and  ( new_n15968_, new_n15967_, new_n15820_ );
or   ( new_n15969_, new_n15968_, new_n15966_ );
and  ( new_n15970_, new_n15969_, new_n15809_ );
or   ( new_n15971_, new_n15970_, new_n15965_ );
or   ( new_n15972_, new_n15971_, new_n15961_ );
and  ( new_n15973_, new_n15972_, new_n15797_ );
and  ( new_n15974_, new_n15973_, new_n15782_ );
and  ( new_n15975_, new_n15773_, new_n15770_ );
and  ( new_n15976_, new_n15780_, new_n15777_ );
and  ( new_n15977_, new_n15976_, new_n15774_ );
or   ( new_n15978_, new_n15977_, new_n15975_ );
and  ( new_n15979_, new_n15788_, new_n15785_ );
and  ( new_n15980_, new_n15795_, new_n15792_ );
and  ( new_n15981_, new_n15980_, new_n15789_ );
or   ( new_n15982_, new_n15981_, new_n15979_ );
and  ( new_n15983_, new_n15982_, new_n15782_ );
or   ( new_n15984_, new_n15983_, new_n15978_ );
or   ( new_n15985_, new_n15984_, new_n15974_ );
and  ( new_n15986_, new_n15985_, new_n15767_ );
or   ( new_n15987_, new_n15986_, new_n15764_ );
and  ( new_n15988_, new_n15987_, new_n15732_ );
and  ( new_n15989_, new_n15988_, new_n15689_ );
or   ( new_n15990_, new_n15989_, new_n15729_ );
or   ( new_n15991_, new_n15641_, new_n15638_ );
and  ( new_n15992_, new_n15991_, new_n15634_ );
and  ( new_n15993_, new_n15992_, new_n15627_ );
and  ( new_n15994_, new_n15993_, new_n15608_ );
and  ( new_n15995_, new_n15994_, new_n15990_ );
or   ( new_n15996_, new_n15995_, new_n15648_ );
and  ( new_n15997_, new_n15996_, new_n15573_ );
or   ( new_n15998_, new_n15997_, new_n15569_ );
and  ( new_n15999_, new_n15998_, new_n15509_ );
or   ( new_n16000_, new_n15999_, new_n15506_ );
xor  ( new_n16001_, new_n506_, new_n491_ );
nand ( new_n16002_, new_n16001_, new_n138_ );
and  ( new_n16003_, new_n16002_, RI2b1c4342baa0_9 );
xor  ( new_n16004_, new_n429_, new_n420_ );
or   ( new_n16005_, new_n16004_, new_n471_ );
xor  ( new_n16006_, new_n499_, new_n488_ );
or   ( new_n16007_, new_n16006_, new_n478_ );
or   ( new_n16008_, new_n16007_, new_n16005_ );
and  ( new_n16009_, new_n16008_, new_n16003_ );
nand ( new_n16010_, new_n16006_, new_n138_ );
and  ( new_n16011_, new_n16010_, RI2b1c4342bb18_10 );
or   ( new_n16012_, new_n16011_, new_n16003_ );
nand ( new_n16013_, new_n16004_, new_n138_ );
and  ( new_n16014_, new_n16013_, RI2b1c4342bb90_11 );
or   ( new_n16015_, new_n16014_, new_n16007_ );
or   ( new_n16016_, new_n16011_, new_n16005_ );
and  ( new_n16017_, new_n16016_, new_n16015_ );
or   ( new_n16018_, new_n16001_, new_n556_ );
or   ( new_n16019_, new_n16018_, new_n16007_ );
and  ( new_n16020_, new_n16019_, new_n16017_ );
and  ( new_n16021_, new_n16020_, new_n16012_ );
and  ( new_n16022_, new_n16021_, RI2b1c4342d648_68 );
or   ( new_n16023_, new_n16014_, new_n16011_ );
and  ( new_n16024_, new_n16023_, new_n16008_ );
and  ( new_n16025_, new_n16024_, RI2b1c4342d5d0_67 );
or   ( new_n16026_, new_n16025_, new_n16022_ );
or   ( new_n16027_, new_n16026_, new_n16009_ );
and  ( new_n16028_, new_n16014_, new_n16011_ );
or   ( new_n16029_, new_n16028_, new_n16018_ );
or   ( new_n16030_, new_n16018_, new_n16011_ );
or   ( new_n16031_, new_n16007_, new_n16003_ );
and  ( new_n16032_, new_n16031_, new_n16030_ );
or   ( new_n16033_, new_n16032_, new_n16024_ );
or   ( new_n16034_, new_n16033_, new_n612_ );
or   ( new_n16035_, new_n16017_, new_n112_ );
and  ( new_n16036_, new_n16035_, new_n16034_ );
or   ( new_n16037_, new_n16036_, new_n16029_ );
and  ( new_n16038_, new_n16037_, new_n16027_ );
xor  ( new_n16039_, new_n258_, new_n257_ );
or   ( new_n16040_, new_n16039_, new_n394_ );
xor  ( new_n16041_, new_n902_, new_n250_ );
nand ( new_n16042_, new_n16041_, new_n138_ );
and  ( new_n16043_, new_n16042_, RI2b1c4342bd70_15 );
xor  ( new_n16044_, new_n907_, new_n255_ );
nand ( new_n16045_, new_n16044_, new_n138_ );
and  ( new_n16046_, new_n16045_, RI2b1c4342bcf8_14 );
and  ( new_n16047_, new_n16046_, new_n16043_ );
or   ( new_n16048_, new_n16047_, new_n16040_ );
xor  ( new_n16049_, new_n392_, new_n391_ );
or   ( new_n16050_, new_n16049_, new_n408_ );
or   ( new_n16051_, new_n16050_, new_n16040_ );
and  ( new_n16052_, new_n16051_, new_n16014_ );
nand ( new_n16053_, new_n16049_, new_n138_ );
and  ( new_n16054_, new_n16053_, RI2b1c4342bc08_12 );
or   ( new_n16055_, new_n16054_, new_n16014_ );
nand ( new_n16056_, new_n16039_, new_n138_ );
and  ( new_n16057_, new_n16056_, RI2b1c4342bc80_13 );
or   ( new_n16058_, new_n16057_, new_n16050_ );
or   ( new_n16059_, new_n16054_, new_n16040_ );
and  ( new_n16060_, new_n16059_, new_n16058_ );
or   ( new_n16061_, new_n16050_, new_n16005_ );
and  ( new_n16062_, new_n16061_, new_n16060_ );
and  ( new_n16063_, new_n16062_, new_n16055_ );
and  ( new_n16064_, new_n16063_, RI2b1c4342d558_66 );
or   ( new_n16065_, new_n16057_, new_n16054_ );
and  ( new_n16066_, new_n16065_, new_n16051_ );
and  ( new_n16067_, new_n16066_, RI2b1c4342d4e0_65 );
or   ( new_n16068_, new_n16067_, new_n16064_ );
or   ( new_n16069_, new_n16068_, new_n16052_ );
and  ( new_n16070_, new_n16057_, new_n16054_ );
or   ( new_n16071_, new_n16070_, new_n16005_ );
or   ( new_n16072_, new_n16054_, new_n16005_ );
or   ( new_n16073_, new_n16050_, new_n16014_ );
and  ( new_n16074_, new_n16073_, new_n16072_ );
or   ( new_n16075_, new_n16074_, new_n16066_ );
or   ( new_n16076_, new_n16075_, new_n526_ );
or   ( new_n16077_, new_n16060_, new_n99_ );
and  ( new_n16078_, new_n16077_, new_n16076_ );
or   ( new_n16079_, new_n16078_, new_n16071_ );
and  ( new_n16080_, new_n16079_, new_n16069_ );
or   ( new_n16081_, new_n16080_, new_n16048_ );
or   ( new_n16082_, new_n16041_, new_n266_ );
or   ( new_n16083_, new_n16044_, new_n263_ );
or   ( new_n16084_, new_n16083_, new_n16082_ );
and  ( new_n16085_, new_n16084_, new_n16057_ );
or   ( new_n16086_, new_n16078_, new_n16052_ );
or   ( new_n16087_, new_n16071_, new_n16068_ );
and  ( new_n16088_, new_n16087_, new_n16086_ );
or   ( new_n16089_, new_n16088_, new_n16085_ );
and  ( new_n16090_, new_n16089_, new_n16081_ );
or   ( new_n16091_, new_n16090_, new_n16038_ );
or   ( new_n16092_, new_n16036_, new_n16009_ );
or   ( new_n16093_, new_n16029_, new_n16026_ );
and  ( new_n16094_, new_n16093_, new_n16092_ );
or   ( new_n16095_, new_n16085_, new_n16080_ );
or   ( new_n16096_, new_n16088_, new_n16048_ );
and  ( new_n16097_, new_n16096_, new_n16095_ );
or   ( new_n16098_, new_n16097_, new_n16094_ );
and  ( new_n16099_, new_n16098_, new_n16091_ );
xor  ( new_n16100_, new_n715_, new_n668_ );
or   ( new_n16101_, new_n16100_, new_n137_ );
and  ( new_n16102_, new_n16101_, RI2b1c4342b6e0_1 );
xor  ( new_n16103_, new_n786_, new_n658_ );
or   ( new_n16104_, new_n16103_, new_n677_ );
xor  ( new_n16105_, new_n832_, new_n663_ );
or   ( new_n16106_, new_n16105_, new_n711_ );
or   ( new_n16107_, new_n16106_, new_n16104_ );
and  ( new_n16108_, new_n16107_, new_n16102_ );
nand ( new_n16109_, new_n16105_, new_n138_ );
and  ( new_n16110_, new_n16109_, RI2b1c4342b758_2 );
nand ( new_n16111_, new_n16103_, new_n138_ );
and  ( new_n16112_, new_n16111_, RI2b1c4342b7d0_3 );
or   ( new_n16113_, new_n16112_, new_n16110_ );
and  ( new_n16114_, new_n16113_, new_n16107_ );
nand ( new_n16115_, new_n16100_, new_n671_ );
or   ( new_n16116_, new_n16115_, new_n16110_ );
or   ( new_n16117_, new_n16106_, new_n16102_ );
and  ( new_n16118_, new_n16117_, new_n16116_ );
or   ( new_n16119_, new_n16118_, new_n16114_ );
or   ( new_n16120_, new_n16119_, new_n886_ );
or   ( new_n16121_, new_n16112_, new_n16106_ );
or   ( new_n16122_, new_n16110_, new_n16104_ );
and  ( new_n16123_, new_n16122_, new_n16121_ );
or   ( new_n16124_, new_n16123_, new_n843_ );
and  ( new_n16125_, new_n16124_, new_n16120_ );
or   ( new_n16126_, new_n16125_, new_n16108_ );
and  ( new_n16127_, new_n16112_, new_n16110_ );
or   ( new_n16128_, new_n16127_, new_n16115_ );
or   ( new_n16129_, new_n16110_, new_n16102_ );
or   ( new_n16130_, new_n16115_, new_n16106_ );
and  ( new_n16131_, new_n16130_, new_n16123_ );
and  ( new_n16132_, new_n16131_, new_n16129_ );
and  ( new_n16133_, new_n16132_, RI2b1c4342da08_76 );
and  ( new_n16134_, new_n16114_, RI2b1c4342d990_75 );
or   ( new_n16135_, new_n16134_, new_n16133_ );
or   ( new_n16136_, new_n16135_, new_n16128_ );
and  ( new_n16137_, new_n16136_, new_n16126_ );
or   ( new_n16138_, new_n16115_, new_n1004_ );
or   ( new_n16139_, new_n16138_, new_n16137_ );
or   ( new_n16140_, new_n16135_, new_n16108_ );
or   ( new_n16141_, new_n16128_, new_n16125_ );
and  ( new_n16142_, new_n16141_, new_n16140_ );
and  ( new_n16143_, new_n16102_, RI2b1c4342da80_77 );
or   ( new_n16144_, new_n16143_, new_n16142_ );
and  ( new_n16145_, new_n16144_, new_n16139_ );
xor  ( new_n16146_, new_n735_, new_n651_ );
or   ( new_n16147_, new_n16146_, new_n685_ );
xor  ( new_n16148_, new_n779_, new_n656_ );
or   ( new_n16149_, new_n16148_, new_n682_ );
or   ( new_n16150_, new_n16149_, new_n16147_ );
and  ( new_n16151_, new_n16150_, new_n16112_ );
nand ( new_n16152_, new_n16148_, new_n138_ );
and  ( new_n16153_, new_n16152_, RI2b1c4342b848_4 );
or   ( new_n16154_, new_n16153_, new_n16112_ );
or   ( new_n16155_, new_n16149_, new_n16104_ );
nand ( new_n16156_, new_n16146_, new_n138_ );
and  ( new_n16157_, new_n16156_, RI2b1c4342b8c0_5 );
or   ( new_n16158_, new_n16157_, new_n16149_ );
or   ( new_n16159_, new_n16153_, new_n16147_ );
and  ( new_n16160_, new_n16159_, new_n16158_ );
and  ( new_n16161_, new_n16160_, new_n16155_ );
and  ( new_n16162_, new_n16161_, new_n16154_ );
and  ( new_n16163_, new_n16162_, RI2b1c4342d918_74 );
or   ( new_n16164_, new_n16157_, new_n16153_ );
and  ( new_n16165_, new_n16164_, new_n16150_ );
and  ( new_n16166_, new_n16165_, RI2b1c4342d8a0_73 );
or   ( new_n16167_, new_n16166_, new_n16163_ );
or   ( new_n16168_, new_n16167_, new_n16151_ );
and  ( new_n16169_, new_n16157_, new_n16153_ );
or   ( new_n16170_, new_n16169_, new_n16104_ );
or   ( new_n16171_, new_n16153_, new_n16104_ );
or   ( new_n16172_, new_n16149_, new_n16112_ );
and  ( new_n16173_, new_n16172_, new_n16171_ );
or   ( new_n16174_, new_n16173_, new_n16165_ );
or   ( new_n16175_, new_n16174_, new_n859_ );
or   ( new_n16176_, new_n16160_, new_n105_ );
and  ( new_n16177_, new_n16176_, new_n16175_ );
or   ( new_n16178_, new_n16177_, new_n16170_ );
and  ( new_n16179_, new_n16178_, new_n16168_ );
xor  ( new_n16180_, new_n592_, new_n576_ );
nand ( new_n16181_, new_n16180_, new_n138_ );
and  ( new_n16182_, new_n16181_, RI2b1c4342b9b0_7 );
xor  ( new_n16183_, new_n584_, new_n573_ );
or   ( new_n16184_, new_n16183_, new_n563_ );
or   ( new_n16185_, new_n16184_, new_n16018_ );
and  ( new_n16186_, new_n16185_, new_n16182_ );
nand ( new_n16187_, new_n16183_, new_n138_ );
and  ( new_n16188_, new_n16187_, RI2b1c4342ba28_8 );
or   ( new_n16189_, new_n16188_, new_n16182_ );
or   ( new_n16190_, new_n16180_, new_n689_ );
or   ( new_n16191_, new_n16190_, new_n16184_ );
or   ( new_n16192_, new_n16184_, new_n16003_ );
or   ( new_n16193_, new_n16188_, new_n16018_ );
and  ( new_n16194_, new_n16193_, new_n16192_ );
and  ( new_n16195_, new_n16194_, new_n16191_ );
and  ( new_n16196_, new_n16195_, new_n16189_ );
and  ( new_n16197_, new_n16196_, RI2b1c4342d738_70 );
or   ( new_n16198_, new_n16188_, new_n16003_ );
and  ( new_n16199_, new_n16198_, new_n16185_ );
and  ( new_n16200_, new_n16199_, RI2b1c4342d6c0_69 );
or   ( new_n16201_, new_n16200_, new_n16197_ );
or   ( new_n16202_, new_n16201_, new_n16186_ );
and  ( new_n16203_, new_n16188_, new_n16003_ );
or   ( new_n16204_, new_n16203_, new_n16190_ );
or   ( new_n16205_, new_n16190_, new_n16188_ );
or   ( new_n16206_, new_n16184_, new_n16182_ );
and  ( new_n16207_, new_n16206_, new_n16205_ );
or   ( new_n16208_, new_n16207_, new_n16199_ );
or   ( new_n16209_, new_n16208_, new_n755_ );
or   ( new_n16210_, new_n16194_, new_n591_ );
and  ( new_n16211_, new_n16210_, new_n16209_ );
or   ( new_n16212_, new_n16211_, new_n16204_ );
and  ( new_n16213_, new_n16212_, new_n16202_ );
xor  ( new_n16214_, new_n728_, new_n646_ );
or   ( new_n16215_, new_n16214_, new_n696_ );
or   ( new_n16216_, new_n16215_, new_n16190_ );
and  ( new_n16217_, new_n16216_, new_n16157_ );
nand ( new_n16218_, new_n16214_, new_n138_ );
and  ( new_n16219_, new_n16218_, RI2b1c4342b938_6 );
or   ( new_n16220_, new_n16219_, new_n16157_ );
or   ( new_n16221_, new_n16215_, new_n16147_ );
or   ( new_n16222_, new_n16215_, new_n16182_ );
or   ( new_n16223_, new_n16219_, new_n16190_ );
and  ( new_n16224_, new_n16223_, new_n16222_ );
and  ( new_n16225_, new_n16224_, new_n16221_ );
and  ( new_n16226_, new_n16225_, new_n16220_ );
and  ( new_n16227_, new_n16226_, RI2b1c4342d828_72 );
or   ( new_n16228_, new_n16219_, new_n16182_ );
and  ( new_n16229_, new_n16228_, new_n16216_ );
and  ( new_n16230_, new_n16229_, RI2b1c4342d7b0_71 );
or   ( new_n16231_, new_n16230_, new_n16227_ );
or   ( new_n16232_, new_n16231_, new_n16217_ );
and  ( new_n16233_, new_n16219_, new_n16182_ );
or   ( new_n16234_, new_n16233_, new_n16147_ );
or   ( new_n16235_, new_n16219_, new_n16147_ );
or   ( new_n16236_, new_n16215_, new_n16157_ );
and  ( new_n16237_, new_n16236_, new_n16235_ );
or   ( new_n16238_, new_n16237_, new_n16229_ );
or   ( new_n16239_, new_n16238_, new_n806_ );
or   ( new_n16240_, new_n16224_, new_n110_ );
and  ( new_n16241_, new_n16240_, new_n16239_ );
or   ( new_n16242_, new_n16241_, new_n16234_ );
and  ( new_n16243_, new_n16242_, new_n16232_ );
or   ( new_n16244_, new_n16243_, new_n16213_ );
or   ( new_n16245_, new_n16211_, new_n16186_ );
or   ( new_n16246_, new_n16204_, new_n16201_ );
and  ( new_n16247_, new_n16246_, new_n16245_ );
or   ( new_n16248_, new_n16241_, new_n16217_ );
or   ( new_n16249_, new_n16234_, new_n16231_ );
and  ( new_n16250_, new_n16249_, new_n16248_ );
or   ( new_n16251_, new_n16250_, new_n16247_ );
and  ( new_n16252_, new_n16251_, new_n16244_ );
or   ( new_n16253_, new_n16252_, new_n16179_ );
or   ( new_n16254_, new_n16177_, new_n16151_ );
or   ( new_n16255_, new_n16170_, new_n16167_ );
and  ( new_n16256_, new_n16255_, new_n16254_ );
or   ( new_n16257_, new_n16247_, new_n16243_ );
or   ( new_n16258_, new_n16250_, new_n16213_ );
and  ( new_n16259_, new_n16258_, new_n16257_ );
or   ( new_n16260_, new_n16259_, new_n16256_ );
and  ( new_n16261_, new_n16260_, new_n16253_ );
or   ( new_n16262_, new_n16261_, new_n16145_ );
or   ( new_n16263_, new_n16143_, new_n16137_ );
or   ( new_n16264_, new_n16142_, new_n16138_ );
and  ( new_n16265_, new_n16264_, new_n16263_ );
or   ( new_n16266_, new_n16259_, new_n16179_ );
or   ( new_n16267_, new_n16256_, new_n16252_ );
and  ( new_n16268_, new_n16267_, new_n16266_ );
or   ( new_n16269_, new_n16268_, new_n16265_ );
and  ( new_n16270_, new_n16269_, new_n16262_ );
or   ( new_n16271_, new_n16270_, new_n16099_ );
or   ( new_n16272_, new_n16097_, new_n16038_ );
or   ( new_n16273_, new_n16094_, new_n16090_ );
and  ( new_n16274_, new_n16273_, new_n16272_ );
or   ( new_n16275_, new_n16265_, new_n16261_ );
or   ( new_n16276_, new_n16268_, new_n16145_ );
and  ( new_n16277_, new_n16276_, new_n16275_ );
or   ( new_n16278_, new_n16277_, new_n16274_ );
and  ( new_n16279_, new_n16278_, new_n16271_ );
and  ( new_n16280_, new_n16102_, RI2b1c4342daf8_78 );
or   ( new_n16281_, new_n16119_, new_n1004_ );
or   ( new_n16282_, new_n16123_, new_n886_ );
and  ( new_n16283_, new_n16282_, new_n16281_ );
or   ( new_n16284_, new_n16283_, new_n16108_ );
and  ( new_n16285_, new_n16132_, RI2b1c4342da80_77 );
and  ( new_n16286_, new_n16114_, RI2b1c4342da08_76 );
or   ( new_n16287_, new_n16286_, new_n16285_ );
or   ( new_n16288_, new_n16287_, new_n16128_ );
and  ( new_n16289_, new_n16288_, new_n16284_ );
or   ( new_n16290_, new_n16289_, new_n16280_ );
or   ( new_n16291_, new_n16287_, new_n16108_ );
or   ( new_n16292_, new_n16283_, new_n16128_ );
and  ( new_n16293_, new_n16292_, new_n16291_ );
or   ( new_n16294_, new_n16115_, new_n1002_ );
or   ( new_n16295_, new_n16294_, new_n16293_ );
and  ( new_n16296_, new_n16295_, new_n16290_ );
and  ( new_n16297_, new_n16162_, RI2b1c4342d990_75 );
and  ( new_n16298_, new_n16165_, RI2b1c4342d918_74 );
or   ( new_n16299_, new_n16298_, new_n16297_ );
or   ( new_n16300_, new_n16299_, new_n16151_ );
or   ( new_n16301_, new_n16174_, new_n843_ );
or   ( new_n16302_, new_n16160_, new_n859_ );
and  ( new_n16303_, new_n16302_, new_n16301_ );
or   ( new_n16304_, new_n16303_, new_n16170_ );
and  ( new_n16305_, new_n16304_, new_n16300_ );
and  ( new_n16306_, new_n16196_, RI2b1c4342d7b0_71 );
and  ( new_n16307_, new_n16199_, RI2b1c4342d738_70 );
or   ( new_n16308_, new_n16307_, new_n16306_ );
or   ( new_n16309_, new_n16308_, new_n16186_ );
or   ( new_n16310_, new_n16208_, new_n110_ );
or   ( new_n16311_, new_n16194_, new_n755_ );
and  ( new_n16312_, new_n16311_, new_n16310_ );
or   ( new_n16313_, new_n16312_, new_n16204_ );
and  ( new_n16314_, new_n16313_, new_n16309_ );
and  ( new_n16315_, new_n16226_, RI2b1c4342d8a0_73 );
and  ( new_n16316_, new_n16229_, RI2b1c4342d828_72 );
or   ( new_n16317_, new_n16316_, new_n16315_ );
or   ( new_n16318_, new_n16317_, new_n16217_ );
or   ( new_n16319_, new_n16238_, new_n105_ );
or   ( new_n16320_, new_n16224_, new_n806_ );
and  ( new_n16321_, new_n16320_, new_n16319_ );
or   ( new_n16322_, new_n16321_, new_n16234_ );
and  ( new_n16323_, new_n16322_, new_n16318_ );
or   ( new_n16324_, new_n16323_, new_n16314_ );
or   ( new_n16325_, new_n16312_, new_n16186_ );
or   ( new_n16326_, new_n16308_, new_n16204_ );
and  ( new_n16327_, new_n16326_, new_n16325_ );
or   ( new_n16328_, new_n16321_, new_n16217_ );
or   ( new_n16329_, new_n16317_, new_n16234_ );
and  ( new_n16330_, new_n16329_, new_n16328_ );
or   ( new_n16331_, new_n16330_, new_n16327_ );
and  ( new_n16332_, new_n16331_, new_n16324_ );
or   ( new_n16333_, new_n16332_, new_n16305_ );
or   ( new_n16334_, new_n16303_, new_n16151_ );
or   ( new_n16335_, new_n16299_, new_n16170_ );
and  ( new_n16336_, new_n16335_, new_n16334_ );
or   ( new_n16337_, new_n16327_, new_n16323_ );
or   ( new_n16338_, new_n16330_, new_n16314_ );
and  ( new_n16339_, new_n16338_, new_n16337_ );
or   ( new_n16340_, new_n16339_, new_n16336_ );
and  ( new_n16341_, new_n16340_, new_n16333_ );
or   ( new_n16342_, new_n16341_, new_n16296_ );
and  ( new_n16343_, new_n16021_, RI2b1c4342d6c0_69 );
and  ( new_n16344_, new_n16024_, RI2b1c4342d648_68 );
or   ( new_n16345_, new_n16344_, new_n16343_ );
or   ( new_n16346_, new_n16345_, new_n16009_ );
or   ( new_n16347_, new_n16033_, new_n591_ );
or   ( new_n16348_, new_n16017_, new_n612_ );
and  ( new_n16349_, new_n16348_, new_n16347_ );
or   ( new_n16350_, new_n16349_, new_n16029_ );
and  ( new_n16351_, new_n16350_, new_n16346_ );
or   ( new_n16352_, new_n16057_, new_n16046_ );
or   ( new_n16353_, new_n16083_, new_n16043_ );
or   ( new_n16354_, new_n16082_, new_n16046_ );
and  ( new_n16355_, new_n16354_, new_n16353_ );
or   ( new_n16356_, new_n16083_, new_n16040_ );
and  ( new_n16357_, new_n16356_, new_n16355_ );
and  ( new_n16358_, new_n16357_, new_n16352_ );
and  ( new_n16359_, new_n16358_, RI2b1c4342d4e0_65 );
or   ( new_n16360_, new_n16359_, new_n16085_ );
or   ( new_n16361_, new_n16046_, new_n16043_ );
and  ( new_n16362_, new_n16361_, new_n16084_ );
or   ( new_n16363_, new_n16046_, new_n16040_ );
or   ( new_n16364_, new_n16083_, new_n16057_ );
and  ( new_n16365_, new_n16364_, new_n16363_ );
or   ( new_n16366_, new_n16365_, new_n16362_ );
or   ( new_n16367_, new_n16366_, new_n99_ );
or   ( new_n16368_, new_n16367_, new_n16048_ );
and  ( new_n16369_, new_n16368_, new_n16360_ );
and  ( new_n16370_, new_n16063_, RI2b1c4342d5d0_67 );
and  ( new_n16371_, new_n16066_, RI2b1c4342d558_66 );
or   ( new_n16372_, new_n16371_, new_n16370_ );
or   ( new_n16373_, new_n16372_, new_n16052_ );
or   ( new_n16374_, new_n16075_, new_n112_ );
or   ( new_n16375_, new_n16060_, new_n526_ );
and  ( new_n16376_, new_n16375_, new_n16374_ );
or   ( new_n16377_, new_n16376_, new_n16071_ );
and  ( new_n16378_, new_n16377_, new_n16373_ );
or   ( new_n16379_, new_n16378_, new_n16369_ );
or   ( new_n16380_, new_n16367_, new_n16085_ );
or   ( new_n16381_, new_n16359_, new_n16048_ );
and  ( new_n16382_, new_n16381_, new_n16380_ );
or   ( new_n16383_, new_n16376_, new_n16052_ );
or   ( new_n16384_, new_n16372_, new_n16071_ );
and  ( new_n16385_, new_n16384_, new_n16383_ );
or   ( new_n16386_, new_n16385_, new_n16382_ );
and  ( new_n16387_, new_n16386_, new_n16379_ );
or   ( new_n16388_, new_n16387_, new_n16351_ );
or   ( new_n16389_, new_n16349_, new_n16009_ );
or   ( new_n16390_, new_n16345_, new_n16029_ );
and  ( new_n16391_, new_n16390_, new_n16389_ );
or   ( new_n16392_, new_n16382_, new_n16378_ );
or   ( new_n16393_, new_n16385_, new_n16369_ );
and  ( new_n16394_, new_n16393_, new_n16392_ );
or   ( new_n16395_, new_n16394_, new_n16391_ );
and  ( new_n16396_, new_n16395_, new_n16388_ );
and  ( new_n16397_, new_n16341_, new_n16296_ );
or   ( new_n16398_, new_n16397_, new_n16396_ );
and  ( new_n16399_, new_n16398_, new_n16342_ );
and  ( new_n16400_, new_n16021_, RI2b1c4342d738_70 );
and  ( new_n16401_, new_n16024_, RI2b1c4342d6c0_69 );
or   ( new_n16402_, new_n16401_, new_n16400_ );
or   ( new_n16403_, new_n16402_, new_n16009_ );
or   ( new_n16404_, new_n16033_, new_n755_ );
or   ( new_n16405_, new_n16017_, new_n591_ );
and  ( new_n16406_, new_n16405_, new_n16404_ );
or   ( new_n16407_, new_n16406_, new_n16029_ );
and  ( new_n16408_, new_n16407_, new_n16403_ );
and  ( new_n16409_, new_n16196_, RI2b1c4342d828_72 );
and  ( new_n16410_, new_n16199_, RI2b1c4342d7b0_71 );
or   ( new_n16411_, new_n16410_, new_n16409_ );
or   ( new_n16412_, new_n16411_, new_n16186_ );
or   ( new_n16413_, new_n16208_, new_n806_ );
or   ( new_n16414_, new_n16194_, new_n110_ );
and  ( new_n16415_, new_n16414_, new_n16413_ );
or   ( new_n16416_, new_n16415_, new_n16204_ );
and  ( new_n16417_, new_n16416_, new_n16412_ );
or   ( new_n16418_, new_n16417_, new_n16408_ );
and  ( new_n16419_, new_n16226_, RI2b1c4342d918_74 );
and  ( new_n16420_, new_n16229_, RI2b1c4342d8a0_73 );
or   ( new_n16421_, new_n16420_, new_n16419_ );
or   ( new_n16422_, new_n16421_, new_n16217_ );
or   ( new_n16423_, new_n16238_, new_n859_ );
or   ( new_n16424_, new_n16224_, new_n105_ );
and  ( new_n16425_, new_n16424_, new_n16423_ );
or   ( new_n16426_, new_n16425_, new_n16234_ );
and  ( new_n16427_, new_n16426_, new_n16422_ );
and  ( new_n16428_, new_n16417_, new_n16408_ );
or   ( new_n16429_, new_n16428_, new_n16427_ );
and  ( new_n16430_, new_n16429_, new_n16418_ );
xor  ( new_n16431_, new_n1345_, new_n246_ );
nand ( new_n16432_, new_n16431_, new_n138_ );
and  ( new_n16433_, new_n16432_, RI2b1c4342be60_17 );
xor  ( new_n16434_, new_n1261_, new_n248_ );
nand ( new_n16435_, new_n16434_, new_n138_ );
and  ( new_n16436_, new_n16435_, RI2b1c4342bde8_16 );
and  ( new_n16437_, new_n16436_, new_n16433_ );
or   ( new_n16438_, new_n16437_, new_n16082_ );
and  ( new_n16439_, new_n16358_, RI2b1c4342d558_66 );
and  ( new_n16440_, new_n16362_, RI2b1c4342d4e0_65 );
or   ( new_n16441_, new_n16440_, new_n16439_ );
or   ( new_n16442_, new_n16441_, new_n16085_ );
or   ( new_n16443_, new_n16366_, new_n526_ );
or   ( new_n16444_, new_n16355_, new_n99_ );
and  ( new_n16445_, new_n16444_, new_n16443_ );
or   ( new_n16446_, new_n16445_, new_n16048_ );
and  ( new_n16447_, new_n16446_, new_n16442_ );
or   ( new_n16448_, new_n16447_, new_n16438_ );
and  ( new_n16449_, new_n16063_, RI2b1c4342d648_68 );
and  ( new_n16450_, new_n16066_, RI2b1c4342d5d0_67 );
or   ( new_n16451_, new_n16450_, new_n16449_ );
or   ( new_n16452_, new_n16451_, new_n16052_ );
or   ( new_n16453_, new_n16075_, new_n612_ );
or   ( new_n16454_, new_n16060_, new_n112_ );
and  ( new_n16455_, new_n16454_, new_n16453_ );
or   ( new_n16456_, new_n16455_, new_n16071_ );
and  ( new_n16457_, new_n16456_, new_n16452_ );
and  ( new_n16458_, new_n16447_, new_n16438_ );
or   ( new_n16459_, new_n16458_, new_n16457_ );
and  ( new_n16460_, new_n16459_, new_n16448_ );
or   ( new_n16461_, new_n16460_, new_n16430_ );
and  ( new_n16462_, new_n16460_, new_n16430_ );
and  ( new_n16463_, new_n16162_, RI2b1c4342da08_76 );
and  ( new_n16464_, new_n16165_, RI2b1c4342d990_75 );
or   ( new_n16465_, new_n16464_, new_n16463_ );
or   ( new_n16466_, new_n16465_, new_n16151_ );
or   ( new_n16467_, new_n16174_, new_n886_ );
or   ( new_n16468_, new_n16160_, new_n843_ );
and  ( new_n16469_, new_n16468_, new_n16467_ );
or   ( new_n16470_, new_n16469_, new_n16170_ );
and  ( new_n16471_, new_n16470_, new_n16466_ );
and  ( new_n16472_, new_n16132_, RI2b1c4342daf8_78 );
and  ( new_n16473_, new_n16114_, RI2b1c4342da80_77 );
or   ( new_n16474_, new_n16473_, new_n16472_ );
or   ( new_n16475_, new_n16474_, new_n16108_ );
or   ( new_n16476_, new_n16119_, new_n1002_ );
or   ( new_n16477_, new_n16123_, new_n1004_ );
and  ( new_n16478_, new_n16477_, new_n16476_ );
or   ( new_n16479_, new_n16478_, new_n16128_ );
and  ( new_n16480_, new_n16479_, new_n16475_ );
or   ( new_n16481_, new_n16480_, new_n16471_ );
and  ( new_n16482_, new_n16102_, RI2b1c4342db70_79 );
and  ( new_n16483_, new_n16480_, new_n16471_ );
or   ( new_n16484_, new_n16483_, new_n16482_ );
and  ( new_n16485_, new_n16484_, new_n16481_ );
or   ( new_n16486_, new_n16485_, new_n16462_ );
and  ( new_n16487_, new_n16486_, new_n16461_ );
or   ( new_n16488_, new_n16487_, new_n16399_ );
or   ( new_n16489_, new_n16293_, new_n16280_ );
or   ( new_n16490_, new_n16294_, new_n16289_ );
and  ( new_n16491_, new_n16490_, new_n16489_ );
or   ( new_n16492_, new_n16339_, new_n16305_ );
or   ( new_n16493_, new_n16336_, new_n16332_ );
and  ( new_n16494_, new_n16493_, new_n16492_ );
or   ( new_n16495_, new_n16494_, new_n16491_ );
or   ( new_n16496_, new_n16394_, new_n16351_ );
or   ( new_n16497_, new_n16391_, new_n16387_ );
and  ( new_n16498_, new_n16497_, new_n16496_ );
and  ( new_n16499_, new_n16494_, new_n16491_ );
or   ( new_n16500_, new_n16499_, new_n16498_ );
and  ( new_n16501_, new_n16500_, new_n16495_ );
or   ( new_n16502_, new_n16431_, new_n274_ );
or   ( new_n16503_, new_n16434_, new_n271_ );
or   ( new_n16504_, new_n16503_, new_n16502_ );
and  ( new_n16505_, new_n16504_, new_n16043_ );
or   ( new_n16506_, new_n16445_, new_n16085_ );
or   ( new_n16507_, new_n16441_, new_n16048_ );
and  ( new_n16508_, new_n16507_, new_n16506_ );
or   ( new_n16509_, new_n16508_, new_n16505_ );
or   ( new_n16510_, new_n16455_, new_n16052_ );
or   ( new_n16511_, new_n16451_, new_n16071_ );
and  ( new_n16512_, new_n16511_, new_n16510_ );
and  ( new_n16513_, new_n16508_, new_n16505_ );
or   ( new_n16514_, new_n16513_, new_n16512_ );
and  ( new_n16515_, new_n16514_, new_n16509_ );
or   ( new_n16516_, new_n16406_, new_n16009_ );
or   ( new_n16517_, new_n16402_, new_n16029_ );
and  ( new_n16518_, new_n16517_, new_n16516_ );
or   ( new_n16519_, new_n16415_, new_n16186_ );
or   ( new_n16520_, new_n16411_, new_n16204_ );
and  ( new_n16521_, new_n16520_, new_n16519_ );
or   ( new_n16522_, new_n16521_, new_n16518_ );
or   ( new_n16523_, new_n16425_, new_n16217_ );
or   ( new_n16524_, new_n16421_, new_n16234_ );
and  ( new_n16525_, new_n16524_, new_n16523_ );
and  ( new_n16526_, new_n16521_, new_n16518_ );
or   ( new_n16527_, new_n16526_, new_n16525_ );
and  ( new_n16528_, new_n16527_, new_n16522_ );
and  ( new_n16529_, new_n16528_, new_n16515_ );
or   ( new_n16530_, new_n16528_, new_n16515_ );
or   ( new_n16531_, new_n16469_, new_n16151_ );
or   ( new_n16532_, new_n16465_, new_n16170_ );
and  ( new_n16533_, new_n16532_, new_n16531_ );
or   ( new_n16534_, new_n16478_, new_n16108_ );
or   ( new_n16535_, new_n16474_, new_n16128_ );
and  ( new_n16536_, new_n16535_, new_n16534_ );
and  ( new_n16537_, new_n16536_, new_n16533_ );
or   ( new_n16538_, new_n16536_, new_n16533_ );
or   ( new_n16539_, new_n16115_, new_n1310_ );
and  ( new_n16540_, new_n16539_, new_n16538_ );
or   ( new_n16541_, new_n16540_, new_n16537_ );
and  ( new_n16542_, new_n16541_, new_n16530_ );
or   ( new_n16543_, new_n16542_, new_n16529_ );
or   ( new_n16544_, new_n16543_, new_n16501_ );
and  ( new_n16545_, new_n16544_, new_n16488_ );
or   ( new_n16546_, new_n16545_, new_n16279_ );
or   ( new_n16547_, new_n16277_, new_n16099_ );
or   ( new_n16548_, new_n16274_, new_n16270_ );
and  ( new_n16549_, new_n16548_, new_n16547_ );
or   ( new_n16550_, new_n16543_, new_n16399_ );
or   ( new_n16551_, new_n16501_, new_n16487_ );
and  ( new_n16552_, new_n16551_, new_n16550_ );
or   ( new_n16553_, new_n16552_, new_n16549_ );
and  ( new_n16554_, new_n16553_, new_n16546_ );
and  ( new_n16555_, new_n16378_, new_n16369_ );
or   ( new_n16556_, new_n16555_, new_n16351_ );
and  ( new_n16557_, new_n16556_, new_n16379_ );
and  ( new_n16558_, new_n16323_, new_n16314_ );
or   ( new_n16559_, new_n16558_, new_n16305_ );
and  ( new_n16560_, new_n16559_, new_n16324_ );
or   ( new_n16561_, new_n16560_, new_n16557_ );
and  ( new_n16562_, new_n16385_, new_n16382_ );
or   ( new_n16563_, new_n16562_, new_n16391_ );
and  ( new_n16564_, new_n16563_, new_n16386_ );
and  ( new_n16565_, new_n16330_, new_n16327_ );
or   ( new_n16566_, new_n16565_, new_n16336_ );
and  ( new_n16567_, new_n16566_, new_n16331_ );
or   ( new_n16568_, new_n16567_, new_n16564_ );
and  ( new_n16569_, new_n16568_, new_n16561_ );
or   ( new_n16570_, new_n16569_, new_n16489_ );
and  ( new_n16571_, new_n16294_, new_n16289_ );
or   ( new_n16572_, new_n16564_, new_n16560_ );
or   ( new_n16573_, new_n16567_, new_n16557_ );
and  ( new_n16574_, new_n16573_, new_n16572_ );
or   ( new_n16575_, new_n16574_, new_n16571_ );
and  ( new_n16576_, new_n16575_, new_n16570_ );
or   ( new_n16577_, new_n16533_, new_n16480_ );
or   ( new_n16578_, new_n16536_, new_n16471_ );
and  ( new_n16579_, new_n16578_, new_n16577_ );
or   ( new_n16580_, new_n16579_, new_n16482_ );
and  ( new_n16581_, new_n16538_, new_n16481_ );
or   ( new_n16582_, new_n16581_, new_n16539_ );
and  ( new_n16583_, new_n16582_, new_n16580_ );
or   ( new_n16584_, new_n16518_, new_n16417_ );
or   ( new_n16585_, new_n16521_, new_n16408_ );
and  ( new_n16586_, new_n16585_, new_n16584_ );
or   ( new_n16587_, new_n16586_, new_n16427_ );
and  ( new_n16588_, new_n16522_, new_n16418_ );
or   ( new_n16589_, new_n16588_, new_n16525_ );
and  ( new_n16590_, new_n16589_, new_n16587_ );
or   ( new_n16591_, new_n16590_, new_n16583_ );
or   ( new_n16592_, new_n16505_, new_n16447_ );
or   ( new_n16593_, new_n16508_, new_n16438_ );
and  ( new_n16594_, new_n16593_, new_n16592_ );
or   ( new_n16595_, new_n16594_, new_n16457_ );
and  ( new_n16596_, new_n16509_, new_n16448_ );
or   ( new_n16597_, new_n16596_, new_n16512_ );
and  ( new_n16598_, new_n16597_, new_n16595_ );
and  ( new_n16599_, new_n16590_, new_n16583_ );
or   ( new_n16600_, new_n16599_, new_n16598_ );
and  ( new_n16601_, new_n16600_, new_n16591_ );
or   ( new_n16602_, new_n16436_, new_n16433_ );
and  ( new_n16603_, new_n16602_, new_n16504_ );
or   ( new_n16604_, new_n16436_, new_n16082_ );
or   ( new_n16605_, new_n16503_, new_n16043_ );
and  ( new_n16606_, new_n16605_, new_n16604_ );
or   ( new_n16607_, new_n16606_, new_n16603_ );
or   ( new_n16608_, new_n16607_, new_n99_ );
or   ( new_n16609_, new_n16608_, new_n16505_ );
or   ( new_n16610_, new_n16436_, new_n16043_ );
or   ( new_n16611_, new_n16503_, new_n16433_ );
or   ( new_n16612_, new_n16502_, new_n16436_ );
and  ( new_n16613_, new_n16612_, new_n16611_ );
or   ( new_n16614_, new_n16503_, new_n16082_ );
and  ( new_n16615_, new_n16614_, new_n16613_ );
and  ( new_n16616_, new_n16615_, new_n16610_ );
and  ( new_n16617_, new_n16616_, RI2b1c4342d4e0_65 );
or   ( new_n16618_, new_n16617_, new_n16438_ );
and  ( new_n16619_, new_n16618_, new_n16609_ );
or   ( new_n16620_, new_n16366_, new_n112_ );
or   ( new_n16621_, new_n16355_, new_n526_ );
and  ( new_n16622_, new_n16621_, new_n16620_ );
or   ( new_n16623_, new_n16622_, new_n16085_ );
and  ( new_n16624_, new_n16358_, RI2b1c4342d5d0_67 );
and  ( new_n16625_, new_n16362_, RI2b1c4342d558_66 );
or   ( new_n16626_, new_n16625_, new_n16624_ );
or   ( new_n16627_, new_n16626_, new_n16048_ );
and  ( new_n16628_, new_n16627_, new_n16623_ );
or   ( new_n16629_, new_n16628_, new_n16619_ );
and  ( new_n16630_, new_n16628_, new_n16619_ );
or   ( new_n16631_, new_n16075_, new_n591_ );
or   ( new_n16632_, new_n16060_, new_n612_ );
and  ( new_n16633_, new_n16632_, new_n16631_ );
or   ( new_n16634_, new_n16633_, new_n16052_ );
and  ( new_n16635_, new_n16063_, RI2b1c4342d6c0_69 );
and  ( new_n16636_, new_n16066_, RI2b1c4342d648_68 );
or   ( new_n16637_, new_n16636_, new_n16635_ );
or   ( new_n16638_, new_n16637_, new_n16071_ );
and  ( new_n16639_, new_n16638_, new_n16634_ );
or   ( new_n16640_, new_n16639_, new_n16630_ );
and  ( new_n16641_, new_n16640_, new_n16629_ );
or   ( new_n16642_, new_n16033_, new_n110_ );
or   ( new_n16643_, new_n16017_, new_n755_ );
and  ( new_n16644_, new_n16643_, new_n16642_ );
or   ( new_n16645_, new_n16644_, new_n16009_ );
and  ( new_n16646_, new_n16021_, RI2b1c4342d7b0_71 );
and  ( new_n16647_, new_n16024_, RI2b1c4342d738_70 );
or   ( new_n16648_, new_n16647_, new_n16646_ );
or   ( new_n16649_, new_n16648_, new_n16029_ );
and  ( new_n16650_, new_n16649_, new_n16645_ );
or   ( new_n16651_, new_n16208_, new_n105_ );
or   ( new_n16652_, new_n16194_, new_n806_ );
and  ( new_n16653_, new_n16652_, new_n16651_ );
or   ( new_n16654_, new_n16653_, new_n16186_ );
and  ( new_n16655_, new_n16196_, RI2b1c4342d8a0_73 );
and  ( new_n16656_, new_n16199_, RI2b1c4342d828_72 );
or   ( new_n16657_, new_n16656_, new_n16655_ );
or   ( new_n16658_, new_n16657_, new_n16204_ );
and  ( new_n16659_, new_n16658_, new_n16654_ );
or   ( new_n16660_, new_n16659_, new_n16650_ );
and  ( new_n16661_, new_n16659_, new_n16650_ );
or   ( new_n16662_, new_n16238_, new_n843_ );
or   ( new_n16663_, new_n16224_, new_n859_ );
and  ( new_n16664_, new_n16663_, new_n16662_ );
or   ( new_n16665_, new_n16664_, new_n16217_ );
and  ( new_n16666_, new_n16226_, RI2b1c4342d990_75 );
and  ( new_n16667_, new_n16229_, RI2b1c4342d918_74 );
or   ( new_n16668_, new_n16667_, new_n16666_ );
or   ( new_n16669_, new_n16668_, new_n16234_ );
and  ( new_n16670_, new_n16669_, new_n16665_ );
or   ( new_n16671_, new_n16670_, new_n16661_ );
and  ( new_n16672_, new_n16671_, new_n16660_ );
and  ( new_n16673_, new_n16672_, new_n16641_ );
or   ( new_n16674_, new_n16672_, new_n16641_ );
or   ( new_n16675_, new_n16174_, new_n1004_ );
or   ( new_n16676_, new_n16160_, new_n886_ );
and  ( new_n16677_, new_n16676_, new_n16675_ );
or   ( new_n16678_, new_n16677_, new_n16151_ );
and  ( new_n16679_, new_n16162_, RI2b1c4342da80_77 );
and  ( new_n16680_, new_n16165_, RI2b1c4342da08_76 );
or   ( new_n16681_, new_n16680_, new_n16679_ );
or   ( new_n16682_, new_n16681_, new_n16170_ );
and  ( new_n16683_, new_n16682_, new_n16678_ );
or   ( new_n16684_, new_n16119_, new_n1310_ );
or   ( new_n16685_, new_n16123_, new_n1002_ );
and  ( new_n16686_, new_n16685_, new_n16684_ );
or   ( new_n16687_, new_n16686_, new_n16108_ );
and  ( new_n16688_, new_n16132_, RI2b1c4342db70_79 );
and  ( new_n16689_, new_n16114_, RI2b1c4342daf8_78 );
or   ( new_n16690_, new_n16689_, new_n16688_ );
or   ( new_n16691_, new_n16690_, new_n16128_ );
and  ( new_n16692_, new_n16691_, new_n16687_ );
and  ( new_n16693_, new_n16692_, new_n16683_ );
or   ( new_n16694_, new_n16692_, new_n16683_ );
or   ( new_n16695_, new_n16115_, new_n1511_ );
and  ( new_n16696_, new_n16695_, new_n16694_ );
or   ( new_n16697_, new_n16696_, new_n16693_ );
and  ( new_n16698_, new_n16697_, new_n16674_ );
or   ( new_n16699_, new_n16698_, new_n16673_ );
and  ( new_n16700_, new_n16699_, new_n16601_ );
or   ( new_n16701_, new_n16699_, new_n16601_ );
or   ( new_n16702_, new_n16491_, new_n16341_ );
or   ( new_n16703_, new_n16494_, new_n16296_ );
and  ( new_n16704_, new_n16703_, new_n16702_ );
or   ( new_n16705_, new_n16704_, new_n16396_ );
and  ( new_n16706_, new_n16495_, new_n16342_ );
or   ( new_n16707_, new_n16706_, new_n16498_ );
and  ( new_n16708_, new_n16707_, new_n16705_ );
and  ( new_n16709_, new_n16708_, new_n16701_ );
or   ( new_n16710_, new_n16709_, new_n16700_ );
or   ( new_n16711_, new_n16710_, new_n16576_ );
or   ( new_n16712_, new_n16617_, new_n16505_ );
or   ( new_n16713_, new_n16608_, new_n16438_ );
and  ( new_n16714_, new_n16713_, new_n16712_ );
or   ( new_n16715_, new_n16626_, new_n16085_ );
or   ( new_n16716_, new_n16622_, new_n16048_ );
and  ( new_n16717_, new_n16716_, new_n16715_ );
or   ( new_n16718_, new_n16717_, new_n16714_ );
and  ( new_n16719_, new_n16717_, new_n16714_ );
or   ( new_n16720_, new_n16637_, new_n16052_ );
or   ( new_n16721_, new_n16633_, new_n16071_ );
and  ( new_n16722_, new_n16721_, new_n16720_ );
or   ( new_n16723_, new_n16722_, new_n16719_ );
and  ( new_n16724_, new_n16723_, new_n16718_ );
or   ( new_n16725_, new_n16648_, new_n16009_ );
or   ( new_n16726_, new_n16644_, new_n16029_ );
and  ( new_n16727_, new_n16726_, new_n16725_ );
or   ( new_n16728_, new_n16657_, new_n16186_ );
or   ( new_n16729_, new_n16653_, new_n16204_ );
and  ( new_n16730_, new_n16729_, new_n16728_ );
or   ( new_n16731_, new_n16730_, new_n16727_ );
and  ( new_n16732_, new_n16730_, new_n16727_ );
or   ( new_n16733_, new_n16668_, new_n16217_ );
or   ( new_n16734_, new_n16664_, new_n16234_ );
and  ( new_n16735_, new_n16734_, new_n16733_ );
or   ( new_n16736_, new_n16735_, new_n16732_ );
and  ( new_n16737_, new_n16736_, new_n16731_ );
or   ( new_n16738_, new_n16737_, new_n16724_ );
and  ( new_n16739_, new_n16737_, new_n16724_ );
or   ( new_n16740_, new_n16690_, new_n16108_ );
or   ( new_n16741_, new_n16686_, new_n16128_ );
and  ( new_n16742_, new_n16741_, new_n16740_ );
or   ( new_n16743_, new_n16681_, new_n16151_ );
or   ( new_n16744_, new_n16677_, new_n16170_ );
and  ( new_n16745_, new_n16744_, new_n16743_ );
or   ( new_n16746_, new_n16745_, new_n16742_ );
and  ( new_n16747_, new_n16745_, new_n16742_ );
and  ( new_n16748_, new_n16102_, RI2b1c4342dbe8_80 );
or   ( new_n16749_, new_n16748_, new_n16747_ );
and  ( new_n16750_, new_n16749_, new_n16746_ );
or   ( new_n16751_, new_n16750_, new_n16739_ );
and  ( new_n16752_, new_n16751_, new_n16738_ );
or   ( new_n16753_, new_n16581_, new_n16482_ );
or   ( new_n16754_, new_n16579_, new_n16539_ );
and  ( new_n16755_, new_n16754_, new_n16753_ );
or   ( new_n16756_, new_n16588_, new_n16427_ );
or   ( new_n16757_, new_n16586_, new_n16525_ );
and  ( new_n16758_, new_n16757_, new_n16756_ );
or   ( new_n16759_, new_n16758_, new_n16755_ );
or   ( new_n16760_, new_n16596_, new_n16457_ );
or   ( new_n16761_, new_n16594_, new_n16512_ );
and  ( new_n16762_, new_n16761_, new_n16760_ );
and  ( new_n16763_, new_n16758_, new_n16755_ );
or   ( new_n16764_, new_n16763_, new_n16762_ );
and  ( new_n16765_, new_n16764_, new_n16759_ );
or   ( new_n16766_, new_n16765_, new_n16752_ );
or   ( new_n16767_, new_n16706_, new_n16396_ );
or   ( new_n16768_, new_n16704_, new_n16498_ );
and  ( new_n16769_, new_n16768_, new_n16767_ );
and  ( new_n16770_, new_n16765_, new_n16752_ );
or   ( new_n16771_, new_n16770_, new_n16769_ );
and  ( new_n16772_, new_n16771_, new_n16766_ );
or   ( new_n16773_, new_n16574_, new_n16489_ );
or   ( new_n16774_, new_n16571_, new_n16569_ );
and  ( new_n16775_, new_n16774_, new_n16773_ );
or   ( new_n16776_, new_n16775_, new_n16772_ );
and  ( new_n16777_, new_n16776_, new_n16711_ );
or   ( new_n16778_, new_n16777_, new_n16554_ );
or   ( new_n16779_, new_n16772_, new_n16576_ );
or   ( new_n16780_, new_n16775_, new_n16710_ );
and  ( new_n16781_, new_n16780_, new_n16779_ );
or   ( new_n16782_, new_n16552_, new_n16279_ );
or   ( new_n16783_, new_n16549_, new_n16545_ );
and  ( new_n16784_, new_n16783_, new_n16782_ );
or   ( new_n16785_, new_n16784_, new_n16781_ );
and  ( new_n16786_, new_n16785_, new_n16778_ );
or   ( new_n16787_, new_n16515_, new_n16430_ );
or   ( new_n16788_, new_n16528_, new_n16460_ );
and  ( new_n16789_, new_n16788_, new_n16787_ );
or   ( new_n16790_, new_n16789_, new_n16485_ );
and  ( new_n16791_, new_n16530_, new_n16461_ );
or   ( new_n16792_, new_n16791_, new_n16541_ );
and  ( new_n16793_, new_n16792_, new_n16790_ );
or   ( new_n16794_, new_n16742_, new_n16683_ );
or   ( new_n16795_, new_n16745_, new_n16692_ );
and  ( new_n16796_, new_n16795_, new_n16794_ );
or   ( new_n16797_, new_n16796_, new_n16748_ );
and  ( new_n16798_, new_n16746_, new_n16694_ );
or   ( new_n16799_, new_n16798_, new_n16695_ );
and  ( new_n16800_, new_n16799_, new_n16797_ );
or   ( new_n16801_, new_n16730_, new_n16650_ );
or   ( new_n16802_, new_n16727_, new_n16659_ );
and  ( new_n16803_, new_n16802_, new_n16801_ );
or   ( new_n16804_, new_n16803_, new_n16735_ );
and  ( new_n16805_, new_n16731_, new_n16660_ );
or   ( new_n16806_, new_n16805_, new_n16670_ );
and  ( new_n16807_, new_n16806_, new_n16804_ );
and  ( new_n16808_, new_n16807_, new_n16800_ );
xor  ( new_n16809_, new_n1711_, new_n1813_ );
or   ( new_n16810_, new_n16809_, new_n282_ );
xor  ( new_n16811_, new_n1704_, new_n1818_ );
or   ( new_n16812_, new_n16811_, new_n279_ );
or   ( new_n16813_, new_n16812_, new_n16810_ );
and  ( new_n16814_, new_n16813_, new_n16433_ );
or   ( new_n16815_, new_n16607_, new_n526_ );
or   ( new_n16816_, new_n16613_, new_n99_ );
and  ( new_n16817_, new_n16816_, new_n16815_ );
or   ( new_n16818_, new_n16817_, new_n16505_ );
and  ( new_n16819_, new_n16616_, RI2b1c4342d558_66 );
and  ( new_n16820_, new_n16603_, RI2b1c4342d4e0_65 );
or   ( new_n16821_, new_n16820_, new_n16819_ );
or   ( new_n16822_, new_n16821_, new_n16438_ );
and  ( new_n16823_, new_n16822_, new_n16818_ );
or   ( new_n16824_, new_n16823_, new_n16814_ );
and  ( new_n16825_, new_n16823_, new_n16814_ );
or   ( new_n16826_, new_n16366_, new_n612_ );
or   ( new_n16827_, new_n16355_, new_n112_ );
and  ( new_n16828_, new_n16827_, new_n16826_ );
or   ( new_n16829_, new_n16828_, new_n16085_ );
and  ( new_n16830_, new_n16358_, RI2b1c4342d648_68 );
and  ( new_n16831_, new_n16362_, RI2b1c4342d5d0_67 );
or   ( new_n16832_, new_n16831_, new_n16830_ );
or   ( new_n16833_, new_n16832_, new_n16048_ );
and  ( new_n16834_, new_n16833_, new_n16829_ );
or   ( new_n16835_, new_n16834_, new_n16825_ );
and  ( new_n16836_, new_n16835_, new_n16824_ );
or   ( new_n16837_, new_n16075_, new_n755_ );
or   ( new_n16838_, new_n16060_, new_n591_ );
and  ( new_n16839_, new_n16838_, new_n16837_ );
or   ( new_n16840_, new_n16839_, new_n16052_ );
and  ( new_n16841_, new_n16063_, RI2b1c4342d738_70 );
and  ( new_n16842_, new_n16066_, RI2b1c4342d6c0_69 );
or   ( new_n16843_, new_n16842_, new_n16841_ );
or   ( new_n16844_, new_n16843_, new_n16071_ );
and  ( new_n16845_, new_n16844_, new_n16840_ );
or   ( new_n16846_, new_n16033_, new_n806_ );
or   ( new_n16847_, new_n16017_, new_n110_ );
and  ( new_n16848_, new_n16847_, new_n16846_ );
or   ( new_n16849_, new_n16848_, new_n16009_ );
and  ( new_n16850_, new_n16021_, RI2b1c4342d828_72 );
and  ( new_n16851_, new_n16024_, RI2b1c4342d7b0_71 );
or   ( new_n16852_, new_n16851_, new_n16850_ );
or   ( new_n16853_, new_n16852_, new_n16029_ );
and  ( new_n16854_, new_n16853_, new_n16849_ );
or   ( new_n16855_, new_n16854_, new_n16845_ );
or   ( new_n16856_, new_n16208_, new_n859_ );
or   ( new_n16857_, new_n16194_, new_n105_ );
and  ( new_n16858_, new_n16857_, new_n16856_ );
or   ( new_n16859_, new_n16858_, new_n16186_ );
and  ( new_n16860_, new_n16196_, RI2b1c4342d918_74 );
and  ( new_n16861_, new_n16199_, RI2b1c4342d8a0_73 );
or   ( new_n16862_, new_n16861_, new_n16860_ );
or   ( new_n16863_, new_n16862_, new_n16204_ );
and  ( new_n16864_, new_n16863_, new_n16859_ );
and  ( new_n16865_, new_n16854_, new_n16845_ );
or   ( new_n16866_, new_n16865_, new_n16864_ );
and  ( new_n16867_, new_n16866_, new_n16855_ );
or   ( new_n16868_, new_n16867_, new_n16836_ );
and  ( new_n16869_, new_n16867_, new_n16836_ );
or   ( new_n16870_, new_n16238_, new_n886_ );
or   ( new_n16871_, new_n16224_, new_n843_ );
and  ( new_n16872_, new_n16871_, new_n16870_ );
or   ( new_n16873_, new_n16872_, new_n16217_ );
and  ( new_n16874_, new_n16226_, RI2b1c4342da08_76 );
and  ( new_n16875_, new_n16229_, RI2b1c4342d990_75 );
or   ( new_n16876_, new_n16875_, new_n16874_ );
or   ( new_n16877_, new_n16876_, new_n16234_ );
and  ( new_n16878_, new_n16877_, new_n16873_ );
or   ( new_n16879_, new_n16174_, new_n1002_ );
or   ( new_n16880_, new_n16160_, new_n1004_ );
and  ( new_n16881_, new_n16880_, new_n16879_ );
or   ( new_n16882_, new_n16881_, new_n16151_ );
and  ( new_n16883_, new_n16162_, RI2b1c4342daf8_78 );
and  ( new_n16884_, new_n16165_, RI2b1c4342da80_77 );
or   ( new_n16885_, new_n16884_, new_n16883_ );
or   ( new_n16886_, new_n16885_, new_n16170_ );
and  ( new_n16887_, new_n16886_, new_n16882_ );
or   ( new_n16888_, new_n16887_, new_n16878_ );
or   ( new_n16889_, new_n16119_, new_n1511_ );
or   ( new_n16890_, new_n16123_, new_n1310_ );
and  ( new_n16891_, new_n16890_, new_n16889_ );
or   ( new_n16892_, new_n16891_, new_n16108_ );
and  ( new_n16893_, new_n16132_, RI2b1c4342dbe8_80 );
and  ( new_n16894_, new_n16114_, RI2b1c4342db70_79 );
or   ( new_n16895_, new_n16894_, new_n16893_ );
or   ( new_n16896_, new_n16895_, new_n16128_ );
and  ( new_n16897_, new_n16896_, new_n16892_ );
and  ( new_n16898_, new_n16887_, new_n16878_ );
or   ( new_n16899_, new_n16898_, new_n16897_ );
and  ( new_n16900_, new_n16899_, new_n16888_ );
or   ( new_n16901_, new_n16900_, new_n16869_ );
and  ( new_n16902_, new_n16901_, new_n16868_ );
or   ( new_n16903_, new_n16902_, new_n16808_ );
or   ( new_n16904_, new_n16758_, new_n16583_ );
or   ( new_n16905_, new_n16755_, new_n16590_ );
and  ( new_n16906_, new_n16905_, new_n16904_ );
or   ( new_n16907_, new_n16906_, new_n16762_ );
and  ( new_n16908_, new_n16759_, new_n16591_ );
or   ( new_n16909_, new_n16908_, new_n16598_ );
and  ( new_n16910_, new_n16909_, new_n16907_ );
and  ( new_n16911_, new_n16902_, new_n16808_ );
or   ( new_n16912_, new_n16911_, new_n16910_ );
and  ( new_n16913_, new_n16912_, new_n16903_ );
or   ( new_n16914_, new_n16913_, new_n16793_ );
or   ( new_n16915_, new_n16765_, new_n16699_ );
or   ( new_n16916_, new_n16752_, new_n16601_ );
and  ( new_n16917_, new_n16916_, new_n16915_ );
or   ( new_n16918_, new_n16917_, new_n16769_ );
and  ( new_n16919_, new_n16766_, new_n16701_ );
or   ( new_n16920_, new_n16919_, new_n16708_ );
and  ( new_n16921_, new_n16920_, new_n16918_ );
and  ( new_n16922_, new_n16913_, new_n16793_ );
or   ( new_n16923_, new_n16922_, new_n16921_ );
and  ( new_n16924_, new_n16923_, new_n16914_ );
or   ( new_n16925_, new_n16924_, new_n16786_ );
and  ( new_n16926_, new_n16196_, RI2b1c4342d6c0_69 );
and  ( new_n16927_, new_n16199_, RI2b1c4342d648_68 );
or   ( new_n16928_, new_n16927_, new_n16926_ );
or   ( new_n16929_, new_n16928_, new_n16186_ );
or   ( new_n16930_, new_n16208_, new_n591_ );
or   ( new_n16931_, new_n16194_, new_n612_ );
and  ( new_n16932_, new_n16931_, new_n16930_ );
or   ( new_n16933_, new_n16932_, new_n16204_ );
and  ( new_n16934_, new_n16933_, new_n16929_ );
and  ( new_n16935_, new_n16063_, RI2b1c4342d4e0_65 );
or   ( new_n16936_, new_n16935_, new_n16052_ );
or   ( new_n16937_, new_n16075_, new_n99_ );
or   ( new_n16938_, new_n16937_, new_n16071_ );
and  ( new_n16939_, new_n16938_, new_n16936_ );
and  ( new_n16940_, new_n16021_, RI2b1c4342d5d0_67 );
and  ( new_n16941_, new_n16024_, RI2b1c4342d558_66 );
or   ( new_n16942_, new_n16941_, new_n16940_ );
or   ( new_n16943_, new_n16942_, new_n16009_ );
or   ( new_n16944_, new_n16033_, new_n112_ );
or   ( new_n16945_, new_n16017_, new_n526_ );
and  ( new_n16946_, new_n16945_, new_n16944_ );
or   ( new_n16947_, new_n16946_, new_n16029_ );
and  ( new_n16948_, new_n16947_, new_n16943_ );
or   ( new_n16949_, new_n16948_, new_n16939_ );
or   ( new_n16950_, new_n16937_, new_n16052_ );
or   ( new_n16951_, new_n16935_, new_n16071_ );
and  ( new_n16952_, new_n16951_, new_n16950_ );
or   ( new_n16953_, new_n16946_, new_n16009_ );
or   ( new_n16954_, new_n16942_, new_n16029_ );
and  ( new_n16955_, new_n16954_, new_n16953_ );
or   ( new_n16956_, new_n16955_, new_n16952_ );
and  ( new_n16957_, new_n16956_, new_n16949_ );
or   ( new_n16958_, new_n16957_, new_n16934_ );
or   ( new_n16959_, new_n16932_, new_n16186_ );
or   ( new_n16960_, new_n16928_, new_n16204_ );
and  ( new_n16961_, new_n16960_, new_n16959_ );
or   ( new_n16962_, new_n16952_, new_n16948_ );
or   ( new_n16963_, new_n16955_, new_n16939_ );
and  ( new_n16964_, new_n16963_, new_n16962_ );
or   ( new_n16965_, new_n16964_, new_n16961_ );
and  ( new_n16966_, new_n16965_, new_n16958_ );
or   ( new_n16967_, new_n16115_, new_n886_ );
and  ( new_n16968_, new_n16132_, RI2b1c4342d990_75 );
and  ( new_n16969_, new_n16114_, RI2b1c4342d918_74 );
or   ( new_n16970_, new_n16969_, new_n16968_ );
or   ( new_n16971_, new_n16970_, new_n16108_ );
or   ( new_n16972_, new_n16119_, new_n843_ );
or   ( new_n16973_, new_n16123_, new_n859_ );
and  ( new_n16974_, new_n16973_, new_n16972_ );
or   ( new_n16975_, new_n16974_, new_n16128_ );
and  ( new_n16976_, new_n16975_, new_n16971_ );
and  ( new_n16977_, new_n16226_, RI2b1c4342d7b0_71 );
and  ( new_n16978_, new_n16229_, RI2b1c4342d738_70 );
or   ( new_n16979_, new_n16978_, new_n16977_ );
or   ( new_n16980_, new_n16979_, new_n16217_ );
or   ( new_n16981_, new_n16238_, new_n110_ );
or   ( new_n16982_, new_n16224_, new_n755_ );
and  ( new_n16983_, new_n16982_, new_n16981_ );
or   ( new_n16984_, new_n16983_, new_n16234_ );
and  ( new_n16985_, new_n16984_, new_n16980_ );
and  ( new_n16986_, new_n16162_, RI2b1c4342d8a0_73 );
and  ( new_n16987_, new_n16165_, RI2b1c4342d828_72 );
or   ( new_n16988_, new_n16987_, new_n16986_ );
or   ( new_n16989_, new_n16988_, new_n16151_ );
or   ( new_n16990_, new_n16174_, new_n105_ );
or   ( new_n16991_, new_n16160_, new_n806_ );
and  ( new_n16992_, new_n16991_, new_n16990_ );
or   ( new_n16993_, new_n16992_, new_n16170_ );
and  ( new_n16994_, new_n16993_, new_n16989_ );
or   ( new_n16995_, new_n16994_, new_n16985_ );
or   ( new_n16996_, new_n16983_, new_n16217_ );
or   ( new_n16997_, new_n16979_, new_n16234_ );
and  ( new_n16998_, new_n16997_, new_n16996_ );
or   ( new_n16999_, new_n16992_, new_n16151_ );
or   ( new_n17000_, new_n16988_, new_n16170_ );
and  ( new_n17001_, new_n17000_, new_n16999_ );
or   ( new_n17002_, new_n17001_, new_n16998_ );
and  ( new_n17003_, new_n17002_, new_n16995_ );
or   ( new_n17004_, new_n17003_, new_n16976_ );
or   ( new_n17005_, new_n16974_, new_n16108_ );
or   ( new_n17006_, new_n16970_, new_n16128_ );
and  ( new_n17007_, new_n17006_, new_n17005_ );
or   ( new_n17008_, new_n16998_, new_n16994_ );
or   ( new_n17009_, new_n17001_, new_n16985_ );
and  ( new_n17010_, new_n17009_, new_n17008_ );
or   ( new_n17011_, new_n17010_, new_n17007_ );
and  ( new_n17012_, new_n17011_, new_n17004_ );
or   ( new_n17013_, new_n17012_, new_n16967_ );
and  ( new_n17014_, new_n16102_, RI2b1c4342da08_76 );
or   ( new_n17015_, new_n17010_, new_n16976_ );
or   ( new_n17016_, new_n17007_, new_n17003_ );
and  ( new_n17017_, new_n17016_, new_n17015_ );
or   ( new_n17018_, new_n17017_, new_n17014_ );
and  ( new_n17019_, new_n17018_, new_n17013_ );
or   ( new_n17020_, new_n17019_, new_n16966_ );
or   ( new_n17021_, new_n16964_, new_n16934_ );
or   ( new_n17022_, new_n16961_, new_n16957_ );
and  ( new_n17023_, new_n17022_, new_n17021_ );
or   ( new_n17024_, new_n17014_, new_n17012_ );
or   ( new_n17025_, new_n17017_, new_n16967_ );
and  ( new_n17026_, new_n17025_, new_n17024_ );
or   ( new_n17027_, new_n17026_, new_n17023_ );
and  ( new_n17028_, new_n17027_, new_n17020_ );
and  ( new_n17029_, new_n16560_, new_n16557_ );
or   ( new_n17030_, new_n17029_, new_n16489_ );
and  ( new_n17031_, new_n17030_, new_n16561_ );
and  ( new_n17032_, new_n16261_, new_n16145_ );
or   ( new_n17033_, new_n17032_, new_n16099_ );
and  ( new_n17034_, new_n17033_, new_n16262_ );
or   ( new_n17035_, new_n17034_, new_n17031_ );
and  ( new_n17036_, new_n16567_, new_n16564_ );
or   ( new_n17037_, new_n17036_, new_n16571_ );
and  ( new_n17038_, new_n17037_, new_n16568_ );
and  ( new_n17039_, new_n16268_, new_n16265_ );
or   ( new_n17040_, new_n17039_, new_n16274_ );
and  ( new_n17041_, new_n17040_, new_n16269_ );
or   ( new_n17042_, new_n17041_, new_n17038_ );
and  ( new_n17043_, new_n17042_, new_n17035_ );
or   ( new_n17044_, new_n17043_, new_n17028_ );
or   ( new_n17045_, new_n17026_, new_n16966_ );
or   ( new_n17046_, new_n17023_, new_n17019_ );
and  ( new_n17047_, new_n17046_, new_n17045_ );
or   ( new_n17048_, new_n17038_, new_n17034_ );
or   ( new_n17049_, new_n17041_, new_n17031_ );
and  ( new_n17050_, new_n17049_, new_n17048_ );
or   ( new_n17051_, new_n17050_, new_n17047_ );
and  ( new_n17052_, new_n17051_, new_n17044_ );
and  ( new_n17053_, new_n16143_, new_n16142_ );
and  ( new_n17054_, new_n16243_, new_n16213_ );
or   ( new_n17055_, new_n17054_, new_n16179_ );
and  ( new_n17056_, new_n17055_, new_n16244_ );
and  ( new_n17057_, new_n16080_, new_n16048_ );
or   ( new_n17058_, new_n17057_, new_n16038_ );
and  ( new_n17059_, new_n17058_, new_n16081_ );
or   ( new_n17060_, new_n17059_, new_n17056_ );
and  ( new_n17061_, new_n16088_, new_n16085_ );
or   ( new_n17062_, new_n17061_, new_n16094_ );
and  ( new_n17063_, new_n17062_, new_n16089_ );
and  ( new_n17064_, new_n16250_, new_n16247_ );
or   ( new_n17065_, new_n17064_, new_n16256_ );
and  ( new_n17066_, new_n17065_, new_n16251_ );
or   ( new_n17067_, new_n17066_, new_n17063_ );
and  ( new_n17068_, new_n17067_, new_n17060_ );
or   ( new_n17069_, new_n17068_, new_n17053_ );
or   ( new_n17070_, new_n17063_, new_n17056_ );
or   ( new_n17071_, new_n17066_, new_n17059_ );
and  ( new_n17072_, new_n17071_, new_n17070_ );
or   ( new_n17073_, new_n17072_, new_n16139_ );
and  ( new_n17074_, new_n17073_, new_n17069_ );
and  ( new_n17075_, new_n16487_, new_n16399_ );
or   ( new_n17076_, new_n17075_, new_n16279_ );
and  ( new_n17077_, new_n17076_, new_n16488_ );
or   ( new_n17078_, new_n17077_, new_n17074_ );
or   ( new_n17079_, new_n17072_, new_n17053_ );
or   ( new_n17080_, new_n17068_, new_n16139_ );
and  ( new_n17081_, new_n17080_, new_n17079_ );
and  ( new_n17082_, new_n16543_, new_n16501_ );
and  ( new_n17083_, new_n16549_, new_n16544_ );
or   ( new_n17084_, new_n17083_, new_n17082_ );
or   ( new_n17085_, new_n17084_, new_n17081_ );
and  ( new_n17086_, new_n17085_, new_n17078_ );
or   ( new_n17087_, new_n17086_, new_n17052_ );
or   ( new_n17088_, new_n17050_, new_n17028_ );
or   ( new_n17089_, new_n17047_, new_n17043_ );
and  ( new_n17090_, new_n17089_, new_n17088_ );
or   ( new_n17091_, new_n17084_, new_n17074_ );
or   ( new_n17092_, new_n17081_, new_n17077_ );
and  ( new_n17093_, new_n17092_, new_n17091_ );
or   ( new_n17094_, new_n17093_, new_n17090_ );
and  ( new_n17095_, new_n17094_, new_n17087_ );
and  ( new_n17096_, new_n16775_, new_n16710_ );
and  ( new_n17097_, new_n16784_, new_n16780_ );
or   ( new_n17098_, new_n17097_, new_n17096_ );
or   ( new_n17099_, new_n17098_, new_n17095_ );
and  ( new_n17100_, new_n16772_, new_n16576_ );
or   ( new_n17101_, new_n17100_, new_n16554_ );
and  ( new_n17102_, new_n17101_, new_n16779_ );
or   ( new_n17103_, new_n17093_, new_n17052_ );
or   ( new_n17104_, new_n17090_, new_n17086_ );
and  ( new_n17105_, new_n17104_, new_n17103_ );
or   ( new_n17106_, new_n17105_, new_n17102_ );
and  ( new_n17107_, new_n17106_, new_n17099_ );
or   ( new_n17108_, new_n17107_, new_n16925_ );
and  ( new_n17109_, new_n17107_, new_n16925_ );
or   ( new_n17110_, new_n16781_, new_n16554_ );
or   ( new_n17111_, new_n16784_, new_n16777_ );
and  ( new_n17112_, new_n17111_, new_n17110_ );
or   ( new_n17113_, new_n17112_, new_n16924_ );
or   ( new_n17114_, new_n16791_, new_n16485_ );
or   ( new_n17115_, new_n16789_, new_n16541_ );
and  ( new_n17116_, new_n17115_, new_n17114_ );
or   ( new_n17117_, new_n16805_, new_n16735_ );
or   ( new_n17118_, new_n16803_, new_n16670_ );
and  ( new_n17119_, new_n17118_, new_n17117_ );
or   ( new_n17120_, new_n16798_, new_n16748_ );
or   ( new_n17121_, new_n16796_, new_n16695_ );
and  ( new_n17122_, new_n17121_, new_n17120_ );
or   ( new_n17123_, new_n17122_, new_n17119_ );
or   ( new_n17124_, new_n16843_, new_n16052_ );
or   ( new_n17125_, new_n16839_, new_n16071_ );
and  ( new_n17126_, new_n17125_, new_n17124_ );
or   ( new_n17127_, new_n16852_, new_n16009_ );
or   ( new_n17128_, new_n16848_, new_n16029_ );
and  ( new_n17129_, new_n17128_, new_n17127_ );
or   ( new_n17130_, new_n17129_, new_n17126_ );
or   ( new_n17131_, new_n16862_, new_n16186_ );
or   ( new_n17132_, new_n16858_, new_n16204_ );
and  ( new_n17133_, new_n17132_, new_n17131_ );
and  ( new_n17134_, new_n17129_, new_n17126_ );
or   ( new_n17135_, new_n17134_, new_n17133_ );
and  ( new_n17136_, new_n17135_, new_n17130_ );
nand ( new_n17137_, new_n16809_, new_n138_ );
and  ( new_n17138_, new_n17137_, RI2b1c4342bf50_19 );
nand ( new_n17139_, new_n16811_, new_n138_ );
and  ( new_n17140_, new_n17139_, RI2b1c4342bed8_18 );
and  ( new_n17141_, new_n17140_, new_n17138_ );
or   ( new_n17142_, new_n17141_, new_n16502_ );
or   ( new_n17143_, new_n16821_, new_n16505_ );
or   ( new_n17144_, new_n16817_, new_n16438_ );
and  ( new_n17145_, new_n17144_, new_n17143_ );
or   ( new_n17146_, new_n17145_, new_n17142_ );
and  ( new_n17147_, new_n17145_, new_n17142_ );
or   ( new_n17148_, new_n16832_, new_n16085_ );
or   ( new_n17149_, new_n16828_, new_n16048_ );
and  ( new_n17150_, new_n17149_, new_n17148_ );
or   ( new_n17151_, new_n17150_, new_n17147_ );
and  ( new_n17152_, new_n17151_, new_n17146_ );
or   ( new_n17153_, new_n17152_, new_n17136_ );
and  ( new_n17154_, new_n17152_, new_n17136_ );
or   ( new_n17155_, new_n16876_, new_n16217_ );
or   ( new_n17156_, new_n16872_, new_n16234_ );
and  ( new_n17157_, new_n17156_, new_n17155_ );
or   ( new_n17158_, new_n16885_, new_n16151_ );
or   ( new_n17159_, new_n16881_, new_n16170_ );
and  ( new_n17160_, new_n17159_, new_n17158_ );
or   ( new_n17161_, new_n17160_, new_n17157_ );
or   ( new_n17162_, new_n16895_, new_n16108_ );
or   ( new_n17163_, new_n16891_, new_n16128_ );
and  ( new_n17164_, new_n17163_, new_n17162_ );
and  ( new_n17165_, new_n17160_, new_n17157_ );
or   ( new_n17166_, new_n17165_, new_n17164_ );
and  ( new_n17167_, new_n17166_, new_n17161_ );
or   ( new_n17168_, new_n17167_, new_n17154_ );
and  ( new_n17169_, new_n17168_, new_n17153_ );
or   ( new_n17170_, new_n17169_, new_n17123_ );
or   ( new_n17171_, new_n16908_, new_n16762_ );
or   ( new_n17172_, new_n16906_, new_n16598_ );
and  ( new_n17173_, new_n17172_, new_n17171_ );
and  ( new_n17174_, new_n17169_, new_n17123_ );
or   ( new_n17175_, new_n17174_, new_n17173_ );
and  ( new_n17176_, new_n17175_, new_n17170_ );
or   ( new_n17177_, new_n17176_, new_n17116_ );
or   ( new_n17178_, new_n16919_, new_n16769_ );
or   ( new_n17179_, new_n16917_, new_n16708_ );
and  ( new_n17180_, new_n17179_, new_n17178_ );
and  ( new_n17181_, new_n17176_, new_n17116_ );
or   ( new_n17182_, new_n17181_, new_n17180_ );
and  ( new_n17183_, new_n17182_, new_n17177_ );
or   ( new_n17184_, new_n17183_, new_n16786_ );
and  ( new_n17185_, new_n17184_, new_n17113_ );
or   ( new_n17186_, new_n16115_, new_n2119_ );
and  ( new_n17187_, new_n16132_, RI2b1c4342dc60_81 );
and  ( new_n17188_, new_n16114_, RI2b1c4342dbe8_80 );
or   ( new_n17189_, new_n17188_, new_n17187_ );
or   ( new_n17190_, new_n17189_, new_n16108_ );
or   ( new_n17191_, new_n16119_, new_n126_ );
or   ( new_n17192_, new_n16123_, new_n1511_ );
and  ( new_n17193_, new_n17192_, new_n17191_ );
or   ( new_n17194_, new_n17193_, new_n16128_ );
and  ( new_n17195_, new_n17194_, new_n17190_ );
and  ( new_n17196_, new_n16162_, RI2b1c4342db70_79 );
and  ( new_n17197_, new_n16165_, RI2b1c4342daf8_78 );
or   ( new_n17198_, new_n17197_, new_n17196_ );
or   ( new_n17199_, new_n17198_, new_n16151_ );
or   ( new_n17200_, new_n16174_, new_n1310_ );
or   ( new_n17201_, new_n16160_, new_n1002_ );
and  ( new_n17202_, new_n17201_, new_n17200_ );
or   ( new_n17203_, new_n17202_, new_n16170_ );
and  ( new_n17204_, new_n17203_, new_n17199_ );
or   ( new_n17205_, new_n16238_, new_n1004_ );
or   ( new_n17206_, new_n16224_, new_n886_ );
and  ( new_n17207_, new_n17206_, new_n17205_ );
or   ( new_n17208_, new_n17207_, new_n16217_ );
and  ( new_n17209_, new_n16226_, RI2b1c4342da80_77 );
and  ( new_n17210_, new_n16229_, RI2b1c4342da08_76 );
or   ( new_n17211_, new_n17210_, new_n17209_ );
or   ( new_n17212_, new_n17211_, new_n16234_ );
and  ( new_n17213_, new_n17212_, new_n17208_ );
or   ( new_n17214_, new_n17213_, new_n17204_ );
or   ( new_n17215_, new_n17211_, new_n16217_ );
or   ( new_n17216_, new_n17207_, new_n16234_ );
and  ( new_n17217_, new_n17216_, new_n17215_ );
or   ( new_n17218_, new_n17202_, new_n16151_ );
or   ( new_n17219_, new_n17198_, new_n16170_ );
and  ( new_n17220_, new_n17219_, new_n17218_ );
or   ( new_n17221_, new_n17220_, new_n17217_ );
and  ( new_n17222_, new_n17221_, new_n17214_ );
or   ( new_n17223_, new_n17222_, new_n17195_ );
or   ( new_n17224_, new_n17193_, new_n16108_ );
or   ( new_n17225_, new_n17189_, new_n16128_ );
and  ( new_n17226_, new_n17225_, new_n17224_ );
or   ( new_n17227_, new_n17217_, new_n17204_ );
or   ( new_n17228_, new_n17220_, new_n17213_ );
and  ( new_n17229_, new_n17228_, new_n17227_ );
or   ( new_n17230_, new_n17229_, new_n17226_ );
and  ( new_n17231_, new_n17230_, new_n17223_ );
and  ( new_n17232_, new_n17231_, new_n17186_ );
xor  ( new_n17233_, new_n2162_, new_n2323_ );
or   ( new_n17234_, new_n17233_, new_n292_ );
xor  ( new_n17235_, new_n2155_, new_n2328_ );
or   ( new_n17236_, new_n17235_, new_n289_ );
or   ( new_n17237_, new_n17236_, new_n17234_ );
and  ( new_n17238_, new_n17237_, new_n17138_ );
or   ( new_n17239_, new_n17140_, new_n17138_ );
and  ( new_n17240_, new_n17239_, new_n16813_ );
or   ( new_n17241_, new_n17140_, new_n16502_ );
or   ( new_n17242_, new_n16812_, new_n16433_ );
and  ( new_n17243_, new_n17242_, new_n17241_ );
or   ( new_n17244_, new_n17243_, new_n17240_ );
or   ( new_n17245_, new_n17244_, new_n526_ );
or   ( new_n17246_, new_n17138_, new_n16812_ );
or   ( new_n17247_, new_n17140_, new_n16810_ );
and  ( new_n17248_, new_n17247_, new_n17246_ );
or   ( new_n17249_, new_n17248_, new_n99_ );
and  ( new_n17250_, new_n17249_, new_n17245_ );
or   ( new_n17251_, new_n17250_, new_n16814_ );
or   ( new_n17252_, new_n17140_, new_n16433_ );
or   ( new_n17253_, new_n16812_, new_n16502_ );
and  ( new_n17254_, new_n17253_, new_n17248_ );
and  ( new_n17255_, new_n17254_, new_n17252_ );
and  ( new_n17256_, new_n17255_, RI2b1c4342d558_66 );
and  ( new_n17257_, new_n17240_, RI2b1c4342d4e0_65 );
or   ( new_n17258_, new_n17257_, new_n17256_ );
or   ( new_n17259_, new_n17258_, new_n17142_ );
and  ( new_n17260_, new_n17259_, new_n17251_ );
or   ( new_n17261_, new_n17260_, new_n17238_ );
or   ( new_n17262_, new_n16607_, new_n612_ );
or   ( new_n17263_, new_n16613_, new_n112_ );
and  ( new_n17264_, new_n17263_, new_n17262_ );
or   ( new_n17265_, new_n17264_, new_n16505_ );
and  ( new_n17266_, new_n16616_, RI2b1c4342d648_68 );
and  ( new_n17267_, new_n16603_, RI2b1c4342d5d0_67 );
or   ( new_n17268_, new_n17267_, new_n17266_ );
or   ( new_n17269_, new_n17268_, new_n16438_ );
and  ( new_n17270_, new_n17269_, new_n17265_ );
and  ( new_n17271_, new_n17260_, new_n17238_ );
or   ( new_n17272_, new_n17271_, new_n17270_ );
and  ( new_n17273_, new_n17272_, new_n17261_ );
or   ( new_n17274_, new_n16366_, new_n755_ );
or   ( new_n17275_, new_n16355_, new_n591_ );
and  ( new_n17276_, new_n17275_, new_n17274_ );
or   ( new_n17277_, new_n17276_, new_n16085_ );
and  ( new_n17278_, new_n16358_, RI2b1c4342d738_70 );
and  ( new_n17279_, new_n16362_, RI2b1c4342d6c0_69 );
or   ( new_n17280_, new_n17279_, new_n17278_ );
or   ( new_n17281_, new_n17280_, new_n16048_ );
and  ( new_n17282_, new_n17281_, new_n17277_ );
or   ( new_n17283_, new_n16075_, new_n806_ );
or   ( new_n17284_, new_n16060_, new_n110_ );
and  ( new_n17285_, new_n17284_, new_n17283_ );
or   ( new_n17286_, new_n17285_, new_n16052_ );
and  ( new_n17287_, new_n16063_, RI2b1c4342d828_72 );
and  ( new_n17288_, new_n16066_, RI2b1c4342d7b0_71 );
or   ( new_n17289_, new_n17288_, new_n17287_ );
or   ( new_n17290_, new_n17289_, new_n16071_ );
and  ( new_n17291_, new_n17290_, new_n17286_ );
or   ( new_n17292_, new_n17291_, new_n17282_ );
or   ( new_n17293_, new_n16033_, new_n859_ );
or   ( new_n17294_, new_n16017_, new_n105_ );
and  ( new_n17295_, new_n17294_, new_n17293_ );
or   ( new_n17296_, new_n17295_, new_n16009_ );
and  ( new_n17297_, new_n16021_, RI2b1c4342d918_74 );
and  ( new_n17298_, new_n16024_, RI2b1c4342d8a0_73 );
or   ( new_n17299_, new_n17298_, new_n17297_ );
or   ( new_n17300_, new_n17299_, new_n16029_ );
and  ( new_n17301_, new_n17300_, new_n17296_ );
and  ( new_n17302_, new_n17291_, new_n17282_ );
or   ( new_n17303_, new_n17302_, new_n17301_ );
and  ( new_n17304_, new_n17303_, new_n17292_ );
or   ( new_n17305_, new_n17304_, new_n17273_ );
or   ( new_n17306_, new_n16208_, new_n886_ );
or   ( new_n17307_, new_n16194_, new_n843_ );
and  ( new_n17308_, new_n17307_, new_n17306_ );
or   ( new_n17309_, new_n17308_, new_n16186_ );
and  ( new_n17310_, new_n16196_, RI2b1c4342da08_76 );
and  ( new_n17311_, new_n16199_, RI2b1c4342d990_75 );
or   ( new_n17312_, new_n17311_, new_n17310_ );
or   ( new_n17313_, new_n17312_, new_n16204_ );
and  ( new_n17314_, new_n17313_, new_n17309_ );
or   ( new_n17315_, new_n16238_, new_n1002_ );
or   ( new_n17316_, new_n16224_, new_n1004_ );
and  ( new_n17317_, new_n17316_, new_n17315_ );
or   ( new_n17318_, new_n17317_, new_n16217_ );
and  ( new_n17319_, new_n16226_, RI2b1c4342daf8_78 );
and  ( new_n17320_, new_n16229_, RI2b1c4342da80_77 );
or   ( new_n17321_, new_n17320_, new_n17319_ );
or   ( new_n17322_, new_n17321_, new_n16234_ );
and  ( new_n17323_, new_n17322_, new_n17318_ );
or   ( new_n17324_, new_n17323_, new_n17314_ );
or   ( new_n17325_, new_n16174_, new_n1511_ );
or   ( new_n17326_, new_n16160_, new_n1310_ );
and  ( new_n17327_, new_n17326_, new_n17325_ );
or   ( new_n17328_, new_n17327_, new_n16151_ );
and  ( new_n17329_, new_n16162_, RI2b1c4342dbe8_80 );
and  ( new_n17330_, new_n16165_, RI2b1c4342db70_79 );
or   ( new_n17331_, new_n17330_, new_n17329_ );
or   ( new_n17332_, new_n17331_, new_n16170_ );
and  ( new_n17333_, new_n17332_, new_n17328_ );
and  ( new_n17334_, new_n17323_, new_n17314_ );
or   ( new_n17335_, new_n17334_, new_n17333_ );
and  ( new_n17336_, new_n17335_, new_n17324_ );
and  ( new_n17337_, new_n17304_, new_n17273_ );
or   ( new_n17338_, new_n17337_, new_n17336_ );
and  ( new_n17339_, new_n17338_, new_n17305_ );
or   ( new_n17340_, new_n17339_, new_n17232_ );
and  ( new_n17341_, new_n16196_, RI2b1c4342d990_75 );
and  ( new_n17342_, new_n16199_, RI2b1c4342d918_74 );
or   ( new_n17343_, new_n17342_, new_n17341_ );
or   ( new_n17344_, new_n17343_, new_n16186_ );
or   ( new_n17345_, new_n16208_, new_n843_ );
or   ( new_n17346_, new_n16194_, new_n859_ );
and  ( new_n17347_, new_n17346_, new_n17345_ );
or   ( new_n17348_, new_n17347_, new_n16204_ );
and  ( new_n17349_, new_n17348_, new_n17344_ );
and  ( new_n17350_, new_n16021_, RI2b1c4342d8a0_73 );
and  ( new_n17351_, new_n16024_, RI2b1c4342d828_72 );
or   ( new_n17352_, new_n17351_, new_n17350_ );
or   ( new_n17353_, new_n17352_, new_n16009_ );
or   ( new_n17354_, new_n16033_, new_n105_ );
or   ( new_n17355_, new_n16017_, new_n806_ );
and  ( new_n17356_, new_n17355_, new_n17354_ );
or   ( new_n17357_, new_n17356_, new_n16029_ );
and  ( new_n17358_, new_n17357_, new_n17353_ );
or   ( new_n17359_, new_n16075_, new_n110_ );
or   ( new_n17360_, new_n16060_, new_n755_ );
and  ( new_n17361_, new_n17360_, new_n17359_ );
or   ( new_n17362_, new_n17361_, new_n16052_ );
and  ( new_n17363_, new_n16063_, RI2b1c4342d7b0_71 );
and  ( new_n17364_, new_n16066_, RI2b1c4342d738_70 );
or   ( new_n17365_, new_n17364_, new_n17363_ );
or   ( new_n17366_, new_n17365_, new_n16071_ );
and  ( new_n17367_, new_n17366_, new_n17362_ );
or   ( new_n17368_, new_n17367_, new_n17358_ );
or   ( new_n17369_, new_n17365_, new_n16052_ );
or   ( new_n17370_, new_n17361_, new_n16071_ );
and  ( new_n17371_, new_n17370_, new_n17369_ );
or   ( new_n17372_, new_n17356_, new_n16009_ );
or   ( new_n17373_, new_n17352_, new_n16029_ );
and  ( new_n17374_, new_n17373_, new_n17372_ );
or   ( new_n17375_, new_n17374_, new_n17371_ );
and  ( new_n17376_, new_n17375_, new_n17368_ );
or   ( new_n17377_, new_n17376_, new_n17349_ );
or   ( new_n17378_, new_n17347_, new_n16186_ );
or   ( new_n17379_, new_n17343_, new_n16204_ );
and  ( new_n17380_, new_n17379_, new_n17378_ );
or   ( new_n17381_, new_n17371_, new_n17358_ );
or   ( new_n17382_, new_n17374_, new_n17367_ );
and  ( new_n17383_, new_n17382_, new_n17381_ );
or   ( new_n17384_, new_n17383_, new_n17380_ );
and  ( new_n17385_, new_n17384_, new_n17377_ );
and  ( new_n17386_, new_n16358_, RI2b1c4342d6c0_69 );
and  ( new_n17387_, new_n16362_, RI2b1c4342d648_68 );
or   ( new_n17388_, new_n17387_, new_n17386_ );
or   ( new_n17389_, new_n17388_, new_n16085_ );
or   ( new_n17390_, new_n16366_, new_n591_ );
or   ( new_n17391_, new_n16355_, new_n612_ );
and  ( new_n17392_, new_n17391_, new_n17390_ );
or   ( new_n17393_, new_n17392_, new_n16048_ );
and  ( new_n17394_, new_n17393_, new_n17389_ );
and  ( new_n17395_, new_n16616_, RI2b1c4342d5d0_67 );
and  ( new_n17396_, new_n16603_, RI2b1c4342d558_66 );
or   ( new_n17397_, new_n17396_, new_n17395_ );
or   ( new_n17398_, new_n17397_, new_n16505_ );
or   ( new_n17399_, new_n16607_, new_n112_ );
or   ( new_n17400_, new_n16613_, new_n526_ );
and  ( new_n17401_, new_n17400_, new_n17399_ );
or   ( new_n17402_, new_n17401_, new_n16438_ );
and  ( new_n17403_, new_n17402_, new_n17398_ );
or   ( new_n17404_, new_n17244_, new_n99_ );
or   ( new_n17405_, new_n17404_, new_n16814_ );
and  ( new_n17406_, new_n17255_, RI2b1c4342d4e0_65 );
or   ( new_n17407_, new_n17406_, new_n17142_ );
and  ( new_n17408_, new_n17407_, new_n17405_ );
or   ( new_n17409_, new_n17408_, new_n17403_ );
or   ( new_n17410_, new_n17406_, new_n16814_ );
or   ( new_n17411_, new_n17404_, new_n17142_ );
and  ( new_n17412_, new_n17411_, new_n17410_ );
or   ( new_n17413_, new_n17401_, new_n16505_ );
or   ( new_n17414_, new_n17397_, new_n16438_ );
and  ( new_n17415_, new_n17414_, new_n17413_ );
or   ( new_n17416_, new_n17415_, new_n17412_ );
and  ( new_n17417_, new_n17416_, new_n17409_ );
or   ( new_n17418_, new_n17417_, new_n17394_ );
or   ( new_n17419_, new_n17392_, new_n16085_ );
or   ( new_n17420_, new_n17388_, new_n16048_ );
and  ( new_n17421_, new_n17420_, new_n17419_ );
or   ( new_n17422_, new_n17412_, new_n17403_ );
or   ( new_n17423_, new_n17415_, new_n17408_ );
and  ( new_n17424_, new_n17423_, new_n17422_ );
or   ( new_n17425_, new_n17424_, new_n17421_ );
and  ( new_n17426_, new_n17425_, new_n17418_ );
or   ( new_n17427_, new_n17426_, new_n17385_ );
and  ( new_n17428_, new_n17339_, new_n17232_ );
or   ( new_n17429_, new_n17428_, new_n17427_ );
and  ( new_n17430_, new_n17429_, new_n17340_ );
or   ( new_n17431_, new_n17145_, new_n16814_ );
or   ( new_n17432_, new_n17142_, new_n16823_ );
and  ( new_n17433_, new_n17432_, new_n17431_ );
or   ( new_n17434_, new_n17433_, new_n17150_ );
and  ( new_n17435_, new_n17146_, new_n16824_ );
or   ( new_n17436_, new_n17435_, new_n16834_ );
and  ( new_n17437_, new_n17436_, new_n17434_ );
and  ( new_n17438_, new_n17130_, new_n16855_ );
or   ( new_n17439_, new_n17438_, new_n17133_ );
or   ( new_n17440_, new_n17129_, new_n16845_ );
or   ( new_n17441_, new_n17126_, new_n16854_ );
and  ( new_n17442_, new_n17441_, new_n17440_ );
or   ( new_n17443_, new_n17442_, new_n16864_ );
and  ( new_n17444_, new_n17443_, new_n17439_ );
and  ( new_n17445_, new_n17161_, new_n16888_ );
or   ( new_n17446_, new_n17445_, new_n17164_ );
or   ( new_n17447_, new_n17160_, new_n16878_ );
or   ( new_n17448_, new_n17157_, new_n16887_ );
and  ( new_n17449_, new_n17448_, new_n17447_ );
or   ( new_n17450_, new_n17449_, new_n16897_ );
and  ( new_n17451_, new_n17450_, new_n17446_ );
or   ( new_n17452_, new_n16115_, new_n126_ );
or   ( new_n17453_, new_n17452_, new_n17451_ );
and  ( new_n17454_, new_n16102_, RI2b1c4342dc60_81 );
or   ( new_n17455_, new_n17449_, new_n17164_ );
or   ( new_n17456_, new_n17445_, new_n16897_ );
and  ( new_n17457_, new_n17456_, new_n17455_ );
or   ( new_n17458_, new_n17457_, new_n17454_ );
and  ( new_n17459_, new_n17458_, new_n17453_ );
or   ( new_n17460_, new_n17459_, new_n17444_ );
or   ( new_n17461_, new_n17442_, new_n17133_ );
or   ( new_n17462_, new_n17438_, new_n16864_ );
and  ( new_n17463_, new_n17462_, new_n17461_ );
or   ( new_n17464_, new_n17454_, new_n17451_ );
or   ( new_n17465_, new_n17457_, new_n17452_ );
and  ( new_n17466_, new_n17465_, new_n17464_ );
or   ( new_n17467_, new_n17466_, new_n17463_ );
and  ( new_n17468_, new_n17467_, new_n17460_ );
or   ( new_n17469_, new_n17468_, new_n17437_ );
and  ( new_n17470_, new_n17468_, new_n17437_ );
and  ( new_n17471_, new_n17217_, new_n17204_ );
or   ( new_n17472_, new_n17471_, new_n17195_ );
and  ( new_n17473_, new_n17472_, new_n17227_ );
and  ( new_n17474_, new_n17371_, new_n17358_ );
or   ( new_n17475_, new_n17474_, new_n17349_ );
and  ( new_n17476_, new_n17475_, new_n17381_ );
and  ( new_n17477_, new_n17415_, new_n17408_ );
or   ( new_n17478_, new_n17477_, new_n17421_ );
and  ( new_n17479_, new_n17478_, new_n17423_ );
or   ( new_n17480_, new_n17479_, new_n17476_ );
and  ( new_n17481_, new_n17412_, new_n17403_ );
or   ( new_n17482_, new_n17481_, new_n17394_ );
and  ( new_n17483_, new_n17482_, new_n17422_ );
and  ( new_n17484_, new_n17374_, new_n17367_ );
or   ( new_n17485_, new_n17484_, new_n17380_ );
and  ( new_n17486_, new_n17485_, new_n17382_ );
or   ( new_n17487_, new_n17486_, new_n17483_ );
and  ( new_n17488_, new_n17487_, new_n17480_ );
or   ( new_n17489_, new_n17488_, new_n17473_ );
and  ( new_n17490_, new_n17220_, new_n17213_ );
or   ( new_n17491_, new_n17490_, new_n17226_ );
and  ( new_n17492_, new_n17491_, new_n17228_ );
or   ( new_n17493_, new_n17483_, new_n17476_ );
or   ( new_n17494_, new_n17486_, new_n17479_ );
and  ( new_n17495_, new_n17494_, new_n17493_ );
or   ( new_n17496_, new_n17495_, new_n17492_ );
and  ( new_n17497_, new_n17496_, new_n17489_ );
or   ( new_n17498_, new_n17497_, new_n17470_ );
and  ( new_n17499_, new_n17498_, new_n17469_ );
or   ( new_n17500_, new_n17499_, new_n17430_ );
and  ( new_n17501_, new_n17499_, new_n17430_ );
or   ( new_n17502_, new_n16807_, new_n16800_ );
and  ( new_n17503_, new_n17502_, new_n17123_ );
or   ( new_n17504_, new_n17503_, new_n17501_ );
and  ( new_n17505_, new_n17504_, new_n17500_ );
or   ( new_n17506_, new_n17136_, new_n16836_ );
or   ( new_n17507_, new_n17152_, new_n16867_ );
and  ( new_n17508_, new_n17507_, new_n17506_ );
or   ( new_n17509_, new_n17508_, new_n17167_ );
and  ( new_n17510_, new_n17153_, new_n16868_ );
or   ( new_n17511_, new_n17510_, new_n16900_ );
and  ( new_n17512_, new_n17511_, new_n17509_ );
and  ( new_n17513_, new_n16718_, new_n16629_ );
or   ( new_n17514_, new_n17513_, new_n16722_ );
or   ( new_n17515_, new_n16717_, new_n16619_ );
or   ( new_n17516_, new_n16714_, new_n16628_ );
and  ( new_n17517_, new_n17516_, new_n17515_ );
or   ( new_n17518_, new_n17517_, new_n16639_ );
and  ( new_n17519_, new_n17518_, new_n17514_ );
and  ( new_n17520_, new_n17454_, new_n17451_ );
or   ( new_n17521_, new_n17520_, new_n17444_ );
and  ( new_n17522_, new_n17521_, new_n17464_ );
and  ( new_n17523_, new_n17486_, new_n17479_ );
or   ( new_n17524_, new_n17523_, new_n17492_ );
and  ( new_n17525_, new_n17524_, new_n17494_ );
or   ( new_n17526_, new_n17525_, new_n17522_ );
and  ( new_n17527_, new_n17483_, new_n17476_ );
or   ( new_n17528_, new_n17527_, new_n17473_ );
and  ( new_n17529_, new_n17528_, new_n17493_ );
and  ( new_n17530_, new_n17457_, new_n17452_ );
or   ( new_n17531_, new_n17530_, new_n17463_ );
and  ( new_n17532_, new_n17531_, new_n17465_ );
or   ( new_n17533_, new_n17532_, new_n17529_ );
and  ( new_n17534_, new_n17533_, new_n17526_ );
or   ( new_n17535_, new_n17534_, new_n17519_ );
or   ( new_n17536_, new_n17529_, new_n17522_ );
or   ( new_n17537_, new_n17532_, new_n17525_ );
and  ( new_n17538_, new_n17537_, new_n17536_ );
or   ( new_n17539_, new_n17517_, new_n16722_ );
or   ( new_n17540_, new_n17513_, new_n16639_ );
and  ( new_n17541_, new_n17540_, new_n17539_ );
or   ( new_n17542_, new_n17541_, new_n17538_ );
and  ( new_n17543_, new_n17542_, new_n17535_ );
or   ( new_n17544_, new_n17543_, new_n17512_ );
and  ( new_n17545_, new_n17544_, new_n17505_ );
and  ( new_n17546_, new_n17170_, new_n16903_ );
or   ( new_n17547_, new_n17546_, new_n17173_ );
or   ( new_n17548_, new_n17123_, new_n16902_ );
or   ( new_n17549_, new_n17169_, new_n16808_ );
and  ( new_n17550_, new_n17549_, new_n17548_ );
or   ( new_n17551_, new_n17550_, new_n16910_ );
and  ( new_n17552_, new_n17551_, new_n17547_ );
and  ( new_n17553_, new_n16738_, new_n16674_ );
or   ( new_n17554_, new_n17553_, new_n16750_ );
or   ( new_n17555_, new_n16737_, new_n16641_ );
or   ( new_n17556_, new_n16724_, new_n16672_ );
and  ( new_n17557_, new_n17556_, new_n17555_ );
or   ( new_n17558_, new_n17557_, new_n16697_ );
and  ( new_n17559_, new_n17558_, new_n17554_ );
and  ( new_n17560_, new_n17532_, new_n17525_ );
or   ( new_n17561_, new_n17560_, new_n17541_ );
and  ( new_n17562_, new_n17561_, new_n17537_ );
or   ( new_n17563_, new_n17562_, new_n17559_ );
and  ( new_n17564_, new_n17529_, new_n17522_ );
or   ( new_n17565_, new_n17564_, new_n17519_ );
and  ( new_n17566_, new_n17565_, new_n17536_ );
or   ( new_n17567_, new_n17557_, new_n16750_ );
or   ( new_n17568_, new_n17553_, new_n16697_ );
and  ( new_n17569_, new_n17568_, new_n17567_ );
or   ( new_n17570_, new_n17569_, new_n17566_ );
and  ( new_n17571_, new_n17570_, new_n17563_ );
or   ( new_n17572_, new_n17571_, new_n17552_ );
or   ( new_n17573_, new_n17566_, new_n17559_ );
or   ( new_n17574_, new_n17569_, new_n17562_ );
and  ( new_n17575_, new_n17574_, new_n17573_ );
or   ( new_n17576_, new_n17550_, new_n17173_ );
or   ( new_n17577_, new_n17546_, new_n16910_ );
and  ( new_n17578_, new_n17577_, new_n17576_ );
or   ( new_n17579_, new_n17578_, new_n17575_ );
and  ( new_n17580_, new_n17579_, new_n17572_ );
or   ( new_n17581_, new_n17544_, new_n17505_ );
and  ( new_n17582_, new_n17581_, new_n17580_ );
or   ( new_n17583_, new_n17582_, new_n17545_ );
and  ( new_n17584_, new_n17569_, new_n17562_ );
or   ( new_n17585_, new_n17584_, new_n17578_ );
and  ( new_n17586_, new_n17585_, new_n17574_ );
or   ( new_n17587_, new_n17586_, new_n17583_ );
or   ( new_n17588_, new_n17116_, new_n16913_ );
or   ( new_n17589_, new_n17176_, new_n16793_ );
and  ( new_n17590_, new_n17589_, new_n17588_ );
or   ( new_n17591_, new_n17590_, new_n17180_ );
and  ( new_n17592_, new_n17177_, new_n16914_ );
or   ( new_n17593_, new_n17592_, new_n16921_ );
and  ( new_n17594_, new_n17593_, new_n17591_ );
and  ( new_n17595_, new_n17586_, new_n17583_ );
or   ( new_n17596_, new_n17595_, new_n17594_ );
and  ( new_n17597_, new_n17596_, new_n17587_ );
or   ( new_n17598_, new_n17597_, new_n17185_ );
or   ( new_n17599_, new_n17598_, new_n17109_ );
and  ( new_n17600_, new_n17599_, new_n17108_ );
and  ( new_n17601_, new_n17597_, new_n17185_ );
or   ( new_n17602_, new_n17601_, new_n17109_ );
or   ( new_n17603_, new_n17575_, new_n17552_ );
or   ( new_n17604_, new_n17578_, new_n17571_ );
and  ( new_n17605_, new_n17604_, new_n17603_ );
or   ( new_n17606_, new_n17510_, new_n17167_ );
or   ( new_n17607_, new_n17508_, new_n16900_ );
and  ( new_n17608_, new_n17607_, new_n17606_ );
or   ( new_n17609_, new_n17538_, new_n17519_ );
or   ( new_n17610_, new_n17541_, new_n17534_ );
and  ( new_n17611_, new_n17610_, new_n17609_ );
and  ( new_n17612_, new_n17611_, new_n17608_ );
or   ( new_n17613_, new_n17612_, new_n17505_ );
or   ( new_n17614_, new_n17435_, new_n17150_ );
or   ( new_n17615_, new_n17433_, new_n16834_ );
and  ( new_n17616_, new_n17615_, new_n17614_ );
or   ( new_n17617_, new_n17466_, new_n17444_ );
or   ( new_n17618_, new_n17463_, new_n17459_ );
and  ( new_n17619_, new_n17618_, new_n17617_ );
or   ( new_n17620_, new_n17619_, new_n17616_ );
and  ( new_n17621_, new_n17619_, new_n17616_ );
or   ( new_n17622_, new_n17495_, new_n17473_ );
or   ( new_n17623_, new_n17492_, new_n17488_ );
and  ( new_n17624_, new_n17623_, new_n17622_ );
or   ( new_n17625_, new_n17624_, new_n17621_ );
and  ( new_n17626_, new_n17625_, new_n17620_ );
or   ( new_n17627_, new_n17229_, new_n17195_ );
or   ( new_n17628_, new_n17226_, new_n17222_ );
and  ( new_n17629_, new_n17628_, new_n17627_ );
and  ( new_n17630_, new_n16102_, RI2b1c4342dcd8_82 );
or   ( new_n17631_, new_n17630_, new_n17629_ );
or   ( new_n17632_, new_n17289_, new_n16052_ );
or   ( new_n17633_, new_n17285_, new_n16071_ );
and  ( new_n17634_, new_n17633_, new_n17632_ );
or   ( new_n17635_, new_n17280_, new_n16085_ );
or   ( new_n17636_, new_n17276_, new_n16048_ );
and  ( new_n17637_, new_n17636_, new_n17635_ );
or   ( new_n17638_, new_n17637_, new_n17634_ );
or   ( new_n17639_, new_n17299_, new_n16009_ );
or   ( new_n17640_, new_n17295_, new_n16029_ );
and  ( new_n17641_, new_n17640_, new_n17639_ );
and  ( new_n17642_, new_n17637_, new_n17634_ );
or   ( new_n17643_, new_n17642_, new_n17641_ );
and  ( new_n17644_, new_n17643_, new_n17638_ );
nand ( new_n17645_, new_n17235_, new_n138_ );
and  ( new_n17646_, new_n17645_, RI2b1c4342bfc8_20 );
nand ( new_n17647_, new_n17233_, new_n138_ );
and  ( new_n17648_, new_n17647_, RI2b1c4342c040_21 );
and  ( new_n17649_, new_n17648_, new_n17646_ );
or   ( new_n17650_, new_n17649_, new_n16810_ );
or   ( new_n17651_, new_n17258_, new_n16814_ );
or   ( new_n17652_, new_n17250_, new_n17142_ );
and  ( new_n17653_, new_n17652_, new_n17651_ );
or   ( new_n17654_, new_n17653_, new_n17650_ );
or   ( new_n17655_, new_n17268_, new_n16505_ );
or   ( new_n17656_, new_n17264_, new_n16438_ );
and  ( new_n17657_, new_n17656_, new_n17655_ );
and  ( new_n17658_, new_n17653_, new_n17650_ );
or   ( new_n17659_, new_n17658_, new_n17657_ );
and  ( new_n17660_, new_n17659_, new_n17654_ );
or   ( new_n17661_, new_n17660_, new_n17644_ );
and  ( new_n17662_, new_n17660_, new_n17644_ );
or   ( new_n17663_, new_n17321_, new_n16217_ );
or   ( new_n17664_, new_n17317_, new_n16234_ );
and  ( new_n17665_, new_n17664_, new_n17663_ );
or   ( new_n17666_, new_n17312_, new_n16186_ );
or   ( new_n17667_, new_n17308_, new_n16204_ );
and  ( new_n17668_, new_n17667_, new_n17666_ );
or   ( new_n17669_, new_n17668_, new_n17665_ );
or   ( new_n17670_, new_n17331_, new_n16151_ );
or   ( new_n17671_, new_n17327_, new_n16170_ );
and  ( new_n17672_, new_n17671_, new_n17670_ );
and  ( new_n17673_, new_n17668_, new_n17665_ );
or   ( new_n17674_, new_n17673_, new_n17672_ );
and  ( new_n17675_, new_n17674_, new_n17669_ );
or   ( new_n17676_, new_n17675_, new_n17662_ );
and  ( new_n17677_, new_n17676_, new_n17661_ );
or   ( new_n17678_, new_n17677_, new_n17631_ );
and  ( new_n17679_, new_n17677_, new_n17631_ );
or   ( new_n17680_, new_n17424_, new_n17394_ );
or   ( new_n17681_, new_n17421_, new_n17417_ );
and  ( new_n17682_, new_n17681_, new_n17680_ );
or   ( new_n17683_, new_n17383_, new_n17349_ );
or   ( new_n17684_, new_n17380_, new_n17376_ );
and  ( new_n17685_, new_n17684_, new_n17683_ );
and  ( new_n17686_, new_n17685_, new_n17682_ );
or   ( new_n17687_, new_n17686_, new_n17679_ );
and  ( new_n17688_, new_n17687_, new_n17678_ );
or   ( new_n17689_, new_n17688_, new_n17626_ );
and  ( new_n17690_, new_n17688_, new_n17626_ );
or   ( new_n17691_, new_n17119_, new_n16800_ );
or   ( new_n17692_, new_n17122_, new_n16807_ );
and  ( new_n17693_, new_n17692_, new_n17691_ );
or   ( new_n17694_, new_n17693_, new_n17690_ );
and  ( new_n17695_, new_n17694_, new_n17689_ );
or   ( new_n17696_, new_n17695_, new_n17544_ );
and  ( new_n17697_, new_n17696_, new_n17613_ );
or   ( new_n17698_, new_n17697_, new_n17605_ );
or   ( new_n17699_, new_n17695_, new_n17612_ );
and  ( new_n17700_, new_n17699_, new_n17581_ );
or   ( new_n17701_, new_n17700_, new_n17580_ );
and  ( new_n17702_, new_n17701_, new_n17698_ );
or   ( new_n17703_, new_n17611_, new_n17512_ );
or   ( new_n17704_, new_n17608_, new_n17543_ );
and  ( new_n17705_, new_n17704_, new_n17703_ );
or   ( new_n17706_, new_n17682_, new_n17385_ );
or   ( new_n17707_, new_n17685_, new_n17426_ );
and  ( new_n17708_, new_n17707_, new_n17706_ );
or   ( new_n17709_, new_n17231_, new_n17186_ );
and  ( new_n17710_, new_n17709_, new_n17631_ );
or   ( new_n17711_, new_n17710_, new_n17708_ );
or   ( new_n17712_, new_n17644_, new_n17273_ );
or   ( new_n17713_, new_n17660_, new_n17304_ );
and  ( new_n17714_, new_n17713_, new_n17712_ );
or   ( new_n17715_, new_n17714_, new_n17675_ );
and  ( new_n17716_, new_n17661_, new_n17305_ );
or   ( new_n17717_, new_n17716_, new_n17336_ );
and  ( new_n17718_, new_n17717_, new_n17715_ );
and  ( new_n17719_, new_n17710_, new_n17708_ );
or   ( new_n17720_, new_n17719_, new_n17718_ );
and  ( new_n17721_, new_n17720_, new_n17711_ );
or   ( new_n17722_, new_n17648_, new_n17646_ );
and  ( new_n17723_, new_n17722_, new_n17237_ );
or   ( new_n17724_, new_n17646_, new_n16810_ );
or   ( new_n17725_, new_n17236_, new_n17138_ );
and  ( new_n17726_, new_n17725_, new_n17724_ );
or   ( new_n17727_, new_n17726_, new_n17723_ );
or   ( new_n17728_, new_n17727_, new_n99_ );
or   ( new_n17729_, new_n17728_, new_n17238_ );
or   ( new_n17730_, new_n17646_, new_n17138_ );
or   ( new_n17731_, new_n17236_, new_n16810_ );
or   ( new_n17732_, new_n17648_, new_n17236_ );
or   ( new_n17733_, new_n17646_, new_n17234_ );
and  ( new_n17734_, new_n17733_, new_n17732_ );
and  ( new_n17735_, new_n17734_, new_n17731_ );
and  ( new_n17736_, new_n17735_, new_n17730_ );
and  ( new_n17737_, new_n17736_, RI2b1c4342d4e0_65 );
or   ( new_n17738_, new_n17737_, new_n17650_ );
and  ( new_n17739_, new_n17738_, new_n17729_ );
or   ( new_n17740_, new_n17244_, new_n112_ );
or   ( new_n17741_, new_n17248_, new_n526_ );
and  ( new_n17742_, new_n17741_, new_n17740_ );
or   ( new_n17743_, new_n17742_, new_n16814_ );
and  ( new_n17744_, new_n17255_, RI2b1c4342d5d0_67 );
and  ( new_n17745_, new_n17240_, RI2b1c4342d558_66 );
or   ( new_n17746_, new_n17745_, new_n17744_ );
or   ( new_n17747_, new_n17746_, new_n17142_ );
and  ( new_n17748_, new_n17747_, new_n17743_ );
or   ( new_n17749_, new_n17748_, new_n17739_ );
and  ( new_n17750_, new_n17748_, new_n17739_ );
or   ( new_n17751_, new_n16607_, new_n591_ );
or   ( new_n17752_, new_n16613_, new_n612_ );
and  ( new_n17753_, new_n17752_, new_n17751_ );
or   ( new_n17754_, new_n17753_, new_n16505_ );
and  ( new_n17755_, new_n16616_, RI2b1c4342d6c0_69 );
and  ( new_n17756_, new_n16603_, RI2b1c4342d648_68 );
or   ( new_n17757_, new_n17756_, new_n17755_ );
or   ( new_n17758_, new_n17757_, new_n16438_ );
and  ( new_n17759_, new_n17758_, new_n17754_ );
or   ( new_n17760_, new_n17759_, new_n17750_ );
and  ( new_n17761_, new_n17760_, new_n17749_ );
or   ( new_n17762_, new_n16366_, new_n110_ );
or   ( new_n17763_, new_n16355_, new_n755_ );
and  ( new_n17764_, new_n17763_, new_n17762_ );
or   ( new_n17765_, new_n17764_, new_n16085_ );
and  ( new_n17766_, new_n16358_, RI2b1c4342d7b0_71 );
and  ( new_n17767_, new_n16362_, RI2b1c4342d738_70 );
or   ( new_n17768_, new_n17767_, new_n17766_ );
or   ( new_n17769_, new_n17768_, new_n16048_ );
and  ( new_n17770_, new_n17769_, new_n17765_ );
or   ( new_n17771_, new_n16075_, new_n105_ );
or   ( new_n17772_, new_n16060_, new_n806_ );
and  ( new_n17773_, new_n17772_, new_n17771_ );
or   ( new_n17774_, new_n17773_, new_n16052_ );
and  ( new_n17775_, new_n16063_, RI2b1c4342d8a0_73 );
and  ( new_n17776_, new_n16066_, RI2b1c4342d828_72 );
or   ( new_n17777_, new_n17776_, new_n17775_ );
or   ( new_n17778_, new_n17777_, new_n16071_ );
and  ( new_n17779_, new_n17778_, new_n17774_ );
or   ( new_n17780_, new_n17779_, new_n17770_ );
and  ( new_n17781_, new_n17779_, new_n17770_ );
or   ( new_n17782_, new_n16033_, new_n843_ );
or   ( new_n17783_, new_n16017_, new_n859_ );
and  ( new_n17784_, new_n17783_, new_n17782_ );
or   ( new_n17785_, new_n17784_, new_n16009_ );
and  ( new_n17786_, new_n16021_, RI2b1c4342d990_75 );
and  ( new_n17787_, new_n16024_, RI2b1c4342d918_74 );
or   ( new_n17788_, new_n17787_, new_n17786_ );
or   ( new_n17789_, new_n17788_, new_n16029_ );
and  ( new_n17790_, new_n17789_, new_n17785_ );
or   ( new_n17791_, new_n17790_, new_n17781_ );
and  ( new_n17792_, new_n17791_, new_n17780_ );
or   ( new_n17793_, new_n17792_, new_n17761_ );
or   ( new_n17794_, new_n16208_, new_n1004_ );
or   ( new_n17795_, new_n16194_, new_n886_ );
and  ( new_n17796_, new_n17795_, new_n17794_ );
or   ( new_n17797_, new_n17796_, new_n16186_ );
and  ( new_n17798_, new_n16196_, RI2b1c4342da80_77 );
and  ( new_n17799_, new_n16199_, RI2b1c4342da08_76 );
or   ( new_n17800_, new_n17799_, new_n17798_ );
or   ( new_n17801_, new_n17800_, new_n16204_ );
and  ( new_n17802_, new_n17801_, new_n17797_ );
or   ( new_n17803_, new_n16238_, new_n1310_ );
or   ( new_n17804_, new_n16224_, new_n1002_ );
and  ( new_n17805_, new_n17804_, new_n17803_ );
or   ( new_n17806_, new_n17805_, new_n16217_ );
and  ( new_n17807_, new_n16226_, RI2b1c4342db70_79 );
and  ( new_n17808_, new_n16229_, RI2b1c4342daf8_78 );
or   ( new_n17809_, new_n17808_, new_n17807_ );
or   ( new_n17810_, new_n17809_, new_n16234_ );
and  ( new_n17811_, new_n17810_, new_n17806_ );
or   ( new_n17812_, new_n17811_, new_n17802_ );
and  ( new_n17813_, new_n17811_, new_n17802_ );
or   ( new_n17814_, new_n16174_, new_n126_ );
or   ( new_n17815_, new_n16160_, new_n1511_ );
and  ( new_n17816_, new_n17815_, new_n17814_ );
or   ( new_n17817_, new_n17816_, new_n16151_ );
and  ( new_n17818_, new_n16162_, RI2b1c4342dc60_81 );
and  ( new_n17819_, new_n16165_, RI2b1c4342dbe8_80 );
or   ( new_n17820_, new_n17819_, new_n17818_ );
or   ( new_n17821_, new_n17820_, new_n16170_ );
and  ( new_n17822_, new_n17821_, new_n17817_ );
or   ( new_n17823_, new_n17822_, new_n17813_ );
and  ( new_n17824_, new_n17823_, new_n17812_ );
and  ( new_n17825_, new_n17792_, new_n17761_ );
or   ( new_n17826_, new_n17825_, new_n17824_ );
and  ( new_n17827_, new_n17826_, new_n17793_ );
or   ( new_n17828_, new_n16119_, new_n121_ );
or   ( new_n17829_, new_n16123_, new_n2119_ );
and  ( new_n17830_, new_n17829_, new_n17828_ );
or   ( new_n17831_, new_n17830_, new_n16108_ );
and  ( new_n17832_, new_n16132_, RI2b1c4342dd50_83 );
and  ( new_n17833_, new_n16114_, RI2b1c4342dcd8_82 );
or   ( new_n17834_, new_n17833_, new_n17832_ );
or   ( new_n17835_, new_n17834_, new_n16128_ );
and  ( new_n17836_, new_n17835_, new_n17831_ );
or   ( new_n17837_, new_n16115_, new_n2541_ );
and  ( new_n17838_, new_n17837_, new_n17836_ );
or   ( new_n17839_, new_n16119_, new_n2119_ );
or   ( new_n17840_, new_n16123_, new_n126_ );
and  ( new_n17841_, new_n17840_, new_n17839_ );
or   ( new_n17842_, new_n17841_, new_n16108_ );
and  ( new_n17843_, new_n16132_, RI2b1c4342dcd8_82 );
and  ( new_n17844_, new_n16114_, RI2b1c4342dc60_81 );
or   ( new_n17845_, new_n17844_, new_n17843_ );
or   ( new_n17846_, new_n17845_, new_n16128_ );
and  ( new_n17847_, new_n17846_, new_n17842_ );
and  ( new_n17848_, new_n17847_, new_n17838_ );
or   ( new_n17849_, new_n17847_, new_n17838_ );
or   ( new_n17850_, new_n16115_, new_n121_ );
and  ( new_n17851_, new_n17850_, new_n17849_ );
or   ( new_n17852_, new_n17851_, new_n17848_ );
and  ( new_n17853_, new_n17852_, new_n17827_ );
or   ( new_n17854_, new_n17852_, new_n17827_ );
or   ( new_n17855_, new_n17665_, new_n17314_ );
or   ( new_n17856_, new_n17668_, new_n17323_ );
and  ( new_n17857_, new_n17856_, new_n17855_ );
or   ( new_n17858_, new_n17857_, new_n17672_ );
and  ( new_n17859_, new_n17669_, new_n17324_ );
or   ( new_n17860_, new_n17859_, new_n17333_ );
and  ( new_n17861_, new_n17860_, new_n17858_ );
or   ( new_n17862_, new_n17634_, new_n17282_ );
or   ( new_n17863_, new_n17637_, new_n17291_ );
and  ( new_n17864_, new_n17863_, new_n17862_ );
or   ( new_n17865_, new_n17864_, new_n17641_ );
and  ( new_n17866_, new_n17638_, new_n17292_ );
or   ( new_n17867_, new_n17866_, new_n17301_ );
and  ( new_n17868_, new_n17867_, new_n17865_ );
or   ( new_n17869_, new_n17868_, new_n17861_ );
or   ( new_n17870_, new_n17653_, new_n17238_ );
or   ( new_n17871_, new_n17650_, new_n17260_ );
and  ( new_n17872_, new_n17871_, new_n17870_ );
or   ( new_n17873_, new_n17872_, new_n17657_ );
and  ( new_n17874_, new_n17654_, new_n17261_ );
or   ( new_n17875_, new_n17874_, new_n17270_ );
and  ( new_n17876_, new_n17875_, new_n17873_ );
and  ( new_n17877_, new_n17868_, new_n17861_ );
or   ( new_n17878_, new_n17877_, new_n17876_ );
and  ( new_n17879_, new_n17878_, new_n17869_ );
and  ( new_n17880_, new_n17879_, new_n17854_ );
or   ( new_n17881_, new_n17880_, new_n17853_ );
and  ( new_n17882_, new_n17881_, new_n17721_ );
or   ( new_n17883_, new_n17881_, new_n17721_ );
or   ( new_n17884_, new_n17619_, new_n17437_ );
or   ( new_n17885_, new_n17616_, new_n17468_ );
and  ( new_n17886_, new_n17885_, new_n17884_ );
or   ( new_n17887_, new_n17886_, new_n17624_ );
and  ( new_n17888_, new_n17620_, new_n17469_ );
or   ( new_n17889_, new_n17888_, new_n17497_ );
and  ( new_n17890_, new_n17889_, new_n17887_ );
and  ( new_n17891_, new_n17890_, new_n17883_ );
or   ( new_n17892_, new_n17891_, new_n17882_ );
and  ( new_n17893_, new_n17892_, new_n17705_ );
or   ( new_n17894_, new_n17892_, new_n17705_ );
or   ( new_n17895_, new_n17626_, new_n17430_ );
or   ( new_n17896_, new_n17688_, new_n17499_ );
and  ( new_n17897_, new_n17896_, new_n17895_ );
or   ( new_n17898_, new_n17897_, new_n17693_ );
and  ( new_n17899_, new_n17689_, new_n17500_ );
or   ( new_n17900_, new_n17899_, new_n17503_ );
and  ( new_n17901_, new_n17900_, new_n17898_ );
and  ( new_n17902_, new_n17901_, new_n17894_ );
or   ( new_n17903_, new_n17902_, new_n17893_ );
or   ( new_n17904_, new_n17903_, new_n17702_ );
or   ( new_n17905_, new_n17592_, new_n17180_ );
or   ( new_n17906_, new_n17590_, new_n16921_ );
and  ( new_n17907_, new_n17906_, new_n17905_ );
and  ( new_n17908_, new_n17566_, new_n17559_ );
or   ( new_n17909_, new_n17908_, new_n17552_ );
and  ( new_n17910_, new_n17909_, new_n17573_ );
or   ( new_n17911_, new_n17910_, new_n17583_ );
and  ( new_n17912_, new_n17695_, new_n17612_ );
or   ( new_n17913_, new_n17912_, new_n17605_ );
and  ( new_n17914_, new_n17913_, new_n17699_ );
or   ( new_n17915_, new_n17914_, new_n17586_ );
and  ( new_n17916_, new_n17915_, new_n17911_ );
or   ( new_n17917_, new_n17916_, new_n17907_ );
or   ( new_n17918_, new_n17914_, new_n17910_ );
and  ( new_n17919_, new_n17918_, new_n17587_ );
or   ( new_n17920_, new_n17919_, new_n17594_ );
and  ( new_n17921_, new_n17920_, new_n17917_ );
or   ( new_n17922_, new_n17921_, new_n17904_ );
and  ( new_n17923_, new_n17921_, new_n17904_ );
or   ( new_n17924_, new_n17899_, new_n17693_ );
or   ( new_n17925_, new_n17897_, new_n17503_ );
and  ( new_n17926_, new_n17925_, new_n17924_ );
or   ( new_n17927_, new_n17611_, new_n17608_ );
and  ( new_n17928_, new_n17927_, new_n17544_ );
or   ( new_n17929_, new_n17928_, new_n17892_ );
or   ( new_n17930_, new_n17746_, new_n16814_ );
or   ( new_n17931_, new_n17742_, new_n17142_ );
and  ( new_n17932_, new_n17931_, new_n17930_ );
or   ( new_n17933_, new_n17737_, new_n17238_ );
or   ( new_n17934_, new_n17728_, new_n17650_ );
and  ( new_n17935_, new_n17934_, new_n17933_ );
or   ( new_n17936_, new_n17935_, new_n17932_ );
and  ( new_n17937_, new_n17935_, new_n17932_ );
or   ( new_n17938_, new_n17757_, new_n16505_ );
or   ( new_n17939_, new_n17753_, new_n16438_ );
and  ( new_n17940_, new_n17939_, new_n17938_ );
or   ( new_n17941_, new_n17940_, new_n17937_ );
and  ( new_n17942_, new_n17941_, new_n17936_ );
or   ( new_n17943_, new_n17777_, new_n16052_ );
or   ( new_n17944_, new_n17773_, new_n16071_ );
and  ( new_n17945_, new_n17944_, new_n17943_ );
or   ( new_n17946_, new_n17768_, new_n16085_ );
or   ( new_n17947_, new_n17764_, new_n16048_ );
and  ( new_n17948_, new_n17947_, new_n17946_ );
or   ( new_n17949_, new_n17948_, new_n17945_ );
and  ( new_n17950_, new_n17948_, new_n17945_ );
or   ( new_n17951_, new_n17788_, new_n16009_ );
or   ( new_n17952_, new_n17784_, new_n16029_ );
and  ( new_n17953_, new_n17952_, new_n17951_ );
or   ( new_n17954_, new_n17953_, new_n17950_ );
and  ( new_n17955_, new_n17954_, new_n17949_ );
or   ( new_n17956_, new_n17955_, new_n17942_ );
or   ( new_n17957_, new_n17800_, new_n16186_ );
or   ( new_n17958_, new_n17796_, new_n16204_ );
and  ( new_n17959_, new_n17958_, new_n17957_ );
or   ( new_n17960_, new_n17809_, new_n16217_ );
or   ( new_n17961_, new_n17805_, new_n16234_ );
and  ( new_n17962_, new_n17961_, new_n17960_ );
or   ( new_n17963_, new_n17962_, new_n17959_ );
and  ( new_n17964_, new_n17962_, new_n17959_ );
or   ( new_n17965_, new_n17820_, new_n16151_ );
or   ( new_n17966_, new_n17816_, new_n16170_ );
and  ( new_n17967_, new_n17966_, new_n17965_ );
or   ( new_n17968_, new_n17967_, new_n17964_ );
and  ( new_n17969_, new_n17968_, new_n17963_ );
and  ( new_n17970_, new_n17955_, new_n17942_ );
or   ( new_n17971_, new_n17970_, new_n17969_ );
and  ( new_n17972_, new_n17971_, new_n17956_ );
and  ( new_n17973_, new_n16102_, RI2b1c4342ddc8_84 );
or   ( new_n17974_, new_n17834_, new_n16108_ );
or   ( new_n17975_, new_n17830_, new_n16128_ );
and  ( new_n17976_, new_n17975_, new_n17974_ );
or   ( new_n17977_, new_n17976_, new_n17973_ );
or   ( new_n17978_, new_n17845_, new_n16108_ );
or   ( new_n17979_, new_n17841_, new_n16128_ );
and  ( new_n17980_, new_n17979_, new_n17978_ );
or   ( new_n17981_, new_n17980_, new_n17977_ );
and  ( new_n17982_, new_n16102_, RI2b1c4342dd50_83 );
and  ( new_n17983_, new_n17980_, new_n17977_ );
or   ( new_n17984_, new_n17983_, new_n17982_ );
and  ( new_n17985_, new_n17984_, new_n17981_ );
or   ( new_n17986_, new_n17985_, new_n17972_ );
or   ( new_n17987_, new_n17859_, new_n17672_ );
or   ( new_n17988_, new_n17857_, new_n17333_ );
and  ( new_n17989_, new_n17988_, new_n17987_ );
or   ( new_n17990_, new_n17866_, new_n17641_ );
or   ( new_n17991_, new_n17864_, new_n17301_ );
and  ( new_n17992_, new_n17991_, new_n17990_ );
or   ( new_n17993_, new_n17992_, new_n17989_ );
or   ( new_n17994_, new_n17874_, new_n17657_ );
or   ( new_n17995_, new_n17872_, new_n17270_ );
and  ( new_n17996_, new_n17995_, new_n17994_ );
and  ( new_n17997_, new_n17992_, new_n17989_ );
or   ( new_n17998_, new_n17997_, new_n17996_ );
and  ( new_n17999_, new_n17998_, new_n17993_ );
and  ( new_n18000_, new_n17985_, new_n17972_ );
or   ( new_n18001_, new_n18000_, new_n17999_ );
and  ( new_n18002_, new_n18001_, new_n17986_ );
or   ( new_n18003_, new_n17685_, new_n17682_ );
and  ( new_n18004_, new_n18003_, new_n17427_ );
or   ( new_n18005_, new_n17629_, new_n17186_ );
or   ( new_n18006_, new_n17630_, new_n17231_ );
and  ( new_n18007_, new_n18006_, new_n18005_ );
or   ( new_n18008_, new_n18007_, new_n18004_ );
or   ( new_n18009_, new_n17716_, new_n17675_ );
or   ( new_n18010_, new_n17714_, new_n17336_ );
and  ( new_n18011_, new_n18010_, new_n18009_ );
and  ( new_n18012_, new_n18007_, new_n18004_ );
or   ( new_n18013_, new_n18012_, new_n18011_ );
and  ( new_n18014_, new_n18013_, new_n18008_ );
or   ( new_n18015_, new_n18014_, new_n18002_ );
and  ( new_n18016_, new_n18014_, new_n18002_ );
or   ( new_n18017_, new_n17888_, new_n17624_ );
or   ( new_n18018_, new_n17886_, new_n17497_ );
and  ( new_n18019_, new_n18018_, new_n18017_ );
or   ( new_n18020_, new_n18019_, new_n18016_ );
and  ( new_n18021_, new_n18020_, new_n18015_ );
or   ( new_n18022_, new_n18021_, new_n17705_ );
and  ( new_n18023_, new_n18022_, new_n17929_ );
or   ( new_n18024_, new_n18023_, new_n17926_ );
or   ( new_n18025_, new_n18021_, new_n17928_ );
and  ( new_n18026_, new_n18025_, new_n17894_ );
or   ( new_n18027_, new_n18026_, new_n17901_ );
and  ( new_n18028_, new_n18027_, new_n18024_ );
or   ( new_n18029_, new_n17631_, new_n17339_ );
or   ( new_n18030_, new_n17677_, new_n17232_ );
and  ( new_n18031_, new_n18030_, new_n18029_ );
or   ( new_n18032_, new_n18031_, new_n17686_ );
and  ( new_n18033_, new_n17678_, new_n17340_ );
or   ( new_n18034_, new_n18033_, new_n17427_ );
and  ( new_n18035_, new_n18034_, new_n18032_ );
or   ( new_n18036_, new_n17992_, new_n17861_ );
or   ( new_n18037_, new_n17989_, new_n17868_ );
and  ( new_n18038_, new_n18037_, new_n18036_ );
or   ( new_n18039_, new_n18038_, new_n17996_ );
and  ( new_n18040_, new_n17993_, new_n17869_ );
or   ( new_n18041_, new_n18040_, new_n17876_ );
and  ( new_n18042_, new_n18041_, new_n18039_ );
or   ( new_n18043_, new_n17980_, new_n17838_ );
or   ( new_n18044_, new_n17977_, new_n17847_ );
and  ( new_n18045_, new_n18044_, new_n18043_ );
or   ( new_n18046_, new_n18045_, new_n17982_ );
and  ( new_n18047_, new_n17981_, new_n17849_ );
or   ( new_n18048_, new_n18047_, new_n17850_ );
and  ( new_n18049_, new_n18048_, new_n18046_ );
or   ( new_n18050_, new_n18049_, new_n18042_ );
or   ( new_n18051_, new_n17955_, new_n17761_ );
or   ( new_n18052_, new_n17942_, new_n17792_ );
and  ( new_n18053_, new_n18052_, new_n18051_ );
or   ( new_n18054_, new_n18053_, new_n17969_ );
and  ( new_n18055_, new_n17956_, new_n17793_ );
or   ( new_n18056_, new_n18055_, new_n17824_ );
and  ( new_n18057_, new_n18056_, new_n18054_ );
and  ( new_n18058_, new_n18049_, new_n18042_ );
or   ( new_n18059_, new_n18058_, new_n18057_ );
and  ( new_n18060_, new_n18059_, new_n18050_ );
xor  ( new_n18061_, new_n2862_, new_n2993_ );
or   ( new_n18062_, new_n18061_, new_n302_ );
xor  ( new_n18063_, new_n2855_, new_n2998_ );
or   ( new_n18064_, new_n18063_, new_n299_ );
or   ( new_n18065_, new_n18064_, new_n18062_ );
and  ( new_n18066_, new_n18065_, new_n17648_ );
or   ( new_n18067_, new_n17727_, new_n526_ );
or   ( new_n18068_, new_n17734_, new_n99_ );
and  ( new_n18069_, new_n18068_, new_n18067_ );
or   ( new_n18070_, new_n18069_, new_n17238_ );
and  ( new_n18071_, new_n17736_, RI2b1c4342d558_66 );
and  ( new_n18072_, new_n17723_, RI2b1c4342d4e0_65 );
or   ( new_n18073_, new_n18072_, new_n18071_ );
or   ( new_n18074_, new_n18073_, new_n17650_ );
and  ( new_n18075_, new_n18074_, new_n18070_ );
or   ( new_n18076_, new_n18075_, new_n18066_ );
or   ( new_n18077_, new_n17244_, new_n612_ );
or   ( new_n18078_, new_n17248_, new_n112_ );
and  ( new_n18079_, new_n18078_, new_n18077_ );
or   ( new_n18080_, new_n18079_, new_n16814_ );
and  ( new_n18081_, new_n17255_, RI2b1c4342d648_68 );
and  ( new_n18082_, new_n17240_, RI2b1c4342d5d0_67 );
or   ( new_n18083_, new_n18082_, new_n18081_ );
or   ( new_n18084_, new_n18083_, new_n17142_ );
and  ( new_n18085_, new_n18084_, new_n18080_ );
and  ( new_n18086_, new_n18075_, new_n18066_ );
or   ( new_n18087_, new_n18086_, new_n18085_ );
and  ( new_n18088_, new_n18087_, new_n18076_ );
or   ( new_n18089_, new_n16607_, new_n755_ );
or   ( new_n18090_, new_n16613_, new_n591_ );
and  ( new_n18091_, new_n18090_, new_n18089_ );
or   ( new_n18092_, new_n18091_, new_n16505_ );
and  ( new_n18093_, new_n16616_, RI2b1c4342d738_70 );
and  ( new_n18094_, new_n16603_, RI2b1c4342d6c0_69 );
or   ( new_n18095_, new_n18094_, new_n18093_ );
or   ( new_n18096_, new_n18095_, new_n16438_ );
and  ( new_n18097_, new_n18096_, new_n18092_ );
or   ( new_n18098_, new_n16366_, new_n806_ );
or   ( new_n18099_, new_n16355_, new_n110_ );
and  ( new_n18100_, new_n18099_, new_n18098_ );
or   ( new_n18101_, new_n18100_, new_n16085_ );
and  ( new_n18102_, new_n16358_, RI2b1c4342d828_72 );
and  ( new_n18103_, new_n16362_, RI2b1c4342d7b0_71 );
or   ( new_n18104_, new_n18103_, new_n18102_ );
or   ( new_n18105_, new_n18104_, new_n16048_ );
and  ( new_n18106_, new_n18105_, new_n18101_ );
or   ( new_n18107_, new_n18106_, new_n18097_ );
or   ( new_n18108_, new_n16075_, new_n859_ );
or   ( new_n18109_, new_n16060_, new_n105_ );
and  ( new_n18110_, new_n18109_, new_n18108_ );
or   ( new_n18111_, new_n18110_, new_n16052_ );
and  ( new_n18112_, new_n16063_, RI2b1c4342d918_74 );
and  ( new_n18113_, new_n16066_, RI2b1c4342d8a0_73 );
or   ( new_n18114_, new_n18113_, new_n18112_ );
or   ( new_n18115_, new_n18114_, new_n16071_ );
and  ( new_n18116_, new_n18115_, new_n18111_ );
and  ( new_n18117_, new_n18106_, new_n18097_ );
or   ( new_n18118_, new_n18117_, new_n18116_ );
and  ( new_n18119_, new_n18118_, new_n18107_ );
or   ( new_n18120_, new_n18119_, new_n18088_ );
or   ( new_n18121_, new_n16033_, new_n886_ );
or   ( new_n18122_, new_n16017_, new_n843_ );
and  ( new_n18123_, new_n18122_, new_n18121_ );
or   ( new_n18124_, new_n18123_, new_n16009_ );
and  ( new_n18125_, new_n16021_, RI2b1c4342da08_76 );
and  ( new_n18126_, new_n16024_, RI2b1c4342d990_75 );
or   ( new_n18127_, new_n18126_, new_n18125_ );
or   ( new_n18128_, new_n18127_, new_n16029_ );
and  ( new_n18129_, new_n18128_, new_n18124_ );
or   ( new_n18130_, new_n16208_, new_n1002_ );
or   ( new_n18131_, new_n16194_, new_n1004_ );
and  ( new_n18132_, new_n18131_, new_n18130_ );
or   ( new_n18133_, new_n18132_, new_n16186_ );
and  ( new_n18134_, new_n16196_, RI2b1c4342daf8_78 );
and  ( new_n18135_, new_n16199_, RI2b1c4342da80_77 );
or   ( new_n18136_, new_n18135_, new_n18134_ );
or   ( new_n18137_, new_n18136_, new_n16204_ );
and  ( new_n18138_, new_n18137_, new_n18133_ );
or   ( new_n18139_, new_n18138_, new_n18129_ );
or   ( new_n18140_, new_n16238_, new_n1511_ );
or   ( new_n18141_, new_n16224_, new_n1310_ );
and  ( new_n18142_, new_n18141_, new_n18140_ );
or   ( new_n18143_, new_n18142_, new_n16217_ );
and  ( new_n18144_, new_n16226_, RI2b1c4342dbe8_80 );
and  ( new_n18145_, new_n16229_, RI2b1c4342db70_79 );
or   ( new_n18146_, new_n18145_, new_n18144_ );
or   ( new_n18147_, new_n18146_, new_n16234_ );
and  ( new_n18148_, new_n18147_, new_n18143_ );
and  ( new_n18149_, new_n18138_, new_n18129_ );
or   ( new_n18150_, new_n18149_, new_n18148_ );
and  ( new_n18151_, new_n18150_, new_n18139_ );
and  ( new_n18152_, new_n18119_, new_n18088_ );
or   ( new_n18153_, new_n18152_, new_n18151_ );
and  ( new_n18154_, new_n18153_, new_n18120_ );
or   ( new_n18155_, new_n17837_, new_n17836_ );
and  ( new_n18156_, new_n18155_, new_n17977_ );
or   ( new_n18157_, new_n16174_, new_n2119_ );
or   ( new_n18158_, new_n16160_, new_n126_ );
and  ( new_n18159_, new_n18158_, new_n18157_ );
or   ( new_n18160_, new_n18159_, new_n16151_ );
and  ( new_n18161_, new_n16162_, RI2b1c4342dcd8_82 );
and  ( new_n18162_, new_n16165_, RI2b1c4342dc60_81 );
or   ( new_n18163_, new_n18162_, new_n18161_ );
or   ( new_n18164_, new_n18163_, new_n16170_ );
and  ( new_n18165_, new_n18164_, new_n18160_ );
or   ( new_n18166_, new_n16119_, new_n2541_ );
or   ( new_n18167_, new_n16123_, new_n121_ );
and  ( new_n18168_, new_n18167_, new_n18166_ );
or   ( new_n18169_, new_n18168_, new_n16108_ );
and  ( new_n18170_, new_n16132_, RI2b1c4342ddc8_84 );
and  ( new_n18171_, new_n16114_, RI2b1c4342dd50_83 );
or   ( new_n18172_, new_n18171_, new_n18170_ );
or   ( new_n18173_, new_n18172_, new_n16128_ );
and  ( new_n18174_, new_n18173_, new_n18169_ );
and  ( new_n18175_, new_n18174_, new_n18165_ );
or   ( new_n18176_, new_n18174_, new_n18165_ );
or   ( new_n18177_, new_n16115_, new_n2806_ );
and  ( new_n18178_, new_n18177_, new_n18176_ );
or   ( new_n18179_, new_n18178_, new_n18175_ );
and  ( new_n18180_, new_n18179_, new_n18156_ );
or   ( new_n18181_, new_n18179_, new_n18156_ );
or   ( new_n18182_, new_n17962_, new_n17802_ );
or   ( new_n18183_, new_n17959_, new_n17811_ );
and  ( new_n18184_, new_n18183_, new_n18182_ );
or   ( new_n18185_, new_n18184_, new_n17967_ );
and  ( new_n18186_, new_n17963_, new_n17812_ );
or   ( new_n18187_, new_n18186_, new_n17822_ );
and  ( new_n18188_, new_n18187_, new_n18185_ );
and  ( new_n18189_, new_n18188_, new_n18181_ );
or   ( new_n18190_, new_n18189_, new_n18180_ );
and  ( new_n18191_, new_n18190_, new_n18154_ );
or   ( new_n18192_, new_n17945_, new_n17770_ );
or   ( new_n18193_, new_n17948_, new_n17779_ );
and  ( new_n18194_, new_n18193_, new_n18192_ );
or   ( new_n18195_, new_n18194_, new_n17953_ );
and  ( new_n18196_, new_n17949_, new_n17780_ );
or   ( new_n18197_, new_n18196_, new_n17790_ );
and  ( new_n18198_, new_n18197_, new_n18195_ );
or   ( new_n18199_, new_n17932_, new_n17739_ );
or   ( new_n18200_, new_n17935_, new_n17748_ );
and  ( new_n18201_, new_n18200_, new_n18199_ );
or   ( new_n18202_, new_n18201_, new_n17940_ );
and  ( new_n18203_, new_n17936_, new_n17749_ );
or   ( new_n18204_, new_n18203_, new_n17759_ );
and  ( new_n18205_, new_n18204_, new_n18202_ );
or   ( new_n18206_, new_n18205_, new_n18198_ );
or   ( new_n18207_, new_n18190_, new_n18154_ );
and  ( new_n18208_, new_n18207_, new_n18206_ );
or   ( new_n18209_, new_n18208_, new_n18191_ );
and  ( new_n18210_, new_n18209_, new_n18060_ );
or   ( new_n18211_, new_n18209_, new_n18060_ );
or   ( new_n18212_, new_n18007_, new_n17708_ );
or   ( new_n18213_, new_n18004_, new_n17710_ );
and  ( new_n18214_, new_n18213_, new_n18212_ );
or   ( new_n18215_, new_n18214_, new_n18011_ );
and  ( new_n18216_, new_n18008_, new_n17711_ );
or   ( new_n18217_, new_n18216_, new_n17718_ );
and  ( new_n18218_, new_n18217_, new_n18215_ );
and  ( new_n18219_, new_n18218_, new_n18211_ );
or   ( new_n18220_, new_n18219_, new_n18210_ );
and  ( new_n18221_, new_n18220_, new_n18035_ );
or   ( new_n18222_, new_n18220_, new_n18035_ );
or   ( new_n18223_, new_n18014_, new_n17881_ );
or   ( new_n18224_, new_n18002_, new_n17721_ );
and  ( new_n18225_, new_n18224_, new_n18223_ );
or   ( new_n18226_, new_n18225_, new_n18019_ );
and  ( new_n18227_, new_n18015_, new_n17883_ );
or   ( new_n18228_, new_n18227_, new_n17890_ );
and  ( new_n18229_, new_n18228_, new_n18226_ );
and  ( new_n18230_, new_n18229_, new_n18222_ );
or   ( new_n18231_, new_n18230_, new_n18221_ );
or   ( new_n18232_, new_n18231_, new_n18028_ );
or   ( new_n18233_, new_n17700_, new_n17605_ );
or   ( new_n18234_, new_n17697_, new_n17580_ );
and  ( new_n18235_, new_n18234_, new_n18233_ );
or   ( new_n18236_, new_n18235_, new_n17903_ );
and  ( new_n18237_, new_n18021_, new_n17928_ );
or   ( new_n18238_, new_n18237_, new_n17926_ );
and  ( new_n18239_, new_n18238_, new_n18025_ );
or   ( new_n18240_, new_n18239_, new_n17702_ );
and  ( new_n18241_, new_n18240_, new_n18236_ );
or   ( new_n18242_, new_n18241_, new_n18232_ );
or   ( new_n18243_, new_n18242_, new_n17923_ );
and  ( new_n18244_, new_n18243_, new_n17922_ );
or   ( new_n18245_, new_n18244_, new_n17602_ );
and  ( new_n18246_, new_n18245_, new_n17600_ );
and  ( new_n18247_, new_n18241_, new_n18232_ );
or   ( new_n18248_, new_n18247_, new_n17923_ );
or   ( new_n18249_, new_n18248_, new_n17602_ );
or   ( new_n18250_, new_n18227_, new_n18019_ );
or   ( new_n18251_, new_n18225_, new_n17890_ );
and  ( new_n18252_, new_n18251_, new_n18250_ );
or   ( new_n18253_, new_n18033_, new_n17686_ );
or   ( new_n18254_, new_n18031_, new_n17427_ );
and  ( new_n18255_, new_n18254_, new_n18253_ );
or   ( new_n18256_, new_n18255_, new_n18220_ );
or   ( new_n18257_, new_n18040_, new_n17996_ );
or   ( new_n18258_, new_n18038_, new_n17876_ );
and  ( new_n18259_, new_n18258_, new_n18257_ );
or   ( new_n18260_, new_n18047_, new_n17982_ );
or   ( new_n18261_, new_n18045_, new_n17850_ );
and  ( new_n18262_, new_n18261_, new_n18260_ );
or   ( new_n18263_, new_n18262_, new_n18259_ );
or   ( new_n18264_, new_n18055_, new_n17969_ );
or   ( new_n18265_, new_n18053_, new_n17824_ );
and  ( new_n18266_, new_n18265_, new_n18264_ );
and  ( new_n18267_, new_n18262_, new_n18259_ );
or   ( new_n18268_, new_n18267_, new_n18266_ );
and  ( new_n18269_, new_n18268_, new_n18263_ );
or   ( new_n18270_, new_n17973_, new_n17836_ );
or   ( new_n18271_, new_n17976_, new_n17837_ );
and  ( new_n18272_, new_n18271_, new_n18270_ );
or   ( new_n18273_, new_n18163_, new_n16151_ );
or   ( new_n18274_, new_n18159_, new_n16170_ );
and  ( new_n18275_, new_n18274_, new_n18273_ );
or   ( new_n18276_, new_n18172_, new_n16108_ );
or   ( new_n18277_, new_n18168_, new_n16128_ );
and  ( new_n18278_, new_n18277_, new_n18276_ );
or   ( new_n18279_, new_n18278_, new_n18275_ );
and  ( new_n18280_, new_n16102_, RI2b1c4342de40_85 );
and  ( new_n18281_, new_n18278_, new_n18275_ );
or   ( new_n18282_, new_n18281_, new_n18280_ );
and  ( new_n18283_, new_n18282_, new_n18279_ );
or   ( new_n18284_, new_n18283_, new_n18272_ );
or   ( new_n18285_, new_n18186_, new_n17967_ );
or   ( new_n18286_, new_n18184_, new_n17822_ );
and  ( new_n18287_, new_n18286_, new_n18285_ );
and  ( new_n18288_, new_n18283_, new_n18272_ );
or   ( new_n18289_, new_n18288_, new_n18287_ );
and  ( new_n18290_, new_n18289_, new_n18284_ );
or   ( new_n18291_, new_n18104_, new_n16085_ );
or   ( new_n18292_, new_n18100_, new_n16048_ );
and  ( new_n18293_, new_n18292_, new_n18291_ );
or   ( new_n18294_, new_n18095_, new_n16505_ );
or   ( new_n18295_, new_n18091_, new_n16438_ );
and  ( new_n18296_, new_n18295_, new_n18294_ );
or   ( new_n18297_, new_n18296_, new_n18293_ );
or   ( new_n18298_, new_n18114_, new_n16052_ );
or   ( new_n18299_, new_n18110_, new_n16071_ );
and  ( new_n18300_, new_n18299_, new_n18298_ );
and  ( new_n18301_, new_n18296_, new_n18293_ );
or   ( new_n18302_, new_n18301_, new_n18300_ );
and  ( new_n18303_, new_n18302_, new_n18297_ );
nand ( new_n18304_, new_n18063_, new_n138_ );
and  ( new_n18305_, new_n18304_, RI2b1c4342c0b8_22 );
nand ( new_n18306_, new_n18061_, new_n138_ );
and  ( new_n18307_, new_n18306_, RI2b1c4342c130_23 );
and  ( new_n18308_, new_n18307_, new_n18305_ );
or   ( new_n18309_, new_n18308_, new_n17234_ );
or   ( new_n18310_, new_n18073_, new_n17238_ );
or   ( new_n18311_, new_n18069_, new_n17650_ );
and  ( new_n18312_, new_n18311_, new_n18310_ );
or   ( new_n18313_, new_n18312_, new_n18309_ );
or   ( new_n18314_, new_n18083_, new_n16814_ );
or   ( new_n18315_, new_n18079_, new_n17142_ );
and  ( new_n18316_, new_n18315_, new_n18314_ );
and  ( new_n18317_, new_n18312_, new_n18309_ );
or   ( new_n18318_, new_n18317_, new_n18316_ );
and  ( new_n18319_, new_n18318_, new_n18313_ );
or   ( new_n18320_, new_n18319_, new_n18303_ );
or   ( new_n18321_, new_n18127_, new_n16009_ );
or   ( new_n18322_, new_n18123_, new_n16029_ );
and  ( new_n18323_, new_n18322_, new_n18321_ );
or   ( new_n18324_, new_n18136_, new_n16186_ );
or   ( new_n18325_, new_n18132_, new_n16204_ );
and  ( new_n18326_, new_n18325_, new_n18324_ );
or   ( new_n18327_, new_n18326_, new_n18323_ );
or   ( new_n18328_, new_n18146_, new_n16217_ );
or   ( new_n18329_, new_n18142_, new_n16234_ );
and  ( new_n18330_, new_n18329_, new_n18328_ );
and  ( new_n18331_, new_n18326_, new_n18323_ );
or   ( new_n18332_, new_n18331_, new_n18330_ );
and  ( new_n18333_, new_n18332_, new_n18327_ );
and  ( new_n18334_, new_n18319_, new_n18303_ );
or   ( new_n18335_, new_n18334_, new_n18333_ );
and  ( new_n18336_, new_n18335_, new_n18320_ );
or   ( new_n18337_, new_n18336_, new_n18290_ );
or   ( new_n18338_, new_n18196_, new_n17953_ );
or   ( new_n18339_, new_n18194_, new_n17790_ );
and  ( new_n18340_, new_n18339_, new_n18338_ );
or   ( new_n18341_, new_n18203_, new_n17940_ );
or   ( new_n18342_, new_n18201_, new_n17759_ );
and  ( new_n18343_, new_n18342_, new_n18341_ );
and  ( new_n18344_, new_n18343_, new_n18340_ );
and  ( new_n18345_, new_n18336_, new_n18290_ );
or   ( new_n18346_, new_n18345_, new_n18344_ );
and  ( new_n18347_, new_n18346_, new_n18337_ );
or   ( new_n18348_, new_n18347_, new_n18269_ );
or   ( new_n18349_, new_n18216_, new_n18011_ );
or   ( new_n18350_, new_n18214_, new_n17718_ );
and  ( new_n18351_, new_n18350_, new_n18349_ );
and  ( new_n18352_, new_n18347_, new_n18269_ );
or   ( new_n18353_, new_n18352_, new_n18351_ );
and  ( new_n18354_, new_n18353_, new_n18348_ );
or   ( new_n18355_, new_n18354_, new_n18035_ );
and  ( new_n18356_, new_n18355_, new_n18256_ );
or   ( new_n18357_, new_n18356_, new_n18252_ );
or   ( new_n18358_, new_n18354_, new_n18255_ );
and  ( new_n18359_, new_n18358_, new_n18222_ );
or   ( new_n18360_, new_n18359_, new_n18229_ );
and  ( new_n18361_, new_n18360_, new_n18357_ );
or   ( new_n18362_, new_n18343_, new_n18198_ );
or   ( new_n18363_, new_n18340_, new_n18205_ );
and  ( new_n18364_, new_n18363_, new_n18362_ );
or   ( new_n18365_, new_n18272_, new_n18179_ );
or   ( new_n18366_, new_n18283_, new_n18156_ );
and  ( new_n18367_, new_n18366_, new_n18365_ );
or   ( new_n18368_, new_n18367_, new_n18287_ );
and  ( new_n18369_, new_n18284_, new_n18181_ );
or   ( new_n18370_, new_n18369_, new_n18188_ );
and  ( new_n18371_, new_n18370_, new_n18368_ );
or   ( new_n18372_, new_n18371_, new_n18364_ );
and  ( new_n18373_, new_n18371_, new_n18364_ );
or   ( new_n18374_, new_n18303_, new_n18088_ );
or   ( new_n18375_, new_n18319_, new_n18119_ );
and  ( new_n18376_, new_n18375_, new_n18374_ );
or   ( new_n18377_, new_n18376_, new_n18333_ );
and  ( new_n18378_, new_n18320_, new_n18120_ );
or   ( new_n18379_, new_n18378_, new_n18151_ );
and  ( new_n18380_, new_n18379_, new_n18377_ );
or   ( new_n18381_, new_n18380_, new_n18373_ );
and  ( new_n18382_, new_n18381_, new_n18372_ );
or   ( new_n18383_, new_n18307_, new_n18305_ );
and  ( new_n18384_, new_n18383_, new_n18065_ );
or   ( new_n18385_, new_n18305_, new_n17234_ );
or   ( new_n18386_, new_n18064_, new_n17648_ );
and  ( new_n18387_, new_n18386_, new_n18385_ );
or   ( new_n18388_, new_n18387_, new_n18384_ );
or   ( new_n18389_, new_n18388_, new_n99_ );
or   ( new_n18390_, new_n18389_, new_n18066_ );
or   ( new_n18391_, new_n18305_, new_n17648_ );
or   ( new_n18392_, new_n18064_, new_n17234_ );
or   ( new_n18393_, new_n18307_, new_n18064_ );
or   ( new_n18394_, new_n18305_, new_n18062_ );
and  ( new_n18395_, new_n18394_, new_n18393_ );
and  ( new_n18396_, new_n18395_, new_n18392_ );
and  ( new_n18397_, new_n18396_, new_n18391_ );
and  ( new_n18398_, new_n18397_, RI2b1c4342d4e0_65 );
or   ( new_n18399_, new_n18398_, new_n18309_ );
and  ( new_n18400_, new_n18399_, new_n18390_ );
or   ( new_n18401_, new_n17727_, new_n112_ );
or   ( new_n18402_, new_n17734_, new_n526_ );
and  ( new_n18403_, new_n18402_, new_n18401_ );
or   ( new_n18404_, new_n18403_, new_n17238_ );
and  ( new_n18405_, new_n17736_, RI2b1c4342d5d0_67 );
and  ( new_n18406_, new_n17723_, RI2b1c4342d558_66 );
or   ( new_n18407_, new_n18406_, new_n18405_ );
or   ( new_n18408_, new_n18407_, new_n17650_ );
and  ( new_n18409_, new_n18408_, new_n18404_ );
or   ( new_n18410_, new_n18409_, new_n18400_ );
and  ( new_n18411_, new_n18409_, new_n18400_ );
or   ( new_n18412_, new_n17244_, new_n591_ );
or   ( new_n18413_, new_n17248_, new_n612_ );
and  ( new_n18414_, new_n18413_, new_n18412_ );
or   ( new_n18415_, new_n18414_, new_n16814_ );
and  ( new_n18416_, new_n17255_, RI2b1c4342d6c0_69 );
and  ( new_n18417_, new_n17240_, RI2b1c4342d648_68 );
or   ( new_n18418_, new_n18417_, new_n18416_ );
or   ( new_n18419_, new_n18418_, new_n17142_ );
and  ( new_n18420_, new_n18419_, new_n18415_ );
or   ( new_n18421_, new_n18420_, new_n18411_ );
and  ( new_n18422_, new_n18421_, new_n18410_ );
or   ( new_n18423_, new_n16607_, new_n110_ );
or   ( new_n18424_, new_n16613_, new_n755_ );
and  ( new_n18425_, new_n18424_, new_n18423_ );
or   ( new_n18426_, new_n18425_, new_n16505_ );
and  ( new_n18427_, new_n16616_, RI2b1c4342d7b0_71 );
and  ( new_n18428_, new_n16603_, RI2b1c4342d738_70 );
or   ( new_n18429_, new_n18428_, new_n18427_ );
or   ( new_n18430_, new_n18429_, new_n16438_ );
and  ( new_n18431_, new_n18430_, new_n18426_ );
or   ( new_n18432_, new_n16366_, new_n105_ );
or   ( new_n18433_, new_n16355_, new_n806_ );
and  ( new_n18434_, new_n18433_, new_n18432_ );
or   ( new_n18435_, new_n18434_, new_n16085_ );
and  ( new_n18436_, new_n16358_, RI2b1c4342d8a0_73 );
and  ( new_n18437_, new_n16362_, RI2b1c4342d828_72 );
or   ( new_n18438_, new_n18437_, new_n18436_ );
or   ( new_n18439_, new_n18438_, new_n16048_ );
and  ( new_n18440_, new_n18439_, new_n18435_ );
or   ( new_n18441_, new_n18440_, new_n18431_ );
and  ( new_n18442_, new_n18440_, new_n18431_ );
or   ( new_n18443_, new_n16075_, new_n843_ );
or   ( new_n18444_, new_n16060_, new_n859_ );
and  ( new_n18445_, new_n18444_, new_n18443_ );
or   ( new_n18446_, new_n18445_, new_n16052_ );
and  ( new_n18447_, new_n16063_, RI2b1c4342d990_75 );
and  ( new_n18448_, new_n16066_, RI2b1c4342d918_74 );
or   ( new_n18449_, new_n18448_, new_n18447_ );
or   ( new_n18450_, new_n18449_, new_n16071_ );
and  ( new_n18451_, new_n18450_, new_n18446_ );
or   ( new_n18452_, new_n18451_, new_n18442_ );
and  ( new_n18453_, new_n18452_, new_n18441_ );
or   ( new_n18454_, new_n18453_, new_n18422_ );
and  ( new_n18455_, new_n18453_, new_n18422_ );
or   ( new_n18456_, new_n16033_, new_n1004_ );
or   ( new_n18457_, new_n16017_, new_n886_ );
and  ( new_n18458_, new_n18457_, new_n18456_ );
or   ( new_n18459_, new_n18458_, new_n16009_ );
and  ( new_n18460_, new_n16021_, RI2b1c4342da80_77 );
and  ( new_n18461_, new_n16024_, RI2b1c4342da08_76 );
or   ( new_n18462_, new_n18461_, new_n18460_ );
or   ( new_n18463_, new_n18462_, new_n16029_ );
and  ( new_n18464_, new_n18463_, new_n18459_ );
or   ( new_n18465_, new_n16208_, new_n1310_ );
or   ( new_n18466_, new_n16194_, new_n1002_ );
and  ( new_n18467_, new_n18466_, new_n18465_ );
or   ( new_n18468_, new_n18467_, new_n16186_ );
and  ( new_n18469_, new_n16196_, RI2b1c4342db70_79 );
and  ( new_n18470_, new_n16199_, RI2b1c4342daf8_78 );
or   ( new_n18471_, new_n18470_, new_n18469_ );
or   ( new_n18472_, new_n18471_, new_n16204_ );
and  ( new_n18473_, new_n18472_, new_n18468_ );
or   ( new_n18474_, new_n18473_, new_n18464_ );
and  ( new_n18475_, new_n18473_, new_n18464_ );
or   ( new_n18476_, new_n16238_, new_n126_ );
or   ( new_n18477_, new_n16224_, new_n1511_ );
and  ( new_n18478_, new_n18477_, new_n18476_ );
or   ( new_n18479_, new_n18478_, new_n16217_ );
and  ( new_n18480_, new_n16226_, RI2b1c4342dc60_81 );
and  ( new_n18481_, new_n16229_, RI2b1c4342dbe8_80 );
or   ( new_n18482_, new_n18481_, new_n18480_ );
or   ( new_n18483_, new_n18482_, new_n16234_ );
and  ( new_n18484_, new_n18483_, new_n18479_ );
or   ( new_n18485_, new_n18484_, new_n18475_ );
and  ( new_n18486_, new_n18485_, new_n18474_ );
or   ( new_n18487_, new_n18486_, new_n18455_ );
and  ( new_n18488_, new_n18487_, new_n18454_ );
or   ( new_n18489_, new_n18278_, new_n18165_ );
or   ( new_n18490_, new_n18275_, new_n18174_ );
and  ( new_n18491_, new_n18490_, new_n18489_ );
or   ( new_n18492_, new_n18491_, new_n18280_ );
and  ( new_n18493_, new_n18279_, new_n18176_ );
or   ( new_n18494_, new_n18493_, new_n18177_ );
and  ( new_n18495_, new_n18494_, new_n18492_ );
or   ( new_n18496_, new_n16174_, new_n121_ );
or   ( new_n18497_, new_n16160_, new_n2119_ );
and  ( new_n18498_, new_n18497_, new_n18496_ );
or   ( new_n18499_, new_n18498_, new_n16151_ );
and  ( new_n18500_, new_n16162_, RI2b1c4342dd50_83 );
and  ( new_n18501_, new_n16165_, RI2b1c4342dcd8_82 );
or   ( new_n18502_, new_n18501_, new_n18500_ );
or   ( new_n18503_, new_n18502_, new_n16170_ );
and  ( new_n18504_, new_n18503_, new_n18499_ );
or   ( new_n18505_, new_n16119_, new_n2806_ );
or   ( new_n18506_, new_n16123_, new_n2541_ );
and  ( new_n18507_, new_n18506_, new_n18505_ );
or   ( new_n18508_, new_n18507_, new_n16108_ );
and  ( new_n18509_, new_n16132_, RI2b1c4342de40_85 );
and  ( new_n18510_, new_n16114_, RI2b1c4342ddc8_84 );
or   ( new_n18511_, new_n18510_, new_n18509_ );
or   ( new_n18512_, new_n18511_, new_n16128_ );
and  ( new_n18513_, new_n18512_, new_n18508_ );
and  ( new_n18514_, new_n18513_, new_n18504_ );
or   ( new_n18515_, new_n18513_, new_n18504_ );
or   ( new_n18516_, new_n16115_, new_n3239_ );
and  ( new_n18517_, new_n18516_, new_n18515_ );
or   ( new_n18518_, new_n18517_, new_n18514_ );
and  ( new_n18519_, new_n18518_, new_n18495_ );
or   ( new_n18520_, new_n18518_, new_n18495_ );
or   ( new_n18521_, new_n18326_, new_n18129_ );
or   ( new_n18522_, new_n18323_, new_n18138_ );
and  ( new_n18523_, new_n18522_, new_n18521_ );
or   ( new_n18524_, new_n18523_, new_n18330_ );
and  ( new_n18525_, new_n18327_, new_n18139_ );
or   ( new_n18526_, new_n18525_, new_n18148_ );
and  ( new_n18527_, new_n18526_, new_n18524_ );
and  ( new_n18528_, new_n18527_, new_n18520_ );
or   ( new_n18529_, new_n18528_, new_n18519_ );
and  ( new_n18530_, new_n18529_, new_n18488_ );
or   ( new_n18531_, new_n18529_, new_n18488_ );
or   ( new_n18532_, new_n18293_, new_n18097_ );
or   ( new_n18533_, new_n18296_, new_n18106_ );
and  ( new_n18534_, new_n18533_, new_n18532_ );
or   ( new_n18535_, new_n18534_, new_n18300_ );
and  ( new_n18536_, new_n18297_, new_n18107_ );
or   ( new_n18537_, new_n18536_, new_n18116_ );
and  ( new_n18538_, new_n18537_, new_n18535_ );
or   ( new_n18539_, new_n18312_, new_n18066_ );
or   ( new_n18540_, new_n18309_, new_n18075_ );
and  ( new_n18541_, new_n18540_, new_n18539_ );
or   ( new_n18542_, new_n18541_, new_n18316_ );
and  ( new_n18543_, new_n18313_, new_n18076_ );
or   ( new_n18544_, new_n18543_, new_n18085_ );
and  ( new_n18545_, new_n18544_, new_n18542_ );
or   ( new_n18546_, new_n18545_, new_n18538_ );
and  ( new_n18547_, new_n18546_, new_n18531_ );
or   ( new_n18548_, new_n18547_, new_n18530_ );
and  ( new_n18549_, new_n18548_, new_n18382_ );
or   ( new_n18550_, new_n18548_, new_n18382_ );
or   ( new_n18551_, new_n18262_, new_n18042_ );
or   ( new_n18552_, new_n18259_, new_n18049_ );
and  ( new_n18553_, new_n18552_, new_n18551_ );
or   ( new_n18554_, new_n18553_, new_n18266_ );
and  ( new_n18555_, new_n18263_, new_n18050_ );
or   ( new_n18556_, new_n18555_, new_n18057_ );
and  ( new_n18557_, new_n18556_, new_n18554_ );
and  ( new_n18558_, new_n18557_, new_n18550_ );
or   ( new_n18559_, new_n18558_, new_n18549_ );
or   ( new_n18560_, new_n17985_, new_n17827_ );
or   ( new_n18561_, new_n17972_, new_n17852_ );
and  ( new_n18562_, new_n18561_, new_n18560_ );
or   ( new_n18563_, new_n18562_, new_n17999_ );
and  ( new_n18564_, new_n17986_, new_n17854_ );
or   ( new_n18565_, new_n18564_, new_n17879_ );
and  ( new_n18566_, new_n18565_, new_n18563_ );
and  ( new_n18567_, new_n18566_, new_n18559_ );
or   ( new_n18568_, new_n18269_, new_n18209_ );
or   ( new_n18569_, new_n18347_, new_n18060_ );
and  ( new_n18570_, new_n18569_, new_n18568_ );
or   ( new_n18571_, new_n18570_, new_n18351_ );
and  ( new_n18572_, new_n18348_, new_n18211_ );
or   ( new_n18573_, new_n18572_, new_n18218_ );
and  ( new_n18574_, new_n18573_, new_n18571_ );
or   ( new_n18575_, new_n18566_, new_n18559_ );
and  ( new_n18576_, new_n18575_, new_n18574_ );
or   ( new_n18577_, new_n18576_, new_n18567_ );
or   ( new_n18578_, new_n18577_, new_n18361_ );
or   ( new_n18579_, new_n18026_, new_n17926_ );
or   ( new_n18580_, new_n18023_, new_n17901_ );
and  ( new_n18581_, new_n18580_, new_n18579_ );
or   ( new_n18582_, new_n18581_, new_n18231_ );
and  ( new_n18583_, new_n18354_, new_n18255_ );
or   ( new_n18584_, new_n18583_, new_n18252_ );
and  ( new_n18585_, new_n18584_, new_n18358_ );
or   ( new_n18586_, new_n18585_, new_n18028_ );
and  ( new_n18587_, new_n18586_, new_n18582_ );
or   ( new_n18588_, new_n18587_, new_n18578_ );
and  ( new_n18589_, new_n18587_, new_n18578_ );
or   ( new_n18590_, new_n18572_, new_n18351_ );
or   ( new_n18591_, new_n18570_, new_n18218_ );
and  ( new_n18592_, new_n18591_, new_n18590_ );
or   ( new_n18593_, new_n18564_, new_n17999_ );
or   ( new_n18594_, new_n18562_, new_n17879_ );
and  ( new_n18595_, new_n18594_, new_n18593_ );
or   ( new_n18596_, new_n18595_, new_n18559_ );
or   ( new_n18597_, new_n18398_, new_n18066_ );
or   ( new_n18598_, new_n18389_, new_n18309_ );
and  ( new_n18599_, new_n18598_, new_n18597_ );
or   ( new_n18600_, new_n18407_, new_n17238_ );
or   ( new_n18601_, new_n18403_, new_n17650_ );
and  ( new_n18602_, new_n18601_, new_n18600_ );
or   ( new_n18603_, new_n18602_, new_n18599_ );
and  ( new_n18604_, new_n18602_, new_n18599_ );
or   ( new_n18605_, new_n18418_, new_n16814_ );
or   ( new_n18606_, new_n18414_, new_n17142_ );
and  ( new_n18607_, new_n18606_, new_n18605_ );
or   ( new_n18608_, new_n18607_, new_n18604_ );
and  ( new_n18609_, new_n18608_, new_n18603_ );
or   ( new_n18610_, new_n18429_, new_n16505_ );
or   ( new_n18611_, new_n18425_, new_n16438_ );
and  ( new_n18612_, new_n18611_, new_n18610_ );
or   ( new_n18613_, new_n18438_, new_n16085_ );
or   ( new_n18614_, new_n18434_, new_n16048_ );
and  ( new_n18615_, new_n18614_, new_n18613_ );
or   ( new_n18616_, new_n18615_, new_n18612_ );
and  ( new_n18617_, new_n18615_, new_n18612_ );
or   ( new_n18618_, new_n18449_, new_n16052_ );
or   ( new_n18619_, new_n18445_, new_n16071_ );
and  ( new_n18620_, new_n18619_, new_n18618_ );
or   ( new_n18621_, new_n18620_, new_n18617_ );
and  ( new_n18622_, new_n18621_, new_n18616_ );
or   ( new_n18623_, new_n18622_, new_n18609_ );
and  ( new_n18624_, new_n18622_, new_n18609_ );
or   ( new_n18625_, new_n18462_, new_n16009_ );
or   ( new_n18626_, new_n18458_, new_n16029_ );
and  ( new_n18627_, new_n18626_, new_n18625_ );
or   ( new_n18628_, new_n18471_, new_n16186_ );
or   ( new_n18629_, new_n18467_, new_n16204_ );
and  ( new_n18630_, new_n18629_, new_n18628_ );
or   ( new_n18631_, new_n18630_, new_n18627_ );
and  ( new_n18632_, new_n18630_, new_n18627_ );
or   ( new_n18633_, new_n18482_, new_n16217_ );
or   ( new_n18634_, new_n18478_, new_n16234_ );
and  ( new_n18635_, new_n18634_, new_n18633_ );
or   ( new_n18636_, new_n18635_, new_n18632_ );
and  ( new_n18637_, new_n18636_, new_n18631_ );
or   ( new_n18638_, new_n18637_, new_n18624_ );
and  ( new_n18639_, new_n18638_, new_n18623_ );
or   ( new_n18640_, new_n18493_, new_n18280_ );
or   ( new_n18641_, new_n18491_, new_n18177_ );
and  ( new_n18642_, new_n18641_, new_n18640_ );
or   ( new_n18643_, new_n18502_, new_n16151_ );
or   ( new_n18644_, new_n18498_, new_n16170_ );
and  ( new_n18645_, new_n18644_, new_n18643_ );
or   ( new_n18646_, new_n18511_, new_n16108_ );
or   ( new_n18647_, new_n18507_, new_n16128_ );
and  ( new_n18648_, new_n18647_, new_n18646_ );
or   ( new_n18649_, new_n18648_, new_n18645_ );
and  ( new_n18650_, new_n18648_, new_n18645_ );
and  ( new_n18651_, new_n16102_, RI2b1c4342deb8_86 );
or   ( new_n18652_, new_n18651_, new_n18650_ );
and  ( new_n18653_, new_n18652_, new_n18649_ );
or   ( new_n18654_, new_n18653_, new_n18642_ );
and  ( new_n18655_, new_n18653_, new_n18642_ );
or   ( new_n18656_, new_n18525_, new_n18330_ );
or   ( new_n18657_, new_n18523_, new_n18148_ );
and  ( new_n18658_, new_n18657_, new_n18656_ );
or   ( new_n18659_, new_n18658_, new_n18655_ );
and  ( new_n18660_, new_n18659_, new_n18654_ );
or   ( new_n18661_, new_n18660_, new_n18639_ );
and  ( new_n18662_, new_n18660_, new_n18639_ );
or   ( new_n18663_, new_n18536_, new_n18300_ );
or   ( new_n18664_, new_n18534_, new_n18116_ );
and  ( new_n18665_, new_n18664_, new_n18663_ );
or   ( new_n18666_, new_n18543_, new_n18316_ );
or   ( new_n18667_, new_n18541_, new_n18085_ );
and  ( new_n18668_, new_n18667_, new_n18666_ );
and  ( new_n18669_, new_n18668_, new_n18665_ );
or   ( new_n18670_, new_n18669_, new_n18662_ );
and  ( new_n18671_, new_n18670_, new_n18661_ );
or   ( new_n18672_, new_n18343_, new_n18340_ );
and  ( new_n18673_, new_n18672_, new_n18206_ );
or   ( new_n18674_, new_n18369_, new_n18287_ );
or   ( new_n18675_, new_n18367_, new_n18188_ );
and  ( new_n18676_, new_n18675_, new_n18674_ );
or   ( new_n18677_, new_n18676_, new_n18673_ );
and  ( new_n18678_, new_n18676_, new_n18673_ );
or   ( new_n18679_, new_n18378_, new_n18333_ );
or   ( new_n18680_, new_n18376_, new_n18151_ );
and  ( new_n18681_, new_n18680_, new_n18679_ );
or   ( new_n18682_, new_n18681_, new_n18678_ );
and  ( new_n18683_, new_n18682_, new_n18677_ );
or   ( new_n18684_, new_n18683_, new_n18671_ );
or   ( new_n18685_, new_n18555_, new_n18266_ );
or   ( new_n18686_, new_n18553_, new_n18057_ );
and  ( new_n18687_, new_n18686_, new_n18685_ );
and  ( new_n18688_, new_n18683_, new_n18671_ );
or   ( new_n18689_, new_n18688_, new_n18687_ );
and  ( new_n18690_, new_n18689_, new_n18684_ );
or   ( new_n18691_, new_n18690_, new_n18566_ );
and  ( new_n18692_, new_n18691_, new_n18596_ );
or   ( new_n18693_, new_n18692_, new_n18592_ );
or   ( new_n18694_, new_n18690_, new_n18595_ );
and  ( new_n18695_, new_n18694_, new_n18575_ );
or   ( new_n18696_, new_n18695_, new_n18574_ );
and  ( new_n18697_, new_n18696_, new_n18693_ );
or   ( new_n18698_, new_n18648_, new_n18504_ );
or   ( new_n18699_, new_n18645_, new_n18513_ );
and  ( new_n18700_, new_n18699_, new_n18698_ );
or   ( new_n18701_, new_n18700_, new_n18651_ );
and  ( new_n18702_, new_n18649_, new_n18515_ );
or   ( new_n18703_, new_n18702_, new_n18516_ );
and  ( new_n18704_, new_n18703_, new_n18701_ );
or   ( new_n18705_, new_n16238_, new_n2119_ );
or   ( new_n18706_, new_n16224_, new_n126_ );
and  ( new_n18707_, new_n18706_, new_n18705_ );
or   ( new_n18708_, new_n18707_, new_n16217_ );
and  ( new_n18709_, new_n16226_, RI2b1c4342dcd8_82 );
and  ( new_n18710_, new_n16229_, RI2b1c4342dc60_81 );
or   ( new_n18711_, new_n18710_, new_n18709_ );
or   ( new_n18712_, new_n18711_, new_n16234_ );
and  ( new_n18713_, new_n18712_, new_n18708_ );
or   ( new_n18714_, new_n16174_, new_n2541_ );
or   ( new_n18715_, new_n16160_, new_n121_ );
and  ( new_n18716_, new_n18715_, new_n18714_ );
or   ( new_n18717_, new_n18716_, new_n16151_ );
and  ( new_n18718_, new_n16162_, RI2b1c4342ddc8_84 );
and  ( new_n18719_, new_n16165_, RI2b1c4342dd50_83 );
or   ( new_n18720_, new_n18719_, new_n18718_ );
or   ( new_n18721_, new_n18720_, new_n16170_ );
and  ( new_n18722_, new_n18721_, new_n18717_ );
or   ( new_n18723_, new_n18722_, new_n18713_ );
and  ( new_n18724_, new_n18722_, new_n18713_ );
or   ( new_n18725_, new_n16119_, new_n3239_ );
or   ( new_n18726_, new_n16123_, new_n2806_ );
and  ( new_n18727_, new_n18726_, new_n18725_ );
or   ( new_n18728_, new_n18727_, new_n16108_ );
and  ( new_n18729_, new_n16132_, RI2b1c4342deb8_86 );
and  ( new_n18730_, new_n16114_, RI2b1c4342de40_85 );
or   ( new_n18731_, new_n18730_, new_n18729_ );
or   ( new_n18732_, new_n18731_, new_n16128_ );
and  ( new_n18733_, new_n18732_, new_n18728_ );
or   ( new_n18734_, new_n18733_, new_n18724_ );
and  ( new_n18735_, new_n18734_, new_n18723_ );
and  ( new_n18736_, new_n18735_, new_n18704_ );
xor  ( new_n18737_, new_n3535_, new_n3685_ );
or   ( new_n18738_, new_n18737_, new_n310_ );
xor  ( new_n18739_, new_n3542_, new_n231_ );
or   ( new_n18740_, new_n18739_, new_n307_ );
or   ( new_n18741_, new_n18740_, new_n18738_ );
and  ( new_n18742_, new_n18741_, new_n18307_ );
or   ( new_n18743_, new_n18388_, new_n526_ );
or   ( new_n18744_, new_n18395_, new_n99_ );
and  ( new_n18745_, new_n18744_, new_n18743_ );
or   ( new_n18746_, new_n18745_, new_n18066_ );
and  ( new_n18747_, new_n18397_, RI2b1c4342d558_66 );
and  ( new_n18748_, new_n18384_, RI2b1c4342d4e0_65 );
or   ( new_n18749_, new_n18748_, new_n18747_ );
or   ( new_n18750_, new_n18749_, new_n18309_ );
and  ( new_n18751_, new_n18750_, new_n18746_ );
or   ( new_n18752_, new_n18751_, new_n18742_ );
and  ( new_n18753_, new_n18751_, new_n18742_ );
or   ( new_n18754_, new_n17727_, new_n612_ );
or   ( new_n18755_, new_n17734_, new_n112_ );
and  ( new_n18756_, new_n18755_, new_n18754_ );
or   ( new_n18757_, new_n18756_, new_n17238_ );
and  ( new_n18758_, new_n17736_, RI2b1c4342d648_68 );
and  ( new_n18759_, new_n17723_, RI2b1c4342d5d0_67 );
or   ( new_n18760_, new_n18759_, new_n18758_ );
or   ( new_n18761_, new_n18760_, new_n17650_ );
and  ( new_n18762_, new_n18761_, new_n18757_ );
or   ( new_n18763_, new_n18762_, new_n18753_ );
and  ( new_n18764_, new_n18763_, new_n18752_ );
or   ( new_n18765_, new_n17244_, new_n755_ );
or   ( new_n18766_, new_n17248_, new_n591_ );
and  ( new_n18767_, new_n18766_, new_n18765_ );
or   ( new_n18768_, new_n18767_, new_n16814_ );
and  ( new_n18769_, new_n17255_, RI2b1c4342d738_70 );
and  ( new_n18770_, new_n17240_, RI2b1c4342d6c0_69 );
or   ( new_n18771_, new_n18770_, new_n18769_ );
or   ( new_n18772_, new_n18771_, new_n17142_ );
and  ( new_n18773_, new_n18772_, new_n18768_ );
or   ( new_n18774_, new_n16607_, new_n806_ );
or   ( new_n18775_, new_n16613_, new_n110_ );
and  ( new_n18776_, new_n18775_, new_n18774_ );
or   ( new_n18777_, new_n18776_, new_n16505_ );
and  ( new_n18778_, new_n16616_, RI2b1c4342d828_72 );
and  ( new_n18779_, new_n16603_, RI2b1c4342d7b0_71 );
or   ( new_n18780_, new_n18779_, new_n18778_ );
or   ( new_n18781_, new_n18780_, new_n16438_ );
and  ( new_n18782_, new_n18781_, new_n18777_ );
or   ( new_n18783_, new_n18782_, new_n18773_ );
and  ( new_n18784_, new_n18782_, new_n18773_ );
or   ( new_n18785_, new_n16366_, new_n859_ );
or   ( new_n18786_, new_n16355_, new_n105_ );
and  ( new_n18787_, new_n18786_, new_n18785_ );
or   ( new_n18788_, new_n18787_, new_n16085_ );
and  ( new_n18789_, new_n16358_, RI2b1c4342d918_74 );
and  ( new_n18790_, new_n16362_, RI2b1c4342d8a0_73 );
or   ( new_n18791_, new_n18790_, new_n18789_ );
or   ( new_n18792_, new_n18791_, new_n16048_ );
and  ( new_n18793_, new_n18792_, new_n18788_ );
or   ( new_n18794_, new_n18793_, new_n18784_ );
and  ( new_n18795_, new_n18794_, new_n18783_ );
or   ( new_n18796_, new_n18795_, new_n18764_ );
and  ( new_n18797_, new_n18795_, new_n18764_ );
or   ( new_n18798_, new_n16075_, new_n886_ );
or   ( new_n18799_, new_n16060_, new_n843_ );
and  ( new_n18800_, new_n18799_, new_n18798_ );
or   ( new_n18801_, new_n18800_, new_n16052_ );
and  ( new_n18802_, new_n16063_, RI2b1c4342da08_76 );
and  ( new_n18803_, new_n16066_, RI2b1c4342d990_75 );
or   ( new_n18804_, new_n18803_, new_n18802_ );
or   ( new_n18805_, new_n18804_, new_n16071_ );
and  ( new_n18806_, new_n18805_, new_n18801_ );
or   ( new_n18807_, new_n16033_, new_n1002_ );
or   ( new_n18808_, new_n16017_, new_n1004_ );
and  ( new_n18809_, new_n18808_, new_n18807_ );
or   ( new_n18810_, new_n18809_, new_n16009_ );
and  ( new_n18811_, new_n16021_, RI2b1c4342daf8_78 );
and  ( new_n18812_, new_n16024_, RI2b1c4342da80_77 );
or   ( new_n18813_, new_n18812_, new_n18811_ );
or   ( new_n18814_, new_n18813_, new_n16029_ );
and  ( new_n18815_, new_n18814_, new_n18810_ );
or   ( new_n18816_, new_n18815_, new_n18806_ );
and  ( new_n18817_, new_n18815_, new_n18806_ );
or   ( new_n18818_, new_n16208_, new_n1511_ );
or   ( new_n18819_, new_n16194_, new_n1310_ );
and  ( new_n18820_, new_n18819_, new_n18818_ );
or   ( new_n18821_, new_n18820_, new_n16186_ );
and  ( new_n18822_, new_n16196_, RI2b1c4342dbe8_80 );
and  ( new_n18823_, new_n16199_, RI2b1c4342db70_79 );
or   ( new_n18824_, new_n18823_, new_n18822_ );
or   ( new_n18825_, new_n18824_, new_n16204_ );
and  ( new_n18826_, new_n18825_, new_n18821_ );
or   ( new_n18827_, new_n18826_, new_n18817_ );
and  ( new_n18828_, new_n18827_, new_n18816_ );
or   ( new_n18829_, new_n18828_, new_n18797_ );
and  ( new_n18830_, new_n18829_, new_n18796_ );
or   ( new_n18831_, new_n18830_, new_n18736_ );
and  ( new_n18832_, new_n18830_, new_n18736_ );
or   ( new_n18833_, new_n18630_, new_n18464_ );
or   ( new_n18834_, new_n18627_, new_n18473_ );
and  ( new_n18835_, new_n18834_, new_n18833_ );
or   ( new_n18836_, new_n18835_, new_n18635_ );
and  ( new_n18837_, new_n18631_, new_n18474_ );
or   ( new_n18838_, new_n18837_, new_n18484_ );
and  ( new_n18839_, new_n18838_, new_n18836_ );
or   ( new_n18840_, new_n18615_, new_n18431_ );
or   ( new_n18841_, new_n18612_, new_n18440_ );
and  ( new_n18842_, new_n18841_, new_n18840_ );
or   ( new_n18843_, new_n18842_, new_n18620_ );
and  ( new_n18844_, new_n18616_, new_n18441_ );
or   ( new_n18845_, new_n18844_, new_n18451_ );
and  ( new_n18846_, new_n18845_, new_n18843_ );
or   ( new_n18847_, new_n18846_, new_n18839_ );
and  ( new_n18848_, new_n18846_, new_n18839_ );
or   ( new_n18849_, new_n18602_, new_n18400_ );
or   ( new_n18850_, new_n18599_, new_n18409_ );
and  ( new_n18851_, new_n18850_, new_n18849_ );
or   ( new_n18852_, new_n18851_, new_n18607_ );
and  ( new_n18853_, new_n18603_, new_n18410_ );
or   ( new_n18854_, new_n18853_, new_n18420_ );
and  ( new_n18855_, new_n18854_, new_n18852_ );
or   ( new_n18856_, new_n18855_, new_n18848_ );
and  ( new_n18857_, new_n18856_, new_n18847_ );
or   ( new_n18858_, new_n18857_, new_n18832_ );
and  ( new_n18859_, new_n18858_, new_n18831_ );
or   ( new_n18860_, new_n18668_, new_n18538_ );
or   ( new_n18861_, new_n18665_, new_n18545_ );
and  ( new_n18862_, new_n18861_, new_n18860_ );
or   ( new_n18863_, new_n18642_, new_n18518_ );
or   ( new_n18864_, new_n18653_, new_n18495_ );
and  ( new_n18865_, new_n18864_, new_n18863_ );
or   ( new_n18866_, new_n18865_, new_n18658_ );
and  ( new_n18867_, new_n18654_, new_n18520_ );
or   ( new_n18868_, new_n18867_, new_n18527_ );
and  ( new_n18869_, new_n18868_, new_n18866_ );
or   ( new_n18870_, new_n18869_, new_n18862_ );
and  ( new_n18871_, new_n18869_, new_n18862_ );
or   ( new_n18872_, new_n18622_, new_n18422_ );
or   ( new_n18873_, new_n18609_, new_n18453_ );
and  ( new_n18874_, new_n18873_, new_n18872_ );
or   ( new_n18875_, new_n18874_, new_n18637_ );
and  ( new_n18876_, new_n18623_, new_n18454_ );
or   ( new_n18877_, new_n18876_, new_n18486_ );
and  ( new_n18878_, new_n18877_, new_n18875_ );
or   ( new_n18879_, new_n18878_, new_n18871_ );
and  ( new_n18880_, new_n18879_, new_n18870_ );
or   ( new_n18881_, new_n18880_, new_n18859_ );
and  ( new_n18882_, new_n18880_, new_n18859_ );
or   ( new_n18883_, new_n18676_, new_n18364_ );
or   ( new_n18884_, new_n18673_, new_n18371_ );
and  ( new_n18885_, new_n18884_, new_n18883_ );
or   ( new_n18886_, new_n18885_, new_n18681_ );
and  ( new_n18887_, new_n18677_, new_n18372_ );
or   ( new_n18888_, new_n18887_, new_n18380_ );
and  ( new_n18889_, new_n18888_, new_n18886_ );
or   ( new_n18890_, new_n18889_, new_n18882_ );
and  ( new_n18891_, new_n18890_, new_n18881_ );
or   ( new_n18892_, new_n18290_, new_n18154_ );
or   ( new_n18893_, new_n18336_, new_n18190_ );
and  ( new_n18894_, new_n18893_, new_n18892_ );
or   ( new_n18895_, new_n18894_, new_n18344_ );
and  ( new_n18896_, new_n18337_, new_n18207_ );
or   ( new_n18897_, new_n18896_, new_n18206_ );
and  ( new_n18898_, new_n18897_, new_n18895_ );
or   ( new_n18899_, new_n18898_, new_n18891_ );
or   ( new_n18900_, new_n18683_, new_n18548_ );
or   ( new_n18901_, new_n18671_, new_n18382_ );
and  ( new_n18902_, new_n18901_, new_n18900_ );
or   ( new_n18903_, new_n18902_, new_n18687_ );
and  ( new_n18904_, new_n18684_, new_n18550_ );
or   ( new_n18905_, new_n18904_, new_n18557_ );
and  ( new_n18906_, new_n18905_, new_n18903_ );
and  ( new_n18907_, new_n18898_, new_n18891_ );
or   ( new_n18908_, new_n18907_, new_n18906_ );
and  ( new_n18909_, new_n18908_, new_n18899_ );
or   ( new_n18910_, new_n18909_, new_n18697_ );
or   ( new_n18911_, new_n18359_, new_n18252_ );
or   ( new_n18912_, new_n18356_, new_n18229_ );
and  ( new_n18913_, new_n18912_, new_n18911_ );
or   ( new_n18914_, new_n18913_, new_n18577_ );
and  ( new_n18915_, new_n18690_, new_n18595_ );
or   ( new_n18916_, new_n18915_, new_n18592_ );
and  ( new_n18917_, new_n18916_, new_n18694_ );
or   ( new_n18918_, new_n18917_, new_n18361_ );
and  ( new_n18919_, new_n18918_, new_n18914_ );
or   ( new_n18920_, new_n18919_, new_n18910_ );
or   ( new_n18921_, new_n18920_, new_n18589_ );
and  ( new_n18922_, new_n18921_, new_n18588_ );
or   ( new_n18923_, new_n18904_, new_n18687_ );
or   ( new_n18924_, new_n18902_, new_n18557_ );
and  ( new_n18925_, new_n18924_, new_n18923_ );
or   ( new_n18926_, new_n18896_, new_n18344_ );
or   ( new_n18927_, new_n18894_, new_n18206_ );
and  ( new_n18928_, new_n18927_, new_n18926_ );
or   ( new_n18929_, new_n18928_, new_n18891_ );
or   ( new_n18930_, new_n18668_, new_n18665_ );
and  ( new_n18931_, new_n18930_, new_n18546_ );
or   ( new_n18932_, new_n18867_, new_n18658_ );
or   ( new_n18933_, new_n18865_, new_n18527_ );
and  ( new_n18934_, new_n18933_, new_n18932_ );
or   ( new_n18935_, new_n18934_, new_n18931_ );
and  ( new_n18936_, new_n18934_, new_n18931_ );
or   ( new_n18937_, new_n18876_, new_n18637_ );
or   ( new_n18938_, new_n18874_, new_n18486_ );
and  ( new_n18939_, new_n18938_, new_n18937_ );
or   ( new_n18940_, new_n18939_, new_n18936_ );
and  ( new_n18941_, new_n18940_, new_n18935_ );
or   ( new_n18942_, new_n18702_, new_n18651_ );
or   ( new_n18943_, new_n18700_, new_n18516_ );
and  ( new_n18944_, new_n18943_, new_n18942_ );
or   ( new_n18945_, new_n18711_, new_n16217_ );
or   ( new_n18946_, new_n18707_, new_n16234_ );
and  ( new_n18947_, new_n18946_, new_n18945_ );
or   ( new_n18948_, new_n18720_, new_n16151_ );
or   ( new_n18949_, new_n18716_, new_n16170_ );
and  ( new_n18950_, new_n18949_, new_n18948_ );
or   ( new_n18951_, new_n18950_, new_n18947_ );
and  ( new_n18952_, new_n18950_, new_n18947_ );
or   ( new_n18953_, new_n18731_, new_n16108_ );
or   ( new_n18954_, new_n18727_, new_n16128_ );
and  ( new_n18955_, new_n18954_, new_n18953_ );
or   ( new_n18956_, new_n18955_, new_n18952_ );
and  ( new_n18957_, new_n18956_, new_n18951_ );
or   ( new_n18958_, new_n18957_, new_n18944_ );
or   ( new_n18959_, new_n18771_, new_n16814_ );
or   ( new_n18960_, new_n18767_, new_n17142_ );
and  ( new_n18961_, new_n18960_, new_n18959_ );
or   ( new_n18962_, new_n18780_, new_n16505_ );
or   ( new_n18963_, new_n18776_, new_n16438_ );
and  ( new_n18964_, new_n18963_, new_n18962_ );
or   ( new_n18965_, new_n18964_, new_n18961_ );
and  ( new_n18966_, new_n18964_, new_n18961_ );
or   ( new_n18967_, new_n18791_, new_n16085_ );
or   ( new_n18968_, new_n18787_, new_n16048_ );
and  ( new_n18969_, new_n18968_, new_n18967_ );
or   ( new_n18970_, new_n18969_, new_n18966_ );
and  ( new_n18971_, new_n18970_, new_n18965_ );
nand ( new_n18972_, new_n18737_, new_n138_ );
and  ( new_n18973_, new_n18972_, RI2b1c4342c220_25 );
nand ( new_n18974_, new_n18739_, new_n138_ );
and  ( new_n18975_, new_n18974_, RI2b1c4342c1a8_24 );
and  ( new_n18976_, new_n18975_, new_n18973_ );
or   ( new_n18977_, new_n18976_, new_n18062_ );
or   ( new_n18978_, new_n18749_, new_n18066_ );
or   ( new_n18979_, new_n18745_, new_n18309_ );
and  ( new_n18980_, new_n18979_, new_n18978_ );
or   ( new_n18981_, new_n18980_, new_n18977_ );
and  ( new_n18982_, new_n18980_, new_n18977_ );
or   ( new_n18983_, new_n18760_, new_n17238_ );
or   ( new_n18984_, new_n18756_, new_n17650_ );
and  ( new_n18985_, new_n18984_, new_n18983_ );
or   ( new_n18986_, new_n18985_, new_n18982_ );
and  ( new_n18987_, new_n18986_, new_n18981_ );
or   ( new_n18988_, new_n18987_, new_n18971_ );
and  ( new_n18989_, new_n18987_, new_n18971_ );
or   ( new_n18990_, new_n18804_, new_n16052_ );
or   ( new_n18991_, new_n18800_, new_n16071_ );
and  ( new_n18992_, new_n18991_, new_n18990_ );
or   ( new_n18993_, new_n18813_, new_n16009_ );
or   ( new_n18994_, new_n18809_, new_n16029_ );
and  ( new_n18995_, new_n18994_, new_n18993_ );
or   ( new_n18996_, new_n18995_, new_n18992_ );
and  ( new_n18997_, new_n18995_, new_n18992_ );
or   ( new_n18998_, new_n18824_, new_n16186_ );
or   ( new_n18999_, new_n18820_, new_n16204_ );
and  ( new_n19000_, new_n18999_, new_n18998_ );
or   ( new_n19001_, new_n19000_, new_n18997_ );
and  ( new_n19002_, new_n19001_, new_n18996_ );
or   ( new_n19003_, new_n19002_, new_n18989_ );
and  ( new_n19004_, new_n19003_, new_n18988_ );
or   ( new_n19005_, new_n19004_, new_n18958_ );
and  ( new_n19006_, new_n19004_, new_n18958_ );
or   ( new_n19007_, new_n18837_, new_n18635_ );
or   ( new_n19008_, new_n18835_, new_n18484_ );
and  ( new_n19009_, new_n19008_, new_n19007_ );
or   ( new_n19010_, new_n18844_, new_n18620_ );
or   ( new_n19011_, new_n18842_, new_n18451_ );
and  ( new_n19012_, new_n19011_, new_n19010_ );
or   ( new_n19013_, new_n19012_, new_n19009_ );
and  ( new_n19014_, new_n19012_, new_n19009_ );
or   ( new_n19015_, new_n18853_, new_n18607_ );
or   ( new_n19016_, new_n18851_, new_n18420_ );
and  ( new_n19017_, new_n19016_, new_n19015_ );
or   ( new_n19018_, new_n19017_, new_n19014_ );
and  ( new_n19019_, new_n19018_, new_n19013_ );
or   ( new_n19020_, new_n19019_, new_n19006_ );
and  ( new_n19021_, new_n19020_, new_n19005_ );
or   ( new_n19022_, new_n19021_, new_n18941_ );
and  ( new_n19023_, new_n19021_, new_n18941_ );
or   ( new_n19024_, new_n18887_, new_n18681_ );
or   ( new_n19025_, new_n18885_, new_n18380_ );
and  ( new_n19026_, new_n19025_, new_n19024_ );
or   ( new_n19027_, new_n19026_, new_n19023_ );
and  ( new_n19028_, new_n19027_, new_n19022_ );
or   ( new_n19029_, new_n19028_, new_n18898_ );
and  ( new_n19030_, new_n19029_, new_n18929_ );
or   ( new_n19031_, new_n19030_, new_n18925_ );
or   ( new_n19032_, new_n19028_, new_n18928_ );
and  ( new_n19033_, new_n19032_, new_n18899_ );
or   ( new_n19034_, new_n19033_, new_n18906_ );
and  ( new_n19035_, new_n19034_, new_n19031_ );
or   ( new_n19036_, new_n18660_, new_n18488_ );
or   ( new_n19037_, new_n18639_, new_n18529_ );
and  ( new_n19038_, new_n19037_, new_n19036_ );
or   ( new_n19039_, new_n19038_, new_n18669_ );
and  ( new_n19040_, new_n18661_, new_n18531_ );
or   ( new_n19041_, new_n19040_, new_n18546_ );
and  ( new_n19042_, new_n19041_, new_n19039_ );
or   ( new_n19043_, new_n18975_, new_n18973_ );
and  ( new_n19044_, new_n19043_, new_n18741_ );
or   ( new_n19045_, new_n18975_, new_n18062_ );
or   ( new_n19046_, new_n18740_, new_n18307_ );
and  ( new_n19047_, new_n19046_, new_n19045_ );
or   ( new_n19048_, new_n19047_, new_n19044_ );
or   ( new_n19049_, new_n19048_, new_n99_ );
or   ( new_n19050_, new_n19049_, new_n18742_ );
or   ( new_n19051_, new_n18975_, new_n18307_ );
or   ( new_n19052_, new_n18740_, new_n18062_ );
or   ( new_n19053_, new_n18973_, new_n18740_ );
or   ( new_n19054_, new_n18975_, new_n18738_ );
and  ( new_n19055_, new_n19054_, new_n19053_ );
and  ( new_n19056_, new_n19055_, new_n19052_ );
and  ( new_n19057_, new_n19056_, new_n19051_ );
and  ( new_n19058_, new_n19057_, RI2b1c4342d4e0_65 );
or   ( new_n19059_, new_n19058_, new_n18977_ );
and  ( new_n19060_, new_n19059_, new_n19050_ );
or   ( new_n19061_, new_n18388_, new_n112_ );
or   ( new_n19062_, new_n18395_, new_n526_ );
and  ( new_n19063_, new_n19062_, new_n19061_ );
or   ( new_n19064_, new_n19063_, new_n18066_ );
and  ( new_n19065_, new_n18397_, RI2b1c4342d5d0_67 );
and  ( new_n19066_, new_n18384_, RI2b1c4342d558_66 );
or   ( new_n19067_, new_n19066_, new_n19065_ );
or   ( new_n19068_, new_n19067_, new_n18309_ );
and  ( new_n19069_, new_n19068_, new_n19064_ );
or   ( new_n19070_, new_n19069_, new_n19060_ );
and  ( new_n19071_, new_n19069_, new_n19060_ );
or   ( new_n19072_, new_n17727_, new_n591_ );
or   ( new_n19073_, new_n17734_, new_n612_ );
and  ( new_n19074_, new_n19073_, new_n19072_ );
or   ( new_n19075_, new_n19074_, new_n17238_ );
and  ( new_n19076_, new_n17736_, RI2b1c4342d6c0_69 );
and  ( new_n19077_, new_n17723_, RI2b1c4342d648_68 );
or   ( new_n19078_, new_n19077_, new_n19076_ );
or   ( new_n19079_, new_n19078_, new_n17650_ );
and  ( new_n19080_, new_n19079_, new_n19075_ );
or   ( new_n19081_, new_n19080_, new_n19071_ );
and  ( new_n19082_, new_n19081_, new_n19070_ );
or   ( new_n19083_, new_n17244_, new_n110_ );
or   ( new_n19084_, new_n17248_, new_n755_ );
and  ( new_n19085_, new_n19084_, new_n19083_ );
or   ( new_n19086_, new_n19085_, new_n16814_ );
and  ( new_n19087_, new_n17255_, RI2b1c4342d7b0_71 );
and  ( new_n19088_, new_n17240_, RI2b1c4342d738_70 );
or   ( new_n19089_, new_n19088_, new_n19087_ );
or   ( new_n19090_, new_n19089_, new_n17142_ );
and  ( new_n19091_, new_n19090_, new_n19086_ );
or   ( new_n19092_, new_n16607_, new_n105_ );
or   ( new_n19093_, new_n16613_, new_n806_ );
and  ( new_n19094_, new_n19093_, new_n19092_ );
or   ( new_n19095_, new_n19094_, new_n16505_ );
and  ( new_n19096_, new_n16616_, RI2b1c4342d8a0_73 );
and  ( new_n19097_, new_n16603_, RI2b1c4342d828_72 );
or   ( new_n19098_, new_n19097_, new_n19096_ );
or   ( new_n19099_, new_n19098_, new_n16438_ );
and  ( new_n19100_, new_n19099_, new_n19095_ );
or   ( new_n19101_, new_n19100_, new_n19091_ );
and  ( new_n19102_, new_n19100_, new_n19091_ );
or   ( new_n19103_, new_n16366_, new_n843_ );
or   ( new_n19104_, new_n16355_, new_n859_ );
and  ( new_n19105_, new_n19104_, new_n19103_ );
or   ( new_n19106_, new_n19105_, new_n16085_ );
and  ( new_n19107_, new_n16358_, RI2b1c4342d990_75 );
and  ( new_n19108_, new_n16362_, RI2b1c4342d918_74 );
or   ( new_n19109_, new_n19108_, new_n19107_ );
or   ( new_n19110_, new_n19109_, new_n16048_ );
and  ( new_n19111_, new_n19110_, new_n19106_ );
or   ( new_n19112_, new_n19111_, new_n19102_ );
and  ( new_n19113_, new_n19112_, new_n19101_ );
or   ( new_n19114_, new_n19113_, new_n19082_ );
and  ( new_n19115_, new_n19113_, new_n19082_ );
or   ( new_n19116_, new_n16075_, new_n1004_ );
or   ( new_n19117_, new_n16060_, new_n886_ );
and  ( new_n19118_, new_n19117_, new_n19116_ );
or   ( new_n19119_, new_n19118_, new_n16052_ );
and  ( new_n19120_, new_n16063_, RI2b1c4342da80_77 );
and  ( new_n19121_, new_n16066_, RI2b1c4342da08_76 );
or   ( new_n19122_, new_n19121_, new_n19120_ );
or   ( new_n19123_, new_n19122_, new_n16071_ );
and  ( new_n19124_, new_n19123_, new_n19119_ );
or   ( new_n19125_, new_n16033_, new_n1310_ );
or   ( new_n19126_, new_n16017_, new_n1002_ );
and  ( new_n19127_, new_n19126_, new_n19125_ );
or   ( new_n19128_, new_n19127_, new_n16009_ );
and  ( new_n19129_, new_n16021_, RI2b1c4342db70_79 );
and  ( new_n19130_, new_n16024_, RI2b1c4342daf8_78 );
or   ( new_n19131_, new_n19130_, new_n19129_ );
or   ( new_n19132_, new_n19131_, new_n16029_ );
and  ( new_n19133_, new_n19132_, new_n19128_ );
or   ( new_n19134_, new_n19133_, new_n19124_ );
and  ( new_n19135_, new_n19133_, new_n19124_ );
or   ( new_n19136_, new_n16208_, new_n126_ );
or   ( new_n19137_, new_n16194_, new_n1511_ );
and  ( new_n19138_, new_n19137_, new_n19136_ );
or   ( new_n19139_, new_n19138_, new_n16186_ );
and  ( new_n19140_, new_n16196_, RI2b1c4342dc60_81 );
and  ( new_n19141_, new_n16199_, RI2b1c4342dbe8_80 );
or   ( new_n19142_, new_n19141_, new_n19140_ );
or   ( new_n19143_, new_n19142_, new_n16204_ );
and  ( new_n19144_, new_n19143_, new_n19139_ );
or   ( new_n19145_, new_n19144_, new_n19135_ );
and  ( new_n19146_, new_n19145_, new_n19134_ );
or   ( new_n19147_, new_n19146_, new_n19115_ );
and  ( new_n19148_, new_n19147_, new_n19114_ );
or   ( new_n19149_, new_n16115_, new_n3902_ );
or   ( new_n19150_, new_n16238_, new_n121_ );
or   ( new_n19151_, new_n16224_, new_n2119_ );
and  ( new_n19152_, new_n19151_, new_n19150_ );
or   ( new_n19153_, new_n19152_, new_n16217_ );
and  ( new_n19154_, new_n16226_, RI2b1c4342dd50_83 );
and  ( new_n19155_, new_n16229_, RI2b1c4342dcd8_82 );
or   ( new_n19156_, new_n19155_, new_n19154_ );
or   ( new_n19157_, new_n19156_, new_n16234_ );
and  ( new_n19158_, new_n19157_, new_n19153_ );
or   ( new_n19159_, new_n16174_, new_n2806_ );
or   ( new_n19160_, new_n16160_, new_n2541_ );
and  ( new_n19161_, new_n19160_, new_n19159_ );
or   ( new_n19162_, new_n19161_, new_n16151_ );
and  ( new_n19163_, new_n16162_, RI2b1c4342de40_85 );
and  ( new_n19164_, new_n16165_, RI2b1c4342ddc8_84 );
or   ( new_n19165_, new_n19164_, new_n19163_ );
or   ( new_n19166_, new_n19165_, new_n16170_ );
and  ( new_n19167_, new_n19166_, new_n19162_ );
or   ( new_n19168_, new_n19167_, new_n19158_ );
and  ( new_n19169_, new_n19167_, new_n19158_ );
or   ( new_n19170_, new_n16119_, new_n3924_ );
or   ( new_n19171_, new_n16123_, new_n3239_ );
and  ( new_n19172_, new_n19171_, new_n19170_ );
or   ( new_n19173_, new_n19172_, new_n16108_ );
and  ( new_n19174_, new_n16132_, RI2b1c4342df30_87 );
and  ( new_n19175_, new_n16114_, RI2b1c4342deb8_86 );
or   ( new_n19176_, new_n19175_, new_n19174_ );
or   ( new_n19177_, new_n19176_, new_n16128_ );
and  ( new_n19178_, new_n19177_, new_n19173_ );
or   ( new_n19179_, new_n19178_, new_n19169_ );
and  ( new_n19180_, new_n19179_, new_n19168_ );
or   ( new_n19181_, new_n19180_, new_n19149_ );
and  ( new_n19182_, new_n19180_, new_n19149_ );
or   ( new_n19183_, new_n16115_, new_n3924_ );
or   ( new_n19184_, new_n19183_, new_n19182_ );
and  ( new_n19185_, new_n19184_, new_n19181_ );
or   ( new_n19186_, new_n19185_, new_n19148_ );
and  ( new_n19187_, new_n19185_, new_n19148_ );
or   ( new_n19188_, new_n18950_, new_n18713_ );
or   ( new_n19189_, new_n18947_, new_n18722_ );
and  ( new_n19190_, new_n19189_, new_n19188_ );
or   ( new_n19191_, new_n19190_, new_n18955_ );
and  ( new_n19192_, new_n18951_, new_n18723_ );
or   ( new_n19193_, new_n19192_, new_n18733_ );
and  ( new_n19194_, new_n19193_, new_n19191_ );
or   ( new_n19195_, new_n18995_, new_n18806_ );
or   ( new_n19196_, new_n18992_, new_n18815_ );
and  ( new_n19197_, new_n19196_, new_n19195_ );
or   ( new_n19198_, new_n19197_, new_n19000_ );
and  ( new_n19199_, new_n18996_, new_n18816_ );
or   ( new_n19200_, new_n19199_, new_n18826_ );
and  ( new_n19201_, new_n19200_, new_n19198_ );
or   ( new_n19202_, new_n19201_, new_n19194_ );
and  ( new_n19203_, new_n19201_, new_n19194_ );
or   ( new_n19204_, new_n18964_, new_n18773_ );
or   ( new_n19205_, new_n18961_, new_n18782_ );
and  ( new_n19206_, new_n19205_, new_n19204_ );
or   ( new_n19207_, new_n19206_, new_n18969_ );
and  ( new_n19208_, new_n18965_, new_n18783_ );
or   ( new_n19209_, new_n19208_, new_n18793_ );
and  ( new_n19210_, new_n19209_, new_n19207_ );
or   ( new_n19211_, new_n19210_, new_n19203_ );
and  ( new_n19212_, new_n19211_, new_n19202_ );
or   ( new_n19213_, new_n19212_, new_n19187_ );
and  ( new_n19214_, new_n19213_, new_n19186_ );
or   ( new_n19215_, new_n19012_, new_n18839_ );
or   ( new_n19216_, new_n19009_, new_n18846_ );
and  ( new_n19217_, new_n19216_, new_n19215_ );
or   ( new_n19218_, new_n19217_, new_n19017_ );
and  ( new_n19219_, new_n19013_, new_n18847_ );
or   ( new_n19220_, new_n19219_, new_n18855_ );
and  ( new_n19221_, new_n19220_, new_n19218_ );
or   ( new_n19222_, new_n18735_, new_n18704_ );
and  ( new_n19223_, new_n19222_, new_n18958_ );
or   ( new_n19224_, new_n19223_, new_n19221_ );
and  ( new_n19225_, new_n19223_, new_n19221_ );
or   ( new_n19226_, new_n18971_, new_n18764_ );
or   ( new_n19227_, new_n18987_, new_n18795_ );
and  ( new_n19228_, new_n19227_, new_n19226_ );
or   ( new_n19229_, new_n19228_, new_n19002_ );
and  ( new_n19230_, new_n18988_, new_n18796_ );
or   ( new_n19231_, new_n19230_, new_n18828_ );
and  ( new_n19232_, new_n19231_, new_n19229_ );
or   ( new_n19233_, new_n19232_, new_n19225_ );
and  ( new_n19234_, new_n19233_, new_n19224_ );
or   ( new_n19235_, new_n19234_, new_n19214_ );
and  ( new_n19236_, new_n19234_, new_n19214_ );
or   ( new_n19237_, new_n18934_, new_n18862_ );
or   ( new_n19238_, new_n18931_, new_n18869_ );
and  ( new_n19239_, new_n19238_, new_n19237_ );
or   ( new_n19240_, new_n19239_, new_n18939_ );
and  ( new_n19241_, new_n18935_, new_n18870_ );
or   ( new_n19242_, new_n19241_, new_n18878_ );
and  ( new_n19243_, new_n19242_, new_n19240_ );
or   ( new_n19244_, new_n19243_, new_n19236_ );
and  ( new_n19245_, new_n19244_, new_n19235_ );
or   ( new_n19246_, new_n19245_, new_n19042_ );
and  ( new_n19247_, new_n19245_, new_n19042_ );
or   ( new_n19248_, new_n18941_, new_n18859_ );
or   ( new_n19249_, new_n19021_, new_n18880_ );
and  ( new_n19250_, new_n19249_, new_n19248_ );
or   ( new_n19251_, new_n19250_, new_n19026_ );
and  ( new_n19252_, new_n19022_, new_n18881_ );
or   ( new_n19253_, new_n19252_, new_n18889_ );
and  ( new_n19254_, new_n19253_, new_n19251_ );
or   ( new_n19255_, new_n19254_, new_n19247_ );
and  ( new_n19256_, new_n19255_, new_n19246_ );
or   ( new_n19257_, new_n19256_, new_n19035_ );
or   ( new_n19258_, new_n18695_, new_n18592_ );
or   ( new_n19259_, new_n18692_, new_n18574_ );
and  ( new_n19260_, new_n19259_, new_n19258_ );
or   ( new_n19261_, new_n19260_, new_n18909_ );
and  ( new_n19262_, new_n19028_, new_n18928_ );
or   ( new_n19263_, new_n19262_, new_n18925_ );
and  ( new_n19264_, new_n19263_, new_n19032_ );
or   ( new_n19265_, new_n19264_, new_n18697_ );
and  ( new_n19266_, new_n19265_, new_n19261_ );
or   ( new_n19267_, new_n19266_, new_n19257_ );
and  ( new_n19268_, new_n19266_, new_n19257_ );
or   ( new_n19269_, new_n19252_, new_n19026_ );
or   ( new_n19270_, new_n19250_, new_n18889_ );
and  ( new_n19271_, new_n19270_, new_n19269_ );
or   ( new_n19272_, new_n19040_, new_n18669_ );
or   ( new_n19273_, new_n19038_, new_n18546_ );
and  ( new_n19274_, new_n19273_, new_n19272_ );
or   ( new_n19275_, new_n19274_, new_n19245_ );
or   ( new_n19276_, new_n19058_, new_n18742_ );
or   ( new_n19277_, new_n19049_, new_n18977_ );
and  ( new_n19278_, new_n19277_, new_n19276_ );
or   ( new_n19279_, new_n19067_, new_n18066_ );
or   ( new_n19280_, new_n19063_, new_n18309_ );
and  ( new_n19281_, new_n19280_, new_n19279_ );
or   ( new_n19282_, new_n19281_, new_n19278_ );
and  ( new_n19283_, new_n19281_, new_n19278_ );
or   ( new_n19284_, new_n19078_, new_n17238_ );
or   ( new_n19285_, new_n19074_, new_n17650_ );
and  ( new_n19286_, new_n19285_, new_n19284_ );
or   ( new_n19287_, new_n19286_, new_n19283_ );
and  ( new_n19288_, new_n19287_, new_n19282_ );
or   ( new_n19289_, new_n19089_, new_n16814_ );
or   ( new_n19290_, new_n19085_, new_n17142_ );
and  ( new_n19291_, new_n19290_, new_n19289_ );
or   ( new_n19292_, new_n19098_, new_n16505_ );
or   ( new_n19293_, new_n19094_, new_n16438_ );
and  ( new_n19294_, new_n19293_, new_n19292_ );
or   ( new_n19295_, new_n19294_, new_n19291_ );
and  ( new_n19296_, new_n19294_, new_n19291_ );
or   ( new_n19297_, new_n19109_, new_n16085_ );
or   ( new_n19298_, new_n19105_, new_n16048_ );
and  ( new_n19299_, new_n19298_, new_n19297_ );
or   ( new_n19300_, new_n19299_, new_n19296_ );
and  ( new_n19301_, new_n19300_, new_n19295_ );
or   ( new_n19302_, new_n19301_, new_n19288_ );
and  ( new_n19303_, new_n19301_, new_n19288_ );
or   ( new_n19304_, new_n19122_, new_n16052_ );
or   ( new_n19305_, new_n19118_, new_n16071_ );
and  ( new_n19306_, new_n19305_, new_n19304_ );
or   ( new_n19307_, new_n19131_, new_n16009_ );
or   ( new_n19308_, new_n19127_, new_n16029_ );
and  ( new_n19309_, new_n19308_, new_n19307_ );
or   ( new_n19310_, new_n19309_, new_n19306_ );
and  ( new_n19311_, new_n19309_, new_n19306_ );
or   ( new_n19312_, new_n19142_, new_n16186_ );
or   ( new_n19313_, new_n19138_, new_n16204_ );
and  ( new_n19314_, new_n19313_, new_n19312_ );
or   ( new_n19315_, new_n19314_, new_n19311_ );
and  ( new_n19316_, new_n19315_, new_n19310_ );
or   ( new_n19317_, new_n19316_, new_n19303_ );
and  ( new_n19318_, new_n19317_, new_n19302_ );
and  ( new_n19319_, new_n16102_, RI2b1c4342dfa8_88 );
or   ( new_n19320_, new_n19156_, new_n16217_ );
or   ( new_n19321_, new_n19152_, new_n16234_ );
and  ( new_n19322_, new_n19321_, new_n19320_ );
or   ( new_n19323_, new_n19165_, new_n16151_ );
or   ( new_n19324_, new_n19161_, new_n16170_ );
and  ( new_n19325_, new_n19324_, new_n19323_ );
or   ( new_n19326_, new_n19325_, new_n19322_ );
and  ( new_n19327_, new_n19325_, new_n19322_ );
or   ( new_n19328_, new_n19176_, new_n16108_ );
or   ( new_n19329_, new_n19172_, new_n16128_ );
and  ( new_n19330_, new_n19329_, new_n19328_ );
or   ( new_n19331_, new_n19330_, new_n19327_ );
and  ( new_n19332_, new_n19331_, new_n19326_ );
or   ( new_n19333_, new_n19332_, new_n19319_ );
and  ( new_n19334_, new_n19332_, new_n19319_ );
and  ( new_n19335_, new_n16102_, RI2b1c4342df30_87 );
or   ( new_n19336_, new_n19335_, new_n19334_ );
and  ( new_n19337_, new_n19336_, new_n19333_ );
or   ( new_n19338_, new_n19337_, new_n19318_ );
and  ( new_n19339_, new_n19337_, new_n19318_ );
or   ( new_n19340_, new_n19192_, new_n18955_ );
or   ( new_n19341_, new_n19190_, new_n18733_ );
and  ( new_n19342_, new_n19341_, new_n19340_ );
or   ( new_n19343_, new_n19199_, new_n19000_ );
or   ( new_n19344_, new_n19197_, new_n18826_ );
and  ( new_n19345_, new_n19344_, new_n19343_ );
or   ( new_n19346_, new_n19345_, new_n19342_ );
and  ( new_n19347_, new_n19345_, new_n19342_ );
or   ( new_n19348_, new_n19208_, new_n18969_ );
or   ( new_n19349_, new_n19206_, new_n18793_ );
and  ( new_n19350_, new_n19349_, new_n19348_ );
or   ( new_n19351_, new_n19350_, new_n19347_ );
and  ( new_n19352_, new_n19351_, new_n19346_ );
or   ( new_n19353_, new_n19352_, new_n19339_ );
and  ( new_n19354_, new_n19353_, new_n19338_ );
or   ( new_n19355_, new_n19219_, new_n19017_ );
or   ( new_n19356_, new_n19217_, new_n18855_ );
and  ( new_n19357_, new_n19356_, new_n19355_ );
or   ( new_n19358_, new_n18944_, new_n18735_ );
or   ( new_n19359_, new_n18957_, new_n18704_ );
and  ( new_n19360_, new_n19359_, new_n19358_ );
or   ( new_n19361_, new_n19360_, new_n19357_ );
and  ( new_n19362_, new_n19360_, new_n19357_ );
or   ( new_n19363_, new_n19230_, new_n19002_ );
or   ( new_n19364_, new_n19228_, new_n18828_ );
and  ( new_n19365_, new_n19364_, new_n19363_ );
or   ( new_n19366_, new_n19365_, new_n19362_ );
and  ( new_n19367_, new_n19366_, new_n19361_ );
or   ( new_n19368_, new_n19367_, new_n19354_ );
and  ( new_n19369_, new_n19367_, new_n19354_ );
or   ( new_n19370_, new_n19241_, new_n18939_ );
or   ( new_n19371_, new_n19239_, new_n18878_ );
and  ( new_n19372_, new_n19371_, new_n19370_ );
or   ( new_n19373_, new_n19372_, new_n19369_ );
and  ( new_n19374_, new_n19373_, new_n19368_ );
or   ( new_n19375_, new_n19374_, new_n19042_ );
and  ( new_n19376_, new_n19375_, new_n19275_ );
or   ( new_n19377_, new_n19376_, new_n19271_ );
or   ( new_n19378_, new_n19374_, new_n19274_ );
and  ( new_n19379_, new_n19378_, new_n19246_ );
or   ( new_n19380_, new_n19379_, new_n19254_ );
and  ( new_n19381_, new_n19380_, new_n19377_ );
or   ( new_n19382_, new_n18958_, new_n18830_ );
or   ( new_n19383_, new_n19004_, new_n18736_ );
and  ( new_n19384_, new_n19383_, new_n19382_ );
or   ( new_n19385_, new_n19384_, new_n19019_ );
and  ( new_n19386_, new_n19005_, new_n18831_ );
or   ( new_n19387_, new_n19386_, new_n18857_ );
and  ( new_n19388_, new_n19387_, new_n19385_ );
xor  ( new_n19389_, new_n4202_, new_n4390_ );
or   ( new_n19390_, new_n19389_, new_n318_ );
xor  ( new_n19391_, new_n4209_, new_n226_ );
or   ( new_n19392_, new_n19391_, new_n315_ );
or   ( new_n19393_, new_n19392_, new_n19390_ );
and  ( new_n19394_, new_n19393_, new_n18973_ );
or   ( new_n19395_, new_n19048_, new_n526_ );
or   ( new_n19396_, new_n19055_, new_n99_ );
and  ( new_n19397_, new_n19396_, new_n19395_ );
or   ( new_n19398_, new_n19397_, new_n18742_ );
and  ( new_n19399_, new_n19057_, RI2b1c4342d558_66 );
and  ( new_n19400_, new_n19044_, RI2b1c4342d4e0_65 );
or   ( new_n19401_, new_n19400_, new_n19399_ );
or   ( new_n19402_, new_n19401_, new_n18977_ );
and  ( new_n19403_, new_n19402_, new_n19398_ );
or   ( new_n19404_, new_n19403_, new_n19394_ );
and  ( new_n19405_, new_n19403_, new_n19394_ );
or   ( new_n19406_, new_n18388_, new_n612_ );
or   ( new_n19407_, new_n18395_, new_n112_ );
and  ( new_n19408_, new_n19407_, new_n19406_ );
or   ( new_n19409_, new_n19408_, new_n18066_ );
and  ( new_n19410_, new_n18397_, RI2b1c4342d648_68 );
and  ( new_n19411_, new_n18384_, RI2b1c4342d5d0_67 );
or   ( new_n19412_, new_n19411_, new_n19410_ );
or   ( new_n19413_, new_n19412_, new_n18309_ );
and  ( new_n19414_, new_n19413_, new_n19409_ );
or   ( new_n19415_, new_n19414_, new_n19405_ );
and  ( new_n19416_, new_n19415_, new_n19404_ );
or   ( new_n19417_, new_n17727_, new_n755_ );
or   ( new_n19418_, new_n17734_, new_n591_ );
and  ( new_n19419_, new_n19418_, new_n19417_ );
or   ( new_n19420_, new_n19419_, new_n17238_ );
and  ( new_n19421_, new_n17736_, RI2b1c4342d738_70 );
and  ( new_n19422_, new_n17723_, RI2b1c4342d6c0_69 );
or   ( new_n19423_, new_n19422_, new_n19421_ );
or   ( new_n19424_, new_n19423_, new_n17650_ );
and  ( new_n19425_, new_n19424_, new_n19420_ );
or   ( new_n19426_, new_n17244_, new_n806_ );
or   ( new_n19427_, new_n17248_, new_n110_ );
and  ( new_n19428_, new_n19427_, new_n19426_ );
or   ( new_n19429_, new_n19428_, new_n16814_ );
and  ( new_n19430_, new_n17255_, RI2b1c4342d828_72 );
and  ( new_n19431_, new_n17240_, RI2b1c4342d7b0_71 );
or   ( new_n19432_, new_n19431_, new_n19430_ );
or   ( new_n19433_, new_n19432_, new_n17142_ );
and  ( new_n19434_, new_n19433_, new_n19429_ );
or   ( new_n19435_, new_n19434_, new_n19425_ );
and  ( new_n19436_, new_n19434_, new_n19425_ );
or   ( new_n19437_, new_n16607_, new_n859_ );
or   ( new_n19438_, new_n16613_, new_n105_ );
and  ( new_n19439_, new_n19438_, new_n19437_ );
or   ( new_n19440_, new_n19439_, new_n16505_ );
and  ( new_n19441_, new_n16616_, RI2b1c4342d918_74 );
and  ( new_n19442_, new_n16603_, RI2b1c4342d8a0_73 );
or   ( new_n19443_, new_n19442_, new_n19441_ );
or   ( new_n19444_, new_n19443_, new_n16438_ );
and  ( new_n19445_, new_n19444_, new_n19440_ );
or   ( new_n19446_, new_n19445_, new_n19436_ );
and  ( new_n19447_, new_n19446_, new_n19435_ );
or   ( new_n19448_, new_n19447_, new_n19416_ );
and  ( new_n19449_, new_n19447_, new_n19416_ );
or   ( new_n19450_, new_n16366_, new_n886_ );
or   ( new_n19451_, new_n16355_, new_n843_ );
and  ( new_n19452_, new_n19451_, new_n19450_ );
or   ( new_n19453_, new_n19452_, new_n16085_ );
and  ( new_n19454_, new_n16358_, RI2b1c4342da08_76 );
and  ( new_n19455_, new_n16362_, RI2b1c4342d990_75 );
or   ( new_n19456_, new_n19455_, new_n19454_ );
or   ( new_n19457_, new_n19456_, new_n16048_ );
and  ( new_n19458_, new_n19457_, new_n19453_ );
or   ( new_n19459_, new_n16075_, new_n1002_ );
or   ( new_n19460_, new_n16060_, new_n1004_ );
and  ( new_n19461_, new_n19460_, new_n19459_ );
or   ( new_n19462_, new_n19461_, new_n16052_ );
and  ( new_n19463_, new_n16063_, RI2b1c4342daf8_78 );
and  ( new_n19464_, new_n16066_, RI2b1c4342da80_77 );
or   ( new_n19465_, new_n19464_, new_n19463_ );
or   ( new_n19466_, new_n19465_, new_n16071_ );
and  ( new_n19467_, new_n19466_, new_n19462_ );
or   ( new_n19468_, new_n19467_, new_n19458_ );
and  ( new_n19469_, new_n19467_, new_n19458_ );
or   ( new_n19470_, new_n16033_, new_n1511_ );
or   ( new_n19471_, new_n16017_, new_n1310_ );
and  ( new_n19472_, new_n19471_, new_n19470_ );
or   ( new_n19473_, new_n19472_, new_n16009_ );
and  ( new_n19474_, new_n16021_, RI2b1c4342dbe8_80 );
and  ( new_n19475_, new_n16024_, RI2b1c4342db70_79 );
or   ( new_n19476_, new_n19475_, new_n19474_ );
or   ( new_n19477_, new_n19476_, new_n16029_ );
and  ( new_n19478_, new_n19477_, new_n19473_ );
or   ( new_n19479_, new_n19478_, new_n19469_ );
and  ( new_n19480_, new_n19479_, new_n19468_ );
or   ( new_n19481_, new_n19480_, new_n19449_ );
and  ( new_n19482_, new_n19481_, new_n19448_ );
or   ( new_n19483_, new_n16208_, new_n2119_ );
or   ( new_n19484_, new_n16194_, new_n126_ );
and  ( new_n19485_, new_n19484_, new_n19483_ );
or   ( new_n19486_, new_n19485_, new_n16186_ );
and  ( new_n19487_, new_n16196_, RI2b1c4342dcd8_82 );
and  ( new_n19488_, new_n16199_, RI2b1c4342dc60_81 );
or   ( new_n19489_, new_n19488_, new_n19487_ );
or   ( new_n19490_, new_n19489_, new_n16204_ );
and  ( new_n19491_, new_n19490_, new_n19486_ );
or   ( new_n19492_, new_n16238_, new_n2541_ );
or   ( new_n19493_, new_n16224_, new_n121_ );
and  ( new_n19494_, new_n19493_, new_n19492_ );
or   ( new_n19495_, new_n19494_, new_n16217_ );
and  ( new_n19496_, new_n16226_, RI2b1c4342ddc8_84 );
and  ( new_n19497_, new_n16229_, RI2b1c4342dd50_83 );
or   ( new_n19498_, new_n19497_, new_n19496_ );
or   ( new_n19499_, new_n19498_, new_n16234_ );
and  ( new_n19500_, new_n19499_, new_n19495_ );
or   ( new_n19501_, new_n19500_, new_n19491_ );
and  ( new_n19502_, new_n19500_, new_n19491_ );
or   ( new_n19503_, new_n16174_, new_n3239_ );
or   ( new_n19504_, new_n16160_, new_n2806_ );
and  ( new_n19505_, new_n19504_, new_n19503_ );
or   ( new_n19506_, new_n19505_, new_n16151_ );
and  ( new_n19507_, new_n16162_, RI2b1c4342deb8_86 );
and  ( new_n19508_, new_n16165_, RI2b1c4342de40_85 );
or   ( new_n19509_, new_n19508_, new_n19507_ );
or   ( new_n19510_, new_n19509_, new_n16170_ );
and  ( new_n19511_, new_n19510_, new_n19506_ );
or   ( new_n19512_, new_n19511_, new_n19502_ );
and  ( new_n19513_, new_n19512_, new_n19501_ );
or   ( new_n19514_, new_n19513_, new_n19319_ );
and  ( new_n19515_, new_n19513_, new_n19319_ );
or   ( new_n19516_, new_n19325_, new_n19158_ );
or   ( new_n19517_, new_n19322_, new_n19167_ );
and  ( new_n19518_, new_n19517_, new_n19516_ );
or   ( new_n19519_, new_n19518_, new_n19330_ );
and  ( new_n19520_, new_n19326_, new_n19168_ );
or   ( new_n19521_, new_n19520_, new_n19178_ );
and  ( new_n19522_, new_n19521_, new_n19519_ );
or   ( new_n19523_, new_n19522_, new_n19515_ );
and  ( new_n19524_, new_n19523_, new_n19514_ );
or   ( new_n19525_, new_n19524_, new_n19482_ );
and  ( new_n19526_, new_n19524_, new_n19482_ );
or   ( new_n19527_, new_n19309_, new_n19124_ );
or   ( new_n19528_, new_n19306_, new_n19133_ );
and  ( new_n19529_, new_n19528_, new_n19527_ );
or   ( new_n19530_, new_n19529_, new_n19314_ );
and  ( new_n19531_, new_n19310_, new_n19134_ );
or   ( new_n19532_, new_n19531_, new_n19144_ );
and  ( new_n19533_, new_n19532_, new_n19530_ );
or   ( new_n19534_, new_n19294_, new_n19091_ );
or   ( new_n19535_, new_n19291_, new_n19100_ );
and  ( new_n19536_, new_n19535_, new_n19534_ );
or   ( new_n19537_, new_n19536_, new_n19299_ );
and  ( new_n19538_, new_n19295_, new_n19101_ );
or   ( new_n19539_, new_n19538_, new_n19111_ );
and  ( new_n19540_, new_n19539_, new_n19537_ );
or   ( new_n19541_, new_n19540_, new_n19533_ );
and  ( new_n19542_, new_n19540_, new_n19533_ );
or   ( new_n19543_, new_n19281_, new_n19060_ );
or   ( new_n19544_, new_n19278_, new_n19069_ );
and  ( new_n19545_, new_n19544_, new_n19543_ );
or   ( new_n19546_, new_n19545_, new_n19286_ );
and  ( new_n19547_, new_n19282_, new_n19070_ );
or   ( new_n19548_, new_n19547_, new_n19080_ );
and  ( new_n19549_, new_n19548_, new_n19546_ );
or   ( new_n19550_, new_n19549_, new_n19542_ );
and  ( new_n19551_, new_n19550_, new_n19541_ );
or   ( new_n19552_, new_n19551_, new_n19526_ );
and  ( new_n19553_, new_n19552_, new_n19525_ );
or   ( new_n19554_, new_n18980_, new_n18742_ );
or   ( new_n19555_, new_n18977_, new_n18751_ );
and  ( new_n19556_, new_n19555_, new_n19554_ );
or   ( new_n19557_, new_n19556_, new_n18985_ );
and  ( new_n19558_, new_n18981_, new_n18752_ );
or   ( new_n19559_, new_n19558_, new_n18762_ );
and  ( new_n19560_, new_n19559_, new_n19557_ );
or   ( new_n19561_, new_n19345_, new_n19194_ );
or   ( new_n19562_, new_n19342_, new_n19201_ );
and  ( new_n19563_, new_n19562_, new_n19561_ );
or   ( new_n19564_, new_n19563_, new_n19350_ );
and  ( new_n19565_, new_n19346_, new_n19202_ );
or   ( new_n19566_, new_n19565_, new_n19210_ );
and  ( new_n19567_, new_n19566_, new_n19564_ );
or   ( new_n19568_, new_n19567_, new_n19560_ );
and  ( new_n19569_, new_n19567_, new_n19560_ );
or   ( new_n19570_, new_n19319_, new_n19180_ );
or   ( new_n19571_, new_n19332_, new_n19149_ );
and  ( new_n19572_, new_n19571_, new_n19570_ );
or   ( new_n19573_, new_n19572_, new_n19335_ );
and  ( new_n19574_, new_n19333_, new_n19181_ );
or   ( new_n19575_, new_n19574_, new_n19183_ );
and  ( new_n19576_, new_n19575_, new_n19573_ );
or   ( new_n19577_, new_n19576_, new_n19569_ );
and  ( new_n19578_, new_n19577_, new_n19568_ );
or   ( new_n19579_, new_n19578_, new_n19553_ );
and  ( new_n19580_, new_n19578_, new_n19553_ );
or   ( new_n19581_, new_n19360_, new_n19221_ );
or   ( new_n19582_, new_n19357_, new_n19223_ );
and  ( new_n19583_, new_n19582_, new_n19581_ );
or   ( new_n19584_, new_n19583_, new_n19365_ );
and  ( new_n19585_, new_n19361_, new_n19224_ );
or   ( new_n19586_, new_n19585_, new_n19232_ );
and  ( new_n19587_, new_n19586_, new_n19584_ );
or   ( new_n19588_, new_n19587_, new_n19580_ );
and  ( new_n19589_, new_n19588_, new_n19579_ );
or   ( new_n19590_, new_n19589_, new_n19388_ );
and  ( new_n19591_, new_n19589_, new_n19388_ );
or   ( new_n19592_, new_n19367_, new_n19214_ );
or   ( new_n19593_, new_n19354_, new_n19234_ );
and  ( new_n19594_, new_n19593_, new_n19592_ );
or   ( new_n19595_, new_n19594_, new_n19372_ );
and  ( new_n19596_, new_n19368_, new_n19235_ );
or   ( new_n19597_, new_n19596_, new_n19243_ );
and  ( new_n19598_, new_n19597_, new_n19595_ );
or   ( new_n19599_, new_n19598_, new_n19591_ );
and  ( new_n19600_, new_n19599_, new_n19590_ );
or   ( new_n19601_, new_n19600_, new_n19381_ );
or   ( new_n19602_, new_n19033_, new_n18925_ );
or   ( new_n19603_, new_n19030_, new_n18906_ );
and  ( new_n19604_, new_n19603_, new_n19602_ );
or   ( new_n19605_, new_n19604_, new_n19256_ );
and  ( new_n19606_, new_n19374_, new_n19274_ );
or   ( new_n19607_, new_n19606_, new_n19271_ );
and  ( new_n19608_, new_n19607_, new_n19378_ );
or   ( new_n19609_, new_n19608_, new_n19035_ );
and  ( new_n19610_, new_n19609_, new_n19605_ );
or   ( new_n19611_, new_n19610_, new_n19601_ );
or   ( new_n19612_, new_n19611_, new_n19268_ );
and  ( new_n19613_, new_n19612_, new_n19267_ );
and  ( new_n19614_, new_n18919_, new_n18910_ );
or   ( new_n19615_, new_n19614_, new_n18589_ );
or   ( new_n19616_, new_n19615_, new_n19613_ );
and  ( new_n19617_, new_n19616_, new_n18922_ );
and  ( new_n19618_, new_n19610_, new_n19601_ );
or   ( new_n19619_, new_n19618_, new_n19268_ );
or   ( new_n19620_, new_n19619_, new_n19615_ );
or   ( new_n19621_, new_n19596_, new_n19372_ );
or   ( new_n19622_, new_n19594_, new_n19243_ );
and  ( new_n19623_, new_n19622_, new_n19621_ );
or   ( new_n19624_, new_n19386_, new_n19019_ );
or   ( new_n19625_, new_n19384_, new_n18857_ );
and  ( new_n19626_, new_n19625_, new_n19624_ );
or   ( new_n19627_, new_n19626_, new_n19589_ );
or   ( new_n19628_, new_n19558_, new_n18985_ );
or   ( new_n19629_, new_n19556_, new_n18762_ );
and  ( new_n19630_, new_n19629_, new_n19628_ );
or   ( new_n19631_, new_n19565_, new_n19350_ );
or   ( new_n19632_, new_n19563_, new_n19210_ );
and  ( new_n19633_, new_n19632_, new_n19631_ );
or   ( new_n19634_, new_n19633_, new_n19630_ );
and  ( new_n19635_, new_n19633_, new_n19630_ );
or   ( new_n19636_, new_n19574_, new_n19335_ );
or   ( new_n19637_, new_n19572_, new_n19183_ );
and  ( new_n19638_, new_n19637_, new_n19636_ );
or   ( new_n19639_, new_n19638_, new_n19635_ );
and  ( new_n19640_, new_n19639_, new_n19634_ );
or   ( new_n19641_, new_n19423_, new_n17238_ );
or   ( new_n19642_, new_n19419_, new_n17650_ );
and  ( new_n19643_, new_n19642_, new_n19641_ );
or   ( new_n19644_, new_n19432_, new_n16814_ );
or   ( new_n19645_, new_n19428_, new_n17142_ );
and  ( new_n19646_, new_n19645_, new_n19644_ );
or   ( new_n19647_, new_n19646_, new_n19643_ );
and  ( new_n19648_, new_n19646_, new_n19643_ );
or   ( new_n19649_, new_n19443_, new_n16505_ );
or   ( new_n19650_, new_n19439_, new_n16438_ );
and  ( new_n19651_, new_n19650_, new_n19649_ );
or   ( new_n19652_, new_n19651_, new_n19648_ );
and  ( new_n19653_, new_n19652_, new_n19647_ );
nand ( new_n19654_, new_n19389_, new_n138_ );
and  ( new_n19655_, new_n19654_, RI2b1c4342c310_27 );
nand ( new_n19656_, new_n19391_, new_n138_ );
and  ( new_n19657_, new_n19656_, RI2b1c4342c298_26 );
and  ( new_n19658_, new_n19657_, new_n19655_ );
or   ( new_n19659_, new_n19658_, new_n18738_ );
or   ( new_n19660_, new_n19401_, new_n18742_ );
or   ( new_n19661_, new_n19397_, new_n18977_ );
and  ( new_n19662_, new_n19661_, new_n19660_ );
or   ( new_n19663_, new_n19662_, new_n19659_ );
and  ( new_n19664_, new_n19662_, new_n19659_ );
or   ( new_n19665_, new_n19412_, new_n18066_ );
or   ( new_n19666_, new_n19408_, new_n18309_ );
and  ( new_n19667_, new_n19666_, new_n19665_ );
or   ( new_n19668_, new_n19667_, new_n19664_ );
and  ( new_n19669_, new_n19668_, new_n19663_ );
or   ( new_n19670_, new_n19669_, new_n19653_ );
and  ( new_n19671_, new_n19669_, new_n19653_ );
or   ( new_n19672_, new_n19456_, new_n16085_ );
or   ( new_n19673_, new_n19452_, new_n16048_ );
and  ( new_n19674_, new_n19673_, new_n19672_ );
or   ( new_n19675_, new_n19465_, new_n16052_ );
or   ( new_n19676_, new_n19461_, new_n16071_ );
and  ( new_n19677_, new_n19676_, new_n19675_ );
or   ( new_n19678_, new_n19677_, new_n19674_ );
and  ( new_n19679_, new_n19677_, new_n19674_ );
or   ( new_n19680_, new_n19476_, new_n16009_ );
or   ( new_n19681_, new_n19472_, new_n16029_ );
and  ( new_n19682_, new_n19681_, new_n19680_ );
or   ( new_n19683_, new_n19682_, new_n19679_ );
and  ( new_n19684_, new_n19683_, new_n19678_ );
or   ( new_n19685_, new_n19684_, new_n19671_ );
and  ( new_n19686_, new_n19685_, new_n19670_ );
or   ( new_n19687_, new_n19489_, new_n16186_ );
or   ( new_n19688_, new_n19485_, new_n16204_ );
and  ( new_n19689_, new_n19688_, new_n19687_ );
or   ( new_n19690_, new_n19498_, new_n16217_ );
or   ( new_n19691_, new_n19494_, new_n16234_ );
and  ( new_n19692_, new_n19691_, new_n19690_ );
or   ( new_n19693_, new_n19692_, new_n19689_ );
and  ( new_n19694_, new_n19692_, new_n19689_ );
or   ( new_n19695_, new_n19509_, new_n16151_ );
or   ( new_n19696_, new_n19505_, new_n16170_ );
and  ( new_n19697_, new_n19696_, new_n19695_ );
or   ( new_n19698_, new_n19697_, new_n19694_ );
and  ( new_n19699_, new_n19698_, new_n19693_ );
and  ( new_n19700_, new_n19699_, new_n19149_ );
or   ( new_n19701_, new_n19699_, new_n19149_ );
or   ( new_n19702_, new_n19520_, new_n19330_ );
or   ( new_n19703_, new_n19518_, new_n19178_ );
and  ( new_n19704_, new_n19703_, new_n19702_ );
and  ( new_n19705_, new_n19704_, new_n19701_ );
or   ( new_n19706_, new_n19705_, new_n19700_ );
or   ( new_n19707_, new_n19706_, new_n19686_ );
and  ( new_n19708_, new_n19706_, new_n19686_ );
or   ( new_n19709_, new_n19531_, new_n19314_ );
or   ( new_n19710_, new_n19529_, new_n19144_ );
and  ( new_n19711_, new_n19710_, new_n19709_ );
or   ( new_n19712_, new_n19538_, new_n19299_ );
or   ( new_n19713_, new_n19536_, new_n19111_ );
and  ( new_n19714_, new_n19713_, new_n19712_ );
or   ( new_n19715_, new_n19714_, new_n19711_ );
and  ( new_n19716_, new_n19714_, new_n19711_ );
or   ( new_n19717_, new_n19547_, new_n19286_ );
or   ( new_n19718_, new_n19545_, new_n19080_ );
and  ( new_n19719_, new_n19718_, new_n19717_ );
or   ( new_n19720_, new_n19719_, new_n19716_ );
and  ( new_n19721_, new_n19720_, new_n19715_ );
or   ( new_n19722_, new_n19721_, new_n19708_ );
and  ( new_n19723_, new_n19722_, new_n19707_ );
or   ( new_n19724_, new_n19723_, new_n19640_ );
and  ( new_n19725_, new_n19723_, new_n19640_ );
or   ( new_n19726_, new_n19585_, new_n19365_ );
or   ( new_n19727_, new_n19583_, new_n19232_ );
and  ( new_n19728_, new_n19727_, new_n19726_ );
or   ( new_n19729_, new_n19728_, new_n19725_ );
and  ( new_n19730_, new_n19729_, new_n19724_ );
or   ( new_n19731_, new_n19730_, new_n19388_ );
and  ( new_n19732_, new_n19731_, new_n19627_ );
or   ( new_n19733_, new_n19732_, new_n19623_ );
or   ( new_n19734_, new_n19730_, new_n19626_ );
and  ( new_n19735_, new_n19734_, new_n19590_ );
or   ( new_n19736_, new_n19735_, new_n19598_ );
and  ( new_n19737_, new_n19736_, new_n19733_ );
or   ( new_n19738_, new_n19633_, new_n19560_ );
or   ( new_n19739_, new_n19630_, new_n19567_ );
and  ( new_n19740_, new_n19739_, new_n19738_ );
or   ( new_n19741_, new_n19740_, new_n19638_ );
and  ( new_n19742_, new_n19634_, new_n19568_ );
or   ( new_n19743_, new_n19742_, new_n19576_ );
and  ( new_n19744_, new_n19743_, new_n19741_ );
or   ( new_n19745_, new_n19706_, new_n19482_ );
or   ( new_n19746_, new_n19686_, new_n19524_ );
and  ( new_n19747_, new_n19746_, new_n19745_ );
or   ( new_n19748_, new_n19747_, new_n19721_ );
and  ( new_n19749_, new_n19707_, new_n19525_ );
or   ( new_n19750_, new_n19749_, new_n19551_ );
and  ( new_n19751_, new_n19750_, new_n19748_ );
or   ( new_n19752_, new_n19751_, new_n19744_ );
or   ( new_n19753_, new_n19657_, new_n19655_ );
and  ( new_n19754_, new_n19753_, new_n19393_ );
or   ( new_n19755_, new_n19657_, new_n18738_ );
or   ( new_n19756_, new_n19392_, new_n18973_ );
and  ( new_n19757_, new_n19756_, new_n19755_ );
or   ( new_n19758_, new_n19757_, new_n19754_ );
or   ( new_n19759_, new_n19758_, new_n99_ );
or   ( new_n19760_, new_n19759_, new_n19394_ );
or   ( new_n19761_, new_n19655_, new_n19392_ );
or   ( new_n19762_, new_n19657_, new_n19390_ );
and  ( new_n19763_, new_n19762_, new_n19761_ );
or   ( new_n19764_, new_n19392_, new_n18738_ );
or   ( new_n19765_, new_n19657_, new_n18973_ );
and  ( new_n19766_, new_n19765_, new_n19764_ );
and  ( new_n19767_, new_n19766_, new_n19763_ );
and  ( new_n19768_, new_n19767_, RI2b1c4342d4e0_65 );
or   ( new_n19769_, new_n19768_, new_n19659_ );
and  ( new_n19770_, new_n19769_, new_n19760_ );
or   ( new_n19771_, new_n19048_, new_n112_ );
or   ( new_n19772_, new_n19055_, new_n526_ );
and  ( new_n19773_, new_n19772_, new_n19771_ );
or   ( new_n19774_, new_n19773_, new_n18742_ );
and  ( new_n19775_, new_n19057_, RI2b1c4342d5d0_67 );
and  ( new_n19776_, new_n19044_, RI2b1c4342d558_66 );
or   ( new_n19777_, new_n19776_, new_n19775_ );
or   ( new_n19778_, new_n19777_, new_n18977_ );
and  ( new_n19779_, new_n19778_, new_n19774_ );
or   ( new_n19780_, new_n19779_, new_n19770_ );
and  ( new_n19781_, new_n19779_, new_n19770_ );
or   ( new_n19782_, new_n18388_, new_n591_ );
or   ( new_n19783_, new_n18395_, new_n612_ );
and  ( new_n19784_, new_n19783_, new_n19782_ );
or   ( new_n19785_, new_n19784_, new_n18066_ );
and  ( new_n19786_, new_n18397_, RI2b1c4342d6c0_69 );
and  ( new_n19787_, new_n18384_, RI2b1c4342d648_68 );
or   ( new_n19788_, new_n19787_, new_n19786_ );
or   ( new_n19789_, new_n19788_, new_n18309_ );
and  ( new_n19790_, new_n19789_, new_n19785_ );
or   ( new_n19791_, new_n19790_, new_n19781_ );
and  ( new_n19792_, new_n19791_, new_n19780_ );
or   ( new_n19793_, new_n17727_, new_n110_ );
or   ( new_n19794_, new_n17734_, new_n755_ );
and  ( new_n19795_, new_n19794_, new_n19793_ );
or   ( new_n19796_, new_n19795_, new_n17238_ );
and  ( new_n19797_, new_n17736_, RI2b1c4342d7b0_71 );
and  ( new_n19798_, new_n17723_, RI2b1c4342d738_70 );
or   ( new_n19799_, new_n19798_, new_n19797_ );
or   ( new_n19800_, new_n19799_, new_n17650_ );
and  ( new_n19801_, new_n19800_, new_n19796_ );
or   ( new_n19802_, new_n17244_, new_n105_ );
or   ( new_n19803_, new_n17248_, new_n806_ );
and  ( new_n19804_, new_n19803_, new_n19802_ );
or   ( new_n19805_, new_n19804_, new_n16814_ );
and  ( new_n19806_, new_n17255_, RI2b1c4342d8a0_73 );
and  ( new_n19807_, new_n17240_, RI2b1c4342d828_72 );
or   ( new_n19808_, new_n19807_, new_n19806_ );
or   ( new_n19809_, new_n19808_, new_n17142_ );
and  ( new_n19810_, new_n19809_, new_n19805_ );
or   ( new_n19811_, new_n19810_, new_n19801_ );
and  ( new_n19812_, new_n19810_, new_n19801_ );
or   ( new_n19813_, new_n16607_, new_n843_ );
or   ( new_n19814_, new_n16613_, new_n859_ );
and  ( new_n19815_, new_n19814_, new_n19813_ );
or   ( new_n19816_, new_n19815_, new_n16505_ );
and  ( new_n19817_, new_n16616_, RI2b1c4342d990_75 );
and  ( new_n19818_, new_n16603_, RI2b1c4342d918_74 );
or   ( new_n19819_, new_n19818_, new_n19817_ );
or   ( new_n19820_, new_n19819_, new_n16438_ );
and  ( new_n19821_, new_n19820_, new_n19816_ );
or   ( new_n19822_, new_n19821_, new_n19812_ );
and  ( new_n19823_, new_n19822_, new_n19811_ );
or   ( new_n19824_, new_n19823_, new_n19792_ );
and  ( new_n19825_, new_n19823_, new_n19792_ );
or   ( new_n19826_, new_n16366_, new_n1004_ );
or   ( new_n19827_, new_n16355_, new_n886_ );
and  ( new_n19828_, new_n19827_, new_n19826_ );
or   ( new_n19829_, new_n19828_, new_n16085_ );
and  ( new_n19830_, new_n16358_, RI2b1c4342da80_77 );
and  ( new_n19831_, new_n16362_, RI2b1c4342da08_76 );
or   ( new_n19832_, new_n19831_, new_n19830_ );
or   ( new_n19833_, new_n19832_, new_n16048_ );
and  ( new_n19834_, new_n19833_, new_n19829_ );
or   ( new_n19835_, new_n16075_, new_n1310_ );
or   ( new_n19836_, new_n16060_, new_n1002_ );
and  ( new_n19837_, new_n19836_, new_n19835_ );
or   ( new_n19838_, new_n19837_, new_n16052_ );
and  ( new_n19839_, new_n16063_, RI2b1c4342db70_79 );
and  ( new_n19840_, new_n16066_, RI2b1c4342daf8_78 );
or   ( new_n19841_, new_n19840_, new_n19839_ );
or   ( new_n19842_, new_n19841_, new_n16071_ );
and  ( new_n19843_, new_n19842_, new_n19838_ );
or   ( new_n19844_, new_n19843_, new_n19834_ );
and  ( new_n19845_, new_n19843_, new_n19834_ );
or   ( new_n19846_, new_n16033_, new_n126_ );
or   ( new_n19847_, new_n16017_, new_n1511_ );
and  ( new_n19848_, new_n19847_, new_n19846_ );
or   ( new_n19849_, new_n19848_, new_n16009_ );
and  ( new_n19850_, new_n16021_, RI2b1c4342dc60_81 );
and  ( new_n19851_, new_n16024_, RI2b1c4342dbe8_80 );
or   ( new_n19852_, new_n19851_, new_n19850_ );
or   ( new_n19853_, new_n19852_, new_n16029_ );
and  ( new_n19854_, new_n19853_, new_n19849_ );
or   ( new_n19855_, new_n19854_, new_n19845_ );
and  ( new_n19856_, new_n19855_, new_n19844_ );
or   ( new_n19857_, new_n19856_, new_n19825_ );
and  ( new_n19858_, new_n19857_, new_n19824_ );
or   ( new_n19859_, new_n16119_, new_n132_ );
or   ( new_n19860_, new_n16123_, new_n3902_ );
and  ( new_n19861_, new_n19860_, new_n19859_ );
or   ( new_n19862_, new_n19861_, new_n16108_ );
and  ( new_n19863_, new_n16132_, RI2b1c4342e020_89 );
and  ( new_n19864_, new_n16114_, RI2b1c4342dfa8_88 );
or   ( new_n19865_, new_n19864_, new_n19863_ );
or   ( new_n19866_, new_n19865_, new_n16128_ );
and  ( new_n19867_, new_n19866_, new_n19862_ );
or   ( new_n19868_, new_n16115_, new_n4635_ );
and  ( new_n19869_, new_n19868_, new_n19867_ );
or   ( new_n19870_, new_n16208_, new_n121_ );
or   ( new_n19871_, new_n16194_, new_n2119_ );
and  ( new_n19872_, new_n19871_, new_n19870_ );
or   ( new_n19873_, new_n19872_, new_n16186_ );
and  ( new_n19874_, new_n16196_, RI2b1c4342dd50_83 );
and  ( new_n19875_, new_n16199_, RI2b1c4342dcd8_82 );
or   ( new_n19876_, new_n19875_, new_n19874_ );
or   ( new_n19877_, new_n19876_, new_n16204_ );
and  ( new_n19878_, new_n19877_, new_n19873_ );
or   ( new_n19879_, new_n16238_, new_n2806_ );
or   ( new_n19880_, new_n16224_, new_n2541_ );
and  ( new_n19881_, new_n19880_, new_n19879_ );
or   ( new_n19882_, new_n19881_, new_n16217_ );
and  ( new_n19883_, new_n16226_, RI2b1c4342de40_85 );
and  ( new_n19884_, new_n16229_, RI2b1c4342ddc8_84 );
or   ( new_n19885_, new_n19884_, new_n19883_ );
or   ( new_n19886_, new_n19885_, new_n16234_ );
and  ( new_n19887_, new_n19886_, new_n19882_ );
or   ( new_n19888_, new_n19887_, new_n19878_ );
and  ( new_n19889_, new_n19887_, new_n19878_ );
or   ( new_n19890_, new_n16174_, new_n3924_ );
or   ( new_n19891_, new_n16160_, new_n3239_ );
and  ( new_n19892_, new_n19891_, new_n19890_ );
or   ( new_n19893_, new_n19892_, new_n16151_ );
and  ( new_n19894_, new_n16162_, RI2b1c4342df30_87 );
and  ( new_n19895_, new_n16165_, RI2b1c4342deb8_86 );
or   ( new_n19896_, new_n19895_, new_n19894_ );
or   ( new_n19897_, new_n19896_, new_n16170_ );
and  ( new_n19898_, new_n19897_, new_n19893_ );
or   ( new_n19899_, new_n19898_, new_n19889_ );
and  ( new_n19900_, new_n19899_, new_n19888_ );
or   ( new_n19901_, new_n19900_, new_n19869_ );
and  ( new_n19902_, new_n19900_, new_n19869_ );
or   ( new_n19903_, new_n16119_, new_n3902_ );
or   ( new_n19904_, new_n16123_, new_n3924_ );
and  ( new_n19905_, new_n19904_, new_n19903_ );
or   ( new_n19906_, new_n19905_, new_n16108_ );
and  ( new_n19907_, new_n16132_, RI2b1c4342dfa8_88 );
and  ( new_n19908_, new_n16114_, RI2b1c4342df30_87 );
or   ( new_n19909_, new_n19908_, new_n19907_ );
or   ( new_n19910_, new_n19909_, new_n16128_ );
and  ( new_n19911_, new_n19910_, new_n19906_ );
or   ( new_n19912_, new_n19911_, new_n19902_ );
and  ( new_n19913_, new_n19912_, new_n19901_ );
or   ( new_n19914_, new_n19913_, new_n19858_ );
and  ( new_n19915_, new_n19913_, new_n19858_ );
or   ( new_n19916_, new_n16115_, new_n132_ );
or   ( new_n19917_, new_n19692_, new_n19491_ );
or   ( new_n19918_, new_n19689_, new_n19500_ );
and  ( new_n19919_, new_n19918_, new_n19917_ );
or   ( new_n19920_, new_n19919_, new_n19697_ );
and  ( new_n19921_, new_n19693_, new_n19501_ );
or   ( new_n19922_, new_n19921_, new_n19511_ );
and  ( new_n19923_, new_n19922_, new_n19920_ );
or   ( new_n19924_, new_n19923_, new_n19916_ );
and  ( new_n19925_, new_n19923_, new_n19916_ );
or   ( new_n19926_, new_n19677_, new_n19458_ );
or   ( new_n19927_, new_n19674_, new_n19467_ );
and  ( new_n19928_, new_n19927_, new_n19926_ );
or   ( new_n19929_, new_n19928_, new_n19682_ );
and  ( new_n19930_, new_n19678_, new_n19468_ );
or   ( new_n19931_, new_n19930_, new_n19478_ );
and  ( new_n19932_, new_n19931_, new_n19929_ );
or   ( new_n19933_, new_n19932_, new_n19925_ );
and  ( new_n19934_, new_n19933_, new_n19924_ );
or   ( new_n19935_, new_n19934_, new_n19915_ );
and  ( new_n19936_, new_n19935_, new_n19914_ );
or   ( new_n19937_, new_n19714_, new_n19533_ );
or   ( new_n19938_, new_n19711_, new_n19540_ );
and  ( new_n19939_, new_n19938_, new_n19937_ );
or   ( new_n19940_, new_n19939_, new_n19719_ );
and  ( new_n19941_, new_n19715_, new_n19541_ );
or   ( new_n19942_, new_n19941_, new_n19549_ );
and  ( new_n19943_, new_n19942_, new_n19940_ );
or   ( new_n19944_, new_n19513_, new_n19149_ );
or   ( new_n19945_, new_n19699_, new_n19319_ );
and  ( new_n19946_, new_n19945_, new_n19944_ );
or   ( new_n19947_, new_n19946_, new_n19704_ );
and  ( new_n19948_, new_n19701_, new_n19514_ );
or   ( new_n19949_, new_n19948_, new_n19522_ );
and  ( new_n19950_, new_n19949_, new_n19947_ );
or   ( new_n19951_, new_n19950_, new_n19943_ );
and  ( new_n19952_, new_n19950_, new_n19943_ );
or   ( new_n19953_, new_n19653_, new_n19416_ );
or   ( new_n19954_, new_n19669_, new_n19447_ );
and  ( new_n19955_, new_n19954_, new_n19953_ );
or   ( new_n19956_, new_n19955_, new_n19684_ );
and  ( new_n19957_, new_n19670_, new_n19448_ );
or   ( new_n19958_, new_n19957_, new_n19480_ );
and  ( new_n19959_, new_n19958_, new_n19956_ );
or   ( new_n19960_, new_n19959_, new_n19952_ );
and  ( new_n19961_, new_n19960_, new_n19951_ );
or   ( new_n19962_, new_n19961_, new_n19936_ );
and  ( new_n19963_, new_n19961_, new_n19936_ );
or   ( new_n19964_, new_n19301_, new_n19082_ );
or   ( new_n19965_, new_n19288_, new_n19113_ );
and  ( new_n19966_, new_n19965_, new_n19964_ );
or   ( new_n19967_, new_n19966_, new_n19316_ );
and  ( new_n19968_, new_n19302_, new_n19114_ );
or   ( new_n19969_, new_n19968_, new_n19146_ );
and  ( new_n19970_, new_n19969_, new_n19967_ );
or   ( new_n19971_, new_n19970_, new_n19963_ );
and  ( new_n19972_, new_n19971_, new_n19962_ );
or   ( new_n19973_, new_n19972_, new_n19752_ );
and  ( new_n19974_, new_n19972_, new_n19752_ );
or   ( new_n19975_, new_n19337_, new_n19148_ );
or   ( new_n19976_, new_n19318_, new_n19185_ );
and  ( new_n19977_, new_n19976_, new_n19975_ );
or   ( new_n19978_, new_n19977_, new_n19352_ );
and  ( new_n19979_, new_n19338_, new_n19186_ );
or   ( new_n19980_, new_n19979_, new_n19212_ );
and  ( new_n19981_, new_n19980_, new_n19978_ );
or   ( new_n19982_, new_n19981_, new_n19974_ );
and  ( new_n19983_, new_n19982_, new_n19973_ );
or   ( new_n19984_, new_n19983_, new_n19737_ );
or   ( new_n19985_, new_n19379_, new_n19271_ );
or   ( new_n19986_, new_n19376_, new_n19254_ );
and  ( new_n19987_, new_n19986_, new_n19985_ );
or   ( new_n19988_, new_n19987_, new_n19600_ );
and  ( new_n19989_, new_n19730_, new_n19626_ );
or   ( new_n19990_, new_n19989_, new_n19623_ );
and  ( new_n19991_, new_n19990_, new_n19734_ );
or   ( new_n19992_, new_n19991_, new_n19381_ );
and  ( new_n19993_, new_n19992_, new_n19988_ );
or   ( new_n19994_, new_n19993_, new_n19984_ );
and  ( new_n19995_, new_n19993_, new_n19984_ );
or   ( new_n19996_, new_n19735_, new_n19623_ );
or   ( new_n19997_, new_n19732_, new_n19598_ );
and  ( new_n19998_, new_n19997_, new_n19996_ );
or   ( new_n19999_, new_n19998_, new_n19983_ );
or   ( new_n20000_, new_n19742_, new_n19638_ );
or   ( new_n20001_, new_n19740_, new_n19576_ );
and  ( new_n20002_, new_n20001_, new_n20000_ );
or   ( new_n20003_, new_n19749_, new_n19721_ );
or   ( new_n20004_, new_n19747_, new_n19551_ );
and  ( new_n20005_, new_n20004_, new_n20003_ );
and  ( new_n20006_, new_n20005_, new_n20002_ );
or   ( new_n20007_, new_n19768_, new_n19394_ );
or   ( new_n20008_, new_n19759_, new_n19659_ );
and  ( new_n20009_, new_n20008_, new_n20007_ );
or   ( new_n20010_, new_n19777_, new_n18742_ );
or   ( new_n20011_, new_n19773_, new_n18977_ );
and  ( new_n20012_, new_n20011_, new_n20010_ );
or   ( new_n20013_, new_n20012_, new_n20009_ );
and  ( new_n20014_, new_n20012_, new_n20009_ );
or   ( new_n20015_, new_n19788_, new_n18066_ );
or   ( new_n20016_, new_n19784_, new_n18309_ );
and  ( new_n20017_, new_n20016_, new_n20015_ );
or   ( new_n20018_, new_n20017_, new_n20014_ );
and  ( new_n20019_, new_n20018_, new_n20013_ );
or   ( new_n20020_, new_n19799_, new_n17238_ );
or   ( new_n20021_, new_n19795_, new_n17650_ );
and  ( new_n20022_, new_n20021_, new_n20020_ );
or   ( new_n20023_, new_n19808_, new_n16814_ );
or   ( new_n20024_, new_n19804_, new_n17142_ );
and  ( new_n20025_, new_n20024_, new_n20023_ );
or   ( new_n20026_, new_n20025_, new_n20022_ );
and  ( new_n20027_, new_n20025_, new_n20022_ );
or   ( new_n20028_, new_n19819_, new_n16505_ );
or   ( new_n20029_, new_n19815_, new_n16438_ );
and  ( new_n20030_, new_n20029_, new_n20028_ );
or   ( new_n20031_, new_n20030_, new_n20027_ );
and  ( new_n20032_, new_n20031_, new_n20026_ );
or   ( new_n20033_, new_n20032_, new_n20019_ );
and  ( new_n20034_, new_n20032_, new_n20019_ );
or   ( new_n20035_, new_n19832_, new_n16085_ );
or   ( new_n20036_, new_n19828_, new_n16048_ );
and  ( new_n20037_, new_n20036_, new_n20035_ );
or   ( new_n20038_, new_n19841_, new_n16052_ );
or   ( new_n20039_, new_n19837_, new_n16071_ );
and  ( new_n20040_, new_n20039_, new_n20038_ );
or   ( new_n20041_, new_n20040_, new_n20037_ );
and  ( new_n20042_, new_n20040_, new_n20037_ );
or   ( new_n20043_, new_n19852_, new_n16009_ );
or   ( new_n20044_, new_n19848_, new_n16029_ );
and  ( new_n20045_, new_n20044_, new_n20043_ );
or   ( new_n20046_, new_n20045_, new_n20042_ );
and  ( new_n20047_, new_n20046_, new_n20041_ );
or   ( new_n20048_, new_n20047_, new_n20034_ );
and  ( new_n20049_, new_n20048_, new_n20033_ );
and  ( new_n20050_, new_n16102_, RI2b1c4342e098_90 );
or   ( new_n20051_, new_n19865_, new_n16108_ );
or   ( new_n20052_, new_n19861_, new_n16128_ );
and  ( new_n20053_, new_n20052_, new_n20051_ );
or   ( new_n20054_, new_n20053_, new_n20050_ );
or   ( new_n20055_, new_n19876_, new_n16186_ );
or   ( new_n20056_, new_n19872_, new_n16204_ );
and  ( new_n20057_, new_n20056_, new_n20055_ );
or   ( new_n20058_, new_n19885_, new_n16217_ );
or   ( new_n20059_, new_n19881_, new_n16234_ );
and  ( new_n20060_, new_n20059_, new_n20058_ );
or   ( new_n20061_, new_n20060_, new_n20057_ );
and  ( new_n20062_, new_n20060_, new_n20057_ );
or   ( new_n20063_, new_n19896_, new_n16151_ );
or   ( new_n20064_, new_n19892_, new_n16170_ );
and  ( new_n20065_, new_n20064_, new_n20063_ );
or   ( new_n20066_, new_n20065_, new_n20062_ );
and  ( new_n20067_, new_n20066_, new_n20061_ );
or   ( new_n20068_, new_n20067_, new_n20054_ );
and  ( new_n20069_, new_n20067_, new_n20054_ );
or   ( new_n20070_, new_n19909_, new_n16108_ );
or   ( new_n20071_, new_n19905_, new_n16128_ );
and  ( new_n20072_, new_n20071_, new_n20070_ );
or   ( new_n20073_, new_n20072_, new_n20069_ );
and  ( new_n20074_, new_n20073_, new_n20068_ );
or   ( new_n20075_, new_n20074_, new_n20049_ );
and  ( new_n20076_, new_n20074_, new_n20049_ );
and  ( new_n20077_, new_n16102_, RI2b1c4342e020_89 );
or   ( new_n20078_, new_n19921_, new_n19697_ );
or   ( new_n20079_, new_n19919_, new_n19511_ );
and  ( new_n20080_, new_n20079_, new_n20078_ );
or   ( new_n20081_, new_n20080_, new_n20077_ );
and  ( new_n20082_, new_n20080_, new_n20077_ );
or   ( new_n20083_, new_n19930_, new_n19682_ );
or   ( new_n20084_, new_n19928_, new_n19478_ );
and  ( new_n20085_, new_n20084_, new_n20083_ );
or   ( new_n20086_, new_n20085_, new_n20082_ );
and  ( new_n20087_, new_n20086_, new_n20081_ );
or   ( new_n20088_, new_n20087_, new_n20076_ );
and  ( new_n20089_, new_n20088_, new_n20075_ );
or   ( new_n20090_, new_n19941_, new_n19719_ );
or   ( new_n20091_, new_n19939_, new_n19549_ );
and  ( new_n20092_, new_n20091_, new_n20090_ );
or   ( new_n20093_, new_n19948_, new_n19704_ );
or   ( new_n20094_, new_n19946_, new_n19522_ );
and  ( new_n20095_, new_n20094_, new_n20093_ );
or   ( new_n20096_, new_n20095_, new_n20092_ );
and  ( new_n20097_, new_n20095_, new_n20092_ );
or   ( new_n20098_, new_n19957_, new_n19684_ );
or   ( new_n20099_, new_n19955_, new_n19480_ );
and  ( new_n20100_, new_n20099_, new_n20098_ );
or   ( new_n20101_, new_n20100_, new_n20097_ );
and  ( new_n20102_, new_n20101_, new_n20096_ );
or   ( new_n20103_, new_n20102_, new_n20089_ );
and  ( new_n20104_, new_n20102_, new_n20089_ );
or   ( new_n20105_, new_n19968_, new_n19316_ );
or   ( new_n20106_, new_n19966_, new_n19146_ );
and  ( new_n20107_, new_n20106_, new_n20105_ );
or   ( new_n20108_, new_n20107_, new_n20104_ );
and  ( new_n20109_, new_n20108_, new_n20103_ );
or   ( new_n20110_, new_n20109_, new_n20006_ );
and  ( new_n20111_, new_n20109_, new_n20006_ );
or   ( new_n20112_, new_n19979_, new_n19352_ );
or   ( new_n20113_, new_n19977_, new_n19212_ );
and  ( new_n20114_, new_n20113_, new_n20112_ );
or   ( new_n20115_, new_n20114_, new_n20111_ );
and  ( new_n20116_, new_n20115_, new_n20110_ );
or   ( new_n20117_, new_n20116_, new_n19737_ );
and  ( new_n20118_, new_n20117_, new_n19999_ );
or   ( new_n20119_, new_n19640_, new_n19553_ );
or   ( new_n20120_, new_n19723_, new_n19578_ );
and  ( new_n20121_, new_n20120_, new_n20119_ );
or   ( new_n20122_, new_n20121_, new_n19728_ );
and  ( new_n20123_, new_n19724_, new_n19579_ );
or   ( new_n20124_, new_n20123_, new_n19587_ );
and  ( new_n20125_, new_n20124_, new_n20122_ );
or   ( new_n20126_, new_n19646_, new_n19425_ );
or   ( new_n20127_, new_n19643_, new_n19434_ );
and  ( new_n20128_, new_n20127_, new_n20126_ );
or   ( new_n20129_, new_n20128_, new_n19651_ );
and  ( new_n20130_, new_n19647_, new_n19435_ );
or   ( new_n20131_, new_n20130_, new_n19445_ );
and  ( new_n20132_, new_n20131_, new_n20129_ );
or   ( new_n20133_, new_n19662_, new_n19394_ );
or   ( new_n20134_, new_n19659_, new_n19403_ );
and  ( new_n20135_, new_n20134_, new_n20133_ );
or   ( new_n20136_, new_n20135_, new_n19667_ );
and  ( new_n20137_, new_n19663_, new_n19404_ );
or   ( new_n20138_, new_n20137_, new_n19414_ );
and  ( new_n20139_, new_n20138_, new_n20136_ );
or   ( new_n20140_, new_n20139_, new_n20132_ );
and  ( new_n20141_, new_n20139_, new_n20132_ );
or   ( new_n20142_, new_n20080_, new_n19916_ );
or   ( new_n20143_, new_n20077_, new_n19923_ );
and  ( new_n20144_, new_n20143_, new_n20142_ );
or   ( new_n20145_, new_n20144_, new_n20085_ );
and  ( new_n20146_, new_n20081_, new_n19924_ );
or   ( new_n20147_, new_n20146_, new_n19932_ );
and  ( new_n20148_, new_n20147_, new_n20145_ );
or   ( new_n20149_, new_n20148_, new_n20141_ );
and  ( new_n20150_, new_n20149_, new_n20140_ );
xor  ( new_n20151_, new_n5015_, new_n5172_ );
or   ( new_n20152_, new_n20151_, new_n326_ );
xor  ( new_n20153_, new_n5022_, new_n221_ );
or   ( new_n20154_, new_n20153_, new_n323_ );
or   ( new_n20155_, new_n20154_, new_n20152_ );
and  ( new_n20156_, new_n20155_, new_n19655_ );
or   ( new_n20157_, new_n19758_, new_n526_ );
or   ( new_n20158_, new_n19763_, new_n99_ );
and  ( new_n20159_, new_n20158_, new_n20157_ );
or   ( new_n20160_, new_n20159_, new_n19394_ );
and  ( new_n20161_, new_n19767_, RI2b1c4342d558_66 );
and  ( new_n20162_, new_n19754_, RI2b1c4342d4e0_65 );
or   ( new_n20163_, new_n20162_, new_n20161_ );
or   ( new_n20164_, new_n20163_, new_n19659_ );
and  ( new_n20165_, new_n20164_, new_n20160_ );
or   ( new_n20166_, new_n20165_, new_n20156_ );
and  ( new_n20167_, new_n20165_, new_n20156_ );
or   ( new_n20168_, new_n19048_, new_n612_ );
or   ( new_n20169_, new_n19055_, new_n112_ );
and  ( new_n20170_, new_n20169_, new_n20168_ );
or   ( new_n20171_, new_n20170_, new_n18742_ );
and  ( new_n20172_, new_n19057_, RI2b1c4342d648_68 );
and  ( new_n20173_, new_n19044_, RI2b1c4342d5d0_67 );
or   ( new_n20174_, new_n20173_, new_n20172_ );
or   ( new_n20175_, new_n20174_, new_n18977_ );
and  ( new_n20176_, new_n20175_, new_n20171_ );
or   ( new_n20177_, new_n20176_, new_n20167_ );
and  ( new_n20178_, new_n20177_, new_n20166_ );
or   ( new_n20179_, new_n18388_, new_n755_ );
or   ( new_n20180_, new_n18395_, new_n591_ );
and  ( new_n20181_, new_n20180_, new_n20179_ );
or   ( new_n20182_, new_n20181_, new_n18066_ );
and  ( new_n20183_, new_n18397_, RI2b1c4342d738_70 );
and  ( new_n20184_, new_n18384_, RI2b1c4342d6c0_69 );
or   ( new_n20185_, new_n20184_, new_n20183_ );
or   ( new_n20186_, new_n20185_, new_n18309_ );
and  ( new_n20187_, new_n20186_, new_n20182_ );
or   ( new_n20188_, new_n17727_, new_n806_ );
or   ( new_n20189_, new_n17734_, new_n110_ );
and  ( new_n20190_, new_n20189_, new_n20188_ );
or   ( new_n20191_, new_n20190_, new_n17238_ );
and  ( new_n20192_, new_n17736_, RI2b1c4342d828_72 );
and  ( new_n20193_, new_n17723_, RI2b1c4342d7b0_71 );
or   ( new_n20194_, new_n20193_, new_n20192_ );
or   ( new_n20195_, new_n20194_, new_n17650_ );
and  ( new_n20196_, new_n20195_, new_n20191_ );
or   ( new_n20197_, new_n20196_, new_n20187_ );
and  ( new_n20198_, new_n20196_, new_n20187_ );
or   ( new_n20199_, new_n17244_, new_n859_ );
or   ( new_n20200_, new_n17248_, new_n105_ );
and  ( new_n20201_, new_n20200_, new_n20199_ );
or   ( new_n20202_, new_n20201_, new_n16814_ );
and  ( new_n20203_, new_n17255_, RI2b1c4342d918_74 );
and  ( new_n20204_, new_n17240_, RI2b1c4342d8a0_73 );
or   ( new_n20205_, new_n20204_, new_n20203_ );
or   ( new_n20206_, new_n20205_, new_n17142_ );
and  ( new_n20207_, new_n20206_, new_n20202_ );
or   ( new_n20208_, new_n20207_, new_n20198_ );
and  ( new_n20209_, new_n20208_, new_n20197_ );
or   ( new_n20210_, new_n20209_, new_n20178_ );
and  ( new_n20211_, new_n20209_, new_n20178_ );
or   ( new_n20212_, new_n16607_, new_n886_ );
or   ( new_n20213_, new_n16613_, new_n843_ );
and  ( new_n20214_, new_n20213_, new_n20212_ );
or   ( new_n20215_, new_n20214_, new_n16505_ );
and  ( new_n20216_, new_n16616_, RI2b1c4342da08_76 );
and  ( new_n20217_, new_n16603_, RI2b1c4342d990_75 );
or   ( new_n20218_, new_n20217_, new_n20216_ );
or   ( new_n20219_, new_n20218_, new_n16438_ );
and  ( new_n20220_, new_n20219_, new_n20215_ );
or   ( new_n20221_, new_n16366_, new_n1002_ );
or   ( new_n20222_, new_n16355_, new_n1004_ );
and  ( new_n20223_, new_n20222_, new_n20221_ );
or   ( new_n20224_, new_n20223_, new_n16085_ );
and  ( new_n20225_, new_n16358_, RI2b1c4342daf8_78 );
and  ( new_n20226_, new_n16362_, RI2b1c4342da80_77 );
or   ( new_n20227_, new_n20226_, new_n20225_ );
or   ( new_n20228_, new_n20227_, new_n16048_ );
and  ( new_n20229_, new_n20228_, new_n20224_ );
or   ( new_n20230_, new_n20229_, new_n20220_ );
and  ( new_n20231_, new_n20229_, new_n20220_ );
or   ( new_n20232_, new_n16075_, new_n1511_ );
or   ( new_n20233_, new_n16060_, new_n1310_ );
and  ( new_n20234_, new_n20233_, new_n20232_ );
or   ( new_n20235_, new_n20234_, new_n16052_ );
and  ( new_n20236_, new_n16063_, RI2b1c4342dbe8_80 );
and  ( new_n20237_, new_n16066_, RI2b1c4342db70_79 );
or   ( new_n20238_, new_n20237_, new_n20236_ );
or   ( new_n20239_, new_n20238_, new_n16071_ );
and  ( new_n20240_, new_n20239_, new_n20235_ );
or   ( new_n20241_, new_n20240_, new_n20231_ );
and  ( new_n20242_, new_n20241_, new_n20230_ );
or   ( new_n20243_, new_n20242_, new_n20211_ );
and  ( new_n20244_, new_n20243_, new_n20210_ );
or   ( new_n20245_, new_n16033_, new_n2119_ );
or   ( new_n20246_, new_n16017_, new_n126_ );
and  ( new_n20247_, new_n20246_, new_n20245_ );
or   ( new_n20248_, new_n20247_, new_n16009_ );
and  ( new_n20249_, new_n16021_, RI2b1c4342dcd8_82 );
and  ( new_n20250_, new_n16024_, RI2b1c4342dc60_81 );
or   ( new_n20251_, new_n20250_, new_n20249_ );
or   ( new_n20252_, new_n20251_, new_n16029_ );
and  ( new_n20253_, new_n20252_, new_n20248_ );
or   ( new_n20254_, new_n16208_, new_n2541_ );
or   ( new_n20255_, new_n16194_, new_n121_ );
and  ( new_n20256_, new_n20255_, new_n20254_ );
or   ( new_n20257_, new_n20256_, new_n16186_ );
and  ( new_n20258_, new_n16196_, RI2b1c4342ddc8_84 );
and  ( new_n20259_, new_n16199_, RI2b1c4342dd50_83 );
or   ( new_n20260_, new_n20259_, new_n20258_ );
or   ( new_n20261_, new_n20260_, new_n16204_ );
and  ( new_n20262_, new_n20261_, new_n20257_ );
or   ( new_n20263_, new_n20262_, new_n20253_ );
and  ( new_n20264_, new_n20262_, new_n20253_ );
or   ( new_n20265_, new_n16238_, new_n3239_ );
or   ( new_n20266_, new_n16224_, new_n2806_ );
and  ( new_n20267_, new_n20266_, new_n20265_ );
or   ( new_n20268_, new_n20267_, new_n16217_ );
and  ( new_n20269_, new_n16226_, RI2b1c4342deb8_86 );
and  ( new_n20270_, new_n16229_, RI2b1c4342de40_85 );
or   ( new_n20271_, new_n20270_, new_n20269_ );
or   ( new_n20272_, new_n20271_, new_n16234_ );
and  ( new_n20273_, new_n20272_, new_n20268_ );
or   ( new_n20274_, new_n20273_, new_n20264_ );
and  ( new_n20275_, new_n20274_, new_n20263_ );
or   ( new_n20276_, new_n16174_, new_n3902_ );
or   ( new_n20277_, new_n16160_, new_n3924_ );
and  ( new_n20278_, new_n20277_, new_n20276_ );
or   ( new_n20279_, new_n20278_, new_n16151_ );
and  ( new_n20280_, new_n16162_, RI2b1c4342dfa8_88 );
and  ( new_n20281_, new_n16165_, RI2b1c4342df30_87 );
or   ( new_n20282_, new_n20281_, new_n20280_ );
or   ( new_n20283_, new_n20282_, new_n16170_ );
and  ( new_n20284_, new_n20283_, new_n20279_ );
or   ( new_n20285_, new_n16119_, new_n4635_ );
or   ( new_n20286_, new_n16123_, new_n132_ );
and  ( new_n20287_, new_n20286_, new_n20285_ );
or   ( new_n20288_, new_n20287_, new_n16108_ );
and  ( new_n20289_, new_n16132_, RI2b1c4342e098_90 );
and  ( new_n20290_, new_n16114_, RI2b1c4342e020_89 );
or   ( new_n20291_, new_n20290_, new_n20289_ );
or   ( new_n20292_, new_n20291_, new_n16128_ );
and  ( new_n20293_, new_n20292_, new_n20288_ );
and  ( new_n20294_, new_n20293_, new_n20284_ );
or   ( new_n20295_, new_n20293_, new_n20284_ );
or   ( new_n20296_, new_n16115_, new_n117_ );
and  ( new_n20297_, new_n20296_, new_n20295_ );
or   ( new_n20298_, new_n20297_, new_n20294_ );
and  ( new_n20299_, new_n20298_, new_n20275_ );
or   ( new_n20300_, new_n20298_, new_n20275_ );
or   ( new_n20301_, new_n19868_, new_n19867_ );
and  ( new_n20302_, new_n20301_, new_n20054_ );
and  ( new_n20303_, new_n20302_, new_n20300_ );
or   ( new_n20304_, new_n20303_, new_n20299_ );
and  ( new_n20305_, new_n20304_, new_n20244_ );
or   ( new_n20306_, new_n20304_, new_n20244_ );
or   ( new_n20307_, new_n20060_, new_n19878_ );
or   ( new_n20308_, new_n20057_, new_n19887_ );
and  ( new_n20309_, new_n20308_, new_n20307_ );
or   ( new_n20310_, new_n20309_, new_n20065_ );
and  ( new_n20311_, new_n20061_, new_n19888_ );
or   ( new_n20312_, new_n20311_, new_n19898_ );
and  ( new_n20313_, new_n20312_, new_n20310_ );
or   ( new_n20314_, new_n20040_, new_n19834_ );
or   ( new_n20315_, new_n20037_, new_n19843_ );
and  ( new_n20316_, new_n20315_, new_n20314_ );
or   ( new_n20317_, new_n20316_, new_n20045_ );
and  ( new_n20318_, new_n20041_, new_n19844_ );
or   ( new_n20319_, new_n20318_, new_n19854_ );
and  ( new_n20320_, new_n20319_, new_n20317_ );
or   ( new_n20321_, new_n20320_, new_n20313_ );
and  ( new_n20322_, new_n20320_, new_n20313_ );
or   ( new_n20323_, new_n20025_, new_n19801_ );
or   ( new_n20324_, new_n20022_, new_n19810_ );
and  ( new_n20325_, new_n20324_, new_n20323_ );
or   ( new_n20326_, new_n20325_, new_n20030_ );
and  ( new_n20327_, new_n20026_, new_n19811_ );
or   ( new_n20328_, new_n20327_, new_n19821_ );
and  ( new_n20329_, new_n20328_, new_n20326_ );
or   ( new_n20330_, new_n20329_, new_n20322_ );
and  ( new_n20331_, new_n20330_, new_n20321_ );
and  ( new_n20332_, new_n20331_, new_n20306_ );
or   ( new_n20333_, new_n20332_, new_n20305_ );
and  ( new_n20334_, new_n20333_, new_n20150_ );
or   ( new_n20335_, new_n20333_, new_n20150_ );
or   ( new_n20336_, new_n20095_, new_n19943_ );
or   ( new_n20337_, new_n20092_, new_n19950_ );
and  ( new_n20338_, new_n20337_, new_n20336_ );
or   ( new_n20339_, new_n20338_, new_n20100_ );
and  ( new_n20340_, new_n20096_, new_n19951_ );
or   ( new_n20341_, new_n20340_, new_n19959_ );
and  ( new_n20342_, new_n20341_, new_n20339_ );
and  ( new_n20343_, new_n20342_, new_n20335_ );
or   ( new_n20344_, new_n20343_, new_n20334_ );
or   ( new_n20345_, new_n20005_, new_n19744_ );
or   ( new_n20346_, new_n20002_, new_n19751_ );
and  ( new_n20347_, new_n20346_, new_n20345_ );
and  ( new_n20348_, new_n20347_, new_n20344_ );
or   ( new_n20349_, new_n20347_, new_n20344_ );
or   ( new_n20350_, new_n20102_, new_n19936_ );
or   ( new_n20351_, new_n20089_, new_n19961_ );
and  ( new_n20352_, new_n20351_, new_n20350_ );
or   ( new_n20353_, new_n20352_, new_n20107_ );
and  ( new_n20354_, new_n20103_, new_n19962_ );
or   ( new_n20355_, new_n20354_, new_n19970_ );
and  ( new_n20356_, new_n20355_, new_n20353_ );
and  ( new_n20357_, new_n20356_, new_n20349_ );
or   ( new_n20358_, new_n20357_, new_n20348_ );
and  ( new_n20359_, new_n20358_, new_n20125_ );
or   ( new_n20360_, new_n20358_, new_n20125_ );
or   ( new_n20361_, new_n20006_, new_n19972_ );
or   ( new_n20362_, new_n20109_, new_n19752_ );
and  ( new_n20363_, new_n20362_, new_n20361_ );
or   ( new_n20364_, new_n20363_, new_n20114_ );
and  ( new_n20365_, new_n20110_, new_n19973_ );
or   ( new_n20366_, new_n20365_, new_n19981_ );
and  ( new_n20367_, new_n20366_, new_n20364_ );
and  ( new_n20368_, new_n20367_, new_n20360_ );
or   ( new_n20369_, new_n20368_, new_n20359_ );
or   ( new_n20370_, new_n20369_, new_n20118_ );
or   ( new_n20371_, new_n20370_, new_n19995_ );
and  ( new_n20372_, new_n20371_, new_n19994_ );
and  ( new_n20373_, new_n20369_, new_n20118_ );
or   ( new_n20374_, new_n20373_, new_n19995_ );
or   ( new_n20375_, new_n20354_, new_n20107_ );
or   ( new_n20376_, new_n20352_, new_n19970_ );
and  ( new_n20377_, new_n20376_, new_n20375_ );
or   ( new_n20378_, new_n20005_, new_n20002_ );
and  ( new_n20379_, new_n20378_, new_n19752_ );
or   ( new_n20380_, new_n20379_, new_n20344_ );
or   ( new_n20381_, new_n20130_, new_n19651_ );
or   ( new_n20382_, new_n20128_, new_n19445_ );
and  ( new_n20383_, new_n20382_, new_n20381_ );
or   ( new_n20384_, new_n20137_, new_n19667_ );
or   ( new_n20385_, new_n20135_, new_n19414_ );
and  ( new_n20386_, new_n20385_, new_n20384_ );
or   ( new_n20387_, new_n20386_, new_n20383_ );
and  ( new_n20388_, new_n20386_, new_n20383_ );
or   ( new_n20389_, new_n20146_, new_n20085_ );
or   ( new_n20390_, new_n20144_, new_n19932_ );
and  ( new_n20391_, new_n20390_, new_n20389_ );
or   ( new_n20392_, new_n20391_, new_n20388_ );
and  ( new_n20393_, new_n20392_, new_n20387_ );
or   ( new_n20394_, new_n20251_, new_n16009_ );
or   ( new_n20395_, new_n20247_, new_n16029_ );
and  ( new_n20396_, new_n20395_, new_n20394_ );
or   ( new_n20397_, new_n20260_, new_n16186_ );
or   ( new_n20398_, new_n20256_, new_n16204_ );
and  ( new_n20399_, new_n20398_, new_n20397_ );
or   ( new_n20400_, new_n20399_, new_n20396_ );
and  ( new_n20401_, new_n20399_, new_n20396_ );
or   ( new_n20402_, new_n20271_, new_n16217_ );
or   ( new_n20403_, new_n20267_, new_n16234_ );
and  ( new_n20404_, new_n20403_, new_n20402_ );
or   ( new_n20405_, new_n20404_, new_n20401_ );
and  ( new_n20406_, new_n20405_, new_n20400_ );
or   ( new_n20407_, new_n20282_, new_n16151_ );
or   ( new_n20408_, new_n20278_, new_n16170_ );
and  ( new_n20409_, new_n20408_, new_n20407_ );
or   ( new_n20410_, new_n20291_, new_n16108_ );
or   ( new_n20411_, new_n20287_, new_n16128_ );
and  ( new_n20412_, new_n20411_, new_n20410_ );
or   ( new_n20413_, new_n20412_, new_n20409_ );
and  ( new_n20414_, new_n20412_, new_n20409_ );
and  ( new_n20415_, new_n16102_, RI2b1c4342e110_91 );
or   ( new_n20416_, new_n20415_, new_n20414_ );
and  ( new_n20417_, new_n20416_, new_n20413_ );
or   ( new_n20418_, new_n20417_, new_n20406_ );
and  ( new_n20419_, new_n20417_, new_n20406_ );
or   ( new_n20420_, new_n20050_, new_n19867_ );
or   ( new_n20421_, new_n20053_, new_n19868_ );
and  ( new_n20422_, new_n20421_, new_n20420_ );
or   ( new_n20423_, new_n20422_, new_n20419_ );
and  ( new_n20424_, new_n20423_, new_n20418_ );
or   ( new_n20425_, new_n20185_, new_n18066_ );
or   ( new_n20426_, new_n20181_, new_n18309_ );
and  ( new_n20427_, new_n20426_, new_n20425_ );
or   ( new_n20428_, new_n20194_, new_n17238_ );
or   ( new_n20429_, new_n20190_, new_n17650_ );
and  ( new_n20430_, new_n20429_, new_n20428_ );
or   ( new_n20431_, new_n20430_, new_n20427_ );
and  ( new_n20432_, new_n20430_, new_n20427_ );
or   ( new_n20433_, new_n20205_, new_n16814_ );
or   ( new_n20434_, new_n20201_, new_n17142_ );
and  ( new_n20435_, new_n20434_, new_n20433_ );
or   ( new_n20436_, new_n20435_, new_n20432_ );
and  ( new_n20437_, new_n20436_, new_n20431_ );
nand ( new_n20438_, new_n20151_, new_n138_ );
and  ( new_n20439_, new_n20438_, RI2b1c4342c400_29 );
nand ( new_n20440_, new_n20153_, new_n138_ );
and  ( new_n20441_, new_n20440_, RI2b1c4342c388_28 );
and  ( new_n20442_, new_n20441_, new_n20439_ );
or   ( new_n20443_, new_n20442_, new_n19390_ );
or   ( new_n20444_, new_n20163_, new_n19394_ );
or   ( new_n20445_, new_n20159_, new_n19659_ );
and  ( new_n20446_, new_n20445_, new_n20444_ );
or   ( new_n20447_, new_n20446_, new_n20443_ );
and  ( new_n20448_, new_n20446_, new_n20443_ );
or   ( new_n20449_, new_n20174_, new_n18742_ );
or   ( new_n20450_, new_n20170_, new_n18977_ );
and  ( new_n20451_, new_n20450_, new_n20449_ );
or   ( new_n20452_, new_n20451_, new_n20448_ );
and  ( new_n20453_, new_n20452_, new_n20447_ );
or   ( new_n20454_, new_n20453_, new_n20437_ );
and  ( new_n20455_, new_n20453_, new_n20437_ );
or   ( new_n20456_, new_n20218_, new_n16505_ );
or   ( new_n20457_, new_n20214_, new_n16438_ );
and  ( new_n20458_, new_n20457_, new_n20456_ );
or   ( new_n20459_, new_n20227_, new_n16085_ );
or   ( new_n20460_, new_n20223_, new_n16048_ );
and  ( new_n20461_, new_n20460_, new_n20459_ );
or   ( new_n20462_, new_n20461_, new_n20458_ );
and  ( new_n20463_, new_n20461_, new_n20458_ );
or   ( new_n20464_, new_n20238_, new_n16052_ );
or   ( new_n20465_, new_n20234_, new_n16071_ );
and  ( new_n20466_, new_n20465_, new_n20464_ );
or   ( new_n20467_, new_n20466_, new_n20463_ );
and  ( new_n20468_, new_n20467_, new_n20462_ );
or   ( new_n20469_, new_n20468_, new_n20455_ );
and  ( new_n20470_, new_n20469_, new_n20454_ );
or   ( new_n20471_, new_n20470_, new_n20424_ );
and  ( new_n20472_, new_n20470_, new_n20424_ );
or   ( new_n20473_, new_n20311_, new_n20065_ );
or   ( new_n20474_, new_n20309_, new_n19898_ );
and  ( new_n20475_, new_n20474_, new_n20473_ );
or   ( new_n20476_, new_n20318_, new_n20045_ );
or   ( new_n20477_, new_n20316_, new_n19854_ );
and  ( new_n20478_, new_n20477_, new_n20476_ );
or   ( new_n20479_, new_n20478_, new_n20475_ );
and  ( new_n20480_, new_n20478_, new_n20475_ );
or   ( new_n20481_, new_n20327_, new_n20030_ );
or   ( new_n20482_, new_n20325_, new_n19821_ );
and  ( new_n20483_, new_n20482_, new_n20481_ );
or   ( new_n20484_, new_n20483_, new_n20480_ );
and  ( new_n20485_, new_n20484_, new_n20479_ );
or   ( new_n20486_, new_n20485_, new_n20472_ );
and  ( new_n20487_, new_n20486_, new_n20471_ );
or   ( new_n20488_, new_n20487_, new_n20393_ );
and  ( new_n20489_, new_n20487_, new_n20393_ );
or   ( new_n20490_, new_n20340_, new_n20100_ );
or   ( new_n20491_, new_n20338_, new_n19959_ );
and  ( new_n20492_, new_n20491_, new_n20490_ );
or   ( new_n20493_, new_n20492_, new_n20489_ );
and  ( new_n20494_, new_n20493_, new_n20488_ );
or   ( new_n20495_, new_n20494_, new_n20347_ );
and  ( new_n20496_, new_n20495_, new_n20380_ );
or   ( new_n20497_, new_n20496_, new_n20377_ );
or   ( new_n20498_, new_n20494_, new_n20379_ );
and  ( new_n20499_, new_n20498_, new_n20349_ );
or   ( new_n20500_, new_n20499_, new_n20356_ );
and  ( new_n20501_, new_n20500_, new_n20497_ );
or   ( new_n20502_, new_n20032_, new_n19792_ );
or   ( new_n20503_, new_n20019_, new_n19823_ );
and  ( new_n20504_, new_n20503_, new_n20502_ );
or   ( new_n20505_, new_n20504_, new_n20047_ );
and  ( new_n20506_, new_n20033_, new_n19824_ );
or   ( new_n20507_, new_n20506_, new_n19856_ );
and  ( new_n20508_, new_n20507_, new_n20505_ );
or   ( new_n20509_, new_n20386_, new_n20132_ );
or   ( new_n20510_, new_n20383_, new_n20139_ );
and  ( new_n20511_, new_n20510_, new_n20509_ );
or   ( new_n20512_, new_n20511_, new_n20391_ );
and  ( new_n20513_, new_n20387_, new_n20140_ );
or   ( new_n20514_, new_n20513_, new_n20148_ );
and  ( new_n20515_, new_n20514_, new_n20512_ );
or   ( new_n20516_, new_n20515_, new_n20508_ );
and  ( new_n20517_, new_n20515_, new_n20508_ );
or   ( new_n20518_, new_n20424_, new_n20244_ );
or   ( new_n20519_, new_n20470_, new_n20304_ );
and  ( new_n20520_, new_n20519_, new_n20518_ );
or   ( new_n20521_, new_n20520_, new_n20485_ );
and  ( new_n20522_, new_n20471_, new_n20306_ );
or   ( new_n20523_, new_n20522_, new_n20331_ );
and  ( new_n20524_, new_n20523_, new_n20521_ );
or   ( new_n20525_, new_n20524_, new_n20517_ );
and  ( new_n20526_, new_n20525_, new_n20516_ );
or   ( new_n20527_, new_n20012_, new_n19770_ );
or   ( new_n20528_, new_n20009_, new_n19779_ );
and  ( new_n20529_, new_n20528_, new_n20527_ );
or   ( new_n20530_, new_n20529_, new_n20017_ );
and  ( new_n20531_, new_n20013_, new_n19780_ );
or   ( new_n20532_, new_n20531_, new_n19790_ );
and  ( new_n20533_, new_n20532_, new_n20530_ );
or   ( new_n20534_, new_n20478_, new_n20313_ );
or   ( new_n20535_, new_n20475_, new_n20320_ );
and  ( new_n20536_, new_n20535_, new_n20534_ );
or   ( new_n20537_, new_n20536_, new_n20483_ );
and  ( new_n20538_, new_n20479_, new_n20321_ );
or   ( new_n20539_, new_n20538_, new_n20329_ );
and  ( new_n20540_, new_n20539_, new_n20537_ );
or   ( new_n20541_, new_n20540_, new_n20533_ );
and  ( new_n20542_, new_n20540_, new_n20533_ );
or   ( new_n20543_, new_n20417_, new_n20275_ );
or   ( new_n20544_, new_n20406_, new_n20298_ );
and  ( new_n20545_, new_n20544_, new_n20543_ );
or   ( new_n20546_, new_n20545_, new_n20422_ );
and  ( new_n20547_, new_n20418_, new_n20300_ );
or   ( new_n20548_, new_n20547_, new_n20302_ );
and  ( new_n20549_, new_n20548_, new_n20546_ );
or   ( new_n20550_, new_n20549_, new_n20542_ );
and  ( new_n20551_, new_n20550_, new_n20541_ );
or   ( new_n20552_, new_n20441_, new_n20439_ );
and  ( new_n20553_, new_n20552_, new_n20155_ );
or   ( new_n20554_, new_n20441_, new_n19390_ );
or   ( new_n20555_, new_n20154_, new_n19655_ );
and  ( new_n20556_, new_n20555_, new_n20554_ );
or   ( new_n20557_, new_n20556_, new_n20553_ );
or   ( new_n20558_, new_n20557_, new_n99_ );
or   ( new_n20559_, new_n20558_, new_n20156_ );
or   ( new_n20560_, new_n20439_, new_n20154_ );
or   ( new_n20561_, new_n20441_, new_n20152_ );
and  ( new_n20562_, new_n20561_, new_n20560_ );
or   ( new_n20563_, new_n20154_, new_n19390_ );
or   ( new_n20564_, new_n20441_, new_n19655_ );
and  ( new_n20565_, new_n20564_, new_n20563_ );
and  ( new_n20566_, new_n20565_, new_n20562_ );
and  ( new_n20567_, new_n20566_, RI2b1c4342d4e0_65 );
or   ( new_n20568_, new_n20567_, new_n20443_ );
and  ( new_n20569_, new_n20568_, new_n20559_ );
or   ( new_n20570_, new_n19758_, new_n112_ );
or   ( new_n20571_, new_n19763_, new_n526_ );
and  ( new_n20572_, new_n20571_, new_n20570_ );
or   ( new_n20573_, new_n20572_, new_n19394_ );
and  ( new_n20574_, new_n19767_, RI2b1c4342d5d0_67 );
and  ( new_n20575_, new_n19754_, RI2b1c4342d558_66 );
or   ( new_n20576_, new_n20575_, new_n20574_ );
or   ( new_n20577_, new_n20576_, new_n19659_ );
and  ( new_n20578_, new_n20577_, new_n20573_ );
or   ( new_n20579_, new_n20578_, new_n20569_ );
and  ( new_n20580_, new_n20578_, new_n20569_ );
or   ( new_n20581_, new_n19048_, new_n591_ );
or   ( new_n20582_, new_n19055_, new_n612_ );
and  ( new_n20583_, new_n20582_, new_n20581_ );
or   ( new_n20584_, new_n20583_, new_n18742_ );
and  ( new_n20585_, new_n19057_, RI2b1c4342d6c0_69 );
and  ( new_n20586_, new_n19044_, RI2b1c4342d648_68 );
or   ( new_n20587_, new_n20586_, new_n20585_ );
or   ( new_n20588_, new_n20587_, new_n18977_ );
and  ( new_n20589_, new_n20588_, new_n20584_ );
or   ( new_n20590_, new_n20589_, new_n20580_ );
and  ( new_n20591_, new_n20590_, new_n20579_ );
or   ( new_n20592_, new_n18388_, new_n110_ );
or   ( new_n20593_, new_n18395_, new_n755_ );
and  ( new_n20594_, new_n20593_, new_n20592_ );
or   ( new_n20595_, new_n20594_, new_n18066_ );
and  ( new_n20596_, new_n18397_, RI2b1c4342d7b0_71 );
and  ( new_n20597_, new_n18384_, RI2b1c4342d738_70 );
or   ( new_n20598_, new_n20597_, new_n20596_ );
or   ( new_n20599_, new_n20598_, new_n18309_ );
and  ( new_n20600_, new_n20599_, new_n20595_ );
or   ( new_n20601_, new_n17727_, new_n105_ );
or   ( new_n20602_, new_n17734_, new_n806_ );
and  ( new_n20603_, new_n20602_, new_n20601_ );
or   ( new_n20604_, new_n20603_, new_n17238_ );
and  ( new_n20605_, new_n17736_, RI2b1c4342d8a0_73 );
and  ( new_n20606_, new_n17723_, RI2b1c4342d828_72 );
or   ( new_n20607_, new_n20606_, new_n20605_ );
or   ( new_n20608_, new_n20607_, new_n17650_ );
and  ( new_n20609_, new_n20608_, new_n20604_ );
or   ( new_n20610_, new_n20609_, new_n20600_ );
and  ( new_n20611_, new_n20609_, new_n20600_ );
or   ( new_n20612_, new_n17244_, new_n843_ );
or   ( new_n20613_, new_n17248_, new_n859_ );
and  ( new_n20614_, new_n20613_, new_n20612_ );
or   ( new_n20615_, new_n20614_, new_n16814_ );
and  ( new_n20616_, new_n17255_, RI2b1c4342d990_75 );
and  ( new_n20617_, new_n17240_, RI2b1c4342d918_74 );
or   ( new_n20618_, new_n20617_, new_n20616_ );
or   ( new_n20619_, new_n20618_, new_n17142_ );
and  ( new_n20620_, new_n20619_, new_n20615_ );
or   ( new_n20621_, new_n20620_, new_n20611_ );
and  ( new_n20622_, new_n20621_, new_n20610_ );
or   ( new_n20623_, new_n20622_, new_n20591_ );
and  ( new_n20624_, new_n20622_, new_n20591_ );
or   ( new_n20625_, new_n16607_, new_n1004_ );
or   ( new_n20626_, new_n16613_, new_n886_ );
and  ( new_n20627_, new_n20626_, new_n20625_ );
or   ( new_n20628_, new_n20627_, new_n16505_ );
and  ( new_n20629_, new_n16616_, RI2b1c4342da80_77 );
and  ( new_n20630_, new_n16603_, RI2b1c4342da08_76 );
or   ( new_n20631_, new_n20630_, new_n20629_ );
or   ( new_n20632_, new_n20631_, new_n16438_ );
and  ( new_n20633_, new_n20632_, new_n20628_ );
or   ( new_n20634_, new_n16366_, new_n1310_ );
or   ( new_n20635_, new_n16355_, new_n1002_ );
and  ( new_n20636_, new_n20635_, new_n20634_ );
or   ( new_n20637_, new_n20636_, new_n16085_ );
and  ( new_n20638_, new_n16358_, RI2b1c4342db70_79 );
and  ( new_n20639_, new_n16362_, RI2b1c4342daf8_78 );
or   ( new_n20640_, new_n20639_, new_n20638_ );
or   ( new_n20641_, new_n20640_, new_n16048_ );
and  ( new_n20642_, new_n20641_, new_n20637_ );
or   ( new_n20643_, new_n20642_, new_n20633_ );
and  ( new_n20644_, new_n20642_, new_n20633_ );
or   ( new_n20645_, new_n16075_, new_n126_ );
or   ( new_n20646_, new_n16060_, new_n1511_ );
and  ( new_n20647_, new_n20646_, new_n20645_ );
or   ( new_n20648_, new_n20647_, new_n16052_ );
and  ( new_n20649_, new_n16063_, RI2b1c4342dc60_81 );
and  ( new_n20650_, new_n16066_, RI2b1c4342dbe8_80 );
or   ( new_n20651_, new_n20650_, new_n20649_ );
or   ( new_n20652_, new_n20651_, new_n16071_ );
and  ( new_n20653_, new_n20652_, new_n20648_ );
or   ( new_n20654_, new_n20653_, new_n20644_ );
and  ( new_n20655_, new_n20654_, new_n20643_ );
or   ( new_n20656_, new_n20655_, new_n20624_ );
and  ( new_n20657_, new_n20656_, new_n20623_ );
or   ( new_n20658_, new_n16033_, new_n121_ );
or   ( new_n20659_, new_n16017_, new_n2119_ );
and  ( new_n20660_, new_n20659_, new_n20658_ );
or   ( new_n20661_, new_n20660_, new_n16009_ );
and  ( new_n20662_, new_n16021_, RI2b1c4342dd50_83 );
and  ( new_n20663_, new_n16024_, RI2b1c4342dcd8_82 );
or   ( new_n20664_, new_n20663_, new_n20662_ );
or   ( new_n20665_, new_n20664_, new_n16029_ );
and  ( new_n20666_, new_n20665_, new_n20661_ );
or   ( new_n20667_, new_n16208_, new_n2806_ );
or   ( new_n20668_, new_n16194_, new_n2541_ );
and  ( new_n20669_, new_n20668_, new_n20667_ );
or   ( new_n20670_, new_n20669_, new_n16186_ );
and  ( new_n20671_, new_n16196_, RI2b1c4342de40_85 );
and  ( new_n20672_, new_n16199_, RI2b1c4342ddc8_84 );
or   ( new_n20673_, new_n20672_, new_n20671_ );
or   ( new_n20674_, new_n20673_, new_n16204_ );
and  ( new_n20675_, new_n20674_, new_n20670_ );
or   ( new_n20676_, new_n20675_, new_n20666_ );
and  ( new_n20677_, new_n20675_, new_n20666_ );
or   ( new_n20678_, new_n16238_, new_n3924_ );
or   ( new_n20679_, new_n16224_, new_n3239_ );
and  ( new_n20680_, new_n20679_, new_n20678_ );
or   ( new_n20681_, new_n20680_, new_n16217_ );
and  ( new_n20682_, new_n16226_, RI2b1c4342df30_87 );
and  ( new_n20683_, new_n16229_, RI2b1c4342deb8_86 );
or   ( new_n20684_, new_n20683_, new_n20682_ );
or   ( new_n20685_, new_n20684_, new_n16234_ );
and  ( new_n20686_, new_n20685_, new_n20681_ );
or   ( new_n20687_, new_n20686_, new_n20677_ );
and  ( new_n20688_, new_n20687_, new_n20676_ );
or   ( new_n20689_, new_n16174_, new_n132_ );
or   ( new_n20690_, new_n16160_, new_n3902_ );
and  ( new_n20691_, new_n20690_, new_n20689_ );
or   ( new_n20692_, new_n20691_, new_n16151_ );
and  ( new_n20693_, new_n16162_, RI2b1c4342e020_89 );
and  ( new_n20694_, new_n16165_, RI2b1c4342dfa8_88 );
or   ( new_n20695_, new_n20694_, new_n20693_ );
or   ( new_n20696_, new_n20695_, new_n16170_ );
and  ( new_n20697_, new_n20696_, new_n20692_ );
or   ( new_n20698_, new_n16119_, new_n117_ );
or   ( new_n20699_, new_n16123_, new_n4635_ );
and  ( new_n20700_, new_n20699_, new_n20698_ );
or   ( new_n20701_, new_n20700_, new_n16108_ );
and  ( new_n20702_, new_n16132_, RI2b1c4342e110_91 );
and  ( new_n20703_, new_n16114_, RI2b1c4342e098_90 );
or   ( new_n20704_, new_n20703_, new_n20702_ );
or   ( new_n20705_, new_n20704_, new_n16128_ );
and  ( new_n20706_, new_n20705_, new_n20701_ );
and  ( new_n20707_, new_n20706_, new_n20697_ );
or   ( new_n20708_, new_n20706_, new_n20697_ );
or   ( new_n20709_, new_n16115_, new_n5459_ );
and  ( new_n20710_, new_n20709_, new_n20708_ );
or   ( new_n20711_, new_n20710_, new_n20707_ );
and  ( new_n20712_, new_n20711_, new_n20688_ );
or   ( new_n20713_, new_n20711_, new_n20688_ );
or   ( new_n20714_, new_n20412_, new_n20284_ );
or   ( new_n20715_, new_n20409_, new_n20293_ );
and  ( new_n20716_, new_n20715_, new_n20714_ );
or   ( new_n20717_, new_n20716_, new_n20415_ );
and  ( new_n20718_, new_n20413_, new_n20295_ );
or   ( new_n20719_, new_n20718_, new_n20296_ );
and  ( new_n20720_, new_n20719_, new_n20717_ );
and  ( new_n20721_, new_n20720_, new_n20713_ );
or   ( new_n20722_, new_n20721_, new_n20712_ );
and  ( new_n20723_, new_n20722_, new_n20657_ );
or   ( new_n20724_, new_n20722_, new_n20657_ );
or   ( new_n20725_, new_n20399_, new_n20253_ );
or   ( new_n20726_, new_n20396_, new_n20262_ );
and  ( new_n20727_, new_n20726_, new_n20725_ );
or   ( new_n20728_, new_n20727_, new_n20404_ );
and  ( new_n20729_, new_n20400_, new_n20263_ );
or   ( new_n20730_, new_n20729_, new_n20273_ );
and  ( new_n20731_, new_n20730_, new_n20728_ );
or   ( new_n20732_, new_n20461_, new_n20220_ );
or   ( new_n20733_, new_n20458_, new_n20229_ );
and  ( new_n20734_, new_n20733_, new_n20732_ );
or   ( new_n20735_, new_n20734_, new_n20466_ );
and  ( new_n20736_, new_n20462_, new_n20230_ );
or   ( new_n20737_, new_n20736_, new_n20240_ );
and  ( new_n20738_, new_n20737_, new_n20735_ );
or   ( new_n20739_, new_n20738_, new_n20731_ );
and  ( new_n20740_, new_n20738_, new_n20731_ );
or   ( new_n20741_, new_n20430_, new_n20187_ );
or   ( new_n20742_, new_n20427_, new_n20196_ );
and  ( new_n20743_, new_n20742_, new_n20741_ );
or   ( new_n20744_, new_n20743_, new_n20435_ );
and  ( new_n20745_, new_n20431_, new_n20197_ );
or   ( new_n20746_, new_n20745_, new_n20207_ );
and  ( new_n20747_, new_n20746_, new_n20744_ );
or   ( new_n20748_, new_n20747_, new_n20740_ );
and  ( new_n20749_, new_n20748_, new_n20739_ );
and  ( new_n20750_, new_n20749_, new_n20724_ );
or   ( new_n20751_, new_n20750_, new_n20723_ );
and  ( new_n20752_, new_n20751_, new_n20551_ );
or   ( new_n20753_, new_n20751_, new_n20551_ );
or   ( new_n20754_, new_n20054_, new_n19900_ );
or   ( new_n20755_, new_n20067_, new_n19869_ );
and  ( new_n20756_, new_n20755_, new_n20754_ );
or   ( new_n20757_, new_n20756_, new_n20072_ );
and  ( new_n20758_, new_n20068_, new_n19901_ );
or   ( new_n20759_, new_n20758_, new_n19911_ );
and  ( new_n20760_, new_n20759_, new_n20757_ );
and  ( new_n20761_, new_n20760_, new_n20753_ );
or   ( new_n20762_, new_n20761_, new_n20752_ );
and  ( new_n20763_, new_n20762_, new_n20526_ );
or   ( new_n20764_, new_n20762_, new_n20526_ );
or   ( new_n20765_, new_n20074_, new_n19858_ );
or   ( new_n20766_, new_n20049_, new_n19913_ );
and  ( new_n20767_, new_n20766_, new_n20765_ );
or   ( new_n20768_, new_n20767_, new_n20087_ );
and  ( new_n20769_, new_n20075_, new_n19914_ );
or   ( new_n20770_, new_n20769_, new_n19934_ );
and  ( new_n20771_, new_n20770_, new_n20768_ );
and  ( new_n20772_, new_n20771_, new_n20764_ );
or   ( new_n20773_, new_n20772_, new_n20763_ );
or   ( new_n20774_, new_n20773_, new_n20501_ );
or   ( new_n20775_, new_n20365_, new_n20114_ );
or   ( new_n20776_, new_n20363_, new_n19981_ );
and  ( new_n20777_, new_n20776_, new_n20775_ );
or   ( new_n20778_, new_n20123_, new_n19728_ );
or   ( new_n20779_, new_n20121_, new_n19587_ );
and  ( new_n20780_, new_n20779_, new_n20778_ );
or   ( new_n20781_, new_n20780_, new_n20358_ );
and  ( new_n20782_, new_n20494_, new_n20379_ );
or   ( new_n20783_, new_n20782_, new_n20377_ );
and  ( new_n20784_, new_n20783_, new_n20498_ );
or   ( new_n20785_, new_n20784_, new_n20125_ );
and  ( new_n20786_, new_n20785_, new_n20781_ );
or   ( new_n20787_, new_n20786_, new_n20777_ );
or   ( new_n20788_, new_n20784_, new_n20780_ );
and  ( new_n20789_, new_n20788_, new_n20360_ );
or   ( new_n20790_, new_n20789_, new_n20367_ );
and  ( new_n20791_, new_n20790_, new_n20787_ );
or   ( new_n20792_, new_n20791_, new_n20774_ );
and  ( new_n20793_, new_n20791_, new_n20774_ );
or   ( new_n20794_, new_n20499_, new_n20377_ );
or   ( new_n20795_, new_n20496_, new_n20356_ );
and  ( new_n20796_, new_n20795_, new_n20794_ );
or   ( new_n20797_, new_n20796_, new_n20773_ );
or   ( new_n20798_, new_n20567_, new_n20156_ );
or   ( new_n20799_, new_n20558_, new_n20443_ );
and  ( new_n20800_, new_n20799_, new_n20798_ );
or   ( new_n20801_, new_n20576_, new_n19394_ );
or   ( new_n20802_, new_n20572_, new_n19659_ );
and  ( new_n20803_, new_n20802_, new_n20801_ );
or   ( new_n20804_, new_n20803_, new_n20800_ );
and  ( new_n20805_, new_n20803_, new_n20800_ );
or   ( new_n20806_, new_n20587_, new_n18742_ );
or   ( new_n20807_, new_n20583_, new_n18977_ );
and  ( new_n20808_, new_n20807_, new_n20806_ );
or   ( new_n20809_, new_n20808_, new_n20805_ );
and  ( new_n20810_, new_n20809_, new_n20804_ );
or   ( new_n20811_, new_n20598_, new_n18066_ );
or   ( new_n20812_, new_n20594_, new_n18309_ );
and  ( new_n20813_, new_n20812_, new_n20811_ );
or   ( new_n20814_, new_n20607_, new_n17238_ );
or   ( new_n20815_, new_n20603_, new_n17650_ );
and  ( new_n20816_, new_n20815_, new_n20814_ );
or   ( new_n20817_, new_n20816_, new_n20813_ );
and  ( new_n20818_, new_n20816_, new_n20813_ );
or   ( new_n20819_, new_n20618_, new_n16814_ );
or   ( new_n20820_, new_n20614_, new_n17142_ );
and  ( new_n20821_, new_n20820_, new_n20819_ );
or   ( new_n20822_, new_n20821_, new_n20818_ );
and  ( new_n20823_, new_n20822_, new_n20817_ );
or   ( new_n20824_, new_n20823_, new_n20810_ );
and  ( new_n20825_, new_n20823_, new_n20810_ );
or   ( new_n20826_, new_n20631_, new_n16505_ );
or   ( new_n20827_, new_n20627_, new_n16438_ );
and  ( new_n20828_, new_n20827_, new_n20826_ );
or   ( new_n20829_, new_n20640_, new_n16085_ );
or   ( new_n20830_, new_n20636_, new_n16048_ );
and  ( new_n20831_, new_n20830_, new_n20829_ );
or   ( new_n20832_, new_n20831_, new_n20828_ );
and  ( new_n20833_, new_n20831_, new_n20828_ );
or   ( new_n20834_, new_n20651_, new_n16052_ );
or   ( new_n20835_, new_n20647_, new_n16071_ );
and  ( new_n20836_, new_n20835_, new_n20834_ );
or   ( new_n20837_, new_n20836_, new_n20833_ );
and  ( new_n20838_, new_n20837_, new_n20832_ );
or   ( new_n20839_, new_n20838_, new_n20825_ );
and  ( new_n20840_, new_n20839_, new_n20824_ );
or   ( new_n20841_, new_n20664_, new_n16009_ );
or   ( new_n20842_, new_n20660_, new_n16029_ );
and  ( new_n20843_, new_n20842_, new_n20841_ );
or   ( new_n20844_, new_n20673_, new_n16186_ );
or   ( new_n20845_, new_n20669_, new_n16204_ );
and  ( new_n20846_, new_n20845_, new_n20844_ );
or   ( new_n20847_, new_n20846_, new_n20843_ );
and  ( new_n20848_, new_n20846_, new_n20843_ );
or   ( new_n20849_, new_n20684_, new_n16217_ );
or   ( new_n20850_, new_n20680_, new_n16234_ );
and  ( new_n20851_, new_n20850_, new_n20849_ );
or   ( new_n20852_, new_n20851_, new_n20848_ );
and  ( new_n20853_, new_n20852_, new_n20847_ );
or   ( new_n20854_, new_n20695_, new_n16151_ );
or   ( new_n20855_, new_n20691_, new_n16170_ );
and  ( new_n20856_, new_n20855_, new_n20854_ );
or   ( new_n20857_, new_n20704_, new_n16108_ );
or   ( new_n20858_, new_n20700_, new_n16128_ );
and  ( new_n20859_, new_n20858_, new_n20857_ );
or   ( new_n20860_, new_n20859_, new_n20856_ );
and  ( new_n20861_, new_n20859_, new_n20856_ );
and  ( new_n20862_, new_n16102_, RI2b1c4342e188_92 );
or   ( new_n20863_, new_n20862_, new_n20861_ );
and  ( new_n20864_, new_n20863_, new_n20860_ );
or   ( new_n20865_, new_n20864_, new_n20853_ );
and  ( new_n20866_, new_n20864_, new_n20853_ );
or   ( new_n20867_, new_n20718_, new_n20415_ );
or   ( new_n20868_, new_n20716_, new_n20296_ );
and  ( new_n20869_, new_n20868_, new_n20867_ );
or   ( new_n20870_, new_n20869_, new_n20866_ );
and  ( new_n20871_, new_n20870_, new_n20865_ );
or   ( new_n20872_, new_n20871_, new_n20840_ );
and  ( new_n20873_, new_n20871_, new_n20840_ );
or   ( new_n20874_, new_n20729_, new_n20404_ );
or   ( new_n20875_, new_n20727_, new_n20273_ );
and  ( new_n20876_, new_n20875_, new_n20874_ );
or   ( new_n20877_, new_n20736_, new_n20466_ );
or   ( new_n20878_, new_n20734_, new_n20240_ );
and  ( new_n20879_, new_n20878_, new_n20877_ );
or   ( new_n20880_, new_n20879_, new_n20876_ );
and  ( new_n20881_, new_n20879_, new_n20876_ );
or   ( new_n20882_, new_n20745_, new_n20435_ );
or   ( new_n20883_, new_n20743_, new_n20207_ );
and  ( new_n20884_, new_n20883_, new_n20882_ );
or   ( new_n20885_, new_n20884_, new_n20881_ );
and  ( new_n20886_, new_n20885_, new_n20880_ );
or   ( new_n20887_, new_n20886_, new_n20873_ );
and  ( new_n20888_, new_n20887_, new_n20872_ );
or   ( new_n20889_, new_n20531_, new_n20017_ );
or   ( new_n20890_, new_n20529_, new_n19790_ );
and  ( new_n20891_, new_n20890_, new_n20889_ );
or   ( new_n20892_, new_n20538_, new_n20483_ );
or   ( new_n20893_, new_n20536_, new_n20329_ );
and  ( new_n20894_, new_n20893_, new_n20892_ );
or   ( new_n20895_, new_n20894_, new_n20891_ );
and  ( new_n20896_, new_n20894_, new_n20891_ );
or   ( new_n20897_, new_n20547_, new_n20422_ );
or   ( new_n20898_, new_n20545_, new_n20302_ );
and  ( new_n20899_, new_n20898_, new_n20897_ );
or   ( new_n20900_, new_n20899_, new_n20896_ );
and  ( new_n20901_, new_n20900_, new_n20895_ );
or   ( new_n20902_, new_n20901_, new_n20888_ );
and  ( new_n20903_, new_n20901_, new_n20888_ );
or   ( new_n20904_, new_n20758_, new_n20072_ );
or   ( new_n20905_, new_n20756_, new_n19911_ );
and  ( new_n20906_, new_n20905_, new_n20904_ );
or   ( new_n20907_, new_n20906_, new_n20903_ );
and  ( new_n20908_, new_n20907_, new_n20902_ );
or   ( new_n20909_, new_n20506_, new_n20047_ );
or   ( new_n20910_, new_n20504_, new_n19856_ );
and  ( new_n20911_, new_n20910_, new_n20909_ );
or   ( new_n20912_, new_n20513_, new_n20391_ );
or   ( new_n20913_, new_n20511_, new_n20148_ );
and  ( new_n20914_, new_n20913_, new_n20912_ );
or   ( new_n20915_, new_n20914_, new_n20911_ );
and  ( new_n20916_, new_n20914_, new_n20911_ );
or   ( new_n20917_, new_n20522_, new_n20485_ );
or   ( new_n20918_, new_n20520_, new_n20331_ );
and  ( new_n20919_, new_n20918_, new_n20917_ );
or   ( new_n20920_, new_n20919_, new_n20916_ );
and  ( new_n20921_, new_n20920_, new_n20915_ );
or   ( new_n20922_, new_n20921_, new_n20908_ );
and  ( new_n20923_, new_n20921_, new_n20908_ );
or   ( new_n20924_, new_n20769_, new_n20087_ );
or   ( new_n20925_, new_n20767_, new_n19934_ );
and  ( new_n20926_, new_n20925_, new_n20924_ );
or   ( new_n20927_, new_n20926_, new_n20923_ );
and  ( new_n20928_, new_n20927_, new_n20922_ );
or   ( new_n20929_, new_n20928_, new_n20501_ );
and  ( new_n20930_, new_n20929_, new_n20797_ );
or   ( new_n20931_, new_n20393_, new_n20333_ );
or   ( new_n20932_, new_n20487_, new_n20150_ );
and  ( new_n20933_, new_n20932_, new_n20931_ );
or   ( new_n20934_, new_n20933_, new_n20492_ );
and  ( new_n20935_, new_n20488_, new_n20335_ );
or   ( new_n20936_, new_n20935_, new_n20342_ );
and  ( new_n20937_, new_n20936_, new_n20934_ );
or   ( new_n20938_, new_n20914_, new_n20508_ );
or   ( new_n20939_, new_n20911_, new_n20515_ );
and  ( new_n20940_, new_n20939_, new_n20938_ );
or   ( new_n20941_, new_n20940_, new_n20919_ );
and  ( new_n20942_, new_n20915_, new_n20516_ );
or   ( new_n20943_, new_n20942_, new_n20524_ );
and  ( new_n20944_, new_n20943_, new_n20941_ );
or   ( new_n20945_, new_n16075_, new_n2119_ );
or   ( new_n20946_, new_n16060_, new_n126_ );
and  ( new_n20947_, new_n20946_, new_n20945_ );
or   ( new_n20948_, new_n20947_, new_n16052_ );
and  ( new_n20949_, new_n16063_, RI2b1c4342dcd8_82 );
and  ( new_n20950_, new_n16066_, RI2b1c4342dc60_81 );
or   ( new_n20951_, new_n20950_, new_n20949_ );
or   ( new_n20952_, new_n20951_, new_n16071_ );
and  ( new_n20953_, new_n20952_, new_n20948_ );
or   ( new_n20954_, new_n16033_, new_n2541_ );
or   ( new_n20955_, new_n16017_, new_n121_ );
and  ( new_n20956_, new_n20955_, new_n20954_ );
or   ( new_n20957_, new_n20956_, new_n16009_ );
and  ( new_n20958_, new_n16021_, RI2b1c4342ddc8_84 );
and  ( new_n20959_, new_n16024_, RI2b1c4342dd50_83 );
or   ( new_n20960_, new_n20959_, new_n20958_ );
or   ( new_n20961_, new_n20960_, new_n16029_ );
and  ( new_n20962_, new_n20961_, new_n20957_ );
or   ( new_n20963_, new_n20962_, new_n20953_ );
and  ( new_n20964_, new_n20962_, new_n20953_ );
or   ( new_n20965_, new_n16208_, new_n3239_ );
or   ( new_n20966_, new_n16194_, new_n2806_ );
and  ( new_n20967_, new_n20966_, new_n20965_ );
or   ( new_n20968_, new_n20967_, new_n16186_ );
and  ( new_n20969_, new_n16196_, RI2b1c4342deb8_86 );
and  ( new_n20970_, new_n16199_, RI2b1c4342de40_85 );
or   ( new_n20971_, new_n20970_, new_n20969_ );
or   ( new_n20972_, new_n20971_, new_n16204_ );
and  ( new_n20973_, new_n20972_, new_n20968_ );
or   ( new_n20974_, new_n20973_, new_n20964_ );
and  ( new_n20975_, new_n20974_, new_n20963_ );
or   ( new_n20976_, new_n16238_, new_n3902_ );
or   ( new_n20977_, new_n16224_, new_n3924_ );
and  ( new_n20978_, new_n20977_, new_n20976_ );
or   ( new_n20979_, new_n20978_, new_n16217_ );
and  ( new_n20980_, new_n16226_, RI2b1c4342dfa8_88 );
and  ( new_n20981_, new_n16229_, RI2b1c4342df30_87 );
or   ( new_n20982_, new_n20981_, new_n20980_ );
or   ( new_n20983_, new_n20982_, new_n16234_ );
and  ( new_n20984_, new_n20983_, new_n20979_ );
or   ( new_n20985_, new_n16174_, new_n4635_ );
or   ( new_n20986_, new_n16160_, new_n132_ );
and  ( new_n20987_, new_n20986_, new_n20985_ );
or   ( new_n20988_, new_n20987_, new_n16151_ );
and  ( new_n20989_, new_n16162_, RI2b1c4342e098_90 );
and  ( new_n20990_, new_n16165_, RI2b1c4342e020_89 );
or   ( new_n20991_, new_n20990_, new_n20989_ );
or   ( new_n20992_, new_n20991_, new_n16170_ );
and  ( new_n20993_, new_n20992_, new_n20988_ );
or   ( new_n20994_, new_n20993_, new_n20984_ );
and  ( new_n20995_, new_n20993_, new_n20984_ );
or   ( new_n20996_, new_n16119_, new_n5459_ );
or   ( new_n20997_, new_n16123_, new_n117_ );
and  ( new_n20998_, new_n20997_, new_n20996_ );
or   ( new_n20999_, new_n20998_, new_n16108_ );
and  ( new_n21000_, new_n16132_, RI2b1c4342e188_92 );
and  ( new_n21001_, new_n16114_, RI2b1c4342e110_91 );
or   ( new_n21002_, new_n21001_, new_n21000_ );
or   ( new_n21003_, new_n21002_, new_n16128_ );
and  ( new_n21004_, new_n21003_, new_n20999_ );
or   ( new_n21005_, new_n21004_, new_n20995_ );
and  ( new_n21006_, new_n21005_, new_n20994_ );
and  ( new_n21007_, new_n21006_, new_n20975_ );
xor  ( new_n21008_, new_n6033_, new_n214_ );
or   ( new_n21009_, new_n21008_, new_n336_ );
xor  ( new_n21010_, new_n5861_, new_n6028_ );
or   ( new_n21011_, new_n21010_, new_n333_ );
or   ( new_n21012_, new_n21011_, new_n21009_ );
and  ( new_n21013_, new_n21012_, new_n20439_ );
or   ( new_n21014_, new_n20557_, new_n526_ );
or   ( new_n21015_, new_n20562_, new_n99_ );
and  ( new_n21016_, new_n21015_, new_n21014_ );
or   ( new_n21017_, new_n21016_, new_n20156_ );
and  ( new_n21018_, new_n20566_, RI2b1c4342d558_66 );
and  ( new_n21019_, new_n20553_, RI2b1c4342d4e0_65 );
or   ( new_n21020_, new_n21019_, new_n21018_ );
or   ( new_n21021_, new_n21020_, new_n20443_ );
and  ( new_n21022_, new_n21021_, new_n21017_ );
or   ( new_n21023_, new_n21022_, new_n21013_ );
and  ( new_n21024_, new_n21022_, new_n21013_ );
or   ( new_n21025_, new_n19758_, new_n612_ );
or   ( new_n21026_, new_n19763_, new_n112_ );
and  ( new_n21027_, new_n21026_, new_n21025_ );
or   ( new_n21028_, new_n21027_, new_n19394_ );
and  ( new_n21029_, new_n19767_, RI2b1c4342d648_68 );
and  ( new_n21030_, new_n19754_, RI2b1c4342d5d0_67 );
or   ( new_n21031_, new_n21030_, new_n21029_ );
or   ( new_n21032_, new_n21031_, new_n19659_ );
and  ( new_n21033_, new_n21032_, new_n21028_ );
or   ( new_n21034_, new_n21033_, new_n21024_ );
and  ( new_n21035_, new_n21034_, new_n21023_ );
or   ( new_n21036_, new_n19048_, new_n755_ );
or   ( new_n21037_, new_n19055_, new_n591_ );
and  ( new_n21038_, new_n21037_, new_n21036_ );
or   ( new_n21039_, new_n21038_, new_n18742_ );
and  ( new_n21040_, new_n19057_, RI2b1c4342d738_70 );
and  ( new_n21041_, new_n19044_, RI2b1c4342d6c0_69 );
or   ( new_n21042_, new_n21041_, new_n21040_ );
or   ( new_n21043_, new_n21042_, new_n18977_ );
and  ( new_n21044_, new_n21043_, new_n21039_ );
or   ( new_n21045_, new_n18388_, new_n806_ );
or   ( new_n21046_, new_n18395_, new_n110_ );
and  ( new_n21047_, new_n21046_, new_n21045_ );
or   ( new_n21048_, new_n21047_, new_n18066_ );
and  ( new_n21049_, new_n18397_, RI2b1c4342d828_72 );
and  ( new_n21050_, new_n18384_, RI2b1c4342d7b0_71 );
or   ( new_n21051_, new_n21050_, new_n21049_ );
or   ( new_n21052_, new_n21051_, new_n18309_ );
and  ( new_n21053_, new_n21052_, new_n21048_ );
or   ( new_n21054_, new_n21053_, new_n21044_ );
and  ( new_n21055_, new_n21053_, new_n21044_ );
or   ( new_n21056_, new_n17727_, new_n859_ );
or   ( new_n21057_, new_n17734_, new_n105_ );
and  ( new_n21058_, new_n21057_, new_n21056_ );
or   ( new_n21059_, new_n21058_, new_n17238_ );
and  ( new_n21060_, new_n17736_, RI2b1c4342d918_74 );
and  ( new_n21061_, new_n17723_, RI2b1c4342d8a0_73 );
or   ( new_n21062_, new_n21061_, new_n21060_ );
or   ( new_n21063_, new_n21062_, new_n17650_ );
and  ( new_n21064_, new_n21063_, new_n21059_ );
or   ( new_n21065_, new_n21064_, new_n21055_ );
and  ( new_n21066_, new_n21065_, new_n21054_ );
or   ( new_n21067_, new_n21066_, new_n21035_ );
and  ( new_n21068_, new_n21066_, new_n21035_ );
or   ( new_n21069_, new_n17244_, new_n886_ );
or   ( new_n21070_, new_n17248_, new_n843_ );
and  ( new_n21071_, new_n21070_, new_n21069_ );
or   ( new_n21072_, new_n21071_, new_n16814_ );
and  ( new_n21073_, new_n17255_, RI2b1c4342da08_76 );
and  ( new_n21074_, new_n17240_, RI2b1c4342d990_75 );
or   ( new_n21075_, new_n21074_, new_n21073_ );
or   ( new_n21076_, new_n21075_, new_n17142_ );
and  ( new_n21077_, new_n21076_, new_n21072_ );
or   ( new_n21078_, new_n16607_, new_n1002_ );
or   ( new_n21079_, new_n16613_, new_n1004_ );
and  ( new_n21080_, new_n21079_, new_n21078_ );
or   ( new_n21081_, new_n21080_, new_n16505_ );
and  ( new_n21082_, new_n16616_, RI2b1c4342daf8_78 );
and  ( new_n21083_, new_n16603_, RI2b1c4342da80_77 );
or   ( new_n21084_, new_n21083_, new_n21082_ );
or   ( new_n21085_, new_n21084_, new_n16438_ );
and  ( new_n21086_, new_n21085_, new_n21081_ );
or   ( new_n21087_, new_n21086_, new_n21077_ );
and  ( new_n21088_, new_n21086_, new_n21077_ );
or   ( new_n21089_, new_n16366_, new_n1511_ );
or   ( new_n21090_, new_n16355_, new_n1310_ );
and  ( new_n21091_, new_n21090_, new_n21089_ );
or   ( new_n21092_, new_n21091_, new_n16085_ );
and  ( new_n21093_, new_n16358_, RI2b1c4342dbe8_80 );
and  ( new_n21094_, new_n16362_, RI2b1c4342db70_79 );
or   ( new_n21095_, new_n21094_, new_n21093_ );
or   ( new_n21096_, new_n21095_, new_n16048_ );
and  ( new_n21097_, new_n21096_, new_n21092_ );
or   ( new_n21098_, new_n21097_, new_n21088_ );
and  ( new_n21099_, new_n21098_, new_n21087_ );
or   ( new_n21100_, new_n21099_, new_n21068_ );
and  ( new_n21101_, new_n21100_, new_n21067_ );
or   ( new_n21102_, new_n21101_, new_n21007_ );
and  ( new_n21103_, new_n21101_, new_n21007_ );
or   ( new_n21104_, new_n20859_, new_n20697_ );
or   ( new_n21105_, new_n20856_, new_n20706_ );
and  ( new_n21106_, new_n21105_, new_n21104_ );
or   ( new_n21107_, new_n21106_, new_n20862_ );
and  ( new_n21108_, new_n20860_, new_n20708_ );
or   ( new_n21109_, new_n21108_, new_n20709_ );
and  ( new_n21110_, new_n21109_, new_n21107_ );
or   ( new_n21111_, new_n20846_, new_n20666_ );
or   ( new_n21112_, new_n20843_, new_n20675_ );
and  ( new_n21113_, new_n21112_, new_n21111_ );
or   ( new_n21114_, new_n21113_, new_n20851_ );
and  ( new_n21115_, new_n20847_, new_n20676_ );
or   ( new_n21116_, new_n21115_, new_n20686_ );
and  ( new_n21117_, new_n21116_, new_n21114_ );
or   ( new_n21118_, new_n21117_, new_n21110_ );
and  ( new_n21119_, new_n21117_, new_n21110_ );
or   ( new_n21120_, new_n20831_, new_n20633_ );
or   ( new_n21121_, new_n20828_, new_n20642_ );
and  ( new_n21122_, new_n21121_, new_n21120_ );
or   ( new_n21123_, new_n21122_, new_n20836_ );
and  ( new_n21124_, new_n20832_, new_n20643_ );
or   ( new_n21125_, new_n21124_, new_n20653_ );
and  ( new_n21126_, new_n21125_, new_n21123_ );
or   ( new_n21127_, new_n21126_, new_n21119_ );
and  ( new_n21128_, new_n21127_, new_n21118_ );
or   ( new_n21129_, new_n21128_, new_n21103_ );
and  ( new_n21130_, new_n21129_, new_n21102_ );
or   ( new_n21131_, new_n20446_, new_n20156_ );
or   ( new_n21132_, new_n20443_, new_n20165_ );
and  ( new_n21133_, new_n21132_, new_n21131_ );
or   ( new_n21134_, new_n21133_, new_n20451_ );
and  ( new_n21135_, new_n20447_, new_n20166_ );
or   ( new_n21136_, new_n21135_, new_n20176_ );
and  ( new_n21137_, new_n21136_, new_n21134_ );
or   ( new_n21138_, new_n20879_, new_n20731_ );
or   ( new_n21139_, new_n20876_, new_n20738_ );
and  ( new_n21140_, new_n21139_, new_n21138_ );
or   ( new_n21141_, new_n21140_, new_n20884_ );
and  ( new_n21142_, new_n20880_, new_n20739_ );
or   ( new_n21143_, new_n21142_, new_n20747_ );
and  ( new_n21144_, new_n21143_, new_n21141_ );
or   ( new_n21145_, new_n21144_, new_n21137_ );
and  ( new_n21146_, new_n21144_, new_n21137_ );
or   ( new_n21147_, new_n20864_, new_n20688_ );
or   ( new_n21148_, new_n20853_, new_n20711_ );
and  ( new_n21149_, new_n21148_, new_n21147_ );
or   ( new_n21150_, new_n21149_, new_n20869_ );
and  ( new_n21151_, new_n20865_, new_n20713_ );
or   ( new_n21152_, new_n21151_, new_n20720_ );
and  ( new_n21153_, new_n21152_, new_n21150_ );
or   ( new_n21154_, new_n21153_, new_n21146_ );
and  ( new_n21155_, new_n21154_, new_n21145_ );
or   ( new_n21156_, new_n21155_, new_n21130_ );
and  ( new_n21157_, new_n21155_, new_n21130_ );
or   ( new_n21158_, new_n20437_, new_n20178_ );
or   ( new_n21159_, new_n20453_, new_n20209_ );
and  ( new_n21160_, new_n21159_, new_n21158_ );
or   ( new_n21161_, new_n21160_, new_n20468_ );
and  ( new_n21162_, new_n20454_, new_n20210_ );
or   ( new_n21163_, new_n21162_, new_n20242_ );
and  ( new_n21164_, new_n21163_, new_n21161_ );
or   ( new_n21165_, new_n21164_, new_n21157_ );
and  ( new_n21166_, new_n21165_, new_n21156_ );
or   ( new_n21167_, new_n21166_, new_n20944_ );
and  ( new_n21168_, new_n21166_, new_n20944_ );
or   ( new_n21169_, new_n20901_, new_n20751_ );
or   ( new_n21170_, new_n20888_, new_n20551_ );
and  ( new_n21171_, new_n21170_, new_n21169_ );
or   ( new_n21172_, new_n21171_, new_n20906_ );
and  ( new_n21173_, new_n20902_, new_n20753_ );
or   ( new_n21174_, new_n21173_, new_n20760_ );
and  ( new_n21175_, new_n21174_, new_n21172_ );
or   ( new_n21176_, new_n21175_, new_n21168_ );
and  ( new_n21177_, new_n21176_, new_n21167_ );
or   ( new_n21178_, new_n21177_, new_n20937_ );
or   ( new_n21179_, new_n20921_, new_n20762_ );
or   ( new_n21180_, new_n20908_, new_n20526_ );
and  ( new_n21181_, new_n21180_, new_n21179_ );
or   ( new_n21182_, new_n21181_, new_n20926_ );
and  ( new_n21183_, new_n20922_, new_n20764_ );
or   ( new_n21184_, new_n21183_, new_n20771_ );
and  ( new_n21185_, new_n21184_, new_n21182_ );
and  ( new_n21186_, new_n21177_, new_n20937_ );
or   ( new_n21187_, new_n21186_, new_n21185_ );
and  ( new_n21188_, new_n21187_, new_n21178_ );
or   ( new_n21189_, new_n21188_, new_n20930_ );
or   ( new_n21190_, new_n21189_, new_n20793_ );
and  ( new_n21191_, new_n21190_, new_n20792_ );
or   ( new_n21192_, new_n21191_, new_n20374_ );
and  ( new_n21193_, new_n21192_, new_n20372_ );
and  ( new_n21194_, new_n21188_, new_n20930_ );
or   ( new_n21195_, new_n21194_, new_n20793_ );
or   ( new_n21196_, new_n21195_, new_n20374_ );
or   ( new_n21197_, new_n21183_, new_n20926_ );
or   ( new_n21198_, new_n21181_, new_n20771_ );
and  ( new_n21199_, new_n21198_, new_n21197_ );
or   ( new_n21200_, new_n20935_, new_n20492_ );
or   ( new_n21201_, new_n20933_, new_n20342_ );
and  ( new_n21202_, new_n21201_, new_n21200_ );
or   ( new_n21203_, new_n21202_, new_n21177_ );
or   ( new_n21204_, new_n20942_, new_n20919_ );
or   ( new_n21205_, new_n20940_, new_n20524_ );
and  ( new_n21206_, new_n21205_, new_n21204_ );
or   ( new_n21207_, new_n21135_, new_n20451_ );
or   ( new_n21208_, new_n21133_, new_n20176_ );
and  ( new_n21209_, new_n21208_, new_n21207_ );
or   ( new_n21210_, new_n21142_, new_n20884_ );
or   ( new_n21211_, new_n21140_, new_n20747_ );
and  ( new_n21212_, new_n21211_, new_n21210_ );
or   ( new_n21213_, new_n21212_, new_n21209_ );
and  ( new_n21214_, new_n21212_, new_n21209_ );
or   ( new_n21215_, new_n21151_, new_n20869_ );
or   ( new_n21216_, new_n21149_, new_n20720_ );
and  ( new_n21217_, new_n21216_, new_n21215_ );
or   ( new_n21218_, new_n21217_, new_n21214_ );
and  ( new_n21219_, new_n21218_, new_n21213_ );
or   ( new_n21220_, new_n20982_, new_n16217_ );
or   ( new_n21221_, new_n20978_, new_n16234_ );
and  ( new_n21222_, new_n21221_, new_n21220_ );
or   ( new_n21223_, new_n20991_, new_n16151_ );
or   ( new_n21224_, new_n20987_, new_n16170_ );
and  ( new_n21225_, new_n21224_, new_n21223_ );
or   ( new_n21226_, new_n21225_, new_n21222_ );
and  ( new_n21227_, new_n21225_, new_n21222_ );
or   ( new_n21228_, new_n21002_, new_n16108_ );
or   ( new_n21229_, new_n20998_, new_n16128_ );
and  ( new_n21230_, new_n21229_, new_n21228_ );
or   ( new_n21231_, new_n21230_, new_n21227_ );
and  ( new_n21232_, new_n21231_, new_n21226_ );
or   ( new_n21233_, new_n20951_, new_n16052_ );
or   ( new_n21234_, new_n20947_, new_n16071_ );
and  ( new_n21235_, new_n21234_, new_n21233_ );
or   ( new_n21236_, new_n20960_, new_n16009_ );
or   ( new_n21237_, new_n20956_, new_n16029_ );
and  ( new_n21238_, new_n21237_, new_n21236_ );
or   ( new_n21239_, new_n21238_, new_n21235_ );
and  ( new_n21240_, new_n21238_, new_n21235_ );
or   ( new_n21241_, new_n20971_, new_n16186_ );
or   ( new_n21242_, new_n20967_, new_n16204_ );
and  ( new_n21243_, new_n21242_, new_n21241_ );
or   ( new_n21244_, new_n21243_, new_n21240_ );
and  ( new_n21245_, new_n21244_, new_n21239_ );
or   ( new_n21246_, new_n21245_, new_n21232_ );
or   ( new_n21247_, new_n21042_, new_n18742_ );
or   ( new_n21248_, new_n21038_, new_n18977_ );
and  ( new_n21249_, new_n21248_, new_n21247_ );
or   ( new_n21250_, new_n21051_, new_n18066_ );
or   ( new_n21251_, new_n21047_, new_n18309_ );
and  ( new_n21252_, new_n21251_, new_n21250_ );
or   ( new_n21253_, new_n21252_, new_n21249_ );
and  ( new_n21254_, new_n21252_, new_n21249_ );
or   ( new_n21255_, new_n21062_, new_n17238_ );
or   ( new_n21256_, new_n21058_, new_n17650_ );
and  ( new_n21257_, new_n21256_, new_n21255_ );
or   ( new_n21258_, new_n21257_, new_n21254_ );
and  ( new_n21259_, new_n21258_, new_n21253_ );
nand ( new_n21260_, new_n21008_, new_n138_ );
and  ( new_n21261_, new_n21260_, RI2b1c4342c4f0_31 );
nand ( new_n21262_, new_n21010_, new_n138_ );
and  ( new_n21263_, new_n21262_, RI2b1c4342c478_30 );
and  ( new_n21264_, new_n21263_, new_n21261_ );
or   ( new_n21265_, new_n21264_, new_n20152_ );
or   ( new_n21266_, new_n21020_, new_n20156_ );
or   ( new_n21267_, new_n21016_, new_n20443_ );
and  ( new_n21268_, new_n21267_, new_n21266_ );
or   ( new_n21269_, new_n21268_, new_n21265_ );
and  ( new_n21270_, new_n21268_, new_n21265_ );
or   ( new_n21271_, new_n21031_, new_n19394_ );
or   ( new_n21272_, new_n21027_, new_n19659_ );
and  ( new_n21273_, new_n21272_, new_n21271_ );
or   ( new_n21274_, new_n21273_, new_n21270_ );
and  ( new_n21275_, new_n21274_, new_n21269_ );
or   ( new_n21276_, new_n21275_, new_n21259_ );
and  ( new_n21277_, new_n21275_, new_n21259_ );
or   ( new_n21278_, new_n21075_, new_n16814_ );
or   ( new_n21279_, new_n21071_, new_n17142_ );
and  ( new_n21280_, new_n21279_, new_n21278_ );
or   ( new_n21281_, new_n21084_, new_n16505_ );
or   ( new_n21282_, new_n21080_, new_n16438_ );
and  ( new_n21283_, new_n21282_, new_n21281_ );
or   ( new_n21284_, new_n21283_, new_n21280_ );
and  ( new_n21285_, new_n21283_, new_n21280_ );
or   ( new_n21286_, new_n21095_, new_n16085_ );
or   ( new_n21287_, new_n21091_, new_n16048_ );
and  ( new_n21288_, new_n21287_, new_n21286_ );
or   ( new_n21289_, new_n21288_, new_n21285_ );
and  ( new_n21290_, new_n21289_, new_n21284_ );
or   ( new_n21291_, new_n21290_, new_n21277_ );
and  ( new_n21292_, new_n21291_, new_n21276_ );
or   ( new_n21293_, new_n21292_, new_n21246_ );
and  ( new_n21294_, new_n21292_, new_n21246_ );
or   ( new_n21295_, new_n21108_, new_n20862_ );
or   ( new_n21296_, new_n21106_, new_n20709_ );
and  ( new_n21297_, new_n21296_, new_n21295_ );
or   ( new_n21298_, new_n21115_, new_n20851_ );
or   ( new_n21299_, new_n21113_, new_n20686_ );
and  ( new_n21300_, new_n21299_, new_n21298_ );
or   ( new_n21301_, new_n21300_, new_n21297_ );
and  ( new_n21302_, new_n21300_, new_n21297_ );
or   ( new_n21303_, new_n21124_, new_n20836_ );
or   ( new_n21304_, new_n21122_, new_n20653_ );
and  ( new_n21305_, new_n21304_, new_n21303_ );
or   ( new_n21306_, new_n21305_, new_n21302_ );
and  ( new_n21307_, new_n21306_, new_n21301_ );
or   ( new_n21308_, new_n21307_, new_n21294_ );
and  ( new_n21309_, new_n21308_, new_n21293_ );
or   ( new_n21310_, new_n21309_, new_n21219_ );
and  ( new_n21311_, new_n21309_, new_n21219_ );
or   ( new_n21312_, new_n21162_, new_n20468_ );
or   ( new_n21313_, new_n21160_, new_n20242_ );
and  ( new_n21314_, new_n21313_, new_n21312_ );
or   ( new_n21315_, new_n21314_, new_n21311_ );
and  ( new_n21316_, new_n21315_, new_n21310_ );
or   ( new_n21317_, new_n21316_, new_n21206_ );
and  ( new_n21318_, new_n21316_, new_n21206_ );
or   ( new_n21319_, new_n21173_, new_n20906_ );
or   ( new_n21320_, new_n21171_, new_n20760_ );
and  ( new_n21321_, new_n21320_, new_n21319_ );
or   ( new_n21322_, new_n21321_, new_n21318_ );
and  ( new_n21323_, new_n21322_, new_n21317_ );
or   ( new_n21324_, new_n21323_, new_n20937_ );
and  ( new_n21325_, new_n21324_, new_n21203_ );
or   ( new_n21326_, new_n21325_, new_n21199_ );
or   ( new_n21327_, new_n21323_, new_n21202_ );
and  ( new_n21328_, new_n21327_, new_n21178_ );
or   ( new_n21329_, new_n21328_, new_n21185_ );
and  ( new_n21330_, new_n21329_, new_n21326_ );
or   ( new_n21331_, new_n20871_, new_n20657_ );
or   ( new_n21332_, new_n20840_, new_n20722_ );
and  ( new_n21333_, new_n21332_, new_n21331_ );
or   ( new_n21334_, new_n21333_, new_n20886_ );
and  ( new_n21335_, new_n20872_, new_n20724_ );
or   ( new_n21336_, new_n21335_, new_n20749_ );
and  ( new_n21337_, new_n21336_, new_n21334_ );
or   ( new_n21338_, new_n21219_, new_n21130_ );
or   ( new_n21339_, new_n21309_, new_n21155_ );
and  ( new_n21340_, new_n21339_, new_n21338_ );
or   ( new_n21341_, new_n21340_, new_n21314_ );
and  ( new_n21342_, new_n21310_, new_n21156_ );
or   ( new_n21343_, new_n21342_, new_n21164_ );
and  ( new_n21344_, new_n21343_, new_n21341_ );
or   ( new_n21345_, new_n21344_, new_n21337_ );
or   ( new_n21346_, new_n20823_, new_n20591_ );
or   ( new_n21347_, new_n20810_, new_n20622_ );
and  ( new_n21348_, new_n21347_, new_n21346_ );
or   ( new_n21349_, new_n21348_, new_n20838_ );
and  ( new_n21350_, new_n20824_, new_n20623_ );
or   ( new_n21351_, new_n21350_, new_n20655_ );
and  ( new_n21352_, new_n21351_, new_n21349_ );
or   ( new_n21353_, new_n21212_, new_n21137_ );
or   ( new_n21354_, new_n21209_, new_n21144_ );
and  ( new_n21355_, new_n21354_, new_n21353_ );
or   ( new_n21356_, new_n21355_, new_n21217_ );
and  ( new_n21357_, new_n21213_, new_n21145_ );
or   ( new_n21358_, new_n21357_, new_n21153_ );
and  ( new_n21359_, new_n21358_, new_n21356_ );
or   ( new_n21360_, new_n21359_, new_n21352_ );
and  ( new_n21361_, new_n21359_, new_n21352_ );
or   ( new_n21362_, new_n21246_, new_n21101_ );
or   ( new_n21363_, new_n21292_, new_n21007_ );
and  ( new_n21364_, new_n21363_, new_n21362_ );
or   ( new_n21365_, new_n21364_, new_n21307_ );
and  ( new_n21366_, new_n21293_, new_n21102_ );
or   ( new_n21367_, new_n21366_, new_n21128_ );
and  ( new_n21368_, new_n21367_, new_n21365_ );
or   ( new_n21369_, new_n21368_, new_n21361_ );
and  ( new_n21370_, new_n21369_, new_n21360_ );
or   ( new_n21371_, new_n20816_, new_n20600_ );
or   ( new_n21372_, new_n20813_, new_n20609_ );
and  ( new_n21373_, new_n21372_, new_n21371_ );
or   ( new_n21374_, new_n21373_, new_n20821_ );
and  ( new_n21375_, new_n20817_, new_n20610_ );
or   ( new_n21376_, new_n21375_, new_n20620_ );
and  ( new_n21377_, new_n21376_, new_n21374_ );
or   ( new_n21378_, new_n21283_, new_n21077_ );
or   ( new_n21379_, new_n21280_, new_n21086_ );
and  ( new_n21380_, new_n21379_, new_n21378_ );
or   ( new_n21381_, new_n21380_, new_n21288_ );
and  ( new_n21382_, new_n21284_, new_n21087_ );
or   ( new_n21383_, new_n21382_, new_n21097_ );
and  ( new_n21384_, new_n21383_, new_n21381_ );
or   ( new_n21385_, new_n21252_, new_n21044_ );
or   ( new_n21386_, new_n21249_, new_n21053_ );
and  ( new_n21387_, new_n21386_, new_n21385_ );
or   ( new_n21388_, new_n21387_, new_n21257_ );
and  ( new_n21389_, new_n21253_, new_n21054_ );
or   ( new_n21390_, new_n21389_, new_n21064_ );
and  ( new_n21391_, new_n21390_, new_n21388_ );
or   ( new_n21392_, new_n21391_, new_n21384_ );
and  ( new_n21393_, new_n21391_, new_n21384_ );
or   ( new_n21394_, new_n21268_, new_n21013_ );
or   ( new_n21395_, new_n21265_, new_n21022_ );
and  ( new_n21396_, new_n21395_, new_n21394_ );
or   ( new_n21397_, new_n21396_, new_n21273_ );
and  ( new_n21398_, new_n21269_, new_n21023_ );
or   ( new_n21399_, new_n21398_, new_n21033_ );
and  ( new_n21400_, new_n21399_, new_n21397_ );
or   ( new_n21401_, new_n21400_, new_n21393_ );
and  ( new_n21402_, new_n21401_, new_n21392_ );
or   ( new_n21403_, new_n21402_, new_n21377_ );
and  ( new_n21404_, new_n21402_, new_n21377_ );
or   ( new_n21405_, new_n20803_, new_n20569_ );
or   ( new_n21406_, new_n20800_, new_n20578_ );
and  ( new_n21407_, new_n21406_, new_n21405_ );
or   ( new_n21408_, new_n21407_, new_n20808_ );
and  ( new_n21409_, new_n20804_, new_n20579_ );
or   ( new_n21410_, new_n21409_, new_n20589_ );
and  ( new_n21411_, new_n21410_, new_n21408_ );
or   ( new_n21412_, new_n21411_, new_n21404_ );
and  ( new_n21413_, new_n21412_, new_n21403_ );
or   ( new_n21414_, new_n21263_, new_n21261_ );
and  ( new_n21415_, new_n21414_, new_n21012_ );
or   ( new_n21416_, new_n21263_, new_n20152_ );
or   ( new_n21417_, new_n21011_, new_n20439_ );
and  ( new_n21418_, new_n21417_, new_n21416_ );
or   ( new_n21419_, new_n21418_, new_n21415_ );
or   ( new_n21420_, new_n21419_, new_n99_ );
or   ( new_n21421_, new_n21420_, new_n21013_ );
or   ( new_n21422_, new_n21261_, new_n21011_ );
or   ( new_n21423_, new_n21263_, new_n21009_ );
and  ( new_n21424_, new_n21423_, new_n21422_ );
or   ( new_n21425_, new_n21011_, new_n20152_ );
or   ( new_n21426_, new_n21263_, new_n20439_ );
and  ( new_n21427_, new_n21426_, new_n21425_ );
and  ( new_n21428_, new_n21427_, new_n21424_ );
and  ( new_n21429_, new_n21428_, RI2b1c4342d4e0_65 );
or   ( new_n21430_, new_n21429_, new_n21265_ );
and  ( new_n21431_, new_n21430_, new_n21421_ );
or   ( new_n21432_, new_n20557_, new_n112_ );
or   ( new_n21433_, new_n20562_, new_n526_ );
and  ( new_n21434_, new_n21433_, new_n21432_ );
or   ( new_n21435_, new_n21434_, new_n20156_ );
and  ( new_n21436_, new_n20566_, RI2b1c4342d5d0_67 );
and  ( new_n21437_, new_n20553_, RI2b1c4342d558_66 );
or   ( new_n21438_, new_n21437_, new_n21436_ );
or   ( new_n21439_, new_n21438_, new_n20443_ );
and  ( new_n21440_, new_n21439_, new_n21435_ );
or   ( new_n21441_, new_n21440_, new_n21431_ );
and  ( new_n21442_, new_n21440_, new_n21431_ );
or   ( new_n21443_, new_n19758_, new_n591_ );
or   ( new_n21444_, new_n19763_, new_n612_ );
and  ( new_n21445_, new_n21444_, new_n21443_ );
or   ( new_n21446_, new_n21445_, new_n19394_ );
and  ( new_n21447_, new_n19767_, RI2b1c4342d6c0_69 );
and  ( new_n21448_, new_n19754_, RI2b1c4342d648_68 );
or   ( new_n21449_, new_n21448_, new_n21447_ );
or   ( new_n21450_, new_n21449_, new_n19659_ );
and  ( new_n21451_, new_n21450_, new_n21446_ );
or   ( new_n21452_, new_n21451_, new_n21442_ );
and  ( new_n21453_, new_n21452_, new_n21441_ );
or   ( new_n21454_, new_n19048_, new_n110_ );
or   ( new_n21455_, new_n19055_, new_n755_ );
and  ( new_n21456_, new_n21455_, new_n21454_ );
or   ( new_n21457_, new_n21456_, new_n18742_ );
and  ( new_n21458_, new_n19057_, RI2b1c4342d7b0_71 );
and  ( new_n21459_, new_n19044_, RI2b1c4342d738_70 );
or   ( new_n21460_, new_n21459_, new_n21458_ );
or   ( new_n21461_, new_n21460_, new_n18977_ );
and  ( new_n21462_, new_n21461_, new_n21457_ );
or   ( new_n21463_, new_n18388_, new_n105_ );
or   ( new_n21464_, new_n18395_, new_n806_ );
and  ( new_n21465_, new_n21464_, new_n21463_ );
or   ( new_n21466_, new_n21465_, new_n18066_ );
and  ( new_n21467_, new_n18397_, RI2b1c4342d8a0_73 );
and  ( new_n21468_, new_n18384_, RI2b1c4342d828_72 );
or   ( new_n21469_, new_n21468_, new_n21467_ );
or   ( new_n21470_, new_n21469_, new_n18309_ );
and  ( new_n21471_, new_n21470_, new_n21466_ );
or   ( new_n21472_, new_n21471_, new_n21462_ );
and  ( new_n21473_, new_n21471_, new_n21462_ );
or   ( new_n21474_, new_n17727_, new_n843_ );
or   ( new_n21475_, new_n17734_, new_n859_ );
and  ( new_n21476_, new_n21475_, new_n21474_ );
or   ( new_n21477_, new_n21476_, new_n17238_ );
and  ( new_n21478_, new_n17736_, RI2b1c4342d990_75 );
and  ( new_n21479_, new_n17723_, RI2b1c4342d918_74 );
or   ( new_n21480_, new_n21479_, new_n21478_ );
or   ( new_n21481_, new_n21480_, new_n17650_ );
and  ( new_n21482_, new_n21481_, new_n21477_ );
or   ( new_n21483_, new_n21482_, new_n21473_ );
and  ( new_n21484_, new_n21483_, new_n21472_ );
or   ( new_n21485_, new_n21484_, new_n21453_ );
and  ( new_n21486_, new_n21484_, new_n21453_ );
or   ( new_n21487_, new_n17244_, new_n1004_ );
or   ( new_n21488_, new_n17248_, new_n886_ );
and  ( new_n21489_, new_n21488_, new_n21487_ );
or   ( new_n21490_, new_n21489_, new_n16814_ );
and  ( new_n21491_, new_n17255_, RI2b1c4342da80_77 );
and  ( new_n21492_, new_n17240_, RI2b1c4342da08_76 );
or   ( new_n21493_, new_n21492_, new_n21491_ );
or   ( new_n21494_, new_n21493_, new_n17142_ );
and  ( new_n21495_, new_n21494_, new_n21490_ );
or   ( new_n21496_, new_n16607_, new_n1310_ );
or   ( new_n21497_, new_n16613_, new_n1002_ );
and  ( new_n21498_, new_n21497_, new_n21496_ );
or   ( new_n21499_, new_n21498_, new_n16505_ );
and  ( new_n21500_, new_n16616_, RI2b1c4342db70_79 );
and  ( new_n21501_, new_n16603_, RI2b1c4342daf8_78 );
or   ( new_n21502_, new_n21501_, new_n21500_ );
or   ( new_n21503_, new_n21502_, new_n16438_ );
and  ( new_n21504_, new_n21503_, new_n21499_ );
or   ( new_n21505_, new_n21504_, new_n21495_ );
and  ( new_n21506_, new_n21504_, new_n21495_ );
or   ( new_n21507_, new_n16366_, new_n126_ );
or   ( new_n21508_, new_n16355_, new_n1511_ );
and  ( new_n21509_, new_n21508_, new_n21507_ );
or   ( new_n21510_, new_n21509_, new_n16085_ );
and  ( new_n21511_, new_n16358_, RI2b1c4342dc60_81 );
and  ( new_n21512_, new_n16362_, RI2b1c4342dbe8_80 );
or   ( new_n21513_, new_n21512_, new_n21511_ );
or   ( new_n21514_, new_n21513_, new_n16048_ );
and  ( new_n21515_, new_n21514_, new_n21510_ );
or   ( new_n21516_, new_n21515_, new_n21506_ );
and  ( new_n21517_, new_n21516_, new_n21505_ );
or   ( new_n21518_, new_n21517_, new_n21486_ );
and  ( new_n21519_, new_n21518_, new_n21485_ );
or   ( new_n21520_, new_n16075_, new_n121_ );
or   ( new_n21521_, new_n16060_, new_n2119_ );
and  ( new_n21522_, new_n21521_, new_n21520_ );
or   ( new_n21523_, new_n21522_, new_n16052_ );
and  ( new_n21524_, new_n16063_, RI2b1c4342dd50_83 );
and  ( new_n21525_, new_n16066_, RI2b1c4342dcd8_82 );
or   ( new_n21526_, new_n21525_, new_n21524_ );
or   ( new_n21527_, new_n21526_, new_n16071_ );
and  ( new_n21528_, new_n21527_, new_n21523_ );
or   ( new_n21529_, new_n16033_, new_n2806_ );
or   ( new_n21530_, new_n16017_, new_n2541_ );
and  ( new_n21531_, new_n21530_, new_n21529_ );
or   ( new_n21532_, new_n21531_, new_n16009_ );
and  ( new_n21533_, new_n16021_, RI2b1c4342de40_85 );
and  ( new_n21534_, new_n16024_, RI2b1c4342ddc8_84 );
or   ( new_n21535_, new_n21534_, new_n21533_ );
or   ( new_n21536_, new_n21535_, new_n16029_ );
and  ( new_n21537_, new_n21536_, new_n21532_ );
or   ( new_n21538_, new_n21537_, new_n21528_ );
and  ( new_n21539_, new_n21537_, new_n21528_ );
or   ( new_n21540_, new_n16208_, new_n3924_ );
or   ( new_n21541_, new_n16194_, new_n3239_ );
and  ( new_n21542_, new_n21541_, new_n21540_ );
or   ( new_n21543_, new_n21542_, new_n16186_ );
and  ( new_n21544_, new_n16196_, RI2b1c4342df30_87 );
and  ( new_n21545_, new_n16199_, RI2b1c4342deb8_86 );
or   ( new_n21546_, new_n21545_, new_n21544_ );
or   ( new_n21547_, new_n21546_, new_n16204_ );
and  ( new_n21548_, new_n21547_, new_n21543_ );
or   ( new_n21549_, new_n21548_, new_n21539_ );
and  ( new_n21550_, new_n21549_, new_n21538_ );
or   ( new_n21551_, new_n16238_, new_n132_ );
or   ( new_n21552_, new_n16224_, new_n3902_ );
and  ( new_n21553_, new_n21552_, new_n21551_ );
or   ( new_n21554_, new_n21553_, new_n16217_ );
and  ( new_n21555_, new_n16226_, RI2b1c4342e020_89 );
and  ( new_n21556_, new_n16229_, RI2b1c4342dfa8_88 );
or   ( new_n21557_, new_n21556_, new_n21555_ );
or   ( new_n21558_, new_n21557_, new_n16234_ );
and  ( new_n21559_, new_n21558_, new_n21554_ );
or   ( new_n21560_, new_n16174_, new_n117_ );
or   ( new_n21561_, new_n16160_, new_n4635_ );
and  ( new_n21562_, new_n21561_, new_n21560_ );
or   ( new_n21563_, new_n21562_, new_n16151_ );
and  ( new_n21564_, new_n16162_, RI2b1c4342e110_91 );
and  ( new_n21565_, new_n16165_, RI2b1c4342e098_90 );
or   ( new_n21566_, new_n21565_, new_n21564_ );
or   ( new_n21567_, new_n21566_, new_n16170_ );
and  ( new_n21568_, new_n21567_, new_n21563_ );
or   ( new_n21569_, new_n21568_, new_n21559_ );
and  ( new_n21570_, new_n21568_, new_n21559_ );
or   ( new_n21571_, new_n16119_, new_n6307_ );
or   ( new_n21572_, new_n16123_, new_n5459_ );
and  ( new_n21573_, new_n21572_, new_n21571_ );
or   ( new_n21574_, new_n21573_, new_n16108_ );
and  ( new_n21575_, new_n16132_, RI2b1c4342e200_93 );
and  ( new_n21576_, new_n16114_, RI2b1c4342e188_92 );
or   ( new_n21577_, new_n21576_, new_n21575_ );
or   ( new_n21578_, new_n21577_, new_n16128_ );
and  ( new_n21579_, new_n21578_, new_n21574_ );
or   ( new_n21580_, new_n21579_, new_n21570_ );
and  ( new_n21581_, new_n21580_, new_n21569_ );
and  ( new_n21582_, new_n21581_, new_n21550_ );
or   ( new_n21583_, new_n21581_, new_n21550_ );
or   ( new_n21584_, new_n16115_, new_n6321_ );
and  ( new_n21585_, new_n21584_, new_n21583_ );
or   ( new_n21586_, new_n21585_, new_n21582_ );
and  ( new_n21587_, new_n21586_, new_n21519_ );
or   ( new_n21588_, new_n21586_, new_n21519_ );
or   ( new_n21589_, new_n16115_, new_n6307_ );
or   ( new_n21590_, new_n21225_, new_n20984_ );
or   ( new_n21591_, new_n21222_, new_n20993_ );
and  ( new_n21592_, new_n21591_, new_n21590_ );
or   ( new_n21593_, new_n21592_, new_n21230_ );
and  ( new_n21594_, new_n21226_, new_n20994_ );
or   ( new_n21595_, new_n21594_, new_n21004_ );
and  ( new_n21596_, new_n21595_, new_n21593_ );
or   ( new_n21597_, new_n21596_, new_n21589_ );
and  ( new_n21598_, new_n21596_, new_n21589_ );
or   ( new_n21599_, new_n21238_, new_n20953_ );
or   ( new_n21600_, new_n21235_, new_n20962_ );
and  ( new_n21601_, new_n21600_, new_n21599_ );
or   ( new_n21602_, new_n21601_, new_n21243_ );
and  ( new_n21603_, new_n21239_, new_n20963_ );
or   ( new_n21604_, new_n21603_, new_n20973_ );
and  ( new_n21605_, new_n21604_, new_n21602_ );
or   ( new_n21606_, new_n21605_, new_n21598_ );
and  ( new_n21607_, new_n21606_, new_n21597_ );
and  ( new_n21608_, new_n21607_, new_n21588_ );
or   ( new_n21609_, new_n21608_, new_n21587_ );
and  ( new_n21610_, new_n21609_, new_n21413_ );
or   ( new_n21611_, new_n21609_, new_n21413_ );
or   ( new_n21612_, new_n21300_, new_n21110_ );
or   ( new_n21613_, new_n21297_, new_n21117_ );
and  ( new_n21614_, new_n21613_, new_n21612_ );
or   ( new_n21615_, new_n21614_, new_n21305_ );
and  ( new_n21616_, new_n21301_, new_n21118_ );
or   ( new_n21617_, new_n21616_, new_n21126_ );
and  ( new_n21618_, new_n21617_, new_n21615_ );
or   ( new_n21619_, new_n21006_, new_n20975_ );
and  ( new_n21620_, new_n21619_, new_n21246_ );
or   ( new_n21621_, new_n21620_, new_n21618_ );
and  ( new_n21622_, new_n21620_, new_n21618_ );
or   ( new_n21623_, new_n21259_, new_n21035_ );
or   ( new_n21624_, new_n21275_, new_n21066_ );
and  ( new_n21625_, new_n21624_, new_n21623_ );
or   ( new_n21626_, new_n21625_, new_n21290_ );
and  ( new_n21627_, new_n21276_, new_n21067_ );
or   ( new_n21628_, new_n21627_, new_n21099_ );
and  ( new_n21629_, new_n21628_, new_n21626_ );
or   ( new_n21630_, new_n21629_, new_n21622_ );
and  ( new_n21631_, new_n21630_, new_n21621_ );
and  ( new_n21632_, new_n21631_, new_n21611_ );
or   ( new_n21633_, new_n21632_, new_n21610_ );
and  ( new_n21634_, new_n21633_, new_n21370_ );
or   ( new_n21635_, new_n21633_, new_n21370_ );
or   ( new_n21636_, new_n20894_, new_n20533_ );
or   ( new_n21637_, new_n20891_, new_n20540_ );
and  ( new_n21638_, new_n21637_, new_n21636_ );
or   ( new_n21639_, new_n21638_, new_n20899_ );
and  ( new_n21640_, new_n20895_, new_n20541_ );
or   ( new_n21641_, new_n21640_, new_n20549_ );
and  ( new_n21642_, new_n21641_, new_n21639_ );
and  ( new_n21643_, new_n21642_, new_n21635_ );
or   ( new_n21644_, new_n21643_, new_n21634_ );
and  ( new_n21645_, new_n21644_, new_n21345_ );
or   ( new_n21646_, new_n21644_, new_n21345_ );
or   ( new_n21647_, new_n21206_, new_n21166_ );
or   ( new_n21648_, new_n21316_, new_n20944_ );
and  ( new_n21649_, new_n21648_, new_n21647_ );
or   ( new_n21650_, new_n21649_, new_n21321_ );
and  ( new_n21651_, new_n21317_, new_n21167_ );
or   ( new_n21652_, new_n21651_, new_n21175_ );
and  ( new_n21653_, new_n21652_, new_n21650_ );
and  ( new_n21654_, new_n21653_, new_n21646_ );
or   ( new_n21655_, new_n21654_, new_n21645_ );
and  ( new_n21656_, new_n21655_, new_n21330_ );
or   ( new_n21657_, new_n21655_, new_n21330_ );
or   ( new_n21658_, new_n21651_, new_n21321_ );
or   ( new_n21659_, new_n21649_, new_n21175_ );
and  ( new_n21660_, new_n21659_, new_n21658_ );
or   ( new_n21661_, new_n21335_, new_n20886_ );
or   ( new_n21662_, new_n21333_, new_n20749_ );
and  ( new_n21663_, new_n21662_, new_n21661_ );
or   ( new_n21664_, new_n21342_, new_n21314_ );
or   ( new_n21665_, new_n21340_, new_n21164_ );
and  ( new_n21666_, new_n21665_, new_n21664_ );
and  ( new_n21667_, new_n21666_, new_n21663_ );
or   ( new_n21668_, new_n21667_, new_n21644_ );
or   ( new_n21669_, new_n21429_, new_n21013_ );
or   ( new_n21670_, new_n21420_, new_n21265_ );
and  ( new_n21671_, new_n21670_, new_n21669_ );
or   ( new_n21672_, new_n21438_, new_n20156_ );
or   ( new_n21673_, new_n21434_, new_n20443_ );
and  ( new_n21674_, new_n21673_, new_n21672_ );
or   ( new_n21675_, new_n21674_, new_n21671_ );
and  ( new_n21676_, new_n21674_, new_n21671_ );
or   ( new_n21677_, new_n21449_, new_n19394_ );
or   ( new_n21678_, new_n21445_, new_n19659_ );
and  ( new_n21679_, new_n21678_, new_n21677_ );
or   ( new_n21680_, new_n21679_, new_n21676_ );
and  ( new_n21681_, new_n21680_, new_n21675_ );
or   ( new_n21682_, new_n21460_, new_n18742_ );
or   ( new_n21683_, new_n21456_, new_n18977_ );
and  ( new_n21684_, new_n21683_, new_n21682_ );
or   ( new_n21685_, new_n21469_, new_n18066_ );
or   ( new_n21686_, new_n21465_, new_n18309_ );
and  ( new_n21687_, new_n21686_, new_n21685_ );
or   ( new_n21688_, new_n21687_, new_n21684_ );
and  ( new_n21689_, new_n21687_, new_n21684_ );
or   ( new_n21690_, new_n21480_, new_n17238_ );
or   ( new_n21691_, new_n21476_, new_n17650_ );
and  ( new_n21692_, new_n21691_, new_n21690_ );
or   ( new_n21693_, new_n21692_, new_n21689_ );
and  ( new_n21694_, new_n21693_, new_n21688_ );
or   ( new_n21695_, new_n21694_, new_n21681_ );
and  ( new_n21696_, new_n21694_, new_n21681_ );
or   ( new_n21697_, new_n21493_, new_n16814_ );
or   ( new_n21698_, new_n21489_, new_n17142_ );
and  ( new_n21699_, new_n21698_, new_n21697_ );
or   ( new_n21700_, new_n21502_, new_n16505_ );
or   ( new_n21701_, new_n21498_, new_n16438_ );
and  ( new_n21702_, new_n21701_, new_n21700_ );
or   ( new_n21703_, new_n21702_, new_n21699_ );
and  ( new_n21704_, new_n21702_, new_n21699_ );
or   ( new_n21705_, new_n21513_, new_n16085_ );
or   ( new_n21706_, new_n21509_, new_n16048_ );
and  ( new_n21707_, new_n21706_, new_n21705_ );
or   ( new_n21708_, new_n21707_, new_n21704_ );
and  ( new_n21709_, new_n21708_, new_n21703_ );
or   ( new_n21710_, new_n21709_, new_n21696_ );
and  ( new_n21711_, new_n21710_, new_n21695_ );
or   ( new_n21712_, new_n21526_, new_n16052_ );
or   ( new_n21713_, new_n21522_, new_n16071_ );
and  ( new_n21714_, new_n21713_, new_n21712_ );
or   ( new_n21715_, new_n21535_, new_n16009_ );
or   ( new_n21716_, new_n21531_, new_n16029_ );
and  ( new_n21717_, new_n21716_, new_n21715_ );
or   ( new_n21718_, new_n21717_, new_n21714_ );
and  ( new_n21719_, new_n21717_, new_n21714_ );
or   ( new_n21720_, new_n21546_, new_n16186_ );
or   ( new_n21721_, new_n21542_, new_n16204_ );
and  ( new_n21722_, new_n21721_, new_n21720_ );
or   ( new_n21723_, new_n21722_, new_n21719_ );
and  ( new_n21724_, new_n21723_, new_n21718_ );
or   ( new_n21725_, new_n21557_, new_n16217_ );
or   ( new_n21726_, new_n21553_, new_n16234_ );
and  ( new_n21727_, new_n21726_, new_n21725_ );
or   ( new_n21728_, new_n21566_, new_n16151_ );
or   ( new_n21729_, new_n21562_, new_n16170_ );
and  ( new_n21730_, new_n21729_, new_n21728_ );
or   ( new_n21731_, new_n21730_, new_n21727_ );
and  ( new_n21732_, new_n21730_, new_n21727_ );
or   ( new_n21733_, new_n21577_, new_n16108_ );
or   ( new_n21734_, new_n21573_, new_n16128_ );
and  ( new_n21735_, new_n21734_, new_n21733_ );
or   ( new_n21736_, new_n21735_, new_n21732_ );
and  ( new_n21737_, new_n21736_, new_n21731_ );
or   ( new_n21738_, new_n21737_, new_n21724_ );
and  ( new_n21739_, new_n21737_, new_n21724_ );
and  ( new_n21740_, new_n16102_, RI2b1c4342e278_94 );
or   ( new_n21741_, new_n21740_, new_n21739_ );
and  ( new_n21742_, new_n21741_, new_n21738_ );
or   ( new_n21743_, new_n21742_, new_n21711_ );
and  ( new_n21744_, new_n21742_, new_n21711_ );
and  ( new_n21745_, new_n16102_, RI2b1c4342e200_93 );
or   ( new_n21746_, new_n21594_, new_n21230_ );
or   ( new_n21747_, new_n21592_, new_n21004_ );
and  ( new_n21748_, new_n21747_, new_n21746_ );
or   ( new_n21749_, new_n21748_, new_n21745_ );
and  ( new_n21750_, new_n21748_, new_n21745_ );
or   ( new_n21751_, new_n21603_, new_n21243_ );
or   ( new_n21752_, new_n21601_, new_n20973_ );
and  ( new_n21753_, new_n21752_, new_n21751_ );
or   ( new_n21754_, new_n21753_, new_n21750_ );
and  ( new_n21755_, new_n21754_, new_n21749_ );
or   ( new_n21756_, new_n21755_, new_n21744_ );
and  ( new_n21757_, new_n21756_, new_n21743_ );
or   ( new_n21758_, new_n21375_, new_n20821_ );
or   ( new_n21759_, new_n21373_, new_n20620_ );
and  ( new_n21760_, new_n21759_, new_n21758_ );
or   ( new_n21761_, new_n21382_, new_n21288_ );
or   ( new_n21762_, new_n21380_, new_n21097_ );
and  ( new_n21763_, new_n21762_, new_n21761_ );
or   ( new_n21764_, new_n21389_, new_n21257_ );
or   ( new_n21765_, new_n21387_, new_n21064_ );
and  ( new_n21766_, new_n21765_, new_n21764_ );
or   ( new_n21767_, new_n21766_, new_n21763_ );
and  ( new_n21768_, new_n21766_, new_n21763_ );
or   ( new_n21769_, new_n21398_, new_n21273_ );
or   ( new_n21770_, new_n21396_, new_n21033_ );
and  ( new_n21771_, new_n21770_, new_n21769_ );
or   ( new_n21772_, new_n21771_, new_n21768_ );
and  ( new_n21773_, new_n21772_, new_n21767_ );
or   ( new_n21774_, new_n21773_, new_n21760_ );
and  ( new_n21775_, new_n21773_, new_n21760_ );
or   ( new_n21776_, new_n21409_, new_n20808_ );
or   ( new_n21777_, new_n21407_, new_n20589_ );
and  ( new_n21778_, new_n21777_, new_n21776_ );
or   ( new_n21779_, new_n21778_, new_n21775_ );
and  ( new_n21780_, new_n21779_, new_n21774_ );
or   ( new_n21781_, new_n21780_, new_n21757_ );
and  ( new_n21782_, new_n21780_, new_n21757_ );
or   ( new_n21783_, new_n21616_, new_n21305_ );
or   ( new_n21784_, new_n21614_, new_n21126_ );
and  ( new_n21785_, new_n21784_, new_n21783_ );
or   ( new_n21786_, new_n21232_, new_n20975_ );
or   ( new_n21787_, new_n21245_, new_n21006_ );
and  ( new_n21788_, new_n21787_, new_n21786_ );
or   ( new_n21789_, new_n21788_, new_n21785_ );
and  ( new_n21790_, new_n21788_, new_n21785_ );
or   ( new_n21791_, new_n21627_, new_n21290_ );
or   ( new_n21792_, new_n21625_, new_n21099_ );
and  ( new_n21793_, new_n21792_, new_n21791_ );
or   ( new_n21794_, new_n21793_, new_n21790_ );
and  ( new_n21795_, new_n21794_, new_n21789_ );
or   ( new_n21796_, new_n21795_, new_n21782_ );
and  ( new_n21797_, new_n21796_, new_n21781_ );
or   ( new_n21798_, new_n21350_, new_n20838_ );
or   ( new_n21799_, new_n21348_, new_n20655_ );
and  ( new_n21800_, new_n21799_, new_n21798_ );
or   ( new_n21801_, new_n21357_, new_n21217_ );
or   ( new_n21802_, new_n21355_, new_n21153_ );
and  ( new_n21803_, new_n21802_, new_n21801_ );
or   ( new_n21804_, new_n21803_, new_n21800_ );
and  ( new_n21805_, new_n21803_, new_n21800_ );
or   ( new_n21806_, new_n21366_, new_n21307_ );
or   ( new_n21807_, new_n21364_, new_n21128_ );
and  ( new_n21808_, new_n21807_, new_n21806_ );
or   ( new_n21809_, new_n21808_, new_n21805_ );
and  ( new_n21810_, new_n21809_, new_n21804_ );
or   ( new_n21811_, new_n21810_, new_n21797_ );
and  ( new_n21812_, new_n21810_, new_n21797_ );
or   ( new_n21813_, new_n21640_, new_n20899_ );
or   ( new_n21814_, new_n21638_, new_n20549_ );
and  ( new_n21815_, new_n21814_, new_n21813_ );
or   ( new_n21816_, new_n21815_, new_n21812_ );
and  ( new_n21817_, new_n21816_, new_n21811_ );
or   ( new_n21818_, new_n21817_, new_n21345_ );
and  ( new_n21819_, new_n21818_, new_n21668_ );
or   ( new_n21820_, new_n21819_, new_n21660_ );
or   ( new_n21821_, new_n21817_, new_n21667_ );
and  ( new_n21822_, new_n21821_, new_n21646_ );
or   ( new_n21823_, new_n21822_, new_n21653_ );
and  ( new_n21824_, new_n21823_, new_n21820_ );
or   ( new_n21825_, new_n21666_, new_n21337_ );
or   ( new_n21826_, new_n21663_, new_n21344_ );
and  ( new_n21827_, new_n21826_, new_n21825_ );
or   ( new_n21828_, new_n21803_, new_n21352_ );
or   ( new_n21829_, new_n21800_, new_n21359_ );
and  ( new_n21830_, new_n21829_, new_n21828_ );
or   ( new_n21831_, new_n21830_, new_n21808_ );
and  ( new_n21832_, new_n21804_, new_n21360_ );
or   ( new_n21833_, new_n21832_, new_n21368_ );
and  ( new_n21834_, new_n21833_, new_n21831_ );
or   ( new_n21835_, new_n21419_, new_n526_ );
or   ( new_n21836_, new_n21424_, new_n99_ );
and  ( new_n21837_, new_n21836_, new_n21835_ );
or   ( new_n21838_, new_n21837_, new_n21013_ );
and  ( new_n21839_, new_n21428_, RI2b1c4342d558_66 );
and  ( new_n21840_, new_n21415_, RI2b1c4342d4e0_65 );
or   ( new_n21841_, new_n21840_, new_n21839_ );
or   ( new_n21842_, new_n21841_, new_n21265_ );
and  ( new_n21843_, new_n21842_, new_n21838_ );
or   ( new_n21844_, new_n21843_, new_n21261_ );
and  ( new_n21845_, new_n21843_, new_n21261_ );
or   ( new_n21846_, new_n20557_, new_n612_ );
or   ( new_n21847_, new_n20562_, new_n112_ );
and  ( new_n21848_, new_n21847_, new_n21846_ );
or   ( new_n21849_, new_n21848_, new_n20156_ );
and  ( new_n21850_, new_n20566_, RI2b1c4342d648_68 );
and  ( new_n21851_, new_n20553_, RI2b1c4342d5d0_67 );
or   ( new_n21852_, new_n21851_, new_n21850_ );
or   ( new_n21853_, new_n21852_, new_n20443_ );
and  ( new_n21854_, new_n21853_, new_n21849_ );
or   ( new_n21855_, new_n21854_, new_n21845_ );
and  ( new_n21856_, new_n21855_, new_n21844_ );
or   ( new_n21857_, new_n19758_, new_n755_ );
or   ( new_n21858_, new_n19763_, new_n591_ );
and  ( new_n21859_, new_n21858_, new_n21857_ );
or   ( new_n21860_, new_n21859_, new_n19394_ );
and  ( new_n21861_, new_n19767_, RI2b1c4342d738_70 );
and  ( new_n21862_, new_n19754_, RI2b1c4342d6c0_69 );
or   ( new_n21863_, new_n21862_, new_n21861_ );
or   ( new_n21864_, new_n21863_, new_n19659_ );
and  ( new_n21865_, new_n21864_, new_n21860_ );
or   ( new_n21866_, new_n19048_, new_n806_ );
or   ( new_n21867_, new_n19055_, new_n110_ );
and  ( new_n21868_, new_n21867_, new_n21866_ );
or   ( new_n21869_, new_n21868_, new_n18742_ );
and  ( new_n21870_, new_n19057_, RI2b1c4342d828_72 );
and  ( new_n21871_, new_n19044_, RI2b1c4342d7b0_71 );
or   ( new_n21872_, new_n21871_, new_n21870_ );
or   ( new_n21873_, new_n21872_, new_n18977_ );
and  ( new_n21874_, new_n21873_, new_n21869_ );
or   ( new_n21875_, new_n21874_, new_n21865_ );
and  ( new_n21876_, new_n21874_, new_n21865_ );
or   ( new_n21877_, new_n18388_, new_n859_ );
or   ( new_n21878_, new_n18395_, new_n105_ );
and  ( new_n21879_, new_n21878_, new_n21877_ );
or   ( new_n21880_, new_n21879_, new_n18066_ );
and  ( new_n21881_, new_n18397_, RI2b1c4342d918_74 );
and  ( new_n21882_, new_n18384_, RI2b1c4342d8a0_73 );
or   ( new_n21883_, new_n21882_, new_n21881_ );
or   ( new_n21884_, new_n21883_, new_n18309_ );
and  ( new_n21885_, new_n21884_, new_n21880_ );
or   ( new_n21886_, new_n21885_, new_n21876_ );
and  ( new_n21887_, new_n21886_, new_n21875_ );
or   ( new_n21888_, new_n21887_, new_n21856_ );
and  ( new_n21889_, new_n21887_, new_n21856_ );
or   ( new_n21890_, new_n17727_, new_n886_ );
or   ( new_n21891_, new_n17734_, new_n843_ );
and  ( new_n21892_, new_n21891_, new_n21890_ );
or   ( new_n21893_, new_n21892_, new_n17238_ );
and  ( new_n21894_, new_n17736_, RI2b1c4342da08_76 );
and  ( new_n21895_, new_n17723_, RI2b1c4342d990_75 );
or   ( new_n21896_, new_n21895_, new_n21894_ );
or   ( new_n21897_, new_n21896_, new_n17650_ );
and  ( new_n21898_, new_n21897_, new_n21893_ );
or   ( new_n21899_, new_n17244_, new_n1002_ );
or   ( new_n21900_, new_n17248_, new_n1004_ );
and  ( new_n21901_, new_n21900_, new_n21899_ );
or   ( new_n21902_, new_n21901_, new_n16814_ );
and  ( new_n21903_, new_n17255_, RI2b1c4342daf8_78 );
and  ( new_n21904_, new_n17240_, RI2b1c4342da80_77 );
or   ( new_n21905_, new_n21904_, new_n21903_ );
or   ( new_n21906_, new_n21905_, new_n17142_ );
and  ( new_n21907_, new_n21906_, new_n21902_ );
or   ( new_n21908_, new_n21907_, new_n21898_ );
and  ( new_n21909_, new_n21907_, new_n21898_ );
or   ( new_n21910_, new_n16607_, new_n1511_ );
or   ( new_n21911_, new_n16613_, new_n1310_ );
and  ( new_n21912_, new_n21911_, new_n21910_ );
or   ( new_n21913_, new_n21912_, new_n16505_ );
and  ( new_n21914_, new_n16616_, RI2b1c4342dbe8_80 );
and  ( new_n21915_, new_n16603_, RI2b1c4342db70_79 );
or   ( new_n21916_, new_n21915_, new_n21914_ );
or   ( new_n21917_, new_n21916_, new_n16438_ );
and  ( new_n21918_, new_n21917_, new_n21913_ );
or   ( new_n21919_, new_n21918_, new_n21909_ );
and  ( new_n21920_, new_n21919_, new_n21908_ );
or   ( new_n21921_, new_n21920_, new_n21889_ );
and  ( new_n21922_, new_n21921_, new_n21888_ );
or   ( new_n21923_, new_n16366_, new_n2119_ );
or   ( new_n21924_, new_n16355_, new_n126_ );
and  ( new_n21925_, new_n21924_, new_n21923_ );
or   ( new_n21926_, new_n21925_, new_n16085_ );
and  ( new_n21927_, new_n16358_, RI2b1c4342dcd8_82 );
and  ( new_n21928_, new_n16362_, RI2b1c4342dc60_81 );
or   ( new_n21929_, new_n21928_, new_n21927_ );
or   ( new_n21930_, new_n21929_, new_n16048_ );
and  ( new_n21931_, new_n21930_, new_n21926_ );
or   ( new_n21932_, new_n16075_, new_n2541_ );
or   ( new_n21933_, new_n16060_, new_n121_ );
and  ( new_n21934_, new_n21933_, new_n21932_ );
or   ( new_n21935_, new_n21934_, new_n16052_ );
and  ( new_n21936_, new_n16063_, RI2b1c4342ddc8_84 );
and  ( new_n21937_, new_n16066_, RI2b1c4342dd50_83 );
or   ( new_n21938_, new_n21937_, new_n21936_ );
or   ( new_n21939_, new_n21938_, new_n16071_ );
and  ( new_n21940_, new_n21939_, new_n21935_ );
or   ( new_n21941_, new_n21940_, new_n21931_ );
and  ( new_n21942_, new_n21940_, new_n21931_ );
or   ( new_n21943_, new_n16033_, new_n3239_ );
or   ( new_n21944_, new_n16017_, new_n2806_ );
and  ( new_n21945_, new_n21944_, new_n21943_ );
or   ( new_n21946_, new_n21945_, new_n16009_ );
and  ( new_n21947_, new_n16021_, RI2b1c4342deb8_86 );
and  ( new_n21948_, new_n16024_, RI2b1c4342de40_85 );
or   ( new_n21949_, new_n21948_, new_n21947_ );
or   ( new_n21950_, new_n21949_, new_n16029_ );
and  ( new_n21951_, new_n21950_, new_n21946_ );
or   ( new_n21952_, new_n21951_, new_n21942_ );
and  ( new_n21953_, new_n21952_, new_n21941_ );
or   ( new_n21954_, new_n16208_, new_n3902_ );
or   ( new_n21955_, new_n16194_, new_n3924_ );
and  ( new_n21956_, new_n21955_, new_n21954_ );
or   ( new_n21957_, new_n21956_, new_n16186_ );
and  ( new_n21958_, new_n16196_, RI2b1c4342dfa8_88 );
and  ( new_n21959_, new_n16199_, RI2b1c4342df30_87 );
or   ( new_n21960_, new_n21959_, new_n21958_ );
or   ( new_n21961_, new_n21960_, new_n16204_ );
and  ( new_n21962_, new_n21961_, new_n21957_ );
or   ( new_n21963_, new_n16238_, new_n4635_ );
or   ( new_n21964_, new_n16224_, new_n132_ );
and  ( new_n21965_, new_n21964_, new_n21963_ );
or   ( new_n21966_, new_n21965_, new_n16217_ );
and  ( new_n21967_, new_n16226_, RI2b1c4342e098_90 );
and  ( new_n21968_, new_n16229_, RI2b1c4342e020_89 );
or   ( new_n21969_, new_n21968_, new_n21967_ );
or   ( new_n21970_, new_n21969_, new_n16234_ );
and  ( new_n21971_, new_n21970_, new_n21966_ );
or   ( new_n21972_, new_n21971_, new_n21962_ );
and  ( new_n21973_, new_n21971_, new_n21962_ );
or   ( new_n21974_, new_n16174_, new_n5459_ );
or   ( new_n21975_, new_n16160_, new_n117_ );
and  ( new_n21976_, new_n21975_, new_n21974_ );
or   ( new_n21977_, new_n21976_, new_n16151_ );
and  ( new_n21978_, new_n16162_, RI2b1c4342e188_92 );
and  ( new_n21979_, new_n16165_, RI2b1c4342e110_91 );
or   ( new_n21980_, new_n21979_, new_n21978_ );
or   ( new_n21981_, new_n21980_, new_n16170_ );
and  ( new_n21982_, new_n21981_, new_n21977_ );
or   ( new_n21983_, new_n21982_, new_n21973_ );
and  ( new_n21984_, new_n21983_, new_n21972_ );
or   ( new_n21985_, new_n21984_, new_n21953_ );
and  ( new_n21986_, new_n21984_, new_n21953_ );
or   ( new_n21987_, new_n16119_, new_n6321_ );
or   ( new_n21988_, new_n16123_, new_n6307_ );
and  ( new_n21989_, new_n21988_, new_n21987_ );
or   ( new_n21990_, new_n21989_, new_n16108_ );
and  ( new_n21991_, new_n16132_, RI2b1c4342e278_94 );
and  ( new_n21992_, new_n16114_, RI2b1c4342e200_93 );
or   ( new_n21993_, new_n21992_, new_n21991_ );
or   ( new_n21994_, new_n21993_, new_n16128_ );
and  ( new_n21995_, new_n21994_, new_n21990_ );
or   ( new_n21996_, new_n16115_, new_n124_ );
and  ( new_n21997_, new_n21996_, new_n21995_ );
or   ( new_n21998_, new_n21997_, new_n21986_ );
and  ( new_n21999_, new_n21998_, new_n21985_ );
or   ( new_n22000_, new_n21999_, new_n21922_ );
and  ( new_n22001_, new_n21999_, new_n21922_ );
or   ( new_n22002_, new_n21730_, new_n21559_ );
or   ( new_n22003_, new_n21727_, new_n21568_ );
and  ( new_n22004_, new_n22003_, new_n22002_ );
or   ( new_n22005_, new_n22004_, new_n21735_ );
and  ( new_n22006_, new_n21731_, new_n21569_ );
or   ( new_n22007_, new_n22006_, new_n21579_ );
and  ( new_n22008_, new_n22007_, new_n22005_ );
or   ( new_n22009_, new_n22008_, new_n21740_ );
and  ( new_n22010_, new_n22008_, new_n21740_ );
or   ( new_n22011_, new_n21717_, new_n21528_ );
or   ( new_n22012_, new_n21714_, new_n21537_ );
and  ( new_n22013_, new_n22012_, new_n22011_ );
or   ( new_n22014_, new_n22013_, new_n21722_ );
and  ( new_n22015_, new_n21718_, new_n21538_ );
or   ( new_n22016_, new_n22015_, new_n21548_ );
and  ( new_n22017_, new_n22016_, new_n22014_ );
or   ( new_n22018_, new_n22017_, new_n22010_ );
and  ( new_n22019_, new_n22018_, new_n22009_ );
or   ( new_n22020_, new_n22019_, new_n22001_ );
and  ( new_n22021_, new_n22020_, new_n22000_ );
or   ( new_n22022_, new_n21766_, new_n21384_ );
or   ( new_n22023_, new_n21763_, new_n21391_ );
and  ( new_n22024_, new_n22023_, new_n22022_ );
or   ( new_n22025_, new_n22024_, new_n21771_ );
and  ( new_n22026_, new_n21767_, new_n21392_ );
or   ( new_n22027_, new_n22026_, new_n21400_ );
and  ( new_n22028_, new_n22027_, new_n22025_ );
or   ( new_n22029_, new_n21702_, new_n21495_ );
or   ( new_n22030_, new_n21699_, new_n21504_ );
and  ( new_n22031_, new_n22030_, new_n22029_ );
or   ( new_n22032_, new_n22031_, new_n21707_ );
and  ( new_n22033_, new_n21703_, new_n21505_ );
or   ( new_n22034_, new_n22033_, new_n21515_ );
and  ( new_n22035_, new_n22034_, new_n22032_ );
or   ( new_n22036_, new_n21687_, new_n21462_ );
or   ( new_n22037_, new_n21684_, new_n21471_ );
and  ( new_n22038_, new_n22037_, new_n22036_ );
or   ( new_n22039_, new_n22038_, new_n21692_ );
and  ( new_n22040_, new_n21688_, new_n21472_ );
or   ( new_n22041_, new_n22040_, new_n21482_ );
and  ( new_n22042_, new_n22041_, new_n22039_ );
or   ( new_n22043_, new_n22042_, new_n22035_ );
and  ( new_n22044_, new_n22042_, new_n22035_ );
or   ( new_n22045_, new_n21674_, new_n21431_ );
or   ( new_n22046_, new_n21671_, new_n21440_ );
and  ( new_n22047_, new_n22046_, new_n22045_ );
or   ( new_n22048_, new_n22047_, new_n21679_ );
and  ( new_n22049_, new_n21675_, new_n21441_ );
or   ( new_n22050_, new_n22049_, new_n21451_ );
and  ( new_n22051_, new_n22050_, new_n22048_ );
or   ( new_n22052_, new_n22051_, new_n22044_ );
and  ( new_n22053_, new_n22052_, new_n22043_ );
or   ( new_n22054_, new_n22053_, new_n22028_ );
and  ( new_n22055_, new_n22053_, new_n22028_ );
or   ( new_n22056_, new_n21748_, new_n21589_ );
or   ( new_n22057_, new_n21745_, new_n21596_ );
and  ( new_n22058_, new_n22057_, new_n22056_ );
or   ( new_n22059_, new_n22058_, new_n21753_ );
and  ( new_n22060_, new_n21749_, new_n21597_ );
or   ( new_n22061_, new_n22060_, new_n21605_ );
and  ( new_n22062_, new_n22061_, new_n22059_ );
or   ( new_n22063_, new_n22062_, new_n22055_ );
and  ( new_n22064_, new_n22063_, new_n22054_ );
or   ( new_n22065_, new_n22064_, new_n22021_ );
and  ( new_n22066_, new_n22064_, new_n22021_ );
or   ( new_n22067_, new_n21788_, new_n21618_ );
or   ( new_n22068_, new_n21785_, new_n21620_ );
and  ( new_n22069_, new_n22068_, new_n22067_ );
or   ( new_n22070_, new_n22069_, new_n21793_ );
and  ( new_n22071_, new_n21789_, new_n21621_ );
or   ( new_n22072_, new_n22071_, new_n21629_ );
and  ( new_n22073_, new_n22072_, new_n22070_ );
or   ( new_n22074_, new_n22073_, new_n22066_ );
and  ( new_n22075_, new_n22074_, new_n22065_ );
or   ( new_n22076_, new_n22075_, new_n21834_ );
or   ( new_n22077_, new_n21780_, new_n21609_ );
or   ( new_n22078_, new_n21757_, new_n21413_ );
and  ( new_n22079_, new_n22078_, new_n22077_ );
or   ( new_n22080_, new_n22079_, new_n21795_ );
and  ( new_n22081_, new_n21781_, new_n21611_ );
or   ( new_n22082_, new_n22081_, new_n21631_ );
and  ( new_n22083_, new_n22082_, new_n22080_ );
and  ( new_n22084_, new_n22075_, new_n21834_ );
or   ( new_n22085_, new_n22084_, new_n22083_ );
and  ( new_n22086_, new_n22085_, new_n22076_ );
or   ( new_n22087_, new_n22086_, new_n21827_ );
or   ( new_n22088_, new_n21810_, new_n21633_ );
or   ( new_n22089_, new_n21797_, new_n21370_ );
and  ( new_n22090_, new_n22089_, new_n22088_ );
or   ( new_n22091_, new_n22090_, new_n21815_ );
and  ( new_n22092_, new_n21811_, new_n21635_ );
or   ( new_n22093_, new_n22092_, new_n21642_ );
and  ( new_n22094_, new_n22093_, new_n22091_ );
and  ( new_n22095_, new_n22086_, new_n21827_ );
or   ( new_n22096_, new_n22095_, new_n22094_ );
and  ( new_n22097_, new_n22096_, new_n22087_ );
or   ( new_n22098_, new_n22097_, new_n21824_ );
and  ( new_n22099_, new_n22098_, new_n21657_ );
or   ( new_n22100_, new_n22099_, new_n21656_ );
and  ( new_n22101_, new_n22097_, new_n21824_ );
or   ( new_n22102_, new_n22101_, new_n21656_ );
or   ( new_n22103_, new_n22092_, new_n21815_ );
or   ( new_n22104_, new_n22090_, new_n21642_ );
and  ( new_n22105_, new_n22104_, new_n22103_ );
or   ( new_n22106_, new_n21666_, new_n21663_ );
and  ( new_n22107_, new_n22106_, new_n21345_ );
or   ( new_n22108_, new_n22107_, new_n22086_ );
or   ( new_n22109_, new_n21832_, new_n21808_ );
or   ( new_n22110_, new_n21830_, new_n21368_ );
and  ( new_n22111_, new_n22110_, new_n22109_ );
or   ( new_n22112_, new_n21929_, new_n16085_ );
or   ( new_n22113_, new_n21925_, new_n16048_ );
and  ( new_n22114_, new_n22113_, new_n22112_ );
or   ( new_n22115_, new_n21938_, new_n16052_ );
or   ( new_n22116_, new_n21934_, new_n16071_ );
and  ( new_n22117_, new_n22116_, new_n22115_ );
or   ( new_n22118_, new_n22117_, new_n22114_ );
and  ( new_n22119_, new_n22117_, new_n22114_ );
or   ( new_n22120_, new_n21949_, new_n16009_ );
or   ( new_n22121_, new_n21945_, new_n16029_ );
and  ( new_n22122_, new_n22121_, new_n22120_ );
or   ( new_n22123_, new_n22122_, new_n22119_ );
and  ( new_n22124_, new_n22123_, new_n22118_ );
or   ( new_n22125_, new_n21960_, new_n16186_ );
or   ( new_n22126_, new_n21956_, new_n16204_ );
and  ( new_n22127_, new_n22126_, new_n22125_ );
or   ( new_n22128_, new_n21969_, new_n16217_ );
or   ( new_n22129_, new_n21965_, new_n16234_ );
and  ( new_n22130_, new_n22129_, new_n22128_ );
or   ( new_n22131_, new_n22130_, new_n22127_ );
and  ( new_n22132_, new_n22130_, new_n22127_ );
or   ( new_n22133_, new_n21980_, new_n16151_ );
or   ( new_n22134_, new_n21976_, new_n16170_ );
and  ( new_n22135_, new_n22134_, new_n22133_ );
or   ( new_n22136_, new_n22135_, new_n22132_ );
and  ( new_n22137_, new_n22136_, new_n22131_ );
or   ( new_n22138_, new_n22137_, new_n22124_ );
and  ( new_n22139_, new_n22137_, new_n22124_ );
and  ( new_n22140_, new_n16102_, RI2b1c4342e2f0_95 );
or   ( new_n22141_, new_n21993_, new_n16108_ );
or   ( new_n22142_, new_n21989_, new_n16128_ );
and  ( new_n22143_, new_n22142_, new_n22141_ );
or   ( new_n22144_, new_n22143_, new_n22140_ );
or   ( new_n22145_, new_n22144_, new_n22139_ );
and  ( new_n22146_, new_n22145_, new_n22138_ );
or   ( new_n22147_, new_n21863_, new_n19394_ );
or   ( new_n22148_, new_n21859_, new_n19659_ );
and  ( new_n22149_, new_n22148_, new_n22147_ );
or   ( new_n22150_, new_n21872_, new_n18742_ );
or   ( new_n22151_, new_n21868_, new_n18977_ );
and  ( new_n22152_, new_n22151_, new_n22150_ );
or   ( new_n22153_, new_n22152_, new_n22149_ );
and  ( new_n22154_, new_n22152_, new_n22149_ );
or   ( new_n22155_, new_n21883_, new_n18066_ );
or   ( new_n22156_, new_n21879_, new_n18309_ );
and  ( new_n22157_, new_n22156_, new_n22155_ );
or   ( new_n22158_, new_n22157_, new_n22154_ );
and  ( new_n22159_, new_n22158_, new_n22153_ );
or   ( new_n22160_, new_n21841_, new_n21013_ );
or   ( new_n22161_, new_n21837_, new_n21265_ );
and  ( new_n22162_, new_n22161_, new_n22160_ );
or   ( new_n22163_, new_n22162_, new_n21009_ );
and  ( new_n22164_, new_n22162_, new_n21009_ );
or   ( new_n22165_, new_n21852_, new_n20156_ );
or   ( new_n22166_, new_n21848_, new_n20443_ );
and  ( new_n22167_, new_n22166_, new_n22165_ );
or   ( new_n22168_, new_n22167_, new_n22164_ );
and  ( new_n22169_, new_n22168_, new_n22163_ );
or   ( new_n22170_, new_n22169_, new_n22159_ );
and  ( new_n22171_, new_n22169_, new_n22159_ );
or   ( new_n22172_, new_n21896_, new_n17238_ );
or   ( new_n22173_, new_n21892_, new_n17650_ );
and  ( new_n22174_, new_n22173_, new_n22172_ );
or   ( new_n22175_, new_n21905_, new_n16814_ );
or   ( new_n22176_, new_n21901_, new_n17142_ );
and  ( new_n22177_, new_n22176_, new_n22175_ );
or   ( new_n22178_, new_n22177_, new_n22174_ );
and  ( new_n22179_, new_n22177_, new_n22174_ );
or   ( new_n22180_, new_n21916_, new_n16505_ );
or   ( new_n22181_, new_n21912_, new_n16438_ );
and  ( new_n22182_, new_n22181_, new_n22180_ );
or   ( new_n22183_, new_n22182_, new_n22179_ );
and  ( new_n22184_, new_n22183_, new_n22178_ );
or   ( new_n22185_, new_n22184_, new_n22171_ );
and  ( new_n22186_, new_n22185_, new_n22170_ );
or   ( new_n22187_, new_n22186_, new_n22146_ );
and  ( new_n22188_, new_n22186_, new_n22146_ );
or   ( new_n22189_, new_n22006_, new_n21735_ );
or   ( new_n22190_, new_n22004_, new_n21579_ );
and  ( new_n22191_, new_n22190_, new_n22189_ );
or   ( new_n22192_, new_n22191_, new_n21584_ );
and  ( new_n22193_, new_n22191_, new_n21584_ );
or   ( new_n22194_, new_n22015_, new_n21722_ );
or   ( new_n22195_, new_n22013_, new_n21548_ );
and  ( new_n22196_, new_n22195_, new_n22194_ );
or   ( new_n22197_, new_n22196_, new_n22193_ );
and  ( new_n22198_, new_n22197_, new_n22192_ );
or   ( new_n22199_, new_n22198_, new_n22188_ );
and  ( new_n22200_, new_n22199_, new_n22187_ );
or   ( new_n22201_, new_n22026_, new_n21771_ );
or   ( new_n22202_, new_n22024_, new_n21400_ );
and  ( new_n22203_, new_n22202_, new_n22201_ );
or   ( new_n22204_, new_n22033_, new_n21707_ );
or   ( new_n22205_, new_n22031_, new_n21515_ );
and  ( new_n22206_, new_n22205_, new_n22204_ );
or   ( new_n22207_, new_n22040_, new_n21692_ );
or   ( new_n22208_, new_n22038_, new_n21482_ );
and  ( new_n22209_, new_n22208_, new_n22207_ );
or   ( new_n22210_, new_n22209_, new_n22206_ );
and  ( new_n22211_, new_n22209_, new_n22206_ );
or   ( new_n22212_, new_n22049_, new_n21679_ );
or   ( new_n22213_, new_n22047_, new_n21451_ );
and  ( new_n22214_, new_n22213_, new_n22212_ );
or   ( new_n22215_, new_n22214_, new_n22211_ );
and  ( new_n22216_, new_n22215_, new_n22210_ );
or   ( new_n22217_, new_n22216_, new_n22203_ );
and  ( new_n22218_, new_n22216_, new_n22203_ );
or   ( new_n22219_, new_n22060_, new_n21753_ );
or   ( new_n22220_, new_n22058_, new_n21605_ );
and  ( new_n22221_, new_n22220_, new_n22219_ );
or   ( new_n22222_, new_n22221_, new_n22218_ );
and  ( new_n22223_, new_n22222_, new_n22217_ );
or   ( new_n22224_, new_n22223_, new_n22200_ );
and  ( new_n22225_, new_n22223_, new_n22200_ );
or   ( new_n22226_, new_n22071_, new_n21793_ );
or   ( new_n22227_, new_n22069_, new_n21629_ );
and  ( new_n22228_, new_n22227_, new_n22226_ );
or   ( new_n22229_, new_n22228_, new_n22225_ );
and  ( new_n22230_, new_n22229_, new_n22224_ );
or   ( new_n22231_, new_n22230_, new_n22111_ );
and  ( new_n22232_, new_n22230_, new_n22111_ );
or   ( new_n22233_, new_n22081_, new_n21795_ );
or   ( new_n22234_, new_n22079_, new_n21631_ );
and  ( new_n22235_, new_n22234_, new_n22233_ );
or   ( new_n22236_, new_n22235_, new_n22232_ );
and  ( new_n22237_, new_n22236_, new_n22231_ );
or   ( new_n22238_, new_n22237_, new_n21827_ );
and  ( new_n22239_, new_n22238_, new_n22108_ );
or   ( new_n22240_, new_n22239_, new_n22105_ );
or   ( new_n22241_, new_n22237_, new_n22107_ );
and  ( new_n22242_, new_n22241_, new_n22087_ );
or   ( new_n22243_, new_n22242_, new_n22094_ );
and  ( new_n22244_, new_n22243_, new_n22240_ );
or   ( new_n22245_, new_n21742_, new_n21519_ );
or   ( new_n22246_, new_n21711_, new_n21586_ );
and  ( new_n22247_, new_n22246_, new_n22245_ );
or   ( new_n22248_, new_n22247_, new_n21755_ );
and  ( new_n22249_, new_n21743_, new_n21588_ );
or   ( new_n22250_, new_n22249_, new_n21607_ );
and  ( new_n22251_, new_n22250_, new_n22248_ );
or   ( new_n22252_, new_n22223_, new_n22021_ );
or   ( new_n22253_, new_n22200_, new_n22064_ );
and  ( new_n22254_, new_n22253_, new_n22252_ );
or   ( new_n22255_, new_n22254_, new_n22228_ );
and  ( new_n22256_, new_n22224_, new_n22065_ );
or   ( new_n22257_, new_n22256_, new_n22073_ );
and  ( new_n22258_, new_n22257_, new_n22255_ );
or   ( new_n22259_, new_n22258_, new_n22251_ );
or   ( new_n22260_, new_n21694_, new_n21453_ );
or   ( new_n22261_, new_n21681_, new_n21484_ );
and  ( new_n22262_, new_n22261_, new_n22260_ );
or   ( new_n22263_, new_n22262_, new_n21709_ );
and  ( new_n22264_, new_n21695_, new_n21485_ );
or   ( new_n22265_, new_n22264_, new_n21517_ );
and  ( new_n22266_, new_n22265_, new_n22263_ );
or   ( new_n22267_, new_n22203_, new_n22053_ );
or   ( new_n22268_, new_n22216_, new_n22028_ );
and  ( new_n22269_, new_n22268_, new_n22267_ );
or   ( new_n22270_, new_n22269_, new_n22221_ );
and  ( new_n22271_, new_n22217_, new_n22054_ );
or   ( new_n22272_, new_n22271_, new_n22062_ );
and  ( new_n22273_, new_n22272_, new_n22270_ );
or   ( new_n22274_, new_n22273_, new_n22266_ );
and  ( new_n22275_, new_n22273_, new_n22266_ );
or   ( new_n22276_, new_n22146_, new_n21922_ );
or   ( new_n22277_, new_n22186_, new_n21999_ );
and  ( new_n22278_, new_n22277_, new_n22276_ );
or   ( new_n22279_, new_n22278_, new_n22198_ );
and  ( new_n22280_, new_n22187_, new_n22000_ );
or   ( new_n22281_, new_n22280_, new_n22019_ );
and  ( new_n22282_, new_n22281_, new_n22279_ );
or   ( new_n22283_, new_n22282_, new_n22275_ );
and  ( new_n22284_, new_n22283_, new_n22274_ );
or   ( new_n22285_, new_n22209_, new_n22035_ );
or   ( new_n22286_, new_n22206_, new_n22042_ );
and  ( new_n22287_, new_n22286_, new_n22285_ );
or   ( new_n22288_, new_n22287_, new_n22214_ );
and  ( new_n22289_, new_n22210_, new_n22043_ );
or   ( new_n22290_, new_n22289_, new_n22051_ );
and  ( new_n22291_, new_n22290_, new_n22288_ );
or   ( new_n22292_, new_n22177_, new_n21898_ );
or   ( new_n22293_, new_n22174_, new_n21907_ );
and  ( new_n22294_, new_n22293_, new_n22292_ );
or   ( new_n22295_, new_n22294_, new_n22182_ );
and  ( new_n22296_, new_n22178_, new_n21908_ );
or   ( new_n22297_, new_n22296_, new_n21918_ );
and  ( new_n22298_, new_n22297_, new_n22295_ );
or   ( new_n22299_, new_n22152_, new_n21865_ );
or   ( new_n22300_, new_n22149_, new_n21874_ );
and  ( new_n22301_, new_n22300_, new_n22299_ );
or   ( new_n22302_, new_n22301_, new_n22157_ );
and  ( new_n22303_, new_n22153_, new_n21875_ );
or   ( new_n22304_, new_n22303_, new_n21885_ );
and  ( new_n22305_, new_n22304_, new_n22302_ );
or   ( new_n22306_, new_n22305_, new_n22298_ );
and  ( new_n22307_, new_n22305_, new_n22298_ );
or   ( new_n22308_, new_n22162_, new_n21261_ );
or   ( new_n22309_, new_n21843_, new_n21009_ );
and  ( new_n22310_, new_n22309_, new_n22308_ );
or   ( new_n22311_, new_n22310_, new_n22167_ );
and  ( new_n22312_, new_n22163_, new_n21844_ );
or   ( new_n22313_, new_n22312_, new_n21854_ );
and  ( new_n22314_, new_n22313_, new_n22311_ );
or   ( new_n22315_, new_n22314_, new_n22307_ );
and  ( new_n22316_, new_n22315_, new_n22306_ );
or   ( new_n22317_, new_n22316_, new_n22291_ );
and  ( new_n22318_, new_n22316_, new_n22291_ );
or   ( new_n22319_, new_n22191_, new_n21740_ );
or   ( new_n22320_, new_n22008_, new_n21584_ );
and  ( new_n22321_, new_n22320_, new_n22319_ );
or   ( new_n22322_, new_n22321_, new_n22196_ );
and  ( new_n22323_, new_n22192_, new_n22009_ );
or   ( new_n22324_, new_n22323_, new_n22017_ );
and  ( new_n22325_, new_n22324_, new_n22322_ );
or   ( new_n22326_, new_n22325_, new_n22318_ );
and  ( new_n22327_, new_n22326_, new_n22317_ );
xor  ( new_n22328_, RI2b1c4342c568_32, RI2b1c4342d468_64 );
or   ( new_n22329_, new_n22328_, new_n137_ );
and  ( new_n22330_, new_n22329_, new_n7097_ );
or   ( new_n22331_, new_n21261_, new_n15246_ );
and  ( new_n22332_, new_n22331_, new_n21009_ );
or   ( new_n22333_, new_n22332_, new_n22330_ );
or   ( new_n22334_, new_n22333_, new_n99_ );
or   ( new_n22335_, new_n22334_, new_n21261_ );
or   ( new_n22336_, new_n22330_, new_n21261_ );
and  ( new_n22337_, new_n22336_, new_n15246_ );
and  ( new_n22338_, new_n22337_, RI2b1c4342d4e0_65 );
or   ( new_n22339_, new_n22338_, new_n21009_ );
and  ( new_n22340_, new_n22339_, new_n22335_ );
or   ( new_n22341_, new_n21419_, new_n112_ );
or   ( new_n22342_, new_n21424_, new_n526_ );
and  ( new_n22343_, new_n22342_, new_n22341_ );
or   ( new_n22344_, new_n22343_, new_n21013_ );
and  ( new_n22345_, new_n21428_, RI2b1c4342d5d0_67 );
and  ( new_n22346_, new_n21415_, RI2b1c4342d558_66 );
or   ( new_n22347_, new_n22346_, new_n22345_ );
or   ( new_n22348_, new_n22347_, new_n21265_ );
and  ( new_n22349_, new_n22348_, new_n22344_ );
or   ( new_n22350_, new_n22349_, new_n22340_ );
or   ( new_n22351_, new_n20557_, new_n591_ );
or   ( new_n22352_, new_n20562_, new_n612_ );
and  ( new_n22353_, new_n22352_, new_n22351_ );
or   ( new_n22354_, new_n22353_, new_n20156_ );
and  ( new_n22355_, new_n20566_, RI2b1c4342d6c0_69 );
and  ( new_n22356_, new_n20553_, RI2b1c4342d648_68 );
or   ( new_n22357_, new_n22356_, new_n22355_ );
or   ( new_n22358_, new_n22357_, new_n20443_ );
and  ( new_n22359_, new_n22358_, new_n22354_ );
or   ( new_n22360_, new_n19758_, new_n110_ );
or   ( new_n22361_, new_n19763_, new_n755_ );
and  ( new_n22362_, new_n22361_, new_n22360_ );
or   ( new_n22363_, new_n22362_, new_n19394_ );
and  ( new_n22364_, new_n19767_, RI2b1c4342d7b0_71 );
and  ( new_n22365_, new_n19754_, RI2b1c4342d738_70 );
or   ( new_n22366_, new_n22365_, new_n22364_ );
or   ( new_n22367_, new_n22366_, new_n19659_ );
and  ( new_n22368_, new_n22367_, new_n22363_ );
or   ( new_n22369_, new_n22368_, new_n22359_ );
and  ( new_n22370_, new_n22368_, new_n22359_ );
or   ( new_n22371_, new_n19048_, new_n105_ );
or   ( new_n22372_, new_n19055_, new_n806_ );
and  ( new_n22373_, new_n22372_, new_n22371_ );
or   ( new_n22374_, new_n22373_, new_n18742_ );
and  ( new_n22375_, new_n19057_, RI2b1c4342d8a0_73 );
and  ( new_n22376_, new_n19044_, RI2b1c4342d828_72 );
or   ( new_n22377_, new_n22376_, new_n22375_ );
or   ( new_n22378_, new_n22377_, new_n18977_ );
and  ( new_n22379_, new_n22378_, new_n22374_ );
or   ( new_n22380_, new_n22379_, new_n22370_ );
and  ( new_n22381_, new_n22380_, new_n22369_ );
or   ( new_n22382_, new_n22381_, new_n22350_ );
and  ( new_n22383_, new_n22381_, new_n22350_ );
or   ( new_n22384_, new_n18388_, new_n843_ );
or   ( new_n22385_, new_n18395_, new_n859_ );
and  ( new_n22386_, new_n22385_, new_n22384_ );
or   ( new_n22387_, new_n22386_, new_n18066_ );
and  ( new_n22388_, new_n18397_, RI2b1c4342d990_75 );
and  ( new_n22389_, new_n18384_, RI2b1c4342d918_74 );
or   ( new_n22390_, new_n22389_, new_n22388_ );
or   ( new_n22391_, new_n22390_, new_n18309_ );
and  ( new_n22392_, new_n22391_, new_n22387_ );
or   ( new_n22393_, new_n17727_, new_n1004_ );
or   ( new_n22394_, new_n17734_, new_n886_ );
and  ( new_n22395_, new_n22394_, new_n22393_ );
or   ( new_n22396_, new_n22395_, new_n17238_ );
and  ( new_n22397_, new_n17736_, RI2b1c4342da80_77 );
and  ( new_n22398_, new_n17723_, RI2b1c4342da08_76 );
or   ( new_n22399_, new_n22398_, new_n22397_ );
or   ( new_n22400_, new_n22399_, new_n17650_ );
and  ( new_n22401_, new_n22400_, new_n22396_ );
or   ( new_n22402_, new_n22401_, new_n22392_ );
and  ( new_n22403_, new_n22401_, new_n22392_ );
or   ( new_n22404_, new_n17244_, new_n1310_ );
or   ( new_n22405_, new_n17248_, new_n1002_ );
and  ( new_n22406_, new_n22405_, new_n22404_ );
or   ( new_n22407_, new_n22406_, new_n16814_ );
and  ( new_n22408_, new_n17255_, RI2b1c4342db70_79 );
and  ( new_n22409_, new_n17240_, RI2b1c4342daf8_78 );
or   ( new_n22410_, new_n22409_, new_n22408_ );
or   ( new_n22411_, new_n22410_, new_n17142_ );
and  ( new_n22412_, new_n22411_, new_n22407_ );
or   ( new_n22413_, new_n22412_, new_n22403_ );
and  ( new_n22414_, new_n22413_, new_n22402_ );
or   ( new_n22415_, new_n22414_, new_n22383_ );
and  ( new_n22416_, new_n22415_, new_n22382_ );
or   ( new_n22417_, new_n16607_, new_n126_ );
or   ( new_n22418_, new_n16613_, new_n1511_ );
and  ( new_n22419_, new_n22418_, new_n22417_ );
or   ( new_n22420_, new_n22419_, new_n16505_ );
and  ( new_n22421_, new_n16616_, RI2b1c4342dc60_81 );
and  ( new_n22422_, new_n16603_, RI2b1c4342dbe8_80 );
or   ( new_n22423_, new_n22422_, new_n22421_ );
or   ( new_n22424_, new_n22423_, new_n16438_ );
and  ( new_n22425_, new_n22424_, new_n22420_ );
or   ( new_n22426_, new_n16366_, new_n121_ );
or   ( new_n22427_, new_n16355_, new_n2119_ );
and  ( new_n22428_, new_n22427_, new_n22426_ );
or   ( new_n22429_, new_n22428_, new_n16085_ );
and  ( new_n22430_, new_n16358_, RI2b1c4342dd50_83 );
and  ( new_n22431_, new_n16362_, RI2b1c4342dcd8_82 );
or   ( new_n22432_, new_n22431_, new_n22430_ );
or   ( new_n22433_, new_n22432_, new_n16048_ );
and  ( new_n22434_, new_n22433_, new_n22429_ );
or   ( new_n22435_, new_n22434_, new_n22425_ );
and  ( new_n22436_, new_n22434_, new_n22425_ );
or   ( new_n22437_, new_n16075_, new_n2806_ );
or   ( new_n22438_, new_n16060_, new_n2541_ );
and  ( new_n22439_, new_n22438_, new_n22437_ );
or   ( new_n22440_, new_n22439_, new_n16052_ );
and  ( new_n22441_, new_n16063_, RI2b1c4342de40_85 );
and  ( new_n22442_, new_n16066_, RI2b1c4342ddc8_84 );
or   ( new_n22443_, new_n22442_, new_n22441_ );
or   ( new_n22444_, new_n22443_, new_n16071_ );
and  ( new_n22445_, new_n22444_, new_n22440_ );
or   ( new_n22446_, new_n22445_, new_n22436_ );
and  ( new_n22447_, new_n22446_, new_n22435_ );
or   ( new_n22448_, new_n16033_, new_n3924_ );
or   ( new_n22449_, new_n16017_, new_n3239_ );
and  ( new_n22450_, new_n22449_, new_n22448_ );
or   ( new_n22451_, new_n22450_, new_n16009_ );
and  ( new_n22452_, new_n16021_, RI2b1c4342df30_87 );
and  ( new_n22453_, new_n16024_, RI2b1c4342deb8_86 );
or   ( new_n22454_, new_n22453_, new_n22452_ );
or   ( new_n22455_, new_n22454_, new_n16029_ );
and  ( new_n22456_, new_n22455_, new_n22451_ );
or   ( new_n22457_, new_n16208_, new_n132_ );
or   ( new_n22458_, new_n16194_, new_n3902_ );
and  ( new_n22459_, new_n22458_, new_n22457_ );
or   ( new_n22460_, new_n22459_, new_n16186_ );
and  ( new_n22461_, new_n16196_, RI2b1c4342e020_89 );
and  ( new_n22462_, new_n16199_, RI2b1c4342dfa8_88 );
or   ( new_n22463_, new_n22462_, new_n22461_ );
or   ( new_n22464_, new_n22463_, new_n16204_ );
and  ( new_n22465_, new_n22464_, new_n22460_ );
or   ( new_n22466_, new_n22465_, new_n22456_ );
and  ( new_n22467_, new_n22465_, new_n22456_ );
or   ( new_n22468_, new_n16238_, new_n117_ );
or   ( new_n22469_, new_n16224_, new_n4635_ );
and  ( new_n22470_, new_n22469_, new_n22468_ );
or   ( new_n22471_, new_n22470_, new_n16217_ );
and  ( new_n22472_, new_n16226_, RI2b1c4342e110_91 );
and  ( new_n22473_, new_n16229_, RI2b1c4342e098_90 );
or   ( new_n22474_, new_n22473_, new_n22472_ );
or   ( new_n22475_, new_n22474_, new_n16234_ );
and  ( new_n22476_, new_n22475_, new_n22471_ );
or   ( new_n22477_, new_n22476_, new_n22467_ );
and  ( new_n22478_, new_n22477_, new_n22466_ );
and  ( new_n22479_, new_n22478_, new_n22447_ );
or   ( new_n22480_, new_n22478_, new_n22447_ );
or   ( new_n22481_, new_n16174_, new_n6307_ );
or   ( new_n22482_, new_n16160_, new_n5459_ );
and  ( new_n22483_, new_n22482_, new_n22481_ );
or   ( new_n22484_, new_n22483_, new_n16151_ );
and  ( new_n22485_, new_n16162_, RI2b1c4342e200_93 );
and  ( new_n22486_, new_n16165_, RI2b1c4342e188_92 );
or   ( new_n22487_, new_n22486_, new_n22485_ );
or   ( new_n22488_, new_n22487_, new_n16170_ );
and  ( new_n22489_, new_n22488_, new_n22484_ );
or   ( new_n22490_, new_n16119_, new_n124_ );
or   ( new_n22491_, new_n16123_, new_n6321_ );
and  ( new_n22492_, new_n22491_, new_n22490_ );
or   ( new_n22493_, new_n22492_, new_n16108_ );
and  ( new_n22494_, new_n16132_, RI2b1c4342e2f0_95 );
and  ( new_n22495_, new_n16114_, RI2b1c4342e278_94 );
or   ( new_n22496_, new_n22495_, new_n22494_ );
or   ( new_n22497_, new_n22496_, new_n16128_ );
and  ( new_n22498_, new_n22497_, new_n22493_ );
and  ( new_n22499_, new_n22498_, new_n22489_ );
or   ( new_n22500_, new_n22498_, new_n22489_ );
or   ( new_n22501_, new_n16115_, new_n7274_ );
and  ( new_n22502_, new_n22501_, new_n22500_ );
or   ( new_n22503_, new_n22502_, new_n22499_ );
and  ( new_n22504_, new_n22503_, new_n22480_ );
or   ( new_n22505_, new_n22504_, new_n22479_ );
and  ( new_n22506_, new_n22505_, new_n22416_ );
or   ( new_n22507_, new_n22505_, new_n22416_ );
or   ( new_n22508_, new_n21996_, new_n21995_ );
and  ( new_n22509_, new_n22508_, new_n22144_ );
or   ( new_n22510_, new_n22130_, new_n21962_ );
or   ( new_n22511_, new_n22127_, new_n21971_ );
and  ( new_n22512_, new_n22511_, new_n22510_ );
or   ( new_n22513_, new_n22512_, new_n22135_ );
and  ( new_n22514_, new_n22131_, new_n21972_ );
or   ( new_n22515_, new_n22514_, new_n21982_ );
and  ( new_n22516_, new_n22515_, new_n22513_ );
or   ( new_n22517_, new_n22516_, new_n22509_ );
and  ( new_n22518_, new_n22516_, new_n22509_ );
or   ( new_n22519_, new_n22117_, new_n21931_ );
or   ( new_n22520_, new_n22114_, new_n21940_ );
and  ( new_n22521_, new_n22520_, new_n22519_ );
or   ( new_n22522_, new_n22521_, new_n22122_ );
and  ( new_n22523_, new_n22118_, new_n21941_ );
or   ( new_n22524_, new_n22523_, new_n21951_ );
and  ( new_n22525_, new_n22524_, new_n22522_ );
or   ( new_n22526_, new_n22525_, new_n22518_ );
and  ( new_n22527_, new_n22526_, new_n22517_ );
and  ( new_n22528_, new_n22527_, new_n22507_ );
or   ( new_n22529_, new_n22528_, new_n22506_ );
and  ( new_n22530_, new_n22529_, new_n22327_ );
or   ( new_n22531_, new_n22529_, new_n22327_ );
or   ( new_n22532_, new_n21737_, new_n21550_ );
or   ( new_n22533_, new_n21724_, new_n21581_ );
and  ( new_n22534_, new_n22533_, new_n22532_ );
or   ( new_n22535_, new_n22534_, new_n21740_ );
and  ( new_n22536_, new_n21738_, new_n21583_ );
or   ( new_n22537_, new_n22536_, new_n21584_ );
and  ( new_n22538_, new_n22537_, new_n22535_ );
and  ( new_n22539_, new_n22538_, new_n22531_ );
or   ( new_n22540_, new_n22539_, new_n22530_ );
and  ( new_n22541_, new_n22540_, new_n22284_ );
or   ( new_n22542_, new_n22540_, new_n22284_ );
or   ( new_n22543_, new_n21760_, new_n21402_ );
or   ( new_n22544_, new_n21773_, new_n21377_ );
and  ( new_n22545_, new_n22544_, new_n22543_ );
or   ( new_n22546_, new_n22545_, new_n21778_ );
and  ( new_n22547_, new_n21774_, new_n21403_ );
or   ( new_n22548_, new_n22547_, new_n21411_ );
and  ( new_n22549_, new_n22548_, new_n22546_ );
and  ( new_n22550_, new_n22549_, new_n22542_ );
or   ( new_n22551_, new_n22550_, new_n22541_ );
and  ( new_n22552_, new_n22551_, new_n22259_ );
or   ( new_n22553_, new_n22551_, new_n22259_ );
or   ( new_n22554_, new_n22111_, new_n22075_ );
or   ( new_n22555_, new_n22230_, new_n21834_ );
and  ( new_n22556_, new_n22555_, new_n22554_ );
or   ( new_n22557_, new_n22556_, new_n22235_ );
and  ( new_n22558_, new_n22231_, new_n22076_ );
or   ( new_n22559_, new_n22558_, new_n22083_ );
and  ( new_n22560_, new_n22559_, new_n22557_ );
and  ( new_n22561_, new_n22560_, new_n22553_ );
or   ( new_n22562_, new_n22561_, new_n22552_ );
and  ( new_n22563_, new_n22562_, new_n22244_ );
or   ( new_n22564_, new_n22562_, new_n22244_ );
or   ( new_n22565_, new_n22558_, new_n22235_ );
or   ( new_n22566_, new_n22556_, new_n22083_ );
and  ( new_n22567_, new_n22566_, new_n22565_ );
or   ( new_n22568_, new_n22249_, new_n21755_ );
or   ( new_n22569_, new_n22247_, new_n21607_ );
and  ( new_n22570_, new_n22569_, new_n22568_ );
or   ( new_n22571_, new_n22256_, new_n22228_ );
or   ( new_n22572_, new_n22254_, new_n22073_ );
and  ( new_n22573_, new_n22572_, new_n22571_ );
and  ( new_n22574_, new_n22573_, new_n22570_ );
or   ( new_n22575_, new_n22574_, new_n22551_ );
or   ( new_n22576_, new_n22338_, new_n21261_ );
or   ( new_n22577_, new_n22334_, new_n21009_ );
and  ( new_n22578_, new_n22577_, new_n22576_ );
or   ( new_n22579_, new_n22347_, new_n21013_ );
or   ( new_n22580_, new_n22343_, new_n21265_ );
and  ( new_n22581_, new_n22580_, new_n22579_ );
and  ( new_n22582_, new_n22581_, new_n22578_ );
or   ( new_n22583_, new_n22357_, new_n20156_ );
or   ( new_n22584_, new_n22353_, new_n20443_ );
and  ( new_n22585_, new_n22584_, new_n22583_ );
or   ( new_n22586_, new_n22366_, new_n19394_ );
or   ( new_n22587_, new_n22362_, new_n19659_ );
and  ( new_n22588_, new_n22587_, new_n22586_ );
or   ( new_n22589_, new_n22588_, new_n22585_ );
and  ( new_n22590_, new_n22588_, new_n22585_ );
or   ( new_n22591_, new_n22377_, new_n18742_ );
or   ( new_n22592_, new_n22373_, new_n18977_ );
and  ( new_n22593_, new_n22592_, new_n22591_ );
or   ( new_n22594_, new_n22593_, new_n22590_ );
and  ( new_n22595_, new_n22594_, new_n22589_ );
or   ( new_n22596_, new_n22595_, new_n22582_ );
and  ( new_n22597_, new_n22595_, new_n22582_ );
or   ( new_n22598_, new_n22390_, new_n18066_ );
or   ( new_n22599_, new_n22386_, new_n18309_ );
and  ( new_n22600_, new_n22599_, new_n22598_ );
or   ( new_n22601_, new_n22399_, new_n17238_ );
or   ( new_n22602_, new_n22395_, new_n17650_ );
and  ( new_n22603_, new_n22602_, new_n22601_ );
or   ( new_n22604_, new_n22603_, new_n22600_ );
and  ( new_n22605_, new_n22603_, new_n22600_ );
or   ( new_n22606_, new_n22410_, new_n16814_ );
or   ( new_n22607_, new_n22406_, new_n17142_ );
and  ( new_n22608_, new_n22607_, new_n22606_ );
or   ( new_n22609_, new_n22608_, new_n22605_ );
and  ( new_n22610_, new_n22609_, new_n22604_ );
or   ( new_n22611_, new_n22610_, new_n22597_ );
and  ( new_n22612_, new_n22611_, new_n22596_ );
or   ( new_n22613_, new_n22423_, new_n16505_ );
or   ( new_n22614_, new_n22419_, new_n16438_ );
and  ( new_n22615_, new_n22614_, new_n22613_ );
or   ( new_n22616_, new_n22432_, new_n16085_ );
or   ( new_n22617_, new_n22428_, new_n16048_ );
and  ( new_n22618_, new_n22617_, new_n22616_ );
or   ( new_n22619_, new_n22618_, new_n22615_ );
and  ( new_n22620_, new_n22618_, new_n22615_ );
or   ( new_n22621_, new_n22443_, new_n16052_ );
or   ( new_n22622_, new_n22439_, new_n16071_ );
and  ( new_n22623_, new_n22622_, new_n22621_ );
or   ( new_n22624_, new_n22623_, new_n22620_ );
and  ( new_n22625_, new_n22624_, new_n22619_ );
or   ( new_n22626_, new_n22454_, new_n16009_ );
or   ( new_n22627_, new_n22450_, new_n16029_ );
and  ( new_n22628_, new_n22627_, new_n22626_ );
or   ( new_n22629_, new_n22463_, new_n16186_ );
or   ( new_n22630_, new_n22459_, new_n16204_ );
and  ( new_n22631_, new_n22630_, new_n22629_ );
or   ( new_n22632_, new_n22631_, new_n22628_ );
and  ( new_n22633_, new_n22631_, new_n22628_ );
or   ( new_n22634_, new_n22474_, new_n16217_ );
or   ( new_n22635_, new_n22470_, new_n16234_ );
and  ( new_n22636_, new_n22635_, new_n22634_ );
or   ( new_n22637_, new_n22636_, new_n22633_ );
and  ( new_n22638_, new_n22637_, new_n22632_ );
or   ( new_n22639_, new_n22638_, new_n22625_ );
and  ( new_n22640_, new_n22638_, new_n22625_ );
or   ( new_n22641_, new_n22487_, new_n16151_ );
or   ( new_n22642_, new_n22483_, new_n16170_ );
and  ( new_n22643_, new_n22642_, new_n22641_ );
or   ( new_n22644_, new_n22496_, new_n16108_ );
or   ( new_n22645_, new_n22492_, new_n16128_ );
and  ( new_n22646_, new_n22645_, new_n22644_ );
or   ( new_n22647_, new_n22646_, new_n22643_ );
and  ( new_n22648_, new_n22646_, new_n22643_ );
and  ( new_n22649_, new_n16102_, RI2b1c4342e368_96 );
or   ( new_n22650_, new_n22649_, new_n22648_ );
and  ( new_n22651_, new_n22650_, new_n22647_ );
or   ( new_n22652_, new_n22651_, new_n22640_ );
and  ( new_n22653_, new_n22652_, new_n22639_ );
or   ( new_n22654_, new_n22653_, new_n22612_ );
and  ( new_n22655_, new_n22653_, new_n22612_ );
or   ( new_n22656_, new_n22140_, new_n21995_ );
or   ( new_n22657_, new_n22143_, new_n21996_ );
and  ( new_n22658_, new_n22657_, new_n22656_ );
or   ( new_n22659_, new_n22514_, new_n22135_ );
or   ( new_n22660_, new_n22512_, new_n21982_ );
and  ( new_n22661_, new_n22660_, new_n22659_ );
or   ( new_n22662_, new_n22661_, new_n22658_ );
and  ( new_n22663_, new_n22661_, new_n22658_ );
or   ( new_n22664_, new_n22523_, new_n22122_ );
or   ( new_n22665_, new_n22521_, new_n21951_ );
and  ( new_n22666_, new_n22665_, new_n22664_ );
or   ( new_n22667_, new_n22666_, new_n22663_ );
and  ( new_n22668_, new_n22667_, new_n22662_ );
or   ( new_n22669_, new_n22668_, new_n22655_ );
and  ( new_n22670_, new_n22669_, new_n22654_ );
or   ( new_n22671_, new_n22289_, new_n22214_ );
or   ( new_n22672_, new_n22287_, new_n22051_ );
and  ( new_n22673_, new_n22672_, new_n22671_ );
or   ( new_n22674_, new_n22296_, new_n22182_ );
or   ( new_n22675_, new_n22294_, new_n21918_ );
and  ( new_n22676_, new_n22675_, new_n22674_ );
or   ( new_n22677_, new_n22303_, new_n22157_ );
or   ( new_n22678_, new_n22301_, new_n21885_ );
and  ( new_n22679_, new_n22678_, new_n22677_ );
or   ( new_n22680_, new_n22679_, new_n22676_ );
and  ( new_n22681_, new_n22679_, new_n22676_ );
or   ( new_n22682_, new_n22312_, new_n22167_ );
or   ( new_n22683_, new_n22310_, new_n21854_ );
and  ( new_n22684_, new_n22683_, new_n22682_ );
or   ( new_n22685_, new_n22684_, new_n22681_ );
and  ( new_n22686_, new_n22685_, new_n22680_ );
or   ( new_n22687_, new_n22686_, new_n22673_ );
and  ( new_n22688_, new_n22686_, new_n22673_ );
or   ( new_n22689_, new_n22323_, new_n22196_ );
or   ( new_n22690_, new_n22321_, new_n22017_ );
and  ( new_n22691_, new_n22690_, new_n22689_ );
or   ( new_n22692_, new_n22691_, new_n22688_ );
and  ( new_n22693_, new_n22692_, new_n22687_ );
or   ( new_n22694_, new_n22693_, new_n22670_ );
and  ( new_n22695_, new_n22693_, new_n22670_ );
or   ( new_n22696_, new_n22536_, new_n21740_ );
or   ( new_n22697_, new_n22534_, new_n21584_ );
and  ( new_n22698_, new_n22697_, new_n22696_ );
or   ( new_n22699_, new_n22698_, new_n22695_ );
and  ( new_n22700_, new_n22699_, new_n22694_ );
or   ( new_n22701_, new_n22264_, new_n21709_ );
or   ( new_n22702_, new_n22262_, new_n21517_ );
and  ( new_n22703_, new_n22702_, new_n22701_ );
or   ( new_n22704_, new_n22271_, new_n22221_ );
or   ( new_n22705_, new_n22269_, new_n22062_ );
and  ( new_n22706_, new_n22705_, new_n22704_ );
or   ( new_n22707_, new_n22706_, new_n22703_ );
and  ( new_n22708_, new_n22706_, new_n22703_ );
or   ( new_n22709_, new_n22280_, new_n22198_ );
or   ( new_n22710_, new_n22278_, new_n22019_ );
and  ( new_n22711_, new_n22710_, new_n22709_ );
or   ( new_n22712_, new_n22711_, new_n22708_ );
and  ( new_n22713_, new_n22712_, new_n22707_ );
or   ( new_n22714_, new_n22713_, new_n22700_ );
and  ( new_n22715_, new_n22713_, new_n22700_ );
or   ( new_n22716_, new_n22547_, new_n21778_ );
or   ( new_n22717_, new_n22545_, new_n21411_ );
and  ( new_n22718_, new_n22717_, new_n22716_ );
or   ( new_n22719_, new_n22718_, new_n22715_ );
and  ( new_n22720_, new_n22719_, new_n22714_ );
or   ( new_n22721_, new_n22720_, new_n22259_ );
and  ( new_n22722_, new_n22721_, new_n22575_ );
or   ( new_n22723_, new_n22722_, new_n22567_ );
or   ( new_n22724_, new_n22720_, new_n22574_ );
and  ( new_n22725_, new_n22724_, new_n22553_ );
or   ( new_n22726_, new_n22725_, new_n22560_ );
and  ( new_n22727_, new_n22726_, new_n22723_ );
or   ( new_n22728_, new_n22573_, new_n22251_ );
or   ( new_n22729_, new_n22570_, new_n22258_ );
and  ( new_n22730_, new_n22729_, new_n22728_ );
nor  ( new_n22731_, new_n22333_, new_n526_ );
nor  ( new_n22732_, new_n22731_, new_n7601_ );
or   ( new_n22733_, new_n22732_, new_n21261_ );
and  ( new_n22734_, new_n22337_, RI2b1c4342d558_66 );
and  ( new_n22735_, new_n22330_, RI2b1c4342d4e0_65 );
or   ( new_n22736_, new_n22735_, new_n22734_ );
or   ( new_n22737_, new_n22736_, new_n21009_ );
and  ( new_n22738_, new_n22737_, new_n22733_ );
or   ( new_n22739_, new_n21419_, new_n612_ );
or   ( new_n22740_, new_n21424_, new_n112_ );
and  ( new_n22741_, new_n22740_, new_n22739_ );
or   ( new_n22742_, new_n22741_, new_n21013_ );
and  ( new_n22743_, new_n21428_, RI2b1c4342d648_68 );
and  ( new_n22744_, new_n21415_, RI2b1c4342d5d0_67 );
or   ( new_n22745_, new_n22744_, new_n22743_ );
or   ( new_n22746_, new_n22745_, new_n21265_ );
and  ( new_n22747_, new_n22746_, new_n22742_ );
or   ( new_n22748_, new_n22747_, new_n22738_ );
and  ( new_n22749_, new_n22747_, new_n22738_ );
or   ( new_n22750_, new_n20557_, new_n755_ );
or   ( new_n22751_, new_n20562_, new_n591_ );
and  ( new_n22752_, new_n22751_, new_n22750_ );
or   ( new_n22753_, new_n22752_, new_n20156_ );
and  ( new_n22754_, new_n20566_, RI2b1c4342d738_70 );
and  ( new_n22755_, new_n20553_, RI2b1c4342d6c0_69 );
or   ( new_n22756_, new_n22755_, new_n22754_ );
or   ( new_n22757_, new_n22756_, new_n20443_ );
and  ( new_n22758_, new_n22757_, new_n22753_ );
or   ( new_n22759_, new_n22758_, new_n22749_ );
and  ( new_n22760_, new_n22759_, new_n22748_ );
or   ( new_n22761_, new_n19758_, new_n806_ );
or   ( new_n22762_, new_n19763_, new_n110_ );
and  ( new_n22763_, new_n22762_, new_n22761_ );
or   ( new_n22764_, new_n22763_, new_n19394_ );
and  ( new_n22765_, new_n19767_, RI2b1c4342d828_72 );
and  ( new_n22766_, new_n19754_, RI2b1c4342d7b0_71 );
or   ( new_n22767_, new_n22766_, new_n22765_ );
or   ( new_n22768_, new_n22767_, new_n19659_ );
and  ( new_n22769_, new_n22768_, new_n22764_ );
or   ( new_n22770_, new_n19048_, new_n859_ );
or   ( new_n22771_, new_n19055_, new_n105_ );
and  ( new_n22772_, new_n22771_, new_n22770_ );
or   ( new_n22773_, new_n22772_, new_n18742_ );
and  ( new_n22774_, new_n19057_, RI2b1c4342d918_74 );
and  ( new_n22775_, new_n19044_, RI2b1c4342d8a0_73 );
or   ( new_n22776_, new_n22775_, new_n22774_ );
or   ( new_n22777_, new_n22776_, new_n18977_ );
and  ( new_n22778_, new_n22777_, new_n22773_ );
or   ( new_n22779_, new_n22778_, new_n22769_ );
and  ( new_n22780_, new_n22778_, new_n22769_ );
or   ( new_n22781_, new_n18388_, new_n886_ );
or   ( new_n22782_, new_n18395_, new_n843_ );
and  ( new_n22783_, new_n22782_, new_n22781_ );
or   ( new_n22784_, new_n22783_, new_n18066_ );
and  ( new_n22785_, new_n18397_, RI2b1c4342da08_76 );
and  ( new_n22786_, new_n18384_, RI2b1c4342d990_75 );
or   ( new_n22787_, new_n22786_, new_n22785_ );
or   ( new_n22788_, new_n22787_, new_n18309_ );
and  ( new_n22789_, new_n22788_, new_n22784_ );
or   ( new_n22790_, new_n22789_, new_n22780_ );
and  ( new_n22791_, new_n22790_, new_n22779_ );
or   ( new_n22792_, new_n22791_, new_n22760_ );
and  ( new_n22793_, new_n22791_, new_n22760_ );
or   ( new_n22794_, new_n17727_, new_n1002_ );
or   ( new_n22795_, new_n17734_, new_n1004_ );
and  ( new_n22796_, new_n22795_, new_n22794_ );
or   ( new_n22797_, new_n22796_, new_n17238_ );
and  ( new_n22798_, new_n17736_, RI2b1c4342daf8_78 );
and  ( new_n22799_, new_n17723_, RI2b1c4342da80_77 );
or   ( new_n22800_, new_n22799_, new_n22798_ );
or   ( new_n22801_, new_n22800_, new_n17650_ );
and  ( new_n22802_, new_n22801_, new_n22797_ );
or   ( new_n22803_, new_n17244_, new_n1511_ );
or   ( new_n22804_, new_n17248_, new_n1310_ );
and  ( new_n22805_, new_n22804_, new_n22803_ );
or   ( new_n22806_, new_n22805_, new_n16814_ );
and  ( new_n22807_, new_n17255_, RI2b1c4342dbe8_80 );
and  ( new_n22808_, new_n17240_, RI2b1c4342db70_79 );
or   ( new_n22809_, new_n22808_, new_n22807_ );
or   ( new_n22810_, new_n22809_, new_n17142_ );
and  ( new_n22811_, new_n22810_, new_n22806_ );
or   ( new_n22812_, new_n22811_, new_n22802_ );
and  ( new_n22813_, new_n22811_, new_n22802_ );
or   ( new_n22814_, new_n16607_, new_n2119_ );
or   ( new_n22815_, new_n16613_, new_n126_ );
and  ( new_n22816_, new_n22815_, new_n22814_ );
or   ( new_n22817_, new_n22816_, new_n16505_ );
and  ( new_n22818_, new_n16616_, RI2b1c4342dcd8_82 );
and  ( new_n22819_, new_n16603_, RI2b1c4342dc60_81 );
or   ( new_n22820_, new_n22819_, new_n22818_ );
or   ( new_n22821_, new_n22820_, new_n16438_ );
and  ( new_n22822_, new_n22821_, new_n22817_ );
or   ( new_n22823_, new_n22822_, new_n22813_ );
and  ( new_n22824_, new_n22823_, new_n22812_ );
or   ( new_n22825_, new_n22824_, new_n22793_ );
and  ( new_n22826_, new_n22825_, new_n22792_ );
or   ( new_n22827_, new_n16366_, new_n2541_ );
or   ( new_n22828_, new_n16355_, new_n121_ );
and  ( new_n22829_, new_n22828_, new_n22827_ );
or   ( new_n22830_, new_n22829_, new_n16085_ );
and  ( new_n22831_, new_n16358_, RI2b1c4342ddc8_84 );
and  ( new_n22832_, new_n16362_, RI2b1c4342dd50_83 );
or   ( new_n22833_, new_n22832_, new_n22831_ );
or   ( new_n22834_, new_n22833_, new_n16048_ );
and  ( new_n22835_, new_n22834_, new_n22830_ );
or   ( new_n22836_, new_n16075_, new_n3239_ );
or   ( new_n22837_, new_n16060_, new_n2806_ );
and  ( new_n22838_, new_n22837_, new_n22836_ );
or   ( new_n22839_, new_n22838_, new_n16052_ );
and  ( new_n22840_, new_n16063_, RI2b1c4342deb8_86 );
and  ( new_n22841_, new_n16066_, RI2b1c4342de40_85 );
or   ( new_n22842_, new_n22841_, new_n22840_ );
or   ( new_n22843_, new_n22842_, new_n16071_ );
and  ( new_n22844_, new_n22843_, new_n22839_ );
or   ( new_n22845_, new_n22844_, new_n22835_ );
and  ( new_n22846_, new_n22844_, new_n22835_ );
or   ( new_n22847_, new_n16033_, new_n3902_ );
or   ( new_n22848_, new_n16017_, new_n3924_ );
and  ( new_n22849_, new_n22848_, new_n22847_ );
or   ( new_n22850_, new_n22849_, new_n16009_ );
and  ( new_n22851_, new_n16021_, RI2b1c4342dfa8_88 );
and  ( new_n22852_, new_n16024_, RI2b1c4342df30_87 );
or   ( new_n22853_, new_n22852_, new_n22851_ );
or   ( new_n22854_, new_n22853_, new_n16029_ );
and  ( new_n22855_, new_n22854_, new_n22850_ );
or   ( new_n22856_, new_n22855_, new_n22846_ );
and  ( new_n22857_, new_n22856_, new_n22845_ );
or   ( new_n22858_, new_n16208_, new_n4635_ );
or   ( new_n22859_, new_n16194_, new_n132_ );
and  ( new_n22860_, new_n22859_, new_n22858_ );
or   ( new_n22861_, new_n22860_, new_n16186_ );
and  ( new_n22862_, new_n16196_, RI2b1c4342e098_90 );
and  ( new_n22863_, new_n16199_, RI2b1c4342e020_89 );
or   ( new_n22864_, new_n22863_, new_n22862_ );
or   ( new_n22865_, new_n22864_, new_n16204_ );
and  ( new_n22866_, new_n22865_, new_n22861_ );
or   ( new_n22867_, new_n16238_, new_n5459_ );
or   ( new_n22868_, new_n16224_, new_n117_ );
and  ( new_n22869_, new_n22868_, new_n22867_ );
or   ( new_n22870_, new_n22869_, new_n16217_ );
and  ( new_n22871_, new_n16226_, RI2b1c4342e188_92 );
and  ( new_n22872_, new_n16229_, RI2b1c4342e110_91 );
or   ( new_n22873_, new_n22872_, new_n22871_ );
or   ( new_n22874_, new_n22873_, new_n16234_ );
and  ( new_n22875_, new_n22874_, new_n22870_ );
or   ( new_n22876_, new_n22875_, new_n22866_ );
and  ( new_n22877_, new_n22875_, new_n22866_ );
or   ( new_n22878_, new_n16174_, new_n6321_ );
or   ( new_n22879_, new_n16160_, new_n6307_ );
and  ( new_n22880_, new_n22879_, new_n22878_ );
or   ( new_n22881_, new_n22880_, new_n16151_ );
and  ( new_n22882_, new_n16162_, RI2b1c4342e278_94 );
and  ( new_n22883_, new_n16165_, RI2b1c4342e200_93 );
or   ( new_n22884_, new_n22883_, new_n22882_ );
or   ( new_n22885_, new_n22884_, new_n16170_ );
and  ( new_n22886_, new_n22885_, new_n22881_ );
or   ( new_n22887_, new_n22886_, new_n22877_ );
and  ( new_n22888_, new_n22887_, new_n22876_ );
or   ( new_n22889_, new_n22888_, new_n22857_ );
and  ( new_n22890_, new_n22888_, new_n22857_ );
or   ( new_n22891_, new_n22646_, new_n22489_ );
or   ( new_n22892_, new_n22643_, new_n22498_ );
and  ( new_n22893_, new_n22892_, new_n22891_ );
or   ( new_n22894_, new_n22893_, new_n22649_ );
and  ( new_n22895_, new_n22647_, new_n22500_ );
or   ( new_n22896_, new_n22895_, new_n22501_ );
and  ( new_n22897_, new_n22896_, new_n22894_ );
or   ( new_n22898_, new_n22897_, new_n22890_ );
and  ( new_n22899_, new_n22898_, new_n22889_ );
or   ( new_n22900_, new_n22899_, new_n22826_ );
and  ( new_n22901_, new_n22899_, new_n22826_ );
or   ( new_n22902_, new_n22631_, new_n22456_ );
or   ( new_n22903_, new_n22628_, new_n22465_ );
and  ( new_n22904_, new_n22903_, new_n22902_ );
or   ( new_n22905_, new_n22904_, new_n22636_ );
and  ( new_n22906_, new_n22632_, new_n22466_ );
or   ( new_n22907_, new_n22906_, new_n22476_ );
and  ( new_n22908_, new_n22907_, new_n22905_ );
or   ( new_n22909_, new_n22618_, new_n22425_ );
or   ( new_n22910_, new_n22615_, new_n22434_ );
and  ( new_n22911_, new_n22910_, new_n22909_ );
or   ( new_n22912_, new_n22911_, new_n22623_ );
and  ( new_n22913_, new_n22619_, new_n22435_ );
or   ( new_n22914_, new_n22913_, new_n22445_ );
and  ( new_n22915_, new_n22914_, new_n22912_ );
or   ( new_n22916_, new_n22915_, new_n22908_ );
and  ( new_n22917_, new_n22915_, new_n22908_ );
or   ( new_n22918_, new_n22603_, new_n22392_ );
or   ( new_n22919_, new_n22600_, new_n22401_ );
and  ( new_n22920_, new_n22919_, new_n22918_ );
or   ( new_n22921_, new_n22920_, new_n22608_ );
and  ( new_n22922_, new_n22604_, new_n22402_ );
or   ( new_n22923_, new_n22922_, new_n22412_ );
and  ( new_n22924_, new_n22923_, new_n22921_ );
or   ( new_n22925_, new_n22924_, new_n22917_ );
and  ( new_n22926_, new_n22925_, new_n22916_ );
or   ( new_n22927_, new_n22926_, new_n22901_ );
and  ( new_n22928_, new_n22927_, new_n22900_ );
or   ( new_n22929_, new_n22679_, new_n22298_ );
or   ( new_n22930_, new_n22676_, new_n22305_ );
and  ( new_n22931_, new_n22930_, new_n22929_ );
or   ( new_n22932_, new_n22931_, new_n22684_ );
and  ( new_n22933_, new_n22680_, new_n22306_ );
or   ( new_n22934_, new_n22933_, new_n22314_ );
and  ( new_n22935_, new_n22934_, new_n22932_ );
or   ( new_n22936_, new_n22661_, new_n22509_ );
or   ( new_n22937_, new_n22658_, new_n22516_ );
and  ( new_n22938_, new_n22937_, new_n22936_ );
or   ( new_n22939_, new_n22938_, new_n22666_ );
and  ( new_n22940_, new_n22662_, new_n22517_ );
or   ( new_n22941_, new_n22940_, new_n22525_ );
and  ( new_n22942_, new_n22941_, new_n22939_ );
or   ( new_n22943_, new_n22942_, new_n22935_ );
and  ( new_n22944_, new_n22942_, new_n22935_ );
or   ( new_n22945_, new_n22638_, new_n22447_ );
or   ( new_n22946_, new_n22625_, new_n22478_ );
and  ( new_n22947_, new_n22946_, new_n22945_ );
or   ( new_n22948_, new_n22947_, new_n22651_ );
and  ( new_n22949_, new_n22639_, new_n22480_ );
or   ( new_n22950_, new_n22949_, new_n22503_ );
and  ( new_n22951_, new_n22950_, new_n22948_ );
or   ( new_n22952_, new_n22951_, new_n22944_ );
and  ( new_n22953_, new_n22952_, new_n22943_ );
or   ( new_n22954_, new_n22953_, new_n22928_ );
and  ( new_n22955_, new_n22953_, new_n22928_ );
or   ( new_n22956_, new_n22137_, new_n21953_ );
or   ( new_n22957_, new_n22124_, new_n21984_ );
and  ( new_n22958_, new_n22957_, new_n22956_ );
or   ( new_n22959_, new_n22958_, new_n22144_ );
and  ( new_n22960_, new_n22138_, new_n21985_ );
or   ( new_n22961_, new_n22960_, new_n21997_ );
and  ( new_n22962_, new_n22961_, new_n22959_ );
or   ( new_n22963_, new_n22962_, new_n22955_ );
and  ( new_n22964_, new_n22963_, new_n22954_ );
or   ( new_n22965_, new_n22159_, new_n21856_ );
or   ( new_n22966_, new_n22169_, new_n21887_ );
and  ( new_n22967_, new_n22966_, new_n22965_ );
or   ( new_n22968_, new_n22967_, new_n22184_ );
and  ( new_n22969_, new_n22170_, new_n21888_ );
or   ( new_n22970_, new_n22969_, new_n21920_ );
and  ( new_n22971_, new_n22970_, new_n22968_ );
or   ( new_n22972_, new_n22673_, new_n22316_ );
or   ( new_n22973_, new_n22686_, new_n22291_ );
and  ( new_n22974_, new_n22973_, new_n22972_ );
or   ( new_n22975_, new_n22974_, new_n22691_ );
and  ( new_n22976_, new_n22687_, new_n22317_ );
or   ( new_n22977_, new_n22976_, new_n22325_ );
and  ( new_n22978_, new_n22977_, new_n22975_ );
or   ( new_n22979_, new_n22978_, new_n22971_ );
and  ( new_n22980_, new_n22978_, new_n22971_ );
or   ( new_n22981_, new_n22653_, new_n22416_ );
or   ( new_n22982_, new_n22612_, new_n22505_ );
and  ( new_n22983_, new_n22982_, new_n22981_ );
or   ( new_n22984_, new_n22983_, new_n22668_ );
and  ( new_n22985_, new_n22654_, new_n22507_ );
or   ( new_n22986_, new_n22985_, new_n22527_ );
and  ( new_n22987_, new_n22986_, new_n22984_ );
or   ( new_n22988_, new_n22987_, new_n22980_ );
and  ( new_n22989_, new_n22988_, new_n22979_ );
or   ( new_n22990_, new_n22989_, new_n22964_ );
and  ( new_n22991_, new_n22989_, new_n22964_ );
or   ( new_n22992_, new_n22706_, new_n22266_ );
or   ( new_n22993_, new_n22703_, new_n22273_ );
and  ( new_n22994_, new_n22993_, new_n22992_ );
or   ( new_n22995_, new_n22994_, new_n22711_ );
and  ( new_n22996_, new_n22707_, new_n22274_ );
or   ( new_n22997_, new_n22996_, new_n22282_ );
and  ( new_n22998_, new_n22997_, new_n22995_ );
or   ( new_n22999_, new_n22998_, new_n22991_ );
and  ( new_n23000_, new_n22999_, new_n22990_ );
or   ( new_n23001_, new_n23000_, new_n22730_ );
or   ( new_n23002_, new_n22713_, new_n22540_ );
or   ( new_n23003_, new_n22700_, new_n22284_ );
and  ( new_n23004_, new_n23003_, new_n23002_ );
or   ( new_n23005_, new_n23004_, new_n22718_ );
and  ( new_n23006_, new_n22714_, new_n22542_ );
or   ( new_n23007_, new_n23006_, new_n22549_ );
and  ( new_n23008_, new_n23007_, new_n23005_ );
and  ( new_n23009_, new_n23000_, new_n22730_ );
or   ( new_n23010_, new_n23009_, new_n23008_ );
and  ( new_n23011_, new_n23010_, new_n23001_ );
or   ( new_n23012_, new_n23011_, new_n22727_ );
and  ( new_n23013_, new_n23012_, new_n22564_ );
or   ( new_n23014_, new_n23013_, new_n22563_ );
or   ( new_n23015_, new_n23014_, new_n22102_ );
and  ( new_n23016_, new_n23015_, new_n22100_ );
and  ( new_n23017_, new_n23011_, new_n22727_ );
or   ( new_n23018_, new_n23017_, new_n22563_ );
or   ( new_n23019_, new_n23018_, new_n22102_ );
or   ( new_n23020_, new_n23006_, new_n22718_ );
or   ( new_n23021_, new_n23004_, new_n22549_ );
and  ( new_n23022_, new_n23021_, new_n23020_ );
or   ( new_n23023_, new_n22573_, new_n22570_ );
and  ( new_n23024_, new_n23023_, new_n22259_ );
or   ( new_n23025_, new_n23024_, new_n23000_ );
or   ( new_n23026_, new_n22969_, new_n22184_ );
or   ( new_n23027_, new_n22967_, new_n21920_ );
and  ( new_n23028_, new_n23027_, new_n23026_ );
or   ( new_n23029_, new_n22976_, new_n22691_ );
or   ( new_n23030_, new_n22974_, new_n22325_ );
and  ( new_n23031_, new_n23030_, new_n23029_ );
or   ( new_n23032_, new_n23031_, new_n23028_ );
and  ( new_n23033_, new_n23031_, new_n23028_ );
or   ( new_n23034_, new_n22985_, new_n22668_ );
or   ( new_n23035_, new_n22983_, new_n22527_ );
and  ( new_n23036_, new_n23035_, new_n23034_ );
or   ( new_n23037_, new_n23036_, new_n23033_ );
and  ( new_n23038_, new_n23037_, new_n23032_ );
or   ( new_n23039_, new_n22736_, new_n21261_ );
or   ( new_n23040_, new_n22732_, new_n21009_ );
and  ( new_n23041_, new_n23040_, new_n23039_ );
or   ( new_n23042_, new_n22745_, new_n21013_ );
or   ( new_n23043_, new_n22741_, new_n21265_ );
and  ( new_n23044_, new_n23043_, new_n23042_ );
or   ( new_n23045_, new_n23044_, new_n23041_ );
and  ( new_n23046_, new_n23044_, new_n23041_ );
or   ( new_n23047_, new_n22756_, new_n20156_ );
or   ( new_n23048_, new_n22752_, new_n20443_ );
and  ( new_n23049_, new_n23048_, new_n23047_ );
or   ( new_n23050_, new_n23049_, new_n23046_ );
and  ( new_n23051_, new_n23050_, new_n23045_ );
or   ( new_n23052_, new_n22767_, new_n19394_ );
or   ( new_n23053_, new_n22763_, new_n19659_ );
and  ( new_n23054_, new_n23053_, new_n23052_ );
or   ( new_n23055_, new_n22776_, new_n18742_ );
or   ( new_n23056_, new_n22772_, new_n18977_ );
and  ( new_n23057_, new_n23056_, new_n23055_ );
or   ( new_n23058_, new_n23057_, new_n23054_ );
and  ( new_n23059_, new_n23057_, new_n23054_ );
or   ( new_n23060_, new_n22787_, new_n18066_ );
or   ( new_n23061_, new_n22783_, new_n18309_ );
and  ( new_n23062_, new_n23061_, new_n23060_ );
or   ( new_n23063_, new_n23062_, new_n23059_ );
and  ( new_n23064_, new_n23063_, new_n23058_ );
or   ( new_n23065_, new_n23064_, new_n23051_ );
and  ( new_n23066_, new_n23064_, new_n23051_ );
or   ( new_n23067_, new_n22800_, new_n17238_ );
or   ( new_n23068_, new_n22796_, new_n17650_ );
and  ( new_n23069_, new_n23068_, new_n23067_ );
or   ( new_n23070_, new_n22809_, new_n16814_ );
or   ( new_n23071_, new_n22805_, new_n17142_ );
and  ( new_n23072_, new_n23071_, new_n23070_ );
or   ( new_n23073_, new_n23072_, new_n23069_ );
and  ( new_n23074_, new_n23072_, new_n23069_ );
or   ( new_n23075_, new_n22820_, new_n16505_ );
or   ( new_n23076_, new_n22816_, new_n16438_ );
and  ( new_n23077_, new_n23076_, new_n23075_ );
or   ( new_n23078_, new_n23077_, new_n23074_ );
and  ( new_n23079_, new_n23078_, new_n23073_ );
or   ( new_n23080_, new_n23079_, new_n23066_ );
and  ( new_n23081_, new_n23080_, new_n23065_ );
or   ( new_n23082_, new_n22833_, new_n16085_ );
or   ( new_n23083_, new_n22829_, new_n16048_ );
and  ( new_n23084_, new_n23083_, new_n23082_ );
or   ( new_n23085_, new_n22842_, new_n16052_ );
or   ( new_n23086_, new_n22838_, new_n16071_ );
and  ( new_n23087_, new_n23086_, new_n23085_ );
or   ( new_n23088_, new_n23087_, new_n23084_ );
and  ( new_n23089_, new_n23087_, new_n23084_ );
or   ( new_n23090_, new_n22853_, new_n16009_ );
or   ( new_n23091_, new_n22849_, new_n16029_ );
and  ( new_n23092_, new_n23091_, new_n23090_ );
or   ( new_n23093_, new_n23092_, new_n23089_ );
and  ( new_n23094_, new_n23093_, new_n23088_ );
or   ( new_n23095_, new_n22864_, new_n16186_ );
or   ( new_n23096_, new_n22860_, new_n16204_ );
and  ( new_n23097_, new_n23096_, new_n23095_ );
or   ( new_n23098_, new_n22873_, new_n16217_ );
or   ( new_n23099_, new_n22869_, new_n16234_ );
and  ( new_n23100_, new_n23099_, new_n23098_ );
or   ( new_n23101_, new_n23100_, new_n23097_ );
and  ( new_n23102_, new_n23100_, new_n23097_ );
or   ( new_n23103_, new_n22884_, new_n16151_ );
or   ( new_n23104_, new_n22880_, new_n16170_ );
and  ( new_n23105_, new_n23104_, new_n23103_ );
or   ( new_n23106_, new_n23105_, new_n23102_ );
and  ( new_n23107_, new_n23106_, new_n23101_ );
or   ( new_n23108_, new_n23107_, new_n23094_ );
and  ( new_n23109_, new_n23107_, new_n23094_ );
or   ( new_n23110_, new_n22895_, new_n22649_ );
or   ( new_n23111_, new_n22893_, new_n22501_ );
and  ( new_n23112_, new_n23111_, new_n23110_ );
or   ( new_n23113_, new_n23112_, new_n23109_ );
and  ( new_n23114_, new_n23113_, new_n23108_ );
or   ( new_n23115_, new_n23114_, new_n23081_ );
and  ( new_n23116_, new_n23114_, new_n23081_ );
or   ( new_n23117_, new_n22906_, new_n22636_ );
or   ( new_n23118_, new_n22904_, new_n22476_ );
and  ( new_n23119_, new_n23118_, new_n23117_ );
or   ( new_n23120_, new_n22913_, new_n22623_ );
or   ( new_n23121_, new_n22911_, new_n22445_ );
and  ( new_n23122_, new_n23121_, new_n23120_ );
or   ( new_n23123_, new_n23122_, new_n23119_ );
and  ( new_n23124_, new_n23122_, new_n23119_ );
or   ( new_n23125_, new_n22922_, new_n22608_ );
or   ( new_n23126_, new_n22920_, new_n22412_ );
and  ( new_n23127_, new_n23126_, new_n23125_ );
or   ( new_n23128_, new_n23127_, new_n23124_ );
and  ( new_n23129_, new_n23128_, new_n23123_ );
or   ( new_n23130_, new_n23129_, new_n23116_ );
and  ( new_n23131_, new_n23130_, new_n23115_ );
or   ( new_n23132_, new_n22933_, new_n22684_ );
or   ( new_n23133_, new_n22931_, new_n22314_ );
and  ( new_n23134_, new_n23133_, new_n23132_ );
or   ( new_n23135_, new_n22940_, new_n22666_ );
or   ( new_n23136_, new_n22938_, new_n22525_ );
and  ( new_n23137_, new_n23136_, new_n23135_ );
or   ( new_n23138_, new_n23137_, new_n23134_ );
and  ( new_n23139_, new_n23137_, new_n23134_ );
or   ( new_n23140_, new_n22949_, new_n22651_ );
or   ( new_n23141_, new_n22947_, new_n22503_ );
and  ( new_n23142_, new_n23141_, new_n23140_ );
or   ( new_n23143_, new_n23142_, new_n23139_ );
and  ( new_n23144_, new_n23143_, new_n23138_ );
or   ( new_n23145_, new_n23144_, new_n23131_ );
and  ( new_n23146_, new_n23144_, new_n23131_ );
or   ( new_n23147_, new_n22960_, new_n22144_ );
or   ( new_n23148_, new_n22958_, new_n21997_ );
and  ( new_n23149_, new_n23148_, new_n23147_ );
or   ( new_n23150_, new_n23149_, new_n23146_ );
and  ( new_n23151_, new_n23150_, new_n23145_ );
or   ( new_n23152_, new_n23151_, new_n23038_ );
and  ( new_n23153_, new_n23151_, new_n23038_ );
or   ( new_n23154_, new_n22996_, new_n22711_ );
or   ( new_n23155_, new_n22994_, new_n22282_ );
and  ( new_n23156_, new_n23155_, new_n23154_ );
or   ( new_n23157_, new_n23156_, new_n23153_ );
and  ( new_n23158_, new_n23157_, new_n23152_ );
or   ( new_n23159_, new_n23158_, new_n22730_ );
and  ( new_n23160_, new_n23159_, new_n23025_ );
or   ( new_n23161_, new_n23160_, new_n23022_ );
or   ( new_n23162_, new_n23158_, new_n23024_ );
and  ( new_n23163_, new_n23162_, new_n23001_ );
or   ( new_n23164_, new_n23163_, new_n23008_ );
and  ( new_n23165_, new_n23164_, new_n23161_ );
or   ( new_n23166_, new_n22693_, new_n22529_ );
or   ( new_n23167_, new_n22670_, new_n22327_ );
and  ( new_n23168_, new_n23167_, new_n23166_ );
or   ( new_n23169_, new_n23168_, new_n22698_ );
and  ( new_n23170_, new_n22694_, new_n22531_ );
or   ( new_n23171_, new_n23170_, new_n22538_ );
and  ( new_n23172_, new_n23171_, new_n23169_ );
or   ( new_n23173_, new_n22595_, new_n22350_ );
or   ( new_n23174_, new_n22582_, new_n22381_ );
and  ( new_n23175_, new_n23174_, new_n23173_ );
or   ( new_n23176_, new_n23175_, new_n22610_ );
and  ( new_n23177_, new_n22596_, new_n22382_ );
or   ( new_n23178_, new_n23177_, new_n22414_ );
and  ( new_n23179_, new_n23178_, new_n23176_ );
or   ( new_n23180_, new_n23137_, new_n22935_ );
or   ( new_n23181_, new_n23134_, new_n22942_ );
and  ( new_n23182_, new_n23181_, new_n23180_ );
or   ( new_n23183_, new_n23182_, new_n23142_ );
and  ( new_n23184_, new_n23138_, new_n22943_ );
or   ( new_n23185_, new_n23184_, new_n22951_ );
and  ( new_n23186_, new_n23185_, new_n23183_ );
or   ( new_n23187_, new_n23186_, new_n23179_ );
and  ( new_n23188_, new_n23186_, new_n23179_ );
or   ( new_n23189_, new_n23114_, new_n22826_ );
or   ( new_n23190_, new_n23081_, new_n22899_ );
and  ( new_n23191_, new_n23190_, new_n23189_ );
or   ( new_n23192_, new_n23191_, new_n23129_ );
and  ( new_n23193_, new_n23115_, new_n22900_ );
or   ( new_n23194_, new_n23193_, new_n22926_ );
and  ( new_n23195_, new_n23194_, new_n23192_ );
or   ( new_n23196_, new_n23195_, new_n23188_ );
and  ( new_n23197_, new_n23196_, new_n23187_ );
or   ( new_n23198_, new_n22588_, new_n22359_ );
or   ( new_n23199_, new_n22585_, new_n22368_ );
and  ( new_n23200_, new_n23199_, new_n23198_ );
or   ( new_n23201_, new_n23200_, new_n22593_ );
and  ( new_n23202_, new_n22589_, new_n22369_ );
or   ( new_n23203_, new_n23202_, new_n22379_ );
and  ( new_n23204_, new_n23203_, new_n23201_ );
or   ( new_n23205_, new_n22581_, new_n22340_ );
or   ( new_n23206_, new_n22578_, new_n22349_ );
and  ( new_n23207_, new_n23206_, new_n23205_ );
or   ( new_n23208_, new_n23207_, new_n23204_ );
and  ( new_n23209_, new_n23207_, new_n23204_ );
or   ( new_n23210_, new_n23122_, new_n22908_ );
or   ( new_n23211_, new_n23119_, new_n22915_ );
and  ( new_n23212_, new_n23211_, new_n23210_ );
or   ( new_n23213_, new_n23212_, new_n23127_ );
and  ( new_n23214_, new_n23123_, new_n22916_ );
or   ( new_n23215_, new_n23214_, new_n22924_ );
and  ( new_n23216_, new_n23215_, new_n23213_ );
or   ( new_n23217_, new_n23216_, new_n23209_ );
and  ( new_n23218_, new_n23217_, new_n23208_ );
or   ( new_n23219_, new_n16607_, new_n121_ );
or   ( new_n23220_, new_n16613_, new_n2119_ );
and  ( new_n23221_, new_n23220_, new_n23219_ );
or   ( new_n23222_, new_n23221_, new_n16505_ );
and  ( new_n23223_, new_n16616_, RI2b1c4342dd50_83 );
and  ( new_n23224_, new_n16603_, RI2b1c4342dcd8_82 );
or   ( new_n23225_, new_n23224_, new_n23223_ );
or   ( new_n23226_, new_n23225_, new_n16438_ );
and  ( new_n23227_, new_n23226_, new_n23222_ );
or   ( new_n23228_, new_n16366_, new_n2806_ );
or   ( new_n23229_, new_n16355_, new_n2541_ );
and  ( new_n23230_, new_n23229_, new_n23228_ );
or   ( new_n23231_, new_n23230_, new_n16085_ );
and  ( new_n23232_, new_n16358_, RI2b1c4342de40_85 );
and  ( new_n23233_, new_n16362_, RI2b1c4342ddc8_84 );
or   ( new_n23234_, new_n23233_, new_n23232_ );
or   ( new_n23235_, new_n23234_, new_n16048_ );
and  ( new_n23236_, new_n23235_, new_n23231_ );
or   ( new_n23237_, new_n23236_, new_n23227_ );
and  ( new_n23238_, new_n23236_, new_n23227_ );
or   ( new_n23239_, new_n16075_, new_n3924_ );
or   ( new_n23240_, new_n16060_, new_n3239_ );
and  ( new_n23241_, new_n23240_, new_n23239_ );
or   ( new_n23242_, new_n23241_, new_n16052_ );
and  ( new_n23243_, new_n16063_, RI2b1c4342df30_87 );
and  ( new_n23244_, new_n16066_, RI2b1c4342deb8_86 );
or   ( new_n23245_, new_n23244_, new_n23243_ );
or   ( new_n23246_, new_n23245_, new_n16071_ );
and  ( new_n23247_, new_n23246_, new_n23242_ );
or   ( new_n23248_, new_n23247_, new_n23238_ );
and  ( new_n23249_, new_n23248_, new_n23237_ );
or   ( new_n23250_, new_n16033_, new_n132_ );
or   ( new_n23251_, new_n16017_, new_n3902_ );
and  ( new_n23252_, new_n23251_, new_n23250_ );
or   ( new_n23253_, new_n23252_, new_n16009_ );
and  ( new_n23254_, new_n16021_, RI2b1c4342e020_89 );
and  ( new_n23255_, new_n16024_, RI2b1c4342dfa8_88 );
or   ( new_n23256_, new_n23255_, new_n23254_ );
or   ( new_n23257_, new_n23256_, new_n16029_ );
and  ( new_n23258_, new_n23257_, new_n23253_ );
or   ( new_n23259_, new_n16208_, new_n117_ );
or   ( new_n23260_, new_n16194_, new_n4635_ );
and  ( new_n23261_, new_n23260_, new_n23259_ );
or   ( new_n23262_, new_n23261_, new_n16186_ );
and  ( new_n23263_, new_n16196_, RI2b1c4342e110_91 );
and  ( new_n23264_, new_n16199_, RI2b1c4342e098_90 );
or   ( new_n23265_, new_n23264_, new_n23263_ );
or   ( new_n23266_, new_n23265_, new_n16204_ );
and  ( new_n23267_, new_n23266_, new_n23262_ );
or   ( new_n23268_, new_n23267_, new_n23258_ );
and  ( new_n23269_, new_n23267_, new_n23258_ );
or   ( new_n23270_, new_n16238_, new_n6307_ );
or   ( new_n23271_, new_n16224_, new_n5459_ );
and  ( new_n23272_, new_n23271_, new_n23270_ );
or   ( new_n23273_, new_n23272_, new_n16217_ );
and  ( new_n23274_, new_n16226_, RI2b1c4342e200_93 );
and  ( new_n23275_, new_n16229_, RI2b1c4342e188_92 );
or   ( new_n23276_, new_n23275_, new_n23274_ );
or   ( new_n23277_, new_n23276_, new_n16234_ );
and  ( new_n23278_, new_n23277_, new_n23273_ );
or   ( new_n23279_, new_n23278_, new_n23269_ );
and  ( new_n23280_, new_n23279_, new_n23268_ );
or   ( new_n23281_, new_n23280_, new_n23249_ );
and  ( new_n23282_, new_n23280_, new_n23249_ );
or   ( new_n23283_, new_n16119_, new_n7274_ );
or   ( new_n23284_, new_n16123_, new_n124_ );
and  ( new_n23285_, new_n23284_, new_n23283_ );
or   ( new_n23286_, new_n23285_, new_n16108_ );
and  ( new_n23287_, new_n16132_, RI2b1c4342e368_96 );
and  ( new_n23288_, new_n16114_, RI2b1c4342e2f0_95 );
or   ( new_n23289_, new_n23288_, new_n23287_ );
or   ( new_n23290_, new_n23289_, new_n16128_ );
and  ( new_n23291_, new_n23290_, new_n23286_ );
or   ( new_n23292_, new_n23291_, new_n23282_ );
and  ( new_n23293_, new_n23292_, new_n23281_ );
or   ( new_n23294_, new_n20557_, new_n110_ );
or   ( new_n23295_, new_n20562_, new_n755_ );
and  ( new_n23296_, new_n23295_, new_n23294_ );
or   ( new_n23297_, new_n23296_, new_n20156_ );
and  ( new_n23298_, new_n20566_, RI2b1c4342d7b0_71 );
and  ( new_n23299_, new_n20553_, RI2b1c4342d738_70 );
or   ( new_n23300_, new_n23299_, new_n23298_ );
or   ( new_n23301_, new_n23300_, new_n20443_ );
and  ( new_n23302_, new_n23301_, new_n23297_ );
or   ( new_n23303_, new_n19758_, new_n105_ );
or   ( new_n23304_, new_n19763_, new_n806_ );
and  ( new_n23305_, new_n23304_, new_n23303_ );
or   ( new_n23306_, new_n23305_, new_n19394_ );
and  ( new_n23307_, new_n19767_, RI2b1c4342d8a0_73 );
and  ( new_n23308_, new_n19754_, RI2b1c4342d828_72 );
or   ( new_n23309_, new_n23308_, new_n23307_ );
or   ( new_n23310_, new_n23309_, new_n19659_ );
and  ( new_n23311_, new_n23310_, new_n23306_ );
or   ( new_n23312_, new_n23311_, new_n23302_ );
and  ( new_n23313_, new_n23311_, new_n23302_ );
or   ( new_n23314_, new_n19048_, new_n843_ );
or   ( new_n23315_, new_n19055_, new_n859_ );
and  ( new_n23316_, new_n23315_, new_n23314_ );
or   ( new_n23317_, new_n23316_, new_n18742_ );
and  ( new_n23318_, new_n19057_, RI2b1c4342d990_75 );
and  ( new_n23319_, new_n19044_, RI2b1c4342d918_74 );
or   ( new_n23320_, new_n23319_, new_n23318_ );
or   ( new_n23321_, new_n23320_, new_n18977_ );
and  ( new_n23322_, new_n23321_, new_n23317_ );
or   ( new_n23323_, new_n23322_, new_n23313_ );
and  ( new_n23324_, new_n23323_, new_n23312_ );
nor  ( new_n23325_, new_n22333_, new_n112_ );
nor  ( new_n23326_, new_n23325_, new_n8170_ );
or   ( new_n23327_, new_n23326_, new_n21261_ );
and  ( new_n23328_, new_n22337_, RI2b1c4342d5d0_67 );
and  ( new_n23329_, new_n22330_, RI2b1c4342d558_66 );
or   ( new_n23330_, new_n23329_, new_n23328_ );
or   ( new_n23331_, new_n23330_, new_n21009_ );
and  ( new_n23332_, new_n23331_, new_n23327_ );
and  ( new_n23333_, new_n23332_, new_n16128_ );
or   ( new_n23334_, new_n23332_, new_n16128_ );
or   ( new_n23335_, new_n21419_, new_n591_ );
or   ( new_n23336_, new_n21424_, new_n612_ );
and  ( new_n23337_, new_n23336_, new_n23335_ );
or   ( new_n23338_, new_n23337_, new_n21013_ );
and  ( new_n23339_, new_n21428_, RI2b1c4342d6c0_69 );
and  ( new_n23340_, new_n21415_, RI2b1c4342d648_68 );
or   ( new_n23341_, new_n23340_, new_n23339_ );
or   ( new_n23342_, new_n23341_, new_n21265_ );
and  ( new_n23343_, new_n23342_, new_n23338_ );
and  ( new_n23344_, new_n23343_, new_n23334_ );
or   ( new_n23345_, new_n23344_, new_n23333_ );
and  ( new_n23346_, new_n23345_, new_n23324_ );
or   ( new_n23347_, new_n23345_, new_n23324_ );
or   ( new_n23348_, new_n18388_, new_n1004_ );
or   ( new_n23349_, new_n18395_, new_n886_ );
and  ( new_n23350_, new_n23349_, new_n23348_ );
or   ( new_n23351_, new_n23350_, new_n18066_ );
and  ( new_n23352_, new_n18397_, RI2b1c4342da80_77 );
and  ( new_n23353_, new_n18384_, RI2b1c4342da08_76 );
or   ( new_n23354_, new_n23353_, new_n23352_ );
or   ( new_n23355_, new_n23354_, new_n18309_ );
and  ( new_n23356_, new_n23355_, new_n23351_ );
or   ( new_n23357_, new_n17727_, new_n1310_ );
or   ( new_n23358_, new_n17734_, new_n1002_ );
and  ( new_n23359_, new_n23358_, new_n23357_ );
or   ( new_n23360_, new_n23359_, new_n17238_ );
and  ( new_n23361_, new_n17736_, RI2b1c4342db70_79 );
and  ( new_n23362_, new_n17723_, RI2b1c4342daf8_78 );
or   ( new_n23363_, new_n23362_, new_n23361_ );
or   ( new_n23364_, new_n23363_, new_n17650_ );
and  ( new_n23365_, new_n23364_, new_n23360_ );
or   ( new_n23366_, new_n23365_, new_n23356_ );
and  ( new_n23367_, new_n23365_, new_n23356_ );
or   ( new_n23368_, new_n17244_, new_n126_ );
or   ( new_n23369_, new_n17248_, new_n1511_ );
and  ( new_n23370_, new_n23369_, new_n23368_ );
or   ( new_n23371_, new_n23370_, new_n16814_ );
and  ( new_n23372_, new_n17255_, RI2b1c4342dc60_81 );
and  ( new_n23373_, new_n17240_, RI2b1c4342dbe8_80 );
or   ( new_n23374_, new_n23373_, new_n23372_ );
or   ( new_n23375_, new_n23374_, new_n17142_ );
and  ( new_n23376_, new_n23375_, new_n23371_ );
or   ( new_n23377_, new_n23376_, new_n23367_ );
and  ( new_n23378_, new_n23377_, new_n23366_ );
and  ( new_n23379_, new_n23378_, new_n23347_ );
or   ( new_n23380_, new_n23379_, new_n23346_ );
and  ( new_n23381_, new_n23380_, new_n23293_ );
or   ( new_n23382_, new_n23380_, new_n23293_ );
or   ( new_n23383_, new_n23100_, new_n22866_ );
or   ( new_n23384_, new_n23097_, new_n22875_ );
and  ( new_n23385_, new_n23384_, new_n23383_ );
or   ( new_n23386_, new_n23385_, new_n23105_ );
and  ( new_n23387_, new_n23101_, new_n22876_ );
or   ( new_n23388_, new_n23387_, new_n22886_ );
and  ( new_n23389_, new_n23388_, new_n23386_ );
or   ( new_n23390_, new_n23087_, new_n22835_ );
or   ( new_n23391_, new_n23084_, new_n22844_ );
and  ( new_n23392_, new_n23391_, new_n23390_ );
or   ( new_n23393_, new_n23392_, new_n23092_ );
and  ( new_n23394_, new_n23088_, new_n22845_ );
or   ( new_n23395_, new_n23394_, new_n22855_ );
and  ( new_n23396_, new_n23395_, new_n23393_ );
or   ( new_n23397_, new_n23396_, new_n23389_ );
and  ( new_n23398_, new_n23396_, new_n23389_ );
or   ( new_n23399_, new_n23072_, new_n22802_ );
or   ( new_n23400_, new_n23069_, new_n22811_ );
and  ( new_n23401_, new_n23400_, new_n23399_ );
or   ( new_n23402_, new_n23401_, new_n23077_ );
and  ( new_n23403_, new_n23073_, new_n22812_ );
or   ( new_n23404_, new_n23403_, new_n22822_ );
and  ( new_n23405_, new_n23404_, new_n23402_ );
or   ( new_n23406_, new_n23405_, new_n23398_ );
and  ( new_n23407_, new_n23406_, new_n23397_ );
and  ( new_n23408_, new_n23407_, new_n23382_ );
or   ( new_n23409_, new_n23408_, new_n23381_ );
and  ( new_n23410_, new_n23409_, new_n23218_ );
or   ( new_n23411_, new_n23409_, new_n23218_ );
or   ( new_n23412_, new_n23107_, new_n22857_ );
or   ( new_n23413_, new_n23094_, new_n22888_ );
and  ( new_n23414_, new_n23413_, new_n23412_ );
or   ( new_n23415_, new_n23414_, new_n23112_ );
and  ( new_n23416_, new_n23108_, new_n22889_ );
or   ( new_n23417_, new_n23416_, new_n22897_ );
and  ( new_n23418_, new_n23417_, new_n23415_ );
or   ( new_n23419_, new_n23064_, new_n22760_ );
or   ( new_n23420_, new_n23051_, new_n22791_ );
and  ( new_n23421_, new_n23420_, new_n23419_ );
or   ( new_n23422_, new_n23421_, new_n23079_ );
and  ( new_n23423_, new_n23065_, new_n22792_ );
or   ( new_n23424_, new_n23423_, new_n22824_ );
and  ( new_n23425_, new_n23424_, new_n23422_ );
or   ( new_n23426_, new_n23425_, new_n23418_ );
and  ( new_n23427_, new_n23426_, new_n23411_ );
or   ( new_n23428_, new_n23427_, new_n23410_ );
and  ( new_n23429_, new_n23428_, new_n23197_ );
or   ( new_n23430_, new_n23428_, new_n23197_ );
or   ( new_n23431_, new_n23031_, new_n22971_ );
or   ( new_n23432_, new_n23028_, new_n22978_ );
and  ( new_n23433_, new_n23432_, new_n23431_ );
or   ( new_n23434_, new_n23433_, new_n23036_ );
and  ( new_n23435_, new_n23032_, new_n22979_ );
or   ( new_n23436_, new_n23435_, new_n22987_ );
and  ( new_n23437_, new_n23436_, new_n23434_ );
and  ( new_n23438_, new_n23437_, new_n23430_ );
or   ( new_n23439_, new_n23438_, new_n23429_ );
and  ( new_n23440_, new_n23439_, new_n23172_ );
or   ( new_n23441_, new_n23439_, new_n23172_ );
or   ( new_n23442_, new_n23038_, new_n22964_ );
or   ( new_n23443_, new_n23151_, new_n22989_ );
and  ( new_n23444_, new_n23443_, new_n23442_ );
or   ( new_n23445_, new_n23444_, new_n23156_ );
and  ( new_n23446_, new_n23152_, new_n22990_ );
or   ( new_n23447_, new_n23446_, new_n22998_ );
and  ( new_n23448_, new_n23447_, new_n23445_ );
and  ( new_n23449_, new_n23448_, new_n23441_ );
or   ( new_n23450_, new_n23449_, new_n23440_ );
and  ( new_n23451_, new_n23450_, new_n23165_ );
or   ( new_n23452_, new_n23450_, new_n23165_ );
or   ( new_n23453_, new_n23446_, new_n23156_ );
or   ( new_n23454_, new_n23444_, new_n22998_ );
and  ( new_n23455_, new_n23454_, new_n23453_ );
or   ( new_n23456_, new_n23170_, new_n22698_ );
or   ( new_n23457_, new_n23168_, new_n22538_ );
and  ( new_n23458_, new_n23457_, new_n23456_ );
or   ( new_n23459_, new_n23458_, new_n23439_ );
or   ( new_n23460_, new_n23177_, new_n22610_ );
or   ( new_n23461_, new_n23175_, new_n22414_ );
and  ( new_n23462_, new_n23461_, new_n23460_ );
or   ( new_n23463_, new_n23184_, new_n23142_ );
or   ( new_n23464_, new_n23182_, new_n22951_ );
and  ( new_n23465_, new_n23464_, new_n23463_ );
or   ( new_n23466_, new_n23465_, new_n23462_ );
and  ( new_n23467_, new_n23465_, new_n23462_ );
or   ( new_n23468_, new_n23193_, new_n23129_ );
or   ( new_n23469_, new_n23191_, new_n22926_ );
and  ( new_n23470_, new_n23469_, new_n23468_ );
or   ( new_n23471_, new_n23470_, new_n23467_ );
and  ( new_n23472_, new_n23471_, new_n23466_ );
or   ( new_n23473_, new_n23202_, new_n22593_ );
or   ( new_n23474_, new_n23200_, new_n22379_ );
and  ( new_n23475_, new_n23474_, new_n23473_ );
or   ( new_n23476_, new_n22581_, new_n22578_ );
and  ( new_n23477_, new_n23476_, new_n22350_ );
or   ( new_n23478_, new_n23477_, new_n23475_ );
and  ( new_n23479_, new_n23477_, new_n23475_ );
or   ( new_n23480_, new_n23214_, new_n23127_ );
or   ( new_n23481_, new_n23212_, new_n22924_ );
and  ( new_n23482_, new_n23481_, new_n23480_ );
or   ( new_n23483_, new_n23482_, new_n23479_ );
and  ( new_n23484_, new_n23483_, new_n23478_ );
or   ( new_n23485_, new_n23225_, new_n16505_ );
or   ( new_n23486_, new_n23221_, new_n16438_ );
and  ( new_n23487_, new_n23486_, new_n23485_ );
or   ( new_n23488_, new_n23234_, new_n16085_ );
or   ( new_n23489_, new_n23230_, new_n16048_ );
and  ( new_n23490_, new_n23489_, new_n23488_ );
or   ( new_n23491_, new_n23490_, new_n23487_ );
and  ( new_n23492_, new_n23490_, new_n23487_ );
or   ( new_n23493_, new_n23245_, new_n16052_ );
or   ( new_n23494_, new_n23241_, new_n16071_ );
and  ( new_n23495_, new_n23494_, new_n23493_ );
or   ( new_n23496_, new_n23495_, new_n23492_ );
and  ( new_n23497_, new_n23496_, new_n23491_ );
or   ( new_n23498_, new_n23256_, new_n16009_ );
or   ( new_n23499_, new_n23252_, new_n16029_ );
and  ( new_n23500_, new_n23499_, new_n23498_ );
or   ( new_n23501_, new_n23265_, new_n16186_ );
or   ( new_n23502_, new_n23261_, new_n16204_ );
and  ( new_n23503_, new_n23502_, new_n23501_ );
or   ( new_n23504_, new_n23503_, new_n23500_ );
and  ( new_n23505_, new_n23503_, new_n23500_ );
or   ( new_n23506_, new_n23276_, new_n16217_ );
or   ( new_n23507_, new_n23272_, new_n16234_ );
and  ( new_n23508_, new_n23507_, new_n23506_ );
or   ( new_n23509_, new_n23508_, new_n23505_ );
and  ( new_n23510_, new_n23509_, new_n23504_ );
or   ( new_n23511_, new_n23510_, new_n23497_ );
and  ( new_n23512_, new_n23510_, new_n23497_ );
or   ( new_n23513_, new_n23289_, new_n16108_ );
or   ( new_n23514_, new_n23285_, new_n16128_ );
and  ( new_n23515_, new_n23514_, new_n23513_ );
or   ( new_n23516_, new_n23515_, new_n23512_ );
and  ( new_n23517_, new_n23516_, new_n23511_ );
or   ( new_n23518_, new_n23300_, new_n20156_ );
or   ( new_n23519_, new_n23296_, new_n20443_ );
and  ( new_n23520_, new_n23519_, new_n23518_ );
or   ( new_n23521_, new_n23309_, new_n19394_ );
or   ( new_n23522_, new_n23305_, new_n19659_ );
and  ( new_n23523_, new_n23522_, new_n23521_ );
or   ( new_n23524_, new_n23523_, new_n23520_ );
and  ( new_n23525_, new_n23523_, new_n23520_ );
or   ( new_n23526_, new_n23320_, new_n18742_ );
or   ( new_n23527_, new_n23316_, new_n18977_ );
and  ( new_n23528_, new_n23527_, new_n23526_ );
or   ( new_n23529_, new_n23528_, new_n23525_ );
and  ( new_n23530_, new_n23529_, new_n23524_ );
or   ( new_n23531_, new_n23330_, new_n21261_ );
or   ( new_n23532_, new_n23326_, new_n21009_ );
and  ( new_n23533_, new_n23532_, new_n23531_ );
or   ( new_n23534_, new_n23533_, new_n16108_ );
and  ( new_n23535_, new_n23533_, new_n16108_ );
or   ( new_n23536_, new_n23341_, new_n21013_ );
or   ( new_n23537_, new_n23337_, new_n21265_ );
and  ( new_n23538_, new_n23537_, new_n23536_ );
or   ( new_n23539_, new_n23538_, new_n23535_ );
and  ( new_n23540_, new_n23539_, new_n23534_ );
or   ( new_n23541_, new_n23540_, new_n23530_ );
and  ( new_n23542_, new_n23540_, new_n23530_ );
or   ( new_n23543_, new_n23354_, new_n18066_ );
or   ( new_n23544_, new_n23350_, new_n18309_ );
and  ( new_n23545_, new_n23544_, new_n23543_ );
or   ( new_n23546_, new_n23363_, new_n17238_ );
or   ( new_n23547_, new_n23359_, new_n17650_ );
and  ( new_n23548_, new_n23547_, new_n23546_ );
or   ( new_n23549_, new_n23548_, new_n23545_ );
and  ( new_n23550_, new_n23548_, new_n23545_ );
or   ( new_n23551_, new_n23374_, new_n16814_ );
or   ( new_n23552_, new_n23370_, new_n17142_ );
and  ( new_n23553_, new_n23552_, new_n23551_ );
or   ( new_n23554_, new_n23553_, new_n23550_ );
and  ( new_n23555_, new_n23554_, new_n23549_ );
or   ( new_n23556_, new_n23555_, new_n23542_ );
and  ( new_n23557_, new_n23556_, new_n23541_ );
or   ( new_n23558_, new_n23557_, new_n23517_ );
and  ( new_n23559_, new_n23557_, new_n23517_ );
or   ( new_n23560_, new_n23387_, new_n23105_ );
or   ( new_n23561_, new_n23385_, new_n22886_ );
and  ( new_n23562_, new_n23561_, new_n23560_ );
or   ( new_n23563_, new_n23394_, new_n23092_ );
or   ( new_n23564_, new_n23392_, new_n22855_ );
and  ( new_n23565_, new_n23564_, new_n23563_ );
or   ( new_n23566_, new_n23565_, new_n23562_ );
and  ( new_n23567_, new_n23565_, new_n23562_ );
or   ( new_n23568_, new_n23403_, new_n23077_ );
or   ( new_n23569_, new_n23401_, new_n22822_ );
and  ( new_n23570_, new_n23569_, new_n23568_ );
or   ( new_n23571_, new_n23570_, new_n23567_ );
and  ( new_n23572_, new_n23571_, new_n23566_ );
or   ( new_n23573_, new_n23572_, new_n23559_ );
and  ( new_n23574_, new_n23573_, new_n23558_ );
or   ( new_n23575_, new_n23574_, new_n23484_ );
and  ( new_n23576_, new_n23574_, new_n23484_ );
or   ( new_n23577_, new_n23416_, new_n23112_ );
or   ( new_n23578_, new_n23414_, new_n22897_ );
and  ( new_n23579_, new_n23578_, new_n23577_ );
or   ( new_n23580_, new_n23423_, new_n23079_ );
or   ( new_n23581_, new_n23421_, new_n22824_ );
and  ( new_n23582_, new_n23581_, new_n23580_ );
and  ( new_n23583_, new_n23582_, new_n23579_ );
or   ( new_n23584_, new_n23583_, new_n23576_ );
and  ( new_n23585_, new_n23584_, new_n23575_ );
or   ( new_n23586_, new_n23585_, new_n23472_ );
and  ( new_n23587_, new_n23585_, new_n23472_ );
or   ( new_n23588_, new_n23435_, new_n23036_ );
or   ( new_n23589_, new_n23433_, new_n22987_ );
and  ( new_n23590_, new_n23589_, new_n23588_ );
or   ( new_n23591_, new_n23590_, new_n23587_ );
and  ( new_n23592_, new_n23591_, new_n23586_ );
or   ( new_n23593_, new_n23592_, new_n23172_ );
and  ( new_n23594_, new_n23593_, new_n23459_ );
or   ( new_n23595_, new_n23594_, new_n23455_ );
or   ( new_n23596_, new_n23592_, new_n23458_ );
and  ( new_n23597_, new_n23596_, new_n23441_ );
or   ( new_n23598_, new_n23597_, new_n23448_ );
and  ( new_n23599_, new_n23598_, new_n23595_ );
or   ( new_n23600_, new_n23144_, new_n22928_ );
or   ( new_n23601_, new_n23131_, new_n22953_ );
and  ( new_n23602_, new_n23601_, new_n23600_ );
or   ( new_n23603_, new_n23602_, new_n23149_ );
and  ( new_n23604_, new_n23145_, new_n22954_ );
or   ( new_n23605_, new_n23604_, new_n22962_ );
and  ( new_n23606_, new_n23605_, new_n23603_ );
nor  ( new_n23607_, new_n22333_, new_n612_ );
nor  ( new_n23608_, new_n23607_, new_n8463_ );
or   ( new_n23609_, new_n23608_, new_n21261_ );
and  ( new_n23610_, new_n22337_, RI2b1c4342d648_68 );
and  ( new_n23611_, new_n22330_, RI2b1c4342d5d0_67 );
or   ( new_n23612_, new_n23611_, new_n23610_ );
or   ( new_n23613_, new_n23612_, new_n21009_ );
and  ( new_n23614_, new_n23613_, new_n23609_ );
or   ( new_n23615_, new_n21419_, new_n755_ );
or   ( new_n23616_, new_n21424_, new_n591_ );
and  ( new_n23617_, new_n23616_, new_n23615_ );
or   ( new_n23618_, new_n23617_, new_n21013_ );
and  ( new_n23619_, new_n21428_, RI2b1c4342d738_70 );
and  ( new_n23620_, new_n21415_, RI2b1c4342d6c0_69 );
or   ( new_n23621_, new_n23620_, new_n23619_ );
or   ( new_n23622_, new_n23621_, new_n21265_ );
and  ( new_n23623_, new_n23622_, new_n23618_ );
or   ( new_n23624_, new_n23623_, new_n23614_ );
and  ( new_n23625_, new_n23623_, new_n23614_ );
or   ( new_n23626_, new_n20557_, new_n806_ );
or   ( new_n23627_, new_n20562_, new_n110_ );
and  ( new_n23628_, new_n23627_, new_n23626_ );
or   ( new_n23629_, new_n23628_, new_n20156_ );
and  ( new_n23630_, new_n20566_, RI2b1c4342d828_72 );
and  ( new_n23631_, new_n20553_, RI2b1c4342d7b0_71 );
or   ( new_n23632_, new_n23631_, new_n23630_ );
or   ( new_n23633_, new_n23632_, new_n20443_ );
and  ( new_n23634_, new_n23633_, new_n23629_ );
or   ( new_n23635_, new_n23634_, new_n23625_ );
and  ( new_n23636_, new_n23635_, new_n23624_ );
or   ( new_n23637_, new_n19758_, new_n859_ );
or   ( new_n23638_, new_n19763_, new_n105_ );
and  ( new_n23639_, new_n23638_, new_n23637_ );
or   ( new_n23640_, new_n23639_, new_n19394_ );
and  ( new_n23641_, new_n19767_, RI2b1c4342d918_74 );
and  ( new_n23642_, new_n19754_, RI2b1c4342d8a0_73 );
or   ( new_n23643_, new_n23642_, new_n23641_ );
or   ( new_n23644_, new_n23643_, new_n19659_ );
and  ( new_n23645_, new_n23644_, new_n23640_ );
or   ( new_n23646_, new_n19048_, new_n886_ );
or   ( new_n23647_, new_n19055_, new_n843_ );
and  ( new_n23648_, new_n23647_, new_n23646_ );
or   ( new_n23649_, new_n23648_, new_n18742_ );
and  ( new_n23650_, new_n19057_, RI2b1c4342da08_76 );
and  ( new_n23651_, new_n19044_, RI2b1c4342d990_75 );
or   ( new_n23652_, new_n23651_, new_n23650_ );
or   ( new_n23653_, new_n23652_, new_n18977_ );
and  ( new_n23654_, new_n23653_, new_n23649_ );
or   ( new_n23655_, new_n23654_, new_n23645_ );
and  ( new_n23656_, new_n23654_, new_n23645_ );
or   ( new_n23657_, new_n18388_, new_n1002_ );
or   ( new_n23658_, new_n18395_, new_n1004_ );
and  ( new_n23659_, new_n23658_, new_n23657_ );
or   ( new_n23660_, new_n23659_, new_n18066_ );
and  ( new_n23661_, new_n18397_, RI2b1c4342daf8_78 );
and  ( new_n23662_, new_n18384_, RI2b1c4342da80_77 );
or   ( new_n23663_, new_n23662_, new_n23661_ );
or   ( new_n23664_, new_n23663_, new_n18309_ );
and  ( new_n23665_, new_n23664_, new_n23660_ );
or   ( new_n23666_, new_n23665_, new_n23656_ );
and  ( new_n23667_, new_n23666_, new_n23655_ );
or   ( new_n23668_, new_n23667_, new_n23636_ );
and  ( new_n23669_, new_n23667_, new_n23636_ );
or   ( new_n23670_, new_n17727_, new_n1511_ );
or   ( new_n23671_, new_n17734_, new_n1310_ );
and  ( new_n23672_, new_n23671_, new_n23670_ );
or   ( new_n23673_, new_n23672_, new_n17238_ );
and  ( new_n23674_, new_n17736_, RI2b1c4342dbe8_80 );
and  ( new_n23675_, new_n17723_, RI2b1c4342db70_79 );
or   ( new_n23676_, new_n23675_, new_n23674_ );
or   ( new_n23677_, new_n23676_, new_n17650_ );
and  ( new_n23678_, new_n23677_, new_n23673_ );
or   ( new_n23679_, new_n17244_, new_n2119_ );
or   ( new_n23680_, new_n17248_, new_n126_ );
and  ( new_n23681_, new_n23680_, new_n23679_ );
or   ( new_n23682_, new_n23681_, new_n16814_ );
and  ( new_n23683_, new_n17255_, RI2b1c4342dcd8_82 );
and  ( new_n23684_, new_n17240_, RI2b1c4342dc60_81 );
or   ( new_n23685_, new_n23684_, new_n23683_ );
or   ( new_n23686_, new_n23685_, new_n17142_ );
and  ( new_n23687_, new_n23686_, new_n23682_ );
or   ( new_n23688_, new_n23687_, new_n23678_ );
and  ( new_n23689_, new_n23687_, new_n23678_ );
or   ( new_n23690_, new_n16607_, new_n2541_ );
or   ( new_n23691_, new_n16613_, new_n121_ );
and  ( new_n23692_, new_n23691_, new_n23690_ );
or   ( new_n23693_, new_n23692_, new_n16505_ );
and  ( new_n23694_, new_n16616_, RI2b1c4342ddc8_84 );
and  ( new_n23695_, new_n16603_, RI2b1c4342dd50_83 );
or   ( new_n23696_, new_n23695_, new_n23694_ );
or   ( new_n23697_, new_n23696_, new_n16438_ );
and  ( new_n23698_, new_n23697_, new_n23693_ );
or   ( new_n23699_, new_n23698_, new_n23689_ );
and  ( new_n23700_, new_n23699_, new_n23688_ );
or   ( new_n23701_, new_n23700_, new_n23669_ );
and  ( new_n23702_, new_n23701_, new_n23668_ );
or   ( new_n23703_, new_n16366_, new_n3239_ );
or   ( new_n23704_, new_n16355_, new_n2806_ );
and  ( new_n23705_, new_n23704_, new_n23703_ );
or   ( new_n23706_, new_n23705_, new_n16085_ );
and  ( new_n23707_, new_n16358_, RI2b1c4342deb8_86 );
and  ( new_n23708_, new_n16362_, RI2b1c4342de40_85 );
or   ( new_n23709_, new_n23708_, new_n23707_ );
or   ( new_n23710_, new_n23709_, new_n16048_ );
and  ( new_n23711_, new_n23710_, new_n23706_ );
or   ( new_n23712_, new_n16075_, new_n3902_ );
or   ( new_n23713_, new_n16060_, new_n3924_ );
and  ( new_n23714_, new_n23713_, new_n23712_ );
or   ( new_n23715_, new_n23714_, new_n16052_ );
and  ( new_n23716_, new_n16063_, RI2b1c4342dfa8_88 );
and  ( new_n23717_, new_n16066_, RI2b1c4342df30_87 );
or   ( new_n23718_, new_n23717_, new_n23716_ );
or   ( new_n23719_, new_n23718_, new_n16071_ );
and  ( new_n23720_, new_n23719_, new_n23715_ );
or   ( new_n23721_, new_n23720_, new_n23711_ );
and  ( new_n23722_, new_n23720_, new_n23711_ );
or   ( new_n23723_, new_n16033_, new_n4635_ );
or   ( new_n23724_, new_n16017_, new_n132_ );
and  ( new_n23725_, new_n23724_, new_n23723_ );
or   ( new_n23726_, new_n23725_, new_n16009_ );
and  ( new_n23727_, new_n16021_, RI2b1c4342e098_90 );
and  ( new_n23728_, new_n16024_, RI2b1c4342e020_89 );
or   ( new_n23729_, new_n23728_, new_n23727_ );
or   ( new_n23730_, new_n23729_, new_n16029_ );
and  ( new_n23731_, new_n23730_, new_n23726_ );
or   ( new_n23732_, new_n23731_, new_n23722_ );
and  ( new_n23733_, new_n23732_, new_n23721_ );
or   ( new_n23734_, new_n16208_, new_n5459_ );
or   ( new_n23735_, new_n16194_, new_n117_ );
and  ( new_n23736_, new_n23735_, new_n23734_ );
or   ( new_n23737_, new_n23736_, new_n16186_ );
and  ( new_n23738_, new_n16196_, RI2b1c4342e188_92 );
and  ( new_n23739_, new_n16199_, RI2b1c4342e110_91 );
or   ( new_n23740_, new_n23739_, new_n23738_ );
or   ( new_n23741_, new_n23740_, new_n16204_ );
and  ( new_n23742_, new_n23741_, new_n23737_ );
or   ( new_n23743_, new_n16238_, new_n6321_ );
or   ( new_n23744_, new_n16224_, new_n6307_ );
and  ( new_n23745_, new_n23744_, new_n23743_ );
or   ( new_n23746_, new_n23745_, new_n16217_ );
and  ( new_n23747_, new_n16226_, RI2b1c4342e278_94 );
and  ( new_n23748_, new_n16229_, RI2b1c4342e200_93 );
or   ( new_n23749_, new_n23748_, new_n23747_ );
or   ( new_n23750_, new_n23749_, new_n16234_ );
and  ( new_n23751_, new_n23750_, new_n23746_ );
or   ( new_n23752_, new_n23751_, new_n23742_ );
and  ( new_n23753_, new_n23751_, new_n23742_ );
or   ( new_n23754_, new_n16174_, new_n7274_ );
or   ( new_n23755_, new_n16160_, new_n124_ );
and  ( new_n23756_, new_n23755_, new_n23754_ );
or   ( new_n23757_, new_n23756_, new_n16151_ );
and  ( new_n23758_, new_n16162_, RI2b1c4342e368_96 );
and  ( new_n23759_, new_n16165_, RI2b1c4342e2f0_95 );
or   ( new_n23760_, new_n23759_, new_n23758_ );
or   ( new_n23761_, new_n23760_, new_n16170_ );
and  ( new_n23762_, new_n23761_, new_n23757_ );
or   ( new_n23763_, new_n23762_, new_n23753_ );
and  ( new_n23764_, new_n23763_, new_n23752_ );
or   ( new_n23765_, new_n23764_, new_n23733_ );
and  ( new_n23766_, new_n23764_, new_n23733_ );
or   ( new_n23767_, new_n16174_, new_n124_ );
or   ( new_n23768_, new_n16160_, new_n6321_ );
and  ( new_n23769_, new_n23768_, new_n23767_ );
or   ( new_n23770_, new_n23769_, new_n16151_ );
and  ( new_n23771_, new_n16162_, RI2b1c4342e2f0_95 );
and  ( new_n23772_, new_n16165_, RI2b1c4342e278_94 );
or   ( new_n23773_, new_n23772_, new_n23771_ );
or   ( new_n23774_, new_n23773_, new_n16170_ );
and  ( new_n23775_, new_n23774_, new_n23770_ );
or   ( new_n23776_, new_n23775_, new_n23766_ );
and  ( new_n23777_, new_n23776_, new_n23765_ );
or   ( new_n23778_, new_n23777_, new_n23702_ );
and  ( new_n23779_, new_n23777_, new_n23702_ );
or   ( new_n23780_, new_n16123_, new_n7274_ );
or   ( new_n23781_, new_n23780_, new_n16108_ );
and  ( new_n23782_, new_n16114_, RI2b1c4342e368_96 );
or   ( new_n23783_, new_n23782_, new_n16128_ );
and  ( new_n23784_, new_n23783_, new_n23781_ );
or   ( new_n23785_, new_n23503_, new_n23258_ );
or   ( new_n23786_, new_n23500_, new_n23267_ );
and  ( new_n23787_, new_n23786_, new_n23785_ );
or   ( new_n23788_, new_n23787_, new_n23508_ );
and  ( new_n23789_, new_n23504_, new_n23268_ );
or   ( new_n23790_, new_n23789_, new_n23278_ );
and  ( new_n23791_, new_n23790_, new_n23788_ );
or   ( new_n23792_, new_n23791_, new_n23784_ );
and  ( new_n23793_, new_n23791_, new_n23784_ );
or   ( new_n23794_, new_n23490_, new_n23227_ );
or   ( new_n23795_, new_n23487_, new_n23236_ );
and  ( new_n23796_, new_n23795_, new_n23794_ );
or   ( new_n23797_, new_n23796_, new_n23495_ );
and  ( new_n23798_, new_n23491_, new_n23237_ );
or   ( new_n23799_, new_n23798_, new_n23247_ );
and  ( new_n23800_, new_n23799_, new_n23797_ );
or   ( new_n23801_, new_n23800_, new_n23793_ );
and  ( new_n23802_, new_n23801_, new_n23792_ );
or   ( new_n23803_, new_n23802_, new_n23779_ );
and  ( new_n23804_, new_n23803_, new_n23778_ );
or   ( new_n23805_, new_n23057_, new_n22769_ );
or   ( new_n23806_, new_n23054_, new_n22778_ );
and  ( new_n23807_, new_n23806_, new_n23805_ );
or   ( new_n23808_, new_n23807_, new_n23062_ );
and  ( new_n23809_, new_n23058_, new_n22779_ );
or   ( new_n23810_, new_n23809_, new_n22789_ );
and  ( new_n23811_, new_n23810_, new_n23808_ );
or   ( new_n23812_, new_n23548_, new_n23356_ );
or   ( new_n23813_, new_n23545_, new_n23365_ );
and  ( new_n23814_, new_n23813_, new_n23812_ );
or   ( new_n23815_, new_n23814_, new_n23553_ );
and  ( new_n23816_, new_n23549_, new_n23366_ );
or   ( new_n23817_, new_n23816_, new_n23376_ );
and  ( new_n23818_, new_n23817_, new_n23815_ );
or   ( new_n23819_, new_n23523_, new_n23302_ );
or   ( new_n23820_, new_n23520_, new_n23311_ );
and  ( new_n23821_, new_n23820_, new_n23819_ );
or   ( new_n23822_, new_n23821_, new_n23528_ );
and  ( new_n23823_, new_n23524_, new_n23312_ );
or   ( new_n23824_, new_n23823_, new_n23322_ );
and  ( new_n23825_, new_n23824_, new_n23822_ );
or   ( new_n23826_, new_n23825_, new_n23818_ );
and  ( new_n23827_, new_n23825_, new_n23818_ );
or   ( new_n23828_, new_n23533_, new_n16128_ );
or   ( new_n23829_, new_n23332_, new_n16108_ );
and  ( new_n23830_, new_n23829_, new_n23828_ );
or   ( new_n23831_, new_n23830_, new_n23538_ );
and  ( new_n23832_, new_n23534_, new_n23334_ );
or   ( new_n23833_, new_n23832_, new_n23343_ );
and  ( new_n23834_, new_n23833_, new_n23831_ );
or   ( new_n23835_, new_n23834_, new_n23827_ );
and  ( new_n23836_, new_n23835_, new_n23826_ );
or   ( new_n23837_, new_n23836_, new_n23811_ );
and  ( new_n23838_, new_n23836_, new_n23811_ );
or   ( new_n23839_, new_n23044_, new_n22738_ );
or   ( new_n23840_, new_n23041_, new_n22747_ );
and  ( new_n23841_, new_n23840_, new_n23839_ );
or   ( new_n23842_, new_n23841_, new_n23049_ );
and  ( new_n23843_, new_n23045_, new_n22748_ );
or   ( new_n23844_, new_n23843_, new_n22758_ );
and  ( new_n23845_, new_n23844_, new_n23842_ );
or   ( new_n23846_, new_n23845_, new_n23838_ );
and  ( new_n23847_, new_n23846_, new_n23837_ );
or   ( new_n23848_, new_n23847_, new_n23804_ );
and  ( new_n23849_, new_n23847_, new_n23804_ );
or   ( new_n23850_, new_n23565_, new_n23389_ );
or   ( new_n23851_, new_n23562_, new_n23396_ );
and  ( new_n23852_, new_n23851_, new_n23850_ );
or   ( new_n23853_, new_n23852_, new_n23570_ );
and  ( new_n23854_, new_n23566_, new_n23397_ );
or   ( new_n23855_, new_n23854_, new_n23405_ );
and  ( new_n23856_, new_n23855_, new_n23853_ );
or   ( new_n23857_, new_n23510_, new_n23249_ );
or   ( new_n23858_, new_n23497_, new_n23280_ );
and  ( new_n23859_, new_n23858_, new_n23857_ );
or   ( new_n23860_, new_n23859_, new_n23515_ );
and  ( new_n23861_, new_n23511_, new_n23281_ );
or   ( new_n23862_, new_n23861_, new_n23291_ );
and  ( new_n23863_, new_n23862_, new_n23860_ );
or   ( new_n23864_, new_n23863_, new_n23856_ );
and  ( new_n23865_, new_n23863_, new_n23856_ );
or   ( new_n23866_, new_n23530_, new_n23345_ );
or   ( new_n23867_, new_n23540_, new_n23324_ );
and  ( new_n23868_, new_n23867_, new_n23866_ );
or   ( new_n23869_, new_n23868_, new_n23555_ );
and  ( new_n23870_, new_n23541_, new_n23347_ );
or   ( new_n23871_, new_n23870_, new_n23378_ );
and  ( new_n23872_, new_n23871_, new_n23869_ );
or   ( new_n23873_, new_n23872_, new_n23865_ );
and  ( new_n23874_, new_n23873_, new_n23864_ );
or   ( new_n23875_, new_n23874_, new_n23849_ );
and  ( new_n23876_, new_n23875_, new_n23848_ );
or   ( new_n23877_, new_n23582_, new_n23418_ );
or   ( new_n23878_, new_n23579_, new_n23425_ );
and  ( new_n23879_, new_n23878_, new_n23877_ );
or   ( new_n23880_, new_n23477_, new_n23204_ );
or   ( new_n23881_, new_n23475_, new_n23207_ );
and  ( new_n23882_, new_n23881_, new_n23880_ );
or   ( new_n23883_, new_n23882_, new_n23482_ );
and  ( new_n23884_, new_n23478_, new_n23208_ );
or   ( new_n23885_, new_n23884_, new_n23216_ );
and  ( new_n23886_, new_n23885_, new_n23883_ );
or   ( new_n23887_, new_n23886_, new_n23879_ );
and  ( new_n23888_, new_n23886_, new_n23879_ );
or   ( new_n23889_, new_n23517_, new_n23380_ );
or   ( new_n23890_, new_n23557_, new_n23293_ );
and  ( new_n23891_, new_n23890_, new_n23889_ );
or   ( new_n23892_, new_n23891_, new_n23572_ );
and  ( new_n23893_, new_n23558_, new_n23382_ );
or   ( new_n23894_, new_n23893_, new_n23407_ );
and  ( new_n23895_, new_n23894_, new_n23892_ );
or   ( new_n23896_, new_n23895_, new_n23888_ );
and  ( new_n23897_, new_n23896_, new_n23887_ );
or   ( new_n23898_, new_n23897_, new_n23876_ );
and  ( new_n23899_, new_n23897_, new_n23876_ );
or   ( new_n23900_, new_n23465_, new_n23179_ );
or   ( new_n23901_, new_n23462_, new_n23186_ );
and  ( new_n23902_, new_n23901_, new_n23900_ );
or   ( new_n23903_, new_n23902_, new_n23470_ );
and  ( new_n23904_, new_n23466_, new_n23187_ );
or   ( new_n23905_, new_n23904_, new_n23195_ );
and  ( new_n23906_, new_n23905_, new_n23903_ );
or   ( new_n23907_, new_n23906_, new_n23899_ );
and  ( new_n23908_, new_n23907_, new_n23898_ );
or   ( new_n23909_, new_n23908_, new_n23606_ );
or   ( new_n23910_, new_n23472_, new_n23428_ );
or   ( new_n23911_, new_n23585_, new_n23197_ );
and  ( new_n23912_, new_n23911_, new_n23910_ );
or   ( new_n23913_, new_n23912_, new_n23590_ );
and  ( new_n23914_, new_n23586_, new_n23430_ );
or   ( new_n23915_, new_n23914_, new_n23437_ );
and  ( new_n23916_, new_n23915_, new_n23913_ );
and  ( new_n23917_, new_n23908_, new_n23606_ );
or   ( new_n23918_, new_n23917_, new_n23916_ );
and  ( new_n23919_, new_n23918_, new_n23909_ );
or   ( new_n23920_, new_n23919_, new_n23599_ );
and  ( new_n23921_, new_n23920_, new_n23452_ );
or   ( new_n23922_, new_n23921_, new_n23451_ );
and  ( new_n23923_, new_n23919_, new_n23599_ );
or   ( new_n23924_, new_n23923_, new_n23451_ );
or   ( new_n23925_, new_n23914_, new_n23590_ );
or   ( new_n23926_, new_n23912_, new_n23437_ );
and  ( new_n23927_, new_n23926_, new_n23925_ );
or   ( new_n23928_, new_n23604_, new_n23149_ );
or   ( new_n23929_, new_n23602_, new_n22962_ );
and  ( new_n23930_, new_n23929_, new_n23928_ );
or   ( new_n23931_, new_n23930_, new_n23908_ );
or   ( new_n23932_, new_n23621_, new_n21013_ );
or   ( new_n23933_, new_n23617_, new_n21265_ );
and  ( new_n23934_, new_n23933_, new_n23932_ );
or   ( new_n23935_, new_n23612_, new_n21261_ );
or   ( new_n23936_, new_n23608_, new_n21009_ );
and  ( new_n23937_, new_n23936_, new_n23935_ );
or   ( new_n23938_, new_n23937_, new_n23934_ );
and  ( new_n23939_, new_n23937_, new_n23934_ );
or   ( new_n23940_, new_n23632_, new_n20156_ );
or   ( new_n23941_, new_n23628_, new_n20443_ );
and  ( new_n23942_, new_n23941_, new_n23940_ );
or   ( new_n23943_, new_n23942_, new_n23939_ );
and  ( new_n23944_, new_n23943_, new_n23938_ );
or   ( new_n23945_, new_n23643_, new_n19394_ );
or   ( new_n23946_, new_n23639_, new_n19659_ );
and  ( new_n23947_, new_n23946_, new_n23945_ );
or   ( new_n23948_, new_n23652_, new_n18742_ );
or   ( new_n23949_, new_n23648_, new_n18977_ );
and  ( new_n23950_, new_n23949_, new_n23948_ );
or   ( new_n23951_, new_n23950_, new_n23947_ );
and  ( new_n23952_, new_n23950_, new_n23947_ );
or   ( new_n23953_, new_n23663_, new_n18066_ );
or   ( new_n23954_, new_n23659_, new_n18309_ );
and  ( new_n23955_, new_n23954_, new_n23953_ );
or   ( new_n23956_, new_n23955_, new_n23952_ );
and  ( new_n23957_, new_n23956_, new_n23951_ );
or   ( new_n23958_, new_n23957_, new_n23944_ );
and  ( new_n23959_, new_n23957_, new_n23944_ );
or   ( new_n23960_, new_n23676_, new_n17238_ );
or   ( new_n23961_, new_n23672_, new_n17650_ );
and  ( new_n23962_, new_n23961_, new_n23960_ );
or   ( new_n23963_, new_n23685_, new_n16814_ );
or   ( new_n23964_, new_n23681_, new_n17142_ );
and  ( new_n23965_, new_n23964_, new_n23963_ );
or   ( new_n23966_, new_n23965_, new_n23962_ );
and  ( new_n23967_, new_n23965_, new_n23962_ );
or   ( new_n23968_, new_n23696_, new_n16505_ );
or   ( new_n23969_, new_n23692_, new_n16438_ );
and  ( new_n23970_, new_n23969_, new_n23968_ );
or   ( new_n23971_, new_n23970_, new_n23967_ );
and  ( new_n23972_, new_n23971_, new_n23966_ );
or   ( new_n23973_, new_n23972_, new_n23959_ );
and  ( new_n23974_, new_n23973_, new_n23958_ );
or   ( new_n23975_, new_n23709_, new_n16085_ );
or   ( new_n23976_, new_n23705_, new_n16048_ );
and  ( new_n23977_, new_n23976_, new_n23975_ );
or   ( new_n23978_, new_n23718_, new_n16052_ );
or   ( new_n23979_, new_n23714_, new_n16071_ );
and  ( new_n23980_, new_n23979_, new_n23978_ );
or   ( new_n23981_, new_n23980_, new_n23977_ );
and  ( new_n23982_, new_n23980_, new_n23977_ );
or   ( new_n23983_, new_n23729_, new_n16009_ );
or   ( new_n23984_, new_n23725_, new_n16029_ );
and  ( new_n23985_, new_n23984_, new_n23983_ );
or   ( new_n23986_, new_n23985_, new_n23982_ );
and  ( new_n23987_, new_n23986_, new_n23981_ );
or   ( new_n23988_, new_n23740_, new_n16186_ );
or   ( new_n23989_, new_n23736_, new_n16204_ );
and  ( new_n23990_, new_n23989_, new_n23988_ );
or   ( new_n23991_, new_n23749_, new_n16217_ );
or   ( new_n23992_, new_n23745_, new_n16234_ );
and  ( new_n23993_, new_n23992_, new_n23991_ );
or   ( new_n23994_, new_n23993_, new_n23990_ );
and  ( new_n23995_, new_n23993_, new_n23990_ );
or   ( new_n23996_, new_n23760_, new_n16151_ );
or   ( new_n23997_, new_n23756_, new_n16170_ );
and  ( new_n23998_, new_n23997_, new_n23996_ );
or   ( new_n23999_, new_n23998_, new_n23995_ );
and  ( new_n24000_, new_n23999_, new_n23994_ );
or   ( new_n24001_, new_n24000_, new_n23987_ );
and  ( new_n24002_, new_n24000_, new_n23987_ );
or   ( new_n24003_, new_n23773_, new_n16151_ );
or   ( new_n24004_, new_n23769_, new_n16170_ );
and  ( new_n24005_, new_n24004_, new_n24003_ );
or   ( new_n24006_, new_n24005_, new_n24002_ );
and  ( new_n24007_, new_n24006_, new_n24001_ );
or   ( new_n24008_, new_n24007_, new_n23974_ );
and  ( new_n24009_, new_n24007_, new_n23974_ );
or   ( new_n24010_, new_n23782_, new_n16108_ );
or   ( new_n24011_, new_n23780_, new_n16128_ );
and  ( new_n24012_, new_n24011_, new_n24010_ );
or   ( new_n24013_, new_n23789_, new_n23508_ );
or   ( new_n24014_, new_n23787_, new_n23278_ );
and  ( new_n24015_, new_n24014_, new_n24013_ );
or   ( new_n24016_, new_n24015_, new_n24012_ );
and  ( new_n24017_, new_n24015_, new_n24012_ );
or   ( new_n24018_, new_n23798_, new_n23495_ );
or   ( new_n24019_, new_n23796_, new_n23247_ );
and  ( new_n24020_, new_n24019_, new_n24018_ );
or   ( new_n24021_, new_n24020_, new_n24017_ );
and  ( new_n24022_, new_n24021_, new_n24016_ );
or   ( new_n24023_, new_n24022_, new_n24009_ );
and  ( new_n24024_, new_n24023_, new_n24008_ );
or   ( new_n24025_, new_n23809_, new_n23062_ );
or   ( new_n24026_, new_n23807_, new_n22789_ );
and  ( new_n24027_, new_n24026_, new_n24025_ );
or   ( new_n24028_, new_n23816_, new_n23553_ );
or   ( new_n24029_, new_n23814_, new_n23376_ );
and  ( new_n24030_, new_n24029_, new_n24028_ );
or   ( new_n24031_, new_n23823_, new_n23528_ );
or   ( new_n24032_, new_n23821_, new_n23322_ );
and  ( new_n24033_, new_n24032_, new_n24031_ );
or   ( new_n24034_, new_n24033_, new_n24030_ );
and  ( new_n24035_, new_n24033_, new_n24030_ );
or   ( new_n24036_, new_n23832_, new_n23538_ );
or   ( new_n24037_, new_n23830_, new_n23343_ );
and  ( new_n24038_, new_n24037_, new_n24036_ );
or   ( new_n24039_, new_n24038_, new_n24035_ );
and  ( new_n24040_, new_n24039_, new_n24034_ );
or   ( new_n24041_, new_n24040_, new_n24027_ );
and  ( new_n24042_, new_n24040_, new_n24027_ );
or   ( new_n24043_, new_n23843_, new_n23049_ );
or   ( new_n24044_, new_n23841_, new_n22758_ );
and  ( new_n24045_, new_n24044_, new_n24043_ );
or   ( new_n24046_, new_n24045_, new_n24042_ );
and  ( new_n24047_, new_n24046_, new_n24041_ );
or   ( new_n24048_, new_n24047_, new_n24024_ );
and  ( new_n24049_, new_n24047_, new_n24024_ );
or   ( new_n24050_, new_n23854_, new_n23570_ );
or   ( new_n24051_, new_n23852_, new_n23405_ );
and  ( new_n24052_, new_n24051_, new_n24050_ );
or   ( new_n24053_, new_n23861_, new_n23515_ );
or   ( new_n24054_, new_n23859_, new_n23291_ );
and  ( new_n24055_, new_n24054_, new_n24053_ );
or   ( new_n24056_, new_n24055_, new_n24052_ );
and  ( new_n24057_, new_n24055_, new_n24052_ );
or   ( new_n24058_, new_n23870_, new_n23555_ );
or   ( new_n24059_, new_n23868_, new_n23378_ );
and  ( new_n24060_, new_n24059_, new_n24058_ );
or   ( new_n24061_, new_n24060_, new_n24057_ );
and  ( new_n24062_, new_n24061_, new_n24056_ );
or   ( new_n24063_, new_n24062_, new_n24049_ );
and  ( new_n24064_, new_n24063_, new_n24048_ );
or   ( new_n24065_, new_n23582_, new_n23579_ );
and  ( new_n24066_, new_n24065_, new_n23426_ );
or   ( new_n24067_, new_n23884_, new_n23482_ );
or   ( new_n24068_, new_n23882_, new_n23216_ );
and  ( new_n24069_, new_n24068_, new_n24067_ );
or   ( new_n24070_, new_n24069_, new_n24066_ );
and  ( new_n24071_, new_n24069_, new_n24066_ );
or   ( new_n24072_, new_n23893_, new_n23572_ );
or   ( new_n24073_, new_n23891_, new_n23407_ );
and  ( new_n24074_, new_n24073_, new_n24072_ );
or   ( new_n24075_, new_n24074_, new_n24071_ );
and  ( new_n24076_, new_n24075_, new_n24070_ );
or   ( new_n24077_, new_n24076_, new_n24064_ );
and  ( new_n24078_, new_n24076_, new_n24064_ );
or   ( new_n24079_, new_n23904_, new_n23470_ );
or   ( new_n24080_, new_n23902_, new_n23195_ );
and  ( new_n24081_, new_n24080_, new_n24079_ );
or   ( new_n24082_, new_n24081_, new_n24078_ );
and  ( new_n24083_, new_n24082_, new_n24077_ );
or   ( new_n24084_, new_n24083_, new_n23606_ );
and  ( new_n24085_, new_n24084_, new_n23931_ );
or   ( new_n24086_, new_n24085_, new_n23927_ );
or   ( new_n24087_, new_n24083_, new_n23930_ );
and  ( new_n24088_, new_n24087_, new_n23909_ );
or   ( new_n24089_, new_n24088_, new_n23916_ );
and  ( new_n24090_, new_n24089_, new_n24086_ );
or   ( new_n24091_, new_n23484_, new_n23409_ );
or   ( new_n24092_, new_n23574_, new_n23218_ );
and  ( new_n24093_, new_n24092_, new_n24091_ );
or   ( new_n24094_, new_n24093_, new_n23583_ );
and  ( new_n24095_, new_n23575_, new_n23411_ );
or   ( new_n24096_, new_n24095_, new_n23426_ );
and  ( new_n24097_, new_n24096_, new_n24094_ );
or   ( new_n24098_, new_n24027_, new_n23836_ );
or   ( new_n24099_, new_n24040_, new_n23811_ );
and  ( new_n24100_, new_n24099_, new_n24098_ );
or   ( new_n24101_, new_n24100_, new_n24045_ );
and  ( new_n24102_, new_n24041_, new_n23837_ );
or   ( new_n24103_, new_n24102_, new_n23845_ );
and  ( new_n24104_, new_n24103_, new_n24101_ );
or   ( new_n24105_, new_n24007_, new_n23702_ );
or   ( new_n24106_, new_n23974_, new_n23777_ );
and  ( new_n24107_, new_n24106_, new_n24105_ );
or   ( new_n24108_, new_n24107_, new_n24022_ );
and  ( new_n24109_, new_n24008_, new_n23778_ );
or   ( new_n24110_, new_n24109_, new_n23802_ );
and  ( new_n24111_, new_n24110_, new_n24108_ );
or   ( new_n24112_, new_n24111_, new_n24104_ );
or   ( new_n24113_, new_n24033_, new_n23818_ );
or   ( new_n24114_, new_n24030_, new_n23825_ );
and  ( new_n24115_, new_n24114_, new_n24113_ );
or   ( new_n24116_, new_n24115_, new_n24038_ );
and  ( new_n24117_, new_n24034_, new_n23826_ );
or   ( new_n24118_, new_n24117_, new_n23834_ );
and  ( new_n24119_, new_n24118_, new_n24116_ );
or   ( new_n24120_, new_n24015_, new_n23784_ );
or   ( new_n24121_, new_n24012_, new_n23791_ );
and  ( new_n24122_, new_n24121_, new_n24120_ );
or   ( new_n24123_, new_n24122_, new_n24020_ );
and  ( new_n24124_, new_n24016_, new_n23792_ );
or   ( new_n24125_, new_n24124_, new_n23800_ );
and  ( new_n24126_, new_n24125_, new_n24123_ );
or   ( new_n24127_, new_n24126_, new_n24119_ );
and  ( new_n24128_, new_n24126_, new_n24119_ );
or   ( new_n24129_, new_n24000_, new_n23733_ );
or   ( new_n24130_, new_n23987_, new_n23764_ );
and  ( new_n24131_, new_n24130_, new_n24129_ );
or   ( new_n24132_, new_n24131_, new_n24005_ );
and  ( new_n24133_, new_n24001_, new_n23765_ );
or   ( new_n24134_, new_n24133_, new_n23775_ );
and  ( new_n24135_, new_n24134_, new_n24132_ );
or   ( new_n24136_, new_n24135_, new_n24128_ );
and  ( new_n24137_, new_n24136_, new_n24127_ );
or   ( new_n24138_, new_n16607_, new_n2806_ );
or   ( new_n24139_, new_n16613_, new_n2541_ );
and  ( new_n24140_, new_n24139_, new_n24138_ );
or   ( new_n24141_, new_n24140_, new_n16505_ );
and  ( new_n24142_, new_n16616_, RI2b1c4342de40_85 );
and  ( new_n24143_, new_n16603_, RI2b1c4342ddc8_84 );
or   ( new_n24144_, new_n24143_, new_n24142_ );
or   ( new_n24145_, new_n24144_, new_n16438_ );
and  ( new_n24146_, new_n24145_, new_n24141_ );
or   ( new_n24147_, new_n16366_, new_n3924_ );
or   ( new_n24148_, new_n16355_, new_n3239_ );
and  ( new_n24149_, new_n24148_, new_n24147_ );
or   ( new_n24150_, new_n24149_, new_n16085_ );
and  ( new_n24151_, new_n16358_, RI2b1c4342df30_87 );
and  ( new_n24152_, new_n16362_, RI2b1c4342deb8_86 );
or   ( new_n24153_, new_n24152_, new_n24151_ );
or   ( new_n24154_, new_n24153_, new_n16048_ );
and  ( new_n24155_, new_n24154_, new_n24150_ );
or   ( new_n24156_, new_n24155_, new_n24146_ );
and  ( new_n24157_, new_n24155_, new_n24146_ );
or   ( new_n24158_, new_n16075_, new_n132_ );
or   ( new_n24159_, new_n16060_, new_n3902_ );
and  ( new_n24160_, new_n24159_, new_n24158_ );
or   ( new_n24161_, new_n24160_, new_n16052_ );
and  ( new_n24162_, new_n16063_, RI2b1c4342e020_89 );
and  ( new_n24163_, new_n16066_, RI2b1c4342dfa8_88 );
or   ( new_n24164_, new_n24163_, new_n24162_ );
or   ( new_n24165_, new_n24164_, new_n16071_ );
and  ( new_n24166_, new_n24165_, new_n24161_ );
or   ( new_n24167_, new_n24166_, new_n24157_ );
and  ( new_n24168_, new_n24167_, new_n24156_ );
or   ( new_n24169_, new_n16033_, new_n117_ );
or   ( new_n24170_, new_n16017_, new_n4635_ );
and  ( new_n24171_, new_n24170_, new_n24169_ );
or   ( new_n24172_, new_n24171_, new_n16009_ );
and  ( new_n24173_, new_n16021_, RI2b1c4342e110_91 );
and  ( new_n24174_, new_n16024_, RI2b1c4342e098_90 );
or   ( new_n24175_, new_n24174_, new_n24173_ );
or   ( new_n24176_, new_n24175_, new_n16029_ );
and  ( new_n24177_, new_n24176_, new_n24172_ );
or   ( new_n24178_, new_n16208_, new_n6307_ );
or   ( new_n24179_, new_n16194_, new_n5459_ );
and  ( new_n24180_, new_n24179_, new_n24178_ );
or   ( new_n24181_, new_n24180_, new_n16186_ );
and  ( new_n24182_, new_n16196_, RI2b1c4342e200_93 );
and  ( new_n24183_, new_n16199_, RI2b1c4342e188_92 );
or   ( new_n24184_, new_n24183_, new_n24182_ );
or   ( new_n24185_, new_n24184_, new_n16204_ );
and  ( new_n24186_, new_n24185_, new_n24181_ );
or   ( new_n24187_, new_n24186_, new_n24177_ );
and  ( new_n24188_, new_n24186_, new_n24177_ );
or   ( new_n24189_, new_n16238_, new_n124_ );
or   ( new_n24190_, new_n16224_, new_n6321_ );
and  ( new_n24191_, new_n24190_, new_n24189_ );
or   ( new_n24192_, new_n24191_, new_n16217_ );
and  ( new_n24193_, new_n16226_, RI2b1c4342e2f0_95 );
and  ( new_n24194_, new_n16229_, RI2b1c4342e278_94 );
or   ( new_n24195_, new_n24194_, new_n24193_ );
or   ( new_n24196_, new_n24195_, new_n16234_ );
and  ( new_n24197_, new_n24196_, new_n24192_ );
or   ( new_n24198_, new_n24197_, new_n24188_ );
and  ( new_n24199_, new_n24198_, new_n24187_ );
or   ( new_n24200_, new_n24199_, new_n24168_ );
and  ( new_n24201_, new_n24199_, new_n24168_ );
or   ( new_n24202_, new_n23993_, new_n23742_ );
or   ( new_n24203_, new_n23990_, new_n23751_ );
and  ( new_n24204_, new_n24203_, new_n24202_ );
or   ( new_n24205_, new_n24204_, new_n23998_ );
and  ( new_n24206_, new_n23994_, new_n23752_ );
or   ( new_n24207_, new_n24206_, new_n23762_ );
and  ( new_n24208_, new_n24207_, new_n24205_ );
or   ( new_n24209_, new_n24208_, new_n24201_ );
and  ( new_n24210_, new_n24209_, new_n24200_ );
or   ( new_n24211_, new_n20557_, new_n105_ );
or   ( new_n24212_, new_n20562_, new_n806_ );
and  ( new_n24213_, new_n24212_, new_n24211_ );
or   ( new_n24214_, new_n24213_, new_n20156_ );
and  ( new_n24215_, new_n20566_, RI2b1c4342d8a0_73 );
and  ( new_n24216_, new_n20553_, RI2b1c4342d828_72 );
or   ( new_n24217_, new_n24216_, new_n24215_ );
or   ( new_n24218_, new_n24217_, new_n20443_ );
and  ( new_n24219_, new_n24218_, new_n24214_ );
or   ( new_n24220_, new_n19758_, new_n843_ );
or   ( new_n24221_, new_n19763_, new_n859_ );
and  ( new_n24222_, new_n24221_, new_n24220_ );
or   ( new_n24223_, new_n24222_, new_n19394_ );
and  ( new_n24224_, new_n19767_, RI2b1c4342d990_75 );
and  ( new_n24225_, new_n19754_, RI2b1c4342d918_74 );
or   ( new_n24226_, new_n24225_, new_n24224_ );
or   ( new_n24227_, new_n24226_, new_n19659_ );
and  ( new_n24228_, new_n24227_, new_n24223_ );
or   ( new_n24229_, new_n24228_, new_n24219_ );
and  ( new_n24230_, new_n24228_, new_n24219_ );
or   ( new_n24231_, new_n19048_, new_n1004_ );
or   ( new_n24232_, new_n19055_, new_n886_ );
and  ( new_n24233_, new_n24232_, new_n24231_ );
or   ( new_n24234_, new_n24233_, new_n18742_ );
and  ( new_n24235_, new_n19057_, RI2b1c4342da80_77 );
and  ( new_n24236_, new_n19044_, RI2b1c4342da08_76 );
or   ( new_n24237_, new_n24236_, new_n24235_ );
or   ( new_n24238_, new_n24237_, new_n18977_ );
and  ( new_n24239_, new_n24238_, new_n24234_ );
or   ( new_n24240_, new_n24239_, new_n24230_ );
and  ( new_n24241_, new_n24240_, new_n24229_ );
nor  ( new_n24242_, new_n22333_, new_n591_ );
nor  ( new_n24243_, new_n24242_, new_n9090_ );
or   ( new_n24244_, new_n24243_, new_n21261_ );
and  ( new_n24245_, new_n22337_, RI2b1c4342d6c0_69 );
and  ( new_n24246_, new_n22330_, RI2b1c4342d648_68 );
or   ( new_n24247_, new_n24246_, new_n24245_ );
or   ( new_n24248_, new_n24247_, new_n21009_ );
and  ( new_n24249_, new_n24248_, new_n24244_ );
and  ( new_n24250_, new_n24249_, new_n16170_ );
or   ( new_n24251_, new_n24249_, new_n16170_ );
or   ( new_n24252_, new_n21419_, new_n110_ );
or   ( new_n24253_, new_n21424_, new_n755_ );
and  ( new_n24254_, new_n24253_, new_n24252_ );
or   ( new_n24255_, new_n24254_, new_n21013_ );
and  ( new_n24256_, new_n21428_, RI2b1c4342d7b0_71 );
and  ( new_n24257_, new_n21415_, RI2b1c4342d738_70 );
or   ( new_n24258_, new_n24257_, new_n24256_ );
or   ( new_n24259_, new_n24258_, new_n21265_ );
and  ( new_n24260_, new_n24259_, new_n24255_ );
and  ( new_n24261_, new_n24260_, new_n24251_ );
or   ( new_n24262_, new_n24261_, new_n24250_ );
and  ( new_n24263_, new_n24262_, new_n24241_ );
or   ( new_n24264_, new_n24262_, new_n24241_ );
or   ( new_n24265_, new_n18388_, new_n1310_ );
or   ( new_n24266_, new_n18395_, new_n1002_ );
and  ( new_n24267_, new_n24266_, new_n24265_ );
or   ( new_n24268_, new_n24267_, new_n18066_ );
and  ( new_n24269_, new_n18397_, RI2b1c4342db70_79 );
and  ( new_n24270_, new_n18384_, RI2b1c4342daf8_78 );
or   ( new_n24271_, new_n24270_, new_n24269_ );
or   ( new_n24272_, new_n24271_, new_n18309_ );
and  ( new_n24273_, new_n24272_, new_n24268_ );
or   ( new_n24274_, new_n17727_, new_n126_ );
or   ( new_n24275_, new_n17734_, new_n1511_ );
and  ( new_n24276_, new_n24275_, new_n24274_ );
or   ( new_n24277_, new_n24276_, new_n17238_ );
and  ( new_n24278_, new_n17736_, RI2b1c4342dc60_81 );
and  ( new_n24279_, new_n17723_, RI2b1c4342dbe8_80 );
or   ( new_n24280_, new_n24279_, new_n24278_ );
or   ( new_n24281_, new_n24280_, new_n17650_ );
and  ( new_n24282_, new_n24281_, new_n24277_ );
or   ( new_n24283_, new_n24282_, new_n24273_ );
and  ( new_n24284_, new_n24282_, new_n24273_ );
or   ( new_n24285_, new_n17244_, new_n121_ );
or   ( new_n24286_, new_n17248_, new_n2119_ );
and  ( new_n24287_, new_n24286_, new_n24285_ );
or   ( new_n24288_, new_n24287_, new_n16814_ );
and  ( new_n24289_, new_n17255_, RI2b1c4342dd50_83 );
and  ( new_n24290_, new_n17240_, RI2b1c4342dcd8_82 );
or   ( new_n24291_, new_n24290_, new_n24289_ );
or   ( new_n24292_, new_n24291_, new_n17142_ );
and  ( new_n24293_, new_n24292_, new_n24288_ );
or   ( new_n24294_, new_n24293_, new_n24284_ );
and  ( new_n24295_, new_n24294_, new_n24283_ );
and  ( new_n24296_, new_n24295_, new_n24264_ );
or   ( new_n24297_, new_n24296_, new_n24263_ );
and  ( new_n24298_, new_n24297_, new_n24210_ );
or   ( new_n24299_, new_n24297_, new_n24210_ );
or   ( new_n24300_, new_n23980_, new_n23711_ );
or   ( new_n24301_, new_n23977_, new_n23720_ );
and  ( new_n24302_, new_n24301_, new_n24300_ );
or   ( new_n24303_, new_n24302_, new_n23985_ );
and  ( new_n24304_, new_n23981_, new_n23721_ );
or   ( new_n24305_, new_n24304_, new_n23731_ );
and  ( new_n24306_, new_n24305_, new_n24303_ );
or   ( new_n24307_, new_n23965_, new_n23678_ );
or   ( new_n24308_, new_n23962_, new_n23687_ );
and  ( new_n24309_, new_n24308_, new_n24307_ );
or   ( new_n24310_, new_n24309_, new_n23970_ );
and  ( new_n24311_, new_n23966_, new_n23688_ );
or   ( new_n24312_, new_n24311_, new_n23698_ );
and  ( new_n24313_, new_n24312_, new_n24310_ );
or   ( new_n24314_, new_n24313_, new_n24306_ );
and  ( new_n24315_, new_n24313_, new_n24306_ );
or   ( new_n24316_, new_n23950_, new_n23645_ );
or   ( new_n24317_, new_n23947_, new_n23654_ );
and  ( new_n24318_, new_n24317_, new_n24316_ );
or   ( new_n24319_, new_n24318_, new_n23955_ );
and  ( new_n24320_, new_n23951_, new_n23655_ );
or   ( new_n24321_, new_n24320_, new_n23665_ );
and  ( new_n24322_, new_n24321_, new_n24319_ );
or   ( new_n24323_, new_n24322_, new_n24315_ );
and  ( new_n24324_, new_n24323_, new_n24314_ );
and  ( new_n24325_, new_n24324_, new_n24299_ );
or   ( new_n24326_, new_n24325_, new_n24298_ );
and  ( new_n24327_, new_n24326_, new_n24137_ );
or   ( new_n24328_, new_n24326_, new_n24137_ );
or   ( new_n24329_, new_n24055_, new_n23856_ );
or   ( new_n24330_, new_n24052_, new_n23863_ );
and  ( new_n24331_, new_n24330_, new_n24329_ );
or   ( new_n24332_, new_n24331_, new_n24060_ );
and  ( new_n24333_, new_n24056_, new_n23864_ );
or   ( new_n24334_, new_n24333_, new_n23872_ );
and  ( new_n24335_, new_n24334_, new_n24332_ );
and  ( new_n24336_, new_n24335_, new_n24328_ );
or   ( new_n24337_, new_n24336_, new_n24327_ );
and  ( new_n24338_, new_n24337_, new_n24112_ );
or   ( new_n24339_, new_n24337_, new_n24112_ );
or   ( new_n24340_, new_n24069_, new_n23879_ );
or   ( new_n24341_, new_n24066_, new_n23886_ );
and  ( new_n24342_, new_n24341_, new_n24340_ );
or   ( new_n24343_, new_n24342_, new_n24074_ );
and  ( new_n24344_, new_n24070_, new_n23887_ );
or   ( new_n24345_, new_n24344_, new_n23895_ );
and  ( new_n24346_, new_n24345_, new_n24343_ );
and  ( new_n24347_, new_n24346_, new_n24339_ );
or   ( new_n24348_, new_n24347_, new_n24338_ );
and  ( new_n24349_, new_n24348_, new_n24097_ );
or   ( new_n24350_, new_n24348_, new_n24097_ );
or   ( new_n24351_, new_n24076_, new_n23876_ );
or   ( new_n24352_, new_n24064_, new_n23897_ );
and  ( new_n24353_, new_n24352_, new_n24351_ );
or   ( new_n24354_, new_n24353_, new_n24081_ );
and  ( new_n24355_, new_n24077_, new_n23898_ );
or   ( new_n24356_, new_n24355_, new_n23906_ );
and  ( new_n24357_, new_n24356_, new_n24354_ );
and  ( new_n24358_, new_n24357_, new_n24350_ );
or   ( new_n24359_, new_n24358_, new_n24349_ );
and  ( new_n24360_, new_n24359_, new_n24090_ );
or   ( new_n24361_, new_n24359_, new_n24090_ );
or   ( new_n24362_, new_n24355_, new_n24081_ );
or   ( new_n24363_, new_n24353_, new_n23906_ );
and  ( new_n24364_, new_n24363_, new_n24362_ );
or   ( new_n24365_, new_n24095_, new_n23583_ );
or   ( new_n24366_, new_n24093_, new_n23426_ );
and  ( new_n24367_, new_n24366_, new_n24365_ );
or   ( new_n24368_, new_n24367_, new_n24348_ );
or   ( new_n24369_, new_n24102_, new_n24045_ );
or   ( new_n24370_, new_n24100_, new_n23845_ );
and  ( new_n24371_, new_n24370_, new_n24369_ );
or   ( new_n24372_, new_n24109_, new_n24022_ );
or   ( new_n24373_, new_n24107_, new_n23802_ );
and  ( new_n24374_, new_n24373_, new_n24372_ );
and  ( new_n24375_, new_n24374_, new_n24371_ );
or   ( new_n24376_, new_n24117_, new_n24038_ );
or   ( new_n24377_, new_n24115_, new_n23834_ );
and  ( new_n24378_, new_n24377_, new_n24376_ );
or   ( new_n24379_, new_n24124_, new_n24020_ );
or   ( new_n24380_, new_n24122_, new_n23800_ );
and  ( new_n24381_, new_n24380_, new_n24379_ );
or   ( new_n24382_, new_n24381_, new_n24378_ );
and  ( new_n24383_, new_n24381_, new_n24378_ );
or   ( new_n24384_, new_n24133_, new_n24005_ );
or   ( new_n24385_, new_n24131_, new_n23775_ );
and  ( new_n24386_, new_n24385_, new_n24384_ );
or   ( new_n24387_, new_n24386_, new_n24383_ );
and  ( new_n24388_, new_n24387_, new_n24382_ );
or   ( new_n24389_, new_n24153_, new_n16085_ );
or   ( new_n24390_, new_n24149_, new_n16048_ );
and  ( new_n24391_, new_n24390_, new_n24389_ );
or   ( new_n24392_, new_n24144_, new_n16505_ );
or   ( new_n24393_, new_n24140_, new_n16438_ );
and  ( new_n24394_, new_n24393_, new_n24392_ );
or   ( new_n24395_, new_n24394_, new_n24391_ );
and  ( new_n24396_, new_n24394_, new_n24391_ );
or   ( new_n24397_, new_n24164_, new_n16052_ );
or   ( new_n24398_, new_n24160_, new_n16071_ );
and  ( new_n24399_, new_n24398_, new_n24397_ );
or   ( new_n24400_, new_n24399_, new_n24396_ );
and  ( new_n24401_, new_n24400_, new_n24395_ );
or   ( new_n24402_, new_n24175_, new_n16009_ );
or   ( new_n24403_, new_n24171_, new_n16029_ );
and  ( new_n24404_, new_n24403_, new_n24402_ );
or   ( new_n24405_, new_n24184_, new_n16186_ );
or   ( new_n24406_, new_n24180_, new_n16204_ );
and  ( new_n24407_, new_n24406_, new_n24405_ );
or   ( new_n24408_, new_n24407_, new_n24404_ );
and  ( new_n24409_, new_n24407_, new_n24404_ );
or   ( new_n24410_, new_n24195_, new_n16217_ );
or   ( new_n24411_, new_n24191_, new_n16234_ );
and  ( new_n24412_, new_n24411_, new_n24410_ );
or   ( new_n24413_, new_n24412_, new_n24409_ );
and  ( new_n24414_, new_n24413_, new_n24408_ );
or   ( new_n24415_, new_n24414_, new_n24401_ );
and  ( new_n24416_, new_n24414_, new_n24401_ );
or   ( new_n24417_, new_n24206_, new_n23998_ );
or   ( new_n24418_, new_n24204_, new_n23762_ );
and  ( new_n24419_, new_n24418_, new_n24417_ );
or   ( new_n24420_, new_n24419_, new_n24416_ );
and  ( new_n24421_, new_n24420_, new_n24415_ );
or   ( new_n24422_, new_n24217_, new_n20156_ );
or   ( new_n24423_, new_n24213_, new_n20443_ );
and  ( new_n24424_, new_n24423_, new_n24422_ );
or   ( new_n24425_, new_n24226_, new_n19394_ );
or   ( new_n24426_, new_n24222_, new_n19659_ );
and  ( new_n24427_, new_n24426_, new_n24425_ );
or   ( new_n24428_, new_n24427_, new_n24424_ );
and  ( new_n24429_, new_n24427_, new_n24424_ );
or   ( new_n24430_, new_n24237_, new_n18742_ );
or   ( new_n24431_, new_n24233_, new_n18977_ );
and  ( new_n24432_, new_n24431_, new_n24430_ );
or   ( new_n24433_, new_n24432_, new_n24429_ );
and  ( new_n24434_, new_n24433_, new_n24428_ );
or   ( new_n24435_, new_n24247_, new_n21261_ );
or   ( new_n24436_, new_n24243_, new_n21009_ );
and  ( new_n24437_, new_n24436_, new_n24435_ );
or   ( new_n24438_, new_n24437_, new_n16151_ );
and  ( new_n24439_, new_n24437_, new_n16151_ );
or   ( new_n24440_, new_n24258_, new_n21013_ );
or   ( new_n24441_, new_n24254_, new_n21265_ );
and  ( new_n24442_, new_n24441_, new_n24440_ );
or   ( new_n24443_, new_n24442_, new_n24439_ );
and  ( new_n24444_, new_n24443_, new_n24438_ );
or   ( new_n24445_, new_n24444_, new_n24434_ );
and  ( new_n24446_, new_n24444_, new_n24434_ );
or   ( new_n24447_, new_n24271_, new_n18066_ );
or   ( new_n24448_, new_n24267_, new_n18309_ );
and  ( new_n24449_, new_n24448_, new_n24447_ );
or   ( new_n24450_, new_n24280_, new_n17238_ );
or   ( new_n24451_, new_n24276_, new_n17650_ );
and  ( new_n24452_, new_n24451_, new_n24450_ );
or   ( new_n24453_, new_n24452_, new_n24449_ );
and  ( new_n24454_, new_n24452_, new_n24449_ );
or   ( new_n24455_, new_n24291_, new_n16814_ );
or   ( new_n24456_, new_n24287_, new_n17142_ );
and  ( new_n24457_, new_n24456_, new_n24455_ );
or   ( new_n24458_, new_n24457_, new_n24454_ );
and  ( new_n24459_, new_n24458_, new_n24453_ );
or   ( new_n24460_, new_n24459_, new_n24446_ );
and  ( new_n24461_, new_n24460_, new_n24445_ );
or   ( new_n24462_, new_n24461_, new_n24421_ );
and  ( new_n24463_, new_n24461_, new_n24421_ );
or   ( new_n24464_, new_n24304_, new_n23985_ );
or   ( new_n24465_, new_n24302_, new_n23731_ );
and  ( new_n24466_, new_n24465_, new_n24464_ );
or   ( new_n24467_, new_n24311_, new_n23970_ );
or   ( new_n24468_, new_n24309_, new_n23698_ );
and  ( new_n24469_, new_n24468_, new_n24467_ );
or   ( new_n24470_, new_n24469_, new_n24466_ );
and  ( new_n24471_, new_n24469_, new_n24466_ );
or   ( new_n24472_, new_n24320_, new_n23955_ );
or   ( new_n24473_, new_n24318_, new_n23665_ );
and  ( new_n24474_, new_n24473_, new_n24472_ );
or   ( new_n24475_, new_n24474_, new_n24471_ );
and  ( new_n24476_, new_n24475_, new_n24470_ );
or   ( new_n24477_, new_n24476_, new_n24463_ );
and  ( new_n24478_, new_n24477_, new_n24462_ );
or   ( new_n24479_, new_n24478_, new_n24388_ );
and  ( new_n24480_, new_n24478_, new_n24388_ );
or   ( new_n24481_, new_n24333_, new_n24060_ );
or   ( new_n24482_, new_n24331_, new_n23872_ );
and  ( new_n24483_, new_n24482_, new_n24481_ );
or   ( new_n24484_, new_n24483_, new_n24480_ );
and  ( new_n24485_, new_n24484_, new_n24479_ );
or   ( new_n24486_, new_n24485_, new_n24375_ );
and  ( new_n24487_, new_n24485_, new_n24375_ );
or   ( new_n24488_, new_n24344_, new_n24074_ );
or   ( new_n24489_, new_n24342_, new_n23895_ );
and  ( new_n24490_, new_n24489_, new_n24488_ );
or   ( new_n24491_, new_n24490_, new_n24487_ );
and  ( new_n24492_, new_n24491_, new_n24486_ );
or   ( new_n24493_, new_n24492_, new_n24097_ );
and  ( new_n24494_, new_n24493_, new_n24368_ );
or   ( new_n24495_, new_n24494_, new_n24364_ );
or   ( new_n24496_, new_n24492_, new_n24367_ );
and  ( new_n24497_, new_n24496_, new_n24350_ );
or   ( new_n24498_, new_n24497_, new_n24357_ );
and  ( new_n24499_, new_n24498_, new_n24495_ );
or   ( new_n24500_, new_n24047_, new_n23804_ );
or   ( new_n24501_, new_n24024_, new_n23847_ );
and  ( new_n24502_, new_n24501_, new_n24500_ );
or   ( new_n24503_, new_n24502_, new_n24062_ );
and  ( new_n24504_, new_n24048_, new_n23848_ );
or   ( new_n24505_, new_n24504_, new_n23874_ );
and  ( new_n24506_, new_n24505_, new_n24503_ );
or   ( new_n24507_, new_n24374_, new_n24104_ );
or   ( new_n24508_, new_n24371_, new_n24111_ );
and  ( new_n24509_, new_n24508_, new_n24507_ );
nor  ( new_n24510_, new_n22333_, new_n755_ );
nor  ( new_n24511_, new_n24510_, new_n9430_ );
or   ( new_n24512_, new_n24511_, new_n21261_ );
and  ( new_n24513_, new_n22337_, RI2b1c4342d738_70 );
and  ( new_n24514_, new_n22330_, RI2b1c4342d6c0_69 );
or   ( new_n24515_, new_n24514_, new_n24513_ );
or   ( new_n24516_, new_n24515_, new_n21009_ );
and  ( new_n24517_, new_n24516_, new_n24512_ );
or   ( new_n24518_, new_n21419_, new_n806_ );
or   ( new_n24519_, new_n21424_, new_n110_ );
and  ( new_n24520_, new_n24519_, new_n24518_ );
or   ( new_n24521_, new_n24520_, new_n21013_ );
and  ( new_n24522_, new_n21428_, RI2b1c4342d828_72 );
and  ( new_n24523_, new_n21415_, RI2b1c4342d7b0_71 );
or   ( new_n24524_, new_n24523_, new_n24522_ );
or   ( new_n24525_, new_n24524_, new_n21265_ );
and  ( new_n24526_, new_n24525_, new_n24521_ );
or   ( new_n24527_, new_n24526_, new_n24517_ );
and  ( new_n24528_, new_n24526_, new_n24517_ );
or   ( new_n24529_, new_n20557_, new_n859_ );
or   ( new_n24530_, new_n20562_, new_n105_ );
and  ( new_n24531_, new_n24530_, new_n24529_ );
or   ( new_n24532_, new_n24531_, new_n20156_ );
and  ( new_n24533_, new_n20566_, RI2b1c4342d918_74 );
and  ( new_n24534_, new_n20553_, RI2b1c4342d8a0_73 );
or   ( new_n24535_, new_n24534_, new_n24533_ );
or   ( new_n24536_, new_n24535_, new_n20443_ );
and  ( new_n24537_, new_n24536_, new_n24532_ );
or   ( new_n24538_, new_n24537_, new_n24528_ );
and  ( new_n24539_, new_n24538_, new_n24527_ );
or   ( new_n24540_, new_n19758_, new_n886_ );
or   ( new_n24541_, new_n19763_, new_n843_ );
and  ( new_n24542_, new_n24541_, new_n24540_ );
or   ( new_n24543_, new_n24542_, new_n19394_ );
and  ( new_n24544_, new_n19767_, RI2b1c4342da08_76 );
and  ( new_n24545_, new_n19754_, RI2b1c4342d990_75 );
or   ( new_n24546_, new_n24545_, new_n24544_ );
or   ( new_n24547_, new_n24546_, new_n19659_ );
and  ( new_n24548_, new_n24547_, new_n24543_ );
or   ( new_n24549_, new_n19048_, new_n1002_ );
or   ( new_n24550_, new_n19055_, new_n1004_ );
and  ( new_n24551_, new_n24550_, new_n24549_ );
or   ( new_n24552_, new_n24551_, new_n18742_ );
and  ( new_n24553_, new_n19057_, RI2b1c4342daf8_78 );
and  ( new_n24554_, new_n19044_, RI2b1c4342da80_77 );
or   ( new_n24555_, new_n24554_, new_n24553_ );
or   ( new_n24556_, new_n24555_, new_n18977_ );
and  ( new_n24557_, new_n24556_, new_n24552_ );
or   ( new_n24558_, new_n24557_, new_n24548_ );
and  ( new_n24559_, new_n24557_, new_n24548_ );
or   ( new_n24560_, new_n18388_, new_n1511_ );
or   ( new_n24561_, new_n18395_, new_n1310_ );
and  ( new_n24562_, new_n24561_, new_n24560_ );
or   ( new_n24563_, new_n24562_, new_n18066_ );
and  ( new_n24564_, new_n18397_, RI2b1c4342dbe8_80 );
and  ( new_n24565_, new_n18384_, RI2b1c4342db70_79 );
or   ( new_n24566_, new_n24565_, new_n24564_ );
or   ( new_n24567_, new_n24566_, new_n18309_ );
and  ( new_n24568_, new_n24567_, new_n24563_ );
or   ( new_n24569_, new_n24568_, new_n24559_ );
and  ( new_n24570_, new_n24569_, new_n24558_ );
or   ( new_n24571_, new_n24570_, new_n24539_ );
and  ( new_n24572_, new_n24570_, new_n24539_ );
or   ( new_n24573_, new_n17727_, new_n2119_ );
or   ( new_n24574_, new_n17734_, new_n126_ );
and  ( new_n24575_, new_n24574_, new_n24573_ );
or   ( new_n24576_, new_n24575_, new_n17238_ );
and  ( new_n24577_, new_n17736_, RI2b1c4342dcd8_82 );
and  ( new_n24578_, new_n17723_, RI2b1c4342dc60_81 );
or   ( new_n24579_, new_n24578_, new_n24577_ );
or   ( new_n24580_, new_n24579_, new_n17650_ );
and  ( new_n24581_, new_n24580_, new_n24576_ );
or   ( new_n24582_, new_n17244_, new_n2541_ );
or   ( new_n24583_, new_n17248_, new_n121_ );
and  ( new_n24584_, new_n24583_, new_n24582_ );
or   ( new_n24585_, new_n24584_, new_n16814_ );
and  ( new_n24586_, new_n17255_, RI2b1c4342ddc8_84 );
and  ( new_n24587_, new_n17240_, RI2b1c4342dd50_83 );
or   ( new_n24588_, new_n24587_, new_n24586_ );
or   ( new_n24589_, new_n24588_, new_n17142_ );
and  ( new_n24590_, new_n24589_, new_n24585_ );
or   ( new_n24591_, new_n24590_, new_n24581_ );
and  ( new_n24592_, new_n24590_, new_n24581_ );
or   ( new_n24593_, new_n16607_, new_n3239_ );
or   ( new_n24594_, new_n16613_, new_n2806_ );
and  ( new_n24595_, new_n24594_, new_n24593_ );
or   ( new_n24596_, new_n24595_, new_n16505_ );
and  ( new_n24597_, new_n16616_, RI2b1c4342deb8_86 );
and  ( new_n24598_, new_n16603_, RI2b1c4342de40_85 );
or   ( new_n24599_, new_n24598_, new_n24597_ );
or   ( new_n24600_, new_n24599_, new_n16438_ );
and  ( new_n24601_, new_n24600_, new_n24596_ );
or   ( new_n24602_, new_n24601_, new_n24592_ );
and  ( new_n24603_, new_n24602_, new_n24591_ );
or   ( new_n24604_, new_n24603_, new_n24572_ );
and  ( new_n24605_, new_n24604_, new_n24571_ );
or   ( new_n24606_, new_n16160_, new_n7274_ );
or   ( new_n24607_, new_n24606_, new_n16151_ );
and  ( new_n24608_, new_n16165_, RI2b1c4342e368_96 );
or   ( new_n24609_, new_n24608_, new_n16170_ );
and  ( new_n24610_, new_n24609_, new_n24607_ );
or   ( new_n24611_, new_n16366_, new_n3902_ );
or   ( new_n24612_, new_n16355_, new_n3924_ );
and  ( new_n24613_, new_n24612_, new_n24611_ );
or   ( new_n24614_, new_n24613_, new_n16085_ );
and  ( new_n24615_, new_n16358_, RI2b1c4342dfa8_88 );
and  ( new_n24616_, new_n16362_, RI2b1c4342df30_87 );
or   ( new_n24617_, new_n24616_, new_n24615_ );
or   ( new_n24618_, new_n24617_, new_n16048_ );
and  ( new_n24619_, new_n24618_, new_n24614_ );
or   ( new_n24620_, new_n16075_, new_n4635_ );
or   ( new_n24621_, new_n16060_, new_n132_ );
and  ( new_n24622_, new_n24621_, new_n24620_ );
or   ( new_n24623_, new_n24622_, new_n16052_ );
and  ( new_n24624_, new_n16063_, RI2b1c4342e098_90 );
and  ( new_n24625_, new_n16066_, RI2b1c4342e020_89 );
or   ( new_n24626_, new_n24625_, new_n24624_ );
or   ( new_n24627_, new_n24626_, new_n16071_ );
and  ( new_n24628_, new_n24627_, new_n24623_ );
or   ( new_n24629_, new_n24628_, new_n24619_ );
and  ( new_n24630_, new_n24628_, new_n24619_ );
or   ( new_n24631_, new_n16033_, new_n5459_ );
or   ( new_n24632_, new_n16017_, new_n117_ );
and  ( new_n24633_, new_n24632_, new_n24631_ );
or   ( new_n24634_, new_n24633_, new_n16009_ );
and  ( new_n24635_, new_n16021_, RI2b1c4342e188_92 );
and  ( new_n24636_, new_n16024_, RI2b1c4342e110_91 );
or   ( new_n24637_, new_n24636_, new_n24635_ );
or   ( new_n24638_, new_n24637_, new_n16029_ );
and  ( new_n24639_, new_n24638_, new_n24634_ );
or   ( new_n24640_, new_n24639_, new_n24630_ );
and  ( new_n24641_, new_n24640_, new_n24629_ );
or   ( new_n24642_, new_n24641_, new_n24610_ );
and  ( new_n24643_, new_n24641_, new_n24610_ );
or   ( new_n24644_, new_n24407_, new_n24177_ );
or   ( new_n24645_, new_n24404_, new_n24186_ );
and  ( new_n24646_, new_n24645_, new_n24644_ );
or   ( new_n24647_, new_n24646_, new_n24412_ );
and  ( new_n24648_, new_n24408_, new_n24187_ );
or   ( new_n24649_, new_n24648_, new_n24197_ );
and  ( new_n24650_, new_n24649_, new_n24647_ );
or   ( new_n24651_, new_n24650_, new_n24643_ );
and  ( new_n24652_, new_n24651_, new_n24642_ );
or   ( new_n24653_, new_n24652_, new_n24605_ );
and  ( new_n24654_, new_n24652_, new_n24605_ );
or   ( new_n24655_, new_n24391_, new_n24146_ );
or   ( new_n24656_, new_n24394_, new_n24155_ );
and  ( new_n24657_, new_n24656_, new_n24655_ );
or   ( new_n24658_, new_n24657_, new_n24399_ );
and  ( new_n24659_, new_n24395_, new_n24156_ );
or   ( new_n24660_, new_n24659_, new_n24166_ );
and  ( new_n24661_, new_n24660_, new_n24658_ );
or   ( new_n24662_, new_n24452_, new_n24273_ );
or   ( new_n24663_, new_n24449_, new_n24282_ );
and  ( new_n24664_, new_n24663_, new_n24662_ );
or   ( new_n24665_, new_n24664_, new_n24457_ );
and  ( new_n24666_, new_n24453_, new_n24283_ );
or   ( new_n24667_, new_n24666_, new_n24293_ );
and  ( new_n24668_, new_n24667_, new_n24665_ );
or   ( new_n24669_, new_n24668_, new_n24661_ );
and  ( new_n24670_, new_n24668_, new_n24661_ );
or   ( new_n24671_, new_n24427_, new_n24219_ );
or   ( new_n24672_, new_n24424_, new_n24228_ );
and  ( new_n24673_, new_n24672_, new_n24671_ );
or   ( new_n24674_, new_n24673_, new_n24432_ );
and  ( new_n24675_, new_n24428_, new_n24229_ );
or   ( new_n24676_, new_n24675_, new_n24239_ );
and  ( new_n24677_, new_n24676_, new_n24674_ );
or   ( new_n24678_, new_n24677_, new_n24670_ );
and  ( new_n24679_, new_n24678_, new_n24669_ );
or   ( new_n24680_, new_n24679_, new_n24654_ );
and  ( new_n24681_, new_n24680_, new_n24653_ );
or   ( new_n24682_, new_n23934_, new_n23614_ );
or   ( new_n24683_, new_n23937_, new_n23623_ );
and  ( new_n24684_, new_n24683_, new_n24682_ );
or   ( new_n24685_, new_n24684_, new_n23942_ );
and  ( new_n24686_, new_n23938_, new_n23624_ );
or   ( new_n24687_, new_n24686_, new_n23634_ );
and  ( new_n24688_, new_n24687_, new_n24685_ );
or   ( new_n24689_, new_n24469_, new_n24306_ );
or   ( new_n24690_, new_n24466_, new_n24313_ );
and  ( new_n24691_, new_n24690_, new_n24689_ );
or   ( new_n24692_, new_n24691_, new_n24474_ );
and  ( new_n24693_, new_n24470_, new_n24314_ );
or   ( new_n24694_, new_n24693_, new_n24322_ );
and  ( new_n24695_, new_n24694_, new_n24692_ );
or   ( new_n24696_, new_n24695_, new_n24688_ );
and  ( new_n24697_, new_n24695_, new_n24688_ );
or   ( new_n24698_, new_n24414_, new_n24168_ );
or   ( new_n24699_, new_n24401_, new_n24199_ );
and  ( new_n24700_, new_n24699_, new_n24698_ );
or   ( new_n24701_, new_n24700_, new_n24419_ );
and  ( new_n24702_, new_n24415_, new_n24200_ );
or   ( new_n24703_, new_n24702_, new_n24208_ );
and  ( new_n24704_, new_n24703_, new_n24701_ );
or   ( new_n24705_, new_n24704_, new_n24697_ );
and  ( new_n24706_, new_n24705_, new_n24696_ );
or   ( new_n24707_, new_n24706_, new_n24681_ );
and  ( new_n24708_, new_n24706_, new_n24681_ );
or   ( new_n24709_, new_n23957_, new_n23636_ );
or   ( new_n24710_, new_n23944_, new_n23667_ );
and  ( new_n24711_, new_n24710_, new_n24709_ );
or   ( new_n24712_, new_n24711_, new_n23972_ );
and  ( new_n24713_, new_n23958_, new_n23668_ );
or   ( new_n24714_, new_n24713_, new_n23700_ );
and  ( new_n24715_, new_n24714_, new_n24712_ );
or   ( new_n24716_, new_n24715_, new_n24708_ );
and  ( new_n24717_, new_n24716_, new_n24707_ );
or   ( new_n24718_, new_n24717_, new_n24509_ );
and  ( new_n24719_, new_n24717_, new_n24509_ );
or   ( new_n24720_, new_n24388_, new_n24326_ );
or   ( new_n24721_, new_n24478_, new_n24137_ );
and  ( new_n24722_, new_n24721_, new_n24720_ );
or   ( new_n24723_, new_n24722_, new_n24483_ );
and  ( new_n24724_, new_n24479_, new_n24328_ );
or   ( new_n24725_, new_n24724_, new_n24335_ );
and  ( new_n24726_, new_n24725_, new_n24723_ );
or   ( new_n24727_, new_n24726_, new_n24719_ );
and  ( new_n24728_, new_n24727_, new_n24718_ );
or   ( new_n24729_, new_n24728_, new_n24506_ );
or   ( new_n24730_, new_n24375_, new_n24337_ );
or   ( new_n24731_, new_n24485_, new_n24112_ );
and  ( new_n24732_, new_n24731_, new_n24730_ );
or   ( new_n24733_, new_n24732_, new_n24490_ );
and  ( new_n24734_, new_n24486_, new_n24339_ );
or   ( new_n24735_, new_n24734_, new_n24346_ );
and  ( new_n24736_, new_n24735_, new_n24733_ );
and  ( new_n24737_, new_n24728_, new_n24506_ );
or   ( new_n24738_, new_n24737_, new_n24736_ );
and  ( new_n24739_, new_n24738_, new_n24729_ );
or   ( new_n24740_, new_n24739_, new_n24499_ );
and  ( new_n24741_, new_n24740_, new_n24361_ );
or   ( new_n24742_, new_n24741_, new_n24360_ );
or   ( new_n24743_, new_n24742_, new_n23924_ );
and  ( new_n24744_, new_n24743_, new_n23922_ );
and  ( new_n24745_, new_n24739_, new_n24499_ );
or   ( new_n24746_, new_n24745_, new_n24360_ );
or   ( new_n24747_, new_n24746_, new_n23924_ );
or   ( new_n24748_, new_n24734_, new_n24490_ );
or   ( new_n24749_, new_n24732_, new_n24346_ );
and  ( new_n24750_, new_n24749_, new_n24748_ );
or   ( new_n24751_, new_n24504_, new_n24062_ );
or   ( new_n24752_, new_n24502_, new_n23874_ );
and  ( new_n24753_, new_n24752_, new_n24751_ );
or   ( new_n24754_, new_n24753_, new_n24728_ );
or   ( new_n24755_, new_n24374_, new_n24371_ );
and  ( new_n24756_, new_n24755_, new_n24112_ );
or   ( new_n24757_, new_n24693_, new_n24474_ );
or   ( new_n24758_, new_n24691_, new_n24322_ );
and  ( new_n24759_, new_n24758_, new_n24757_ );
or   ( new_n24760_, new_n24686_, new_n23942_ );
or   ( new_n24761_, new_n24684_, new_n23634_ );
and  ( new_n24762_, new_n24761_, new_n24760_ );
or   ( new_n24763_, new_n24762_, new_n24759_ );
and  ( new_n24764_, new_n24762_, new_n24759_ );
or   ( new_n24765_, new_n24702_, new_n24419_ );
or   ( new_n24766_, new_n24700_, new_n24208_ );
and  ( new_n24767_, new_n24766_, new_n24765_ );
or   ( new_n24768_, new_n24767_, new_n24764_ );
and  ( new_n24769_, new_n24768_, new_n24763_ );
or   ( new_n24770_, new_n24608_, new_n16151_ );
or   ( new_n24771_, new_n24606_, new_n16170_ );
and  ( new_n24772_, new_n24771_, new_n24770_ );
or   ( new_n24773_, new_n24626_, new_n16052_ );
or   ( new_n24774_, new_n24622_, new_n16071_ );
and  ( new_n24775_, new_n24774_, new_n24773_ );
or   ( new_n24776_, new_n24617_, new_n16085_ );
or   ( new_n24777_, new_n24613_, new_n16048_ );
and  ( new_n24778_, new_n24777_, new_n24776_ );
or   ( new_n24779_, new_n24778_, new_n24775_ );
and  ( new_n24780_, new_n24778_, new_n24775_ );
or   ( new_n24781_, new_n24637_, new_n16009_ );
or   ( new_n24782_, new_n24633_, new_n16029_ );
and  ( new_n24783_, new_n24782_, new_n24781_ );
or   ( new_n24784_, new_n24783_, new_n24780_ );
and  ( new_n24785_, new_n24784_, new_n24779_ );
or   ( new_n24786_, new_n24785_, new_n24772_ );
and  ( new_n24787_, new_n24785_, new_n24772_ );
or   ( new_n24788_, new_n24648_, new_n24412_ );
or   ( new_n24789_, new_n24646_, new_n24197_ );
and  ( new_n24790_, new_n24789_, new_n24788_ );
or   ( new_n24791_, new_n24790_, new_n24787_ );
and  ( new_n24792_, new_n24791_, new_n24786_ );
or   ( new_n24793_, new_n24515_, new_n21261_ );
or   ( new_n24794_, new_n24511_, new_n21009_ );
and  ( new_n24795_, new_n24794_, new_n24793_ );
or   ( new_n24796_, new_n24524_, new_n21013_ );
or   ( new_n24797_, new_n24520_, new_n21265_ );
and  ( new_n24798_, new_n24797_, new_n24796_ );
or   ( new_n24799_, new_n24798_, new_n24795_ );
and  ( new_n24800_, new_n24798_, new_n24795_ );
or   ( new_n24801_, new_n24535_, new_n20156_ );
or   ( new_n24802_, new_n24531_, new_n20443_ );
and  ( new_n24803_, new_n24802_, new_n24801_ );
or   ( new_n24804_, new_n24803_, new_n24800_ );
and  ( new_n24805_, new_n24804_, new_n24799_ );
or   ( new_n24806_, new_n24546_, new_n19394_ );
or   ( new_n24807_, new_n24542_, new_n19659_ );
and  ( new_n24808_, new_n24807_, new_n24806_ );
or   ( new_n24809_, new_n24555_, new_n18742_ );
or   ( new_n24810_, new_n24551_, new_n18977_ );
and  ( new_n24811_, new_n24810_, new_n24809_ );
or   ( new_n24812_, new_n24811_, new_n24808_ );
and  ( new_n24813_, new_n24811_, new_n24808_ );
or   ( new_n24814_, new_n24566_, new_n18066_ );
or   ( new_n24815_, new_n24562_, new_n18309_ );
and  ( new_n24816_, new_n24815_, new_n24814_ );
or   ( new_n24817_, new_n24816_, new_n24813_ );
and  ( new_n24818_, new_n24817_, new_n24812_ );
or   ( new_n24819_, new_n24818_, new_n24805_ );
and  ( new_n24820_, new_n24818_, new_n24805_ );
or   ( new_n24821_, new_n24579_, new_n17238_ );
or   ( new_n24822_, new_n24575_, new_n17650_ );
and  ( new_n24823_, new_n24822_, new_n24821_ );
or   ( new_n24824_, new_n24588_, new_n16814_ );
or   ( new_n24825_, new_n24584_, new_n17142_ );
and  ( new_n24826_, new_n24825_, new_n24824_ );
or   ( new_n24827_, new_n24826_, new_n24823_ );
and  ( new_n24828_, new_n24826_, new_n24823_ );
or   ( new_n24829_, new_n24599_, new_n16505_ );
or   ( new_n24830_, new_n24595_, new_n16438_ );
and  ( new_n24831_, new_n24830_, new_n24829_ );
or   ( new_n24832_, new_n24831_, new_n24828_ );
and  ( new_n24833_, new_n24832_, new_n24827_ );
or   ( new_n24834_, new_n24833_, new_n24820_ );
and  ( new_n24835_, new_n24834_, new_n24819_ );
or   ( new_n24836_, new_n24835_, new_n24792_ );
and  ( new_n24837_, new_n24835_, new_n24792_ );
or   ( new_n24838_, new_n24666_, new_n24457_ );
or   ( new_n24839_, new_n24664_, new_n24293_ );
and  ( new_n24840_, new_n24839_, new_n24838_ );
or   ( new_n24841_, new_n24659_, new_n24399_ );
or   ( new_n24842_, new_n24657_, new_n24166_ );
and  ( new_n24843_, new_n24842_, new_n24841_ );
or   ( new_n24844_, new_n24843_, new_n24840_ );
and  ( new_n24845_, new_n24843_, new_n24840_ );
or   ( new_n24846_, new_n24675_, new_n24432_ );
or   ( new_n24847_, new_n24673_, new_n24239_ );
and  ( new_n24848_, new_n24847_, new_n24846_ );
or   ( new_n24849_, new_n24848_, new_n24845_ );
and  ( new_n24850_, new_n24849_, new_n24844_ );
or   ( new_n24851_, new_n24850_, new_n24837_ );
and  ( new_n24852_, new_n24851_, new_n24836_ );
or   ( new_n24853_, new_n24852_, new_n24769_ );
and  ( new_n24854_, new_n24852_, new_n24769_ );
or   ( new_n24855_, new_n24713_, new_n23972_ );
or   ( new_n24856_, new_n24711_, new_n23700_ );
and  ( new_n24857_, new_n24856_, new_n24855_ );
or   ( new_n24858_, new_n24857_, new_n24854_ );
and  ( new_n24859_, new_n24858_, new_n24853_ );
or   ( new_n24860_, new_n24859_, new_n24756_ );
and  ( new_n24861_, new_n24859_, new_n24756_ );
or   ( new_n24862_, new_n24724_, new_n24483_ );
or   ( new_n24863_, new_n24722_, new_n24335_ );
and  ( new_n24864_, new_n24863_, new_n24862_ );
or   ( new_n24865_, new_n24864_, new_n24861_ );
and  ( new_n24866_, new_n24865_, new_n24860_ );
or   ( new_n24867_, new_n24866_, new_n24506_ );
and  ( new_n24868_, new_n24867_, new_n24754_ );
or   ( new_n24869_, new_n24868_, new_n24750_ );
or   ( new_n24870_, new_n24866_, new_n24753_ );
and  ( new_n24871_, new_n24870_, new_n24729_ );
or   ( new_n24872_, new_n24871_, new_n24736_ );
and  ( new_n24873_, new_n24872_, new_n24869_ );
or   ( new_n24874_, new_n24421_, new_n24297_ );
or   ( new_n24875_, new_n24461_, new_n24210_ );
and  ( new_n24876_, new_n24875_, new_n24874_ );
or   ( new_n24877_, new_n24876_, new_n24476_ );
and  ( new_n24878_, new_n24462_, new_n24299_ );
or   ( new_n24879_, new_n24878_, new_n24324_ );
and  ( new_n24880_, new_n24879_, new_n24877_ );
or   ( new_n24881_, new_n24769_, new_n24681_ );
or   ( new_n24882_, new_n24852_, new_n24706_ );
and  ( new_n24883_, new_n24882_, new_n24881_ );
or   ( new_n24884_, new_n24883_, new_n24857_ );
and  ( new_n24885_, new_n24853_, new_n24707_ );
or   ( new_n24886_, new_n24885_, new_n24715_ );
and  ( new_n24887_, new_n24886_, new_n24884_ );
or   ( new_n24888_, new_n24887_, new_n24880_ );
or   ( new_n24889_, new_n24759_, new_n24688_ );
or   ( new_n24890_, new_n24762_, new_n24695_ );
and  ( new_n24891_, new_n24890_, new_n24889_ );
or   ( new_n24892_, new_n24891_, new_n24767_ );
and  ( new_n24893_, new_n24763_, new_n24696_ );
or   ( new_n24894_, new_n24893_, new_n24704_ );
and  ( new_n24895_, new_n24894_, new_n24892_ );
or   ( new_n24896_, new_n24792_, new_n24605_ );
or   ( new_n24897_, new_n24835_, new_n24652_ );
and  ( new_n24898_, new_n24897_, new_n24896_ );
or   ( new_n24899_, new_n24898_, new_n24850_ );
and  ( new_n24900_, new_n24836_, new_n24653_ );
or   ( new_n24901_, new_n24900_, new_n24679_ );
and  ( new_n24902_, new_n24901_, new_n24899_ );
or   ( new_n24903_, new_n24902_, new_n24895_ );
or   ( new_n24904_, new_n24437_, new_n16170_ );
or   ( new_n24905_, new_n24249_, new_n16151_ );
and  ( new_n24906_, new_n24905_, new_n24904_ );
or   ( new_n24907_, new_n24906_, new_n24442_ );
and  ( new_n24908_, new_n24438_, new_n24251_ );
or   ( new_n24909_, new_n24908_, new_n24260_ );
and  ( new_n24910_, new_n24909_, new_n24907_ );
or   ( new_n24911_, new_n24840_, new_n24661_ );
or   ( new_n24912_, new_n24843_, new_n24668_ );
and  ( new_n24913_, new_n24912_, new_n24911_ );
or   ( new_n24914_, new_n24913_, new_n24848_ );
and  ( new_n24915_, new_n24844_, new_n24669_ );
or   ( new_n24916_, new_n24915_, new_n24677_ );
and  ( new_n24917_, new_n24916_, new_n24914_ );
or   ( new_n24918_, new_n24917_, new_n24910_ );
and  ( new_n24919_, new_n24917_, new_n24910_ );
or   ( new_n24920_, new_n24772_, new_n24641_ );
or   ( new_n24921_, new_n24785_, new_n24610_ );
and  ( new_n24922_, new_n24921_, new_n24920_ );
or   ( new_n24923_, new_n24922_, new_n24790_ );
and  ( new_n24924_, new_n24786_, new_n24642_ );
or   ( new_n24925_, new_n24924_, new_n24650_ );
and  ( new_n24926_, new_n24925_, new_n24923_ );
or   ( new_n24927_, new_n24926_, new_n24919_ );
and  ( new_n24928_, new_n24927_, new_n24918_ );
or   ( new_n24929_, new_n16607_, new_n3924_ );
or   ( new_n24930_, new_n16613_, new_n3239_ );
and  ( new_n24931_, new_n24930_, new_n24929_ );
or   ( new_n24932_, new_n24931_, new_n16505_ );
and  ( new_n24933_, new_n16616_, RI2b1c4342df30_87 );
and  ( new_n24934_, new_n16603_, RI2b1c4342deb8_86 );
or   ( new_n24935_, new_n24934_, new_n24933_ );
or   ( new_n24936_, new_n24935_, new_n16438_ );
and  ( new_n24937_, new_n24936_, new_n24932_ );
or   ( new_n24938_, new_n16366_, new_n132_ );
or   ( new_n24939_, new_n16355_, new_n3902_ );
and  ( new_n24940_, new_n24939_, new_n24938_ );
or   ( new_n24941_, new_n24940_, new_n16085_ );
and  ( new_n24942_, new_n16358_, RI2b1c4342e020_89 );
and  ( new_n24943_, new_n16362_, RI2b1c4342dfa8_88 );
or   ( new_n24944_, new_n24943_, new_n24942_ );
or   ( new_n24945_, new_n24944_, new_n16048_ );
and  ( new_n24946_, new_n24945_, new_n24941_ );
or   ( new_n24947_, new_n24946_, new_n24937_ );
and  ( new_n24948_, new_n24946_, new_n24937_ );
or   ( new_n24949_, new_n16075_, new_n117_ );
or   ( new_n24950_, new_n16060_, new_n4635_ );
and  ( new_n24951_, new_n24950_, new_n24949_ );
or   ( new_n24952_, new_n24951_, new_n16052_ );
and  ( new_n24953_, new_n16063_, RI2b1c4342e110_91 );
and  ( new_n24954_, new_n16066_, RI2b1c4342e098_90 );
or   ( new_n24955_, new_n24954_, new_n24953_ );
or   ( new_n24956_, new_n24955_, new_n16071_ );
and  ( new_n24957_, new_n24956_, new_n24952_ );
or   ( new_n24958_, new_n24957_, new_n24948_ );
and  ( new_n24959_, new_n24958_, new_n24947_ );
or   ( new_n24960_, new_n16033_, new_n6307_ );
or   ( new_n24961_, new_n16017_, new_n5459_ );
and  ( new_n24962_, new_n24961_, new_n24960_ );
or   ( new_n24963_, new_n24962_, new_n16009_ );
and  ( new_n24964_, new_n16021_, RI2b1c4342e200_93 );
and  ( new_n24965_, new_n16024_, RI2b1c4342e188_92 );
or   ( new_n24966_, new_n24965_, new_n24964_ );
or   ( new_n24967_, new_n24966_, new_n16029_ );
and  ( new_n24968_, new_n24967_, new_n24963_ );
or   ( new_n24969_, new_n16208_, new_n124_ );
or   ( new_n24970_, new_n16194_, new_n6321_ );
and  ( new_n24971_, new_n24970_, new_n24969_ );
or   ( new_n24972_, new_n24971_, new_n16186_ );
and  ( new_n24973_, new_n16196_, RI2b1c4342e2f0_95 );
and  ( new_n24974_, new_n16199_, RI2b1c4342e278_94 );
or   ( new_n24975_, new_n24974_, new_n24973_ );
or   ( new_n24976_, new_n24975_, new_n16204_ );
and  ( new_n24977_, new_n24976_, new_n24972_ );
or   ( new_n24978_, new_n24977_, new_n24968_ );
and  ( new_n24979_, new_n24977_, new_n24968_ );
or   ( new_n24980_, new_n16224_, new_n7274_ );
or   ( new_n24981_, new_n24980_, new_n16217_ );
and  ( new_n24982_, new_n16229_, RI2b1c4342e368_96 );
or   ( new_n24983_, new_n24982_, new_n16234_ );
and  ( new_n24984_, new_n24983_, new_n24981_ );
or   ( new_n24985_, new_n24984_, new_n24979_ );
and  ( new_n24986_, new_n24985_, new_n24978_ );
or   ( new_n24987_, new_n24986_, new_n24959_ );
and  ( new_n24988_, new_n24986_, new_n24959_ );
or   ( new_n24989_, new_n16208_, new_n6321_ );
or   ( new_n24990_, new_n16194_, new_n6307_ );
and  ( new_n24991_, new_n24990_, new_n24989_ );
or   ( new_n24992_, new_n24991_, new_n16186_ );
and  ( new_n24993_, new_n16196_, RI2b1c4342e278_94 );
and  ( new_n24994_, new_n16199_, RI2b1c4342e200_93 );
or   ( new_n24995_, new_n24994_, new_n24993_ );
or   ( new_n24996_, new_n24995_, new_n16204_ );
and  ( new_n24997_, new_n24996_, new_n24992_ );
or   ( new_n24998_, new_n24997_, new_n24988_ );
and  ( new_n24999_, new_n24998_, new_n24987_ );
or   ( new_n25000_, new_n20557_, new_n843_ );
or   ( new_n25001_, new_n20562_, new_n859_ );
and  ( new_n25002_, new_n25001_, new_n25000_ );
or   ( new_n25003_, new_n25002_, new_n20156_ );
and  ( new_n25004_, new_n20566_, RI2b1c4342d990_75 );
and  ( new_n25005_, new_n20553_, RI2b1c4342d918_74 );
or   ( new_n25006_, new_n25005_, new_n25004_ );
or   ( new_n25007_, new_n25006_, new_n20443_ );
and  ( new_n25008_, new_n25007_, new_n25003_ );
or   ( new_n25009_, new_n19758_, new_n1004_ );
or   ( new_n25010_, new_n19763_, new_n886_ );
and  ( new_n25011_, new_n25010_, new_n25009_ );
or   ( new_n25012_, new_n25011_, new_n19394_ );
and  ( new_n25013_, new_n19767_, RI2b1c4342da80_77 );
and  ( new_n25014_, new_n19754_, RI2b1c4342da08_76 );
or   ( new_n25015_, new_n25014_, new_n25013_ );
or   ( new_n25016_, new_n25015_, new_n19659_ );
and  ( new_n25017_, new_n25016_, new_n25012_ );
or   ( new_n25018_, new_n25017_, new_n25008_ );
and  ( new_n25019_, new_n25017_, new_n25008_ );
or   ( new_n25020_, new_n19048_, new_n1310_ );
or   ( new_n25021_, new_n19055_, new_n1002_ );
and  ( new_n25022_, new_n25021_, new_n25020_ );
or   ( new_n25023_, new_n25022_, new_n18742_ );
and  ( new_n25024_, new_n19057_, RI2b1c4342db70_79 );
and  ( new_n25025_, new_n19044_, RI2b1c4342daf8_78 );
or   ( new_n25026_, new_n25025_, new_n25024_ );
or   ( new_n25027_, new_n25026_, new_n18977_ );
and  ( new_n25028_, new_n25027_, new_n25023_ );
or   ( new_n25029_, new_n25028_, new_n25019_ );
and  ( new_n25030_, new_n25029_, new_n25018_ );
nor  ( new_n25031_, new_n22333_, new_n110_ );
nor  ( new_n25032_, new_n25031_, new_n9881_ );
or   ( new_n25033_, new_n25032_, new_n21261_ );
and  ( new_n25034_, new_n22337_, RI2b1c4342d7b0_71 );
and  ( new_n25035_, new_n22330_, RI2b1c4342d738_70 );
or   ( new_n25036_, new_n25035_, new_n25034_ );
or   ( new_n25037_, new_n25036_, new_n21009_ );
and  ( new_n25038_, new_n25037_, new_n25033_ );
and  ( new_n25039_, new_n25038_, new_n16234_ );
or   ( new_n25040_, new_n25038_, new_n16234_ );
or   ( new_n25041_, new_n21419_, new_n105_ );
or   ( new_n25042_, new_n21424_, new_n806_ );
and  ( new_n25043_, new_n25042_, new_n25041_ );
or   ( new_n25044_, new_n25043_, new_n21013_ );
and  ( new_n25045_, new_n21428_, RI2b1c4342d8a0_73 );
and  ( new_n25046_, new_n21415_, RI2b1c4342d828_72 );
or   ( new_n25047_, new_n25046_, new_n25045_ );
or   ( new_n25048_, new_n25047_, new_n21265_ );
and  ( new_n25049_, new_n25048_, new_n25044_ );
and  ( new_n25050_, new_n25049_, new_n25040_ );
or   ( new_n25051_, new_n25050_, new_n25039_ );
and  ( new_n25052_, new_n25051_, new_n25030_ );
or   ( new_n25053_, new_n25051_, new_n25030_ );
or   ( new_n25054_, new_n18388_, new_n126_ );
or   ( new_n25055_, new_n18395_, new_n1511_ );
and  ( new_n25056_, new_n25055_, new_n25054_ );
or   ( new_n25057_, new_n25056_, new_n18066_ );
and  ( new_n25058_, new_n18397_, RI2b1c4342dc60_81 );
and  ( new_n25059_, new_n18384_, RI2b1c4342dbe8_80 );
or   ( new_n25060_, new_n25059_, new_n25058_ );
or   ( new_n25061_, new_n25060_, new_n18309_ );
and  ( new_n25062_, new_n25061_, new_n25057_ );
or   ( new_n25063_, new_n17727_, new_n121_ );
or   ( new_n25064_, new_n17734_, new_n2119_ );
and  ( new_n25065_, new_n25064_, new_n25063_ );
or   ( new_n25066_, new_n25065_, new_n17238_ );
and  ( new_n25067_, new_n17736_, RI2b1c4342dd50_83 );
and  ( new_n25068_, new_n17723_, RI2b1c4342dcd8_82 );
or   ( new_n25069_, new_n25068_, new_n25067_ );
or   ( new_n25070_, new_n25069_, new_n17650_ );
and  ( new_n25071_, new_n25070_, new_n25066_ );
or   ( new_n25072_, new_n25071_, new_n25062_ );
and  ( new_n25073_, new_n25071_, new_n25062_ );
or   ( new_n25074_, new_n17244_, new_n2806_ );
or   ( new_n25075_, new_n17248_, new_n2541_ );
and  ( new_n25076_, new_n25075_, new_n25074_ );
or   ( new_n25077_, new_n25076_, new_n16814_ );
and  ( new_n25078_, new_n17255_, RI2b1c4342de40_85 );
and  ( new_n25079_, new_n17240_, RI2b1c4342ddc8_84 );
or   ( new_n25080_, new_n25079_, new_n25078_ );
or   ( new_n25081_, new_n25080_, new_n17142_ );
and  ( new_n25082_, new_n25081_, new_n25077_ );
or   ( new_n25083_, new_n25082_, new_n25073_ );
and  ( new_n25084_, new_n25083_, new_n25072_ );
and  ( new_n25085_, new_n25084_, new_n25053_ );
or   ( new_n25086_, new_n25085_, new_n25052_ );
and  ( new_n25087_, new_n25086_, new_n24999_ );
or   ( new_n25088_, new_n25086_, new_n24999_ );
or   ( new_n25089_, new_n16238_, new_n7274_ );
or   ( new_n25090_, new_n16224_, new_n124_ );
and  ( new_n25091_, new_n25090_, new_n25089_ );
or   ( new_n25092_, new_n25091_, new_n16217_ );
and  ( new_n25093_, new_n16226_, RI2b1c4342e368_96 );
and  ( new_n25094_, new_n16229_, RI2b1c4342e2f0_95 );
or   ( new_n25095_, new_n25094_, new_n25093_ );
or   ( new_n25096_, new_n25095_, new_n16234_ );
and  ( new_n25097_, new_n25096_, new_n25092_ );
or   ( new_n25098_, new_n24775_, new_n24619_ );
or   ( new_n25099_, new_n24778_, new_n24628_ );
and  ( new_n25100_, new_n25099_, new_n25098_ );
or   ( new_n25101_, new_n25100_, new_n24783_ );
and  ( new_n25102_, new_n24779_, new_n24629_ );
or   ( new_n25103_, new_n25102_, new_n24639_ );
and  ( new_n25104_, new_n25103_, new_n25101_ );
or   ( new_n25105_, new_n25104_, new_n25097_ );
and  ( new_n25106_, new_n25104_, new_n25097_ );
or   ( new_n25107_, new_n24826_, new_n24581_ );
or   ( new_n25108_, new_n24823_, new_n24590_ );
and  ( new_n25109_, new_n25108_, new_n25107_ );
or   ( new_n25110_, new_n25109_, new_n24831_ );
and  ( new_n25111_, new_n24827_, new_n24591_ );
or   ( new_n25112_, new_n25111_, new_n24601_ );
and  ( new_n25113_, new_n25112_, new_n25110_ );
or   ( new_n25114_, new_n25113_, new_n25106_ );
and  ( new_n25115_, new_n25114_, new_n25105_ );
and  ( new_n25116_, new_n25115_, new_n25088_ );
or   ( new_n25117_, new_n25116_, new_n25087_ );
and  ( new_n25118_, new_n25117_, new_n24928_ );
or   ( new_n25119_, new_n25117_, new_n24928_ );
or   ( new_n25120_, new_n24434_, new_n24262_ );
or   ( new_n25121_, new_n24444_, new_n24241_ );
and  ( new_n25122_, new_n25121_, new_n25120_ );
or   ( new_n25123_, new_n25122_, new_n24459_ );
and  ( new_n25124_, new_n24445_, new_n24264_ );
or   ( new_n25125_, new_n25124_, new_n24295_ );
and  ( new_n25126_, new_n25125_, new_n25123_ );
and  ( new_n25127_, new_n25126_, new_n25119_ );
or   ( new_n25128_, new_n25127_, new_n25118_ );
and  ( new_n25129_, new_n25128_, new_n24903_ );
or   ( new_n25130_, new_n25128_, new_n24903_ );
or   ( new_n25131_, new_n24381_, new_n24119_ );
or   ( new_n25132_, new_n24378_, new_n24126_ );
and  ( new_n25133_, new_n25132_, new_n25131_ );
or   ( new_n25134_, new_n25133_, new_n24386_ );
and  ( new_n25135_, new_n24382_, new_n24127_ );
or   ( new_n25136_, new_n25135_, new_n24135_ );
and  ( new_n25137_, new_n25136_, new_n25134_ );
and  ( new_n25138_, new_n25137_, new_n25130_ );
or   ( new_n25139_, new_n25138_, new_n25129_ );
and  ( new_n25140_, new_n25139_, new_n24888_ );
or   ( new_n25141_, new_n25139_, new_n24888_ );
or   ( new_n25142_, new_n24756_, new_n24717_ );
or   ( new_n25143_, new_n24859_, new_n24509_ );
and  ( new_n25144_, new_n25143_, new_n25142_ );
or   ( new_n25145_, new_n25144_, new_n24864_ );
and  ( new_n25146_, new_n24860_, new_n24718_ );
or   ( new_n25147_, new_n25146_, new_n24726_ );
and  ( new_n25148_, new_n25147_, new_n25145_ );
and  ( new_n25149_, new_n25148_, new_n25141_ );
or   ( new_n25150_, new_n25149_, new_n25140_ );
and  ( new_n25151_, new_n25150_, new_n24873_ );
or   ( new_n25152_, new_n25150_, new_n24873_ );
or   ( new_n25153_, new_n25146_, new_n24864_ );
or   ( new_n25154_, new_n25144_, new_n24726_ );
and  ( new_n25155_, new_n25154_, new_n25153_ );
or   ( new_n25156_, new_n24878_, new_n24476_ );
or   ( new_n25157_, new_n24876_, new_n24324_ );
and  ( new_n25158_, new_n25157_, new_n25156_ );
or   ( new_n25159_, new_n24885_, new_n24857_ );
or   ( new_n25160_, new_n24883_, new_n24715_ );
and  ( new_n25161_, new_n25160_, new_n25159_ );
and  ( new_n25162_, new_n25161_, new_n25158_ );
or   ( new_n25163_, new_n25162_, new_n25139_ );
or   ( new_n25164_, new_n24893_, new_n24767_ );
or   ( new_n25165_, new_n24891_, new_n24704_ );
and  ( new_n25166_, new_n25165_, new_n25164_ );
or   ( new_n25167_, new_n24900_, new_n24850_ );
or   ( new_n25168_, new_n24898_, new_n24679_ );
and  ( new_n25169_, new_n25168_, new_n25167_ );
and  ( new_n25170_, new_n25169_, new_n25166_ );
or   ( new_n25171_, new_n24908_, new_n24442_ );
or   ( new_n25172_, new_n24906_, new_n24260_ );
and  ( new_n25173_, new_n25172_, new_n25171_ );
or   ( new_n25174_, new_n24915_, new_n24848_ );
or   ( new_n25175_, new_n24913_, new_n24677_ );
and  ( new_n25176_, new_n25175_, new_n25174_ );
or   ( new_n25177_, new_n25176_, new_n25173_ );
and  ( new_n25178_, new_n25176_, new_n25173_ );
or   ( new_n25179_, new_n24924_, new_n24790_ );
or   ( new_n25180_, new_n24922_, new_n24650_ );
and  ( new_n25181_, new_n25180_, new_n25179_ );
or   ( new_n25182_, new_n25181_, new_n25178_ );
and  ( new_n25183_, new_n25182_, new_n25177_ );
or   ( new_n25184_, new_n24935_, new_n16505_ );
or   ( new_n25185_, new_n24931_, new_n16438_ );
and  ( new_n25186_, new_n25185_, new_n25184_ );
or   ( new_n25187_, new_n24944_, new_n16085_ );
or   ( new_n25188_, new_n24940_, new_n16048_ );
and  ( new_n25189_, new_n25188_, new_n25187_ );
or   ( new_n25190_, new_n25189_, new_n25186_ );
and  ( new_n25191_, new_n25189_, new_n25186_ );
or   ( new_n25192_, new_n24955_, new_n16052_ );
or   ( new_n25193_, new_n24951_, new_n16071_ );
and  ( new_n25194_, new_n25193_, new_n25192_ );
or   ( new_n25195_, new_n25194_, new_n25191_ );
and  ( new_n25196_, new_n25195_, new_n25190_ );
or   ( new_n25197_, new_n24966_, new_n16009_ );
or   ( new_n25198_, new_n24962_, new_n16029_ );
and  ( new_n25199_, new_n25198_, new_n25197_ );
or   ( new_n25200_, new_n24975_, new_n16186_ );
or   ( new_n25201_, new_n24971_, new_n16204_ );
and  ( new_n25202_, new_n25201_, new_n25200_ );
or   ( new_n25203_, new_n25202_, new_n25199_ );
and  ( new_n25204_, new_n25202_, new_n25199_ );
or   ( new_n25205_, new_n24982_, new_n16217_ );
or   ( new_n25206_, new_n24980_, new_n16234_ );
and  ( new_n25207_, new_n25206_, new_n25205_ );
or   ( new_n25208_, new_n25207_, new_n25204_ );
and  ( new_n25209_, new_n25208_, new_n25203_ );
or   ( new_n25210_, new_n25209_, new_n25196_ );
and  ( new_n25211_, new_n25209_, new_n25196_ );
or   ( new_n25212_, new_n24995_, new_n16186_ );
or   ( new_n25213_, new_n24991_, new_n16204_ );
and  ( new_n25214_, new_n25213_, new_n25212_ );
or   ( new_n25215_, new_n25214_, new_n25211_ );
and  ( new_n25216_, new_n25215_, new_n25210_ );
or   ( new_n25217_, new_n25006_, new_n20156_ );
or   ( new_n25218_, new_n25002_, new_n20443_ );
and  ( new_n25219_, new_n25218_, new_n25217_ );
or   ( new_n25220_, new_n25015_, new_n19394_ );
or   ( new_n25221_, new_n25011_, new_n19659_ );
and  ( new_n25222_, new_n25221_, new_n25220_ );
or   ( new_n25223_, new_n25222_, new_n25219_ );
and  ( new_n25224_, new_n25222_, new_n25219_ );
or   ( new_n25225_, new_n25026_, new_n18742_ );
or   ( new_n25226_, new_n25022_, new_n18977_ );
and  ( new_n25227_, new_n25226_, new_n25225_ );
or   ( new_n25228_, new_n25227_, new_n25224_ );
and  ( new_n25229_, new_n25228_, new_n25223_ );
or   ( new_n25230_, new_n25036_, new_n21261_ );
or   ( new_n25231_, new_n25032_, new_n21009_ );
and  ( new_n25232_, new_n25231_, new_n25230_ );
or   ( new_n25233_, new_n25232_, new_n16217_ );
and  ( new_n25234_, new_n25232_, new_n16217_ );
or   ( new_n25235_, new_n25047_, new_n21013_ );
or   ( new_n25236_, new_n25043_, new_n21265_ );
and  ( new_n25237_, new_n25236_, new_n25235_ );
or   ( new_n25238_, new_n25237_, new_n25234_ );
and  ( new_n25239_, new_n25238_, new_n25233_ );
or   ( new_n25240_, new_n25239_, new_n25229_ );
and  ( new_n25241_, new_n25239_, new_n25229_ );
or   ( new_n25242_, new_n25060_, new_n18066_ );
or   ( new_n25243_, new_n25056_, new_n18309_ );
and  ( new_n25244_, new_n25243_, new_n25242_ );
or   ( new_n25245_, new_n25069_, new_n17238_ );
or   ( new_n25246_, new_n25065_, new_n17650_ );
and  ( new_n25247_, new_n25246_, new_n25245_ );
or   ( new_n25248_, new_n25247_, new_n25244_ );
and  ( new_n25249_, new_n25247_, new_n25244_ );
or   ( new_n25250_, new_n25080_, new_n16814_ );
or   ( new_n25251_, new_n25076_, new_n17142_ );
and  ( new_n25252_, new_n25251_, new_n25250_ );
or   ( new_n25253_, new_n25252_, new_n25249_ );
and  ( new_n25254_, new_n25253_, new_n25248_ );
or   ( new_n25255_, new_n25254_, new_n25241_ );
and  ( new_n25256_, new_n25255_, new_n25240_ );
or   ( new_n25257_, new_n25256_, new_n25216_ );
and  ( new_n25258_, new_n25256_, new_n25216_ );
or   ( new_n25259_, new_n25095_, new_n16217_ );
or   ( new_n25260_, new_n25091_, new_n16234_ );
and  ( new_n25261_, new_n25260_, new_n25259_ );
or   ( new_n25262_, new_n25102_, new_n24783_ );
or   ( new_n25263_, new_n25100_, new_n24639_ );
and  ( new_n25264_, new_n25263_, new_n25262_ );
or   ( new_n25265_, new_n25264_, new_n25261_ );
and  ( new_n25266_, new_n25264_, new_n25261_ );
or   ( new_n25267_, new_n25111_, new_n24831_ );
or   ( new_n25268_, new_n25109_, new_n24601_ );
and  ( new_n25269_, new_n25268_, new_n25267_ );
or   ( new_n25270_, new_n25269_, new_n25266_ );
and  ( new_n25271_, new_n25270_, new_n25265_ );
or   ( new_n25272_, new_n25271_, new_n25258_ );
and  ( new_n25273_, new_n25272_, new_n25257_ );
or   ( new_n25274_, new_n25273_, new_n25183_ );
and  ( new_n25275_, new_n25273_, new_n25183_ );
or   ( new_n25276_, new_n25124_, new_n24459_ );
or   ( new_n25277_, new_n25122_, new_n24295_ );
and  ( new_n25278_, new_n25277_, new_n25276_ );
or   ( new_n25279_, new_n25278_, new_n25275_ );
and  ( new_n25280_, new_n25279_, new_n25274_ );
or   ( new_n25281_, new_n25280_, new_n25170_ );
and  ( new_n25282_, new_n25280_, new_n25170_ );
or   ( new_n25283_, new_n25135_, new_n24386_ );
or   ( new_n25284_, new_n25133_, new_n24135_ );
and  ( new_n25285_, new_n25284_, new_n25283_ );
or   ( new_n25286_, new_n25285_, new_n25282_ );
and  ( new_n25287_, new_n25286_, new_n25281_ );
or   ( new_n25288_, new_n25287_, new_n24888_ );
and  ( new_n25289_, new_n25288_, new_n25163_ );
or   ( new_n25290_, new_n25289_, new_n25155_ );
or   ( new_n25291_, new_n25287_, new_n25162_ );
and  ( new_n25292_, new_n25291_, new_n25141_ );
or   ( new_n25293_, new_n25292_, new_n25148_ );
and  ( new_n25294_, new_n25293_, new_n25290_ );
or   ( new_n25295_, new_n25161_, new_n24880_ );
or   ( new_n25296_, new_n25158_, new_n24887_ );
and  ( new_n25297_, new_n25296_, new_n25295_ );
or   ( new_n25298_, new_n25169_, new_n24895_ );
or   ( new_n25299_, new_n25166_, new_n24902_ );
and  ( new_n25300_, new_n25299_, new_n25298_ );
nor  ( new_n25301_, new_n22333_, new_n806_ );
nor  ( new_n25302_, new_n25301_, new_n10150_ );
or   ( new_n25303_, new_n25302_, new_n21261_ );
and  ( new_n25304_, new_n22337_, RI2b1c4342d828_72 );
and  ( new_n25305_, new_n22330_, RI2b1c4342d7b0_71 );
or   ( new_n25306_, new_n25305_, new_n25304_ );
or   ( new_n25307_, new_n25306_, new_n21009_ );
and  ( new_n25308_, new_n25307_, new_n25303_ );
or   ( new_n25309_, new_n21419_, new_n859_ );
or   ( new_n25310_, new_n21424_, new_n105_ );
and  ( new_n25311_, new_n25310_, new_n25309_ );
or   ( new_n25312_, new_n25311_, new_n21013_ );
and  ( new_n25313_, new_n21428_, RI2b1c4342d918_74 );
and  ( new_n25314_, new_n21415_, RI2b1c4342d8a0_73 );
or   ( new_n25315_, new_n25314_, new_n25313_ );
or   ( new_n25316_, new_n25315_, new_n21265_ );
and  ( new_n25317_, new_n25316_, new_n25312_ );
or   ( new_n25318_, new_n25317_, new_n25308_ );
and  ( new_n25319_, new_n25317_, new_n25308_ );
or   ( new_n25320_, new_n20557_, new_n886_ );
or   ( new_n25321_, new_n20562_, new_n843_ );
and  ( new_n25322_, new_n25321_, new_n25320_ );
or   ( new_n25323_, new_n25322_, new_n20156_ );
and  ( new_n25324_, new_n20566_, RI2b1c4342da08_76 );
and  ( new_n25325_, new_n20553_, RI2b1c4342d990_75 );
or   ( new_n25326_, new_n25325_, new_n25324_ );
or   ( new_n25327_, new_n25326_, new_n20443_ );
and  ( new_n25328_, new_n25327_, new_n25323_ );
or   ( new_n25329_, new_n25328_, new_n25319_ );
and  ( new_n25330_, new_n25329_, new_n25318_ );
or   ( new_n25331_, new_n19758_, new_n1002_ );
or   ( new_n25332_, new_n19763_, new_n1004_ );
and  ( new_n25333_, new_n25332_, new_n25331_ );
or   ( new_n25334_, new_n25333_, new_n19394_ );
and  ( new_n25335_, new_n19767_, RI2b1c4342daf8_78 );
and  ( new_n25336_, new_n19754_, RI2b1c4342da80_77 );
or   ( new_n25337_, new_n25336_, new_n25335_ );
or   ( new_n25338_, new_n25337_, new_n19659_ );
and  ( new_n25339_, new_n25338_, new_n25334_ );
or   ( new_n25340_, new_n19048_, new_n1511_ );
or   ( new_n25341_, new_n19055_, new_n1310_ );
and  ( new_n25342_, new_n25341_, new_n25340_ );
or   ( new_n25343_, new_n25342_, new_n18742_ );
and  ( new_n25344_, new_n19057_, RI2b1c4342dbe8_80 );
and  ( new_n25345_, new_n19044_, RI2b1c4342db70_79 );
or   ( new_n25346_, new_n25345_, new_n25344_ );
or   ( new_n25347_, new_n25346_, new_n18977_ );
and  ( new_n25348_, new_n25347_, new_n25343_ );
or   ( new_n25349_, new_n25348_, new_n25339_ );
and  ( new_n25350_, new_n25348_, new_n25339_ );
or   ( new_n25351_, new_n18388_, new_n2119_ );
or   ( new_n25352_, new_n18395_, new_n126_ );
and  ( new_n25353_, new_n25352_, new_n25351_ );
or   ( new_n25354_, new_n25353_, new_n18066_ );
and  ( new_n25355_, new_n18397_, RI2b1c4342dcd8_82 );
and  ( new_n25356_, new_n18384_, RI2b1c4342dc60_81 );
or   ( new_n25357_, new_n25356_, new_n25355_ );
or   ( new_n25358_, new_n25357_, new_n18309_ );
and  ( new_n25359_, new_n25358_, new_n25354_ );
or   ( new_n25360_, new_n25359_, new_n25350_ );
and  ( new_n25361_, new_n25360_, new_n25349_ );
or   ( new_n25362_, new_n25361_, new_n25330_ );
and  ( new_n25363_, new_n25361_, new_n25330_ );
or   ( new_n25364_, new_n17727_, new_n2541_ );
or   ( new_n25365_, new_n17734_, new_n121_ );
and  ( new_n25366_, new_n25365_, new_n25364_ );
or   ( new_n25367_, new_n25366_, new_n17238_ );
and  ( new_n25368_, new_n17736_, RI2b1c4342ddc8_84 );
and  ( new_n25369_, new_n17723_, RI2b1c4342dd50_83 );
or   ( new_n25370_, new_n25369_, new_n25368_ );
or   ( new_n25371_, new_n25370_, new_n17650_ );
and  ( new_n25372_, new_n25371_, new_n25367_ );
or   ( new_n25373_, new_n17244_, new_n3239_ );
or   ( new_n25374_, new_n17248_, new_n2806_ );
and  ( new_n25375_, new_n25374_, new_n25373_ );
or   ( new_n25376_, new_n25375_, new_n16814_ );
and  ( new_n25377_, new_n17255_, RI2b1c4342deb8_86 );
and  ( new_n25378_, new_n17240_, RI2b1c4342de40_85 );
or   ( new_n25379_, new_n25378_, new_n25377_ );
or   ( new_n25380_, new_n25379_, new_n17142_ );
and  ( new_n25381_, new_n25380_, new_n25376_ );
or   ( new_n25382_, new_n25381_, new_n25372_ );
and  ( new_n25383_, new_n25381_, new_n25372_ );
or   ( new_n25384_, new_n16607_, new_n3902_ );
or   ( new_n25385_, new_n16613_, new_n3924_ );
and  ( new_n25386_, new_n25385_, new_n25384_ );
or   ( new_n25387_, new_n25386_, new_n16505_ );
and  ( new_n25388_, new_n16616_, RI2b1c4342dfa8_88 );
and  ( new_n25389_, new_n16603_, RI2b1c4342df30_87 );
or   ( new_n25390_, new_n25389_, new_n25388_ );
or   ( new_n25391_, new_n25390_, new_n16438_ );
and  ( new_n25392_, new_n25391_, new_n25387_ );
or   ( new_n25393_, new_n25392_, new_n25383_ );
and  ( new_n25394_, new_n25393_, new_n25382_ );
or   ( new_n25395_, new_n25394_, new_n25363_ );
and  ( new_n25396_, new_n25395_, new_n25362_ );
or   ( new_n25397_, new_n25202_, new_n24968_ );
or   ( new_n25398_, new_n25199_, new_n24977_ );
and  ( new_n25399_, new_n25398_, new_n25397_ );
or   ( new_n25400_, new_n25399_, new_n25207_ );
and  ( new_n25401_, new_n25203_, new_n24978_ );
or   ( new_n25402_, new_n25401_, new_n24984_ );
and  ( new_n25403_, new_n25402_, new_n25400_ );
or   ( new_n25404_, new_n16366_, new_n4635_ );
or   ( new_n25405_, new_n16355_, new_n132_ );
and  ( new_n25406_, new_n25405_, new_n25404_ );
or   ( new_n25407_, new_n25406_, new_n16085_ );
and  ( new_n25408_, new_n16358_, RI2b1c4342e098_90 );
and  ( new_n25409_, new_n16362_, RI2b1c4342e020_89 );
or   ( new_n25410_, new_n25409_, new_n25408_ );
or   ( new_n25411_, new_n25410_, new_n16048_ );
and  ( new_n25412_, new_n25411_, new_n25407_ );
or   ( new_n25413_, new_n16075_, new_n5459_ );
or   ( new_n25414_, new_n16060_, new_n117_ );
and  ( new_n25415_, new_n25414_, new_n25413_ );
or   ( new_n25416_, new_n25415_, new_n16052_ );
and  ( new_n25417_, new_n16063_, RI2b1c4342e188_92 );
and  ( new_n25418_, new_n16066_, RI2b1c4342e110_91 );
or   ( new_n25419_, new_n25418_, new_n25417_ );
or   ( new_n25420_, new_n25419_, new_n16071_ );
and  ( new_n25421_, new_n25420_, new_n25416_ );
or   ( new_n25422_, new_n25421_, new_n25412_ );
and  ( new_n25423_, new_n25421_, new_n25412_ );
or   ( new_n25424_, new_n16033_, new_n6321_ );
or   ( new_n25425_, new_n16017_, new_n6307_ );
and  ( new_n25426_, new_n25425_, new_n25424_ );
or   ( new_n25427_, new_n25426_, new_n16009_ );
and  ( new_n25428_, new_n16021_, RI2b1c4342e278_94 );
and  ( new_n25429_, new_n16024_, RI2b1c4342e200_93 );
or   ( new_n25430_, new_n25429_, new_n25428_ );
or   ( new_n25431_, new_n25430_, new_n16029_ );
and  ( new_n25432_, new_n25431_, new_n25427_ );
or   ( new_n25433_, new_n25432_, new_n25423_ );
and  ( new_n25434_, new_n25433_, new_n25422_ );
or   ( new_n25435_, new_n25434_, new_n25403_ );
and  ( new_n25436_, new_n25434_, new_n25403_ );
or   ( new_n25437_, new_n25189_, new_n24937_ );
or   ( new_n25438_, new_n25186_, new_n24946_ );
and  ( new_n25439_, new_n25438_, new_n25437_ );
or   ( new_n25440_, new_n25439_, new_n25194_ );
and  ( new_n25441_, new_n25190_, new_n24947_ );
or   ( new_n25442_, new_n25441_, new_n24957_ );
and  ( new_n25443_, new_n25442_, new_n25440_ );
or   ( new_n25444_, new_n25443_, new_n25436_ );
and  ( new_n25445_, new_n25444_, new_n25435_ );
or   ( new_n25446_, new_n25445_, new_n25396_ );
and  ( new_n25447_, new_n25445_, new_n25396_ );
or   ( new_n25448_, new_n25247_, new_n25062_ );
or   ( new_n25449_, new_n25244_, new_n25071_ );
and  ( new_n25450_, new_n25449_, new_n25448_ );
or   ( new_n25451_, new_n25450_, new_n25252_ );
and  ( new_n25452_, new_n25248_, new_n25072_ );
or   ( new_n25453_, new_n25452_, new_n25082_ );
and  ( new_n25454_, new_n25453_, new_n25451_ );
or   ( new_n25455_, new_n25222_, new_n25008_ );
or   ( new_n25456_, new_n25219_, new_n25017_ );
and  ( new_n25457_, new_n25456_, new_n25455_ );
or   ( new_n25458_, new_n25457_, new_n25227_ );
and  ( new_n25459_, new_n25223_, new_n25018_ );
or   ( new_n25460_, new_n25459_, new_n25028_ );
and  ( new_n25461_, new_n25460_, new_n25458_ );
or   ( new_n25462_, new_n25461_, new_n25454_ );
and  ( new_n25463_, new_n25461_, new_n25454_ );
or   ( new_n25464_, new_n25232_, new_n16234_ );
or   ( new_n25465_, new_n25038_, new_n16217_ );
and  ( new_n25466_, new_n25465_, new_n25464_ );
or   ( new_n25467_, new_n25466_, new_n25237_ );
and  ( new_n25468_, new_n25233_, new_n25040_ );
or   ( new_n25469_, new_n25468_, new_n25049_ );
and  ( new_n25470_, new_n25469_, new_n25467_ );
or   ( new_n25471_, new_n25470_, new_n25463_ );
and  ( new_n25472_, new_n25471_, new_n25462_ );
or   ( new_n25473_, new_n25472_, new_n25447_ );
and  ( new_n25474_, new_n25473_, new_n25446_ );
or   ( new_n25475_, new_n24811_, new_n24548_ );
or   ( new_n25476_, new_n24808_, new_n24557_ );
and  ( new_n25477_, new_n25476_, new_n25475_ );
or   ( new_n25478_, new_n25477_, new_n24816_ );
and  ( new_n25479_, new_n24812_, new_n24558_ );
or   ( new_n25480_, new_n25479_, new_n24568_ );
and  ( new_n25481_, new_n25480_, new_n25478_ );
or   ( new_n25482_, new_n24798_, new_n24517_ );
or   ( new_n25483_, new_n24795_, new_n24526_ );
and  ( new_n25484_, new_n25483_, new_n25482_ );
or   ( new_n25485_, new_n25484_, new_n24803_ );
and  ( new_n25486_, new_n24799_, new_n24527_ );
or   ( new_n25487_, new_n25486_, new_n24537_ );
and  ( new_n25488_, new_n25487_, new_n25485_ );
or   ( new_n25489_, new_n25488_, new_n25481_ );
and  ( new_n25490_, new_n25488_, new_n25481_ );
or   ( new_n25491_, new_n25264_, new_n25097_ );
or   ( new_n25492_, new_n25261_, new_n25104_ );
and  ( new_n25493_, new_n25492_, new_n25491_ );
or   ( new_n25494_, new_n25493_, new_n25269_ );
and  ( new_n25495_, new_n25265_, new_n25105_ );
or   ( new_n25496_, new_n25495_, new_n25113_ );
and  ( new_n25497_, new_n25496_, new_n25494_ );
or   ( new_n25498_, new_n25497_, new_n25490_ );
and  ( new_n25499_, new_n25498_, new_n25489_ );
or   ( new_n25500_, new_n25499_, new_n25474_ );
and  ( new_n25501_, new_n25499_, new_n25474_ );
or   ( new_n25502_, new_n24818_, new_n24539_ );
or   ( new_n25503_, new_n24805_, new_n24570_ );
and  ( new_n25504_, new_n25503_, new_n25502_ );
or   ( new_n25505_, new_n25504_, new_n24833_ );
and  ( new_n25506_, new_n24819_, new_n24571_ );
or   ( new_n25507_, new_n25506_, new_n24603_ );
and  ( new_n25508_, new_n25507_, new_n25505_ );
or   ( new_n25509_, new_n25508_, new_n25501_ );
and  ( new_n25510_, new_n25509_, new_n25500_ );
or   ( new_n25511_, new_n25510_, new_n25300_ );
and  ( new_n25512_, new_n25510_, new_n25300_ );
or   ( new_n25513_, new_n25183_, new_n25117_ );
or   ( new_n25514_, new_n25273_, new_n24928_ );
and  ( new_n25515_, new_n25514_, new_n25513_ );
or   ( new_n25516_, new_n25515_, new_n25278_ );
and  ( new_n25517_, new_n25274_, new_n25119_ );
or   ( new_n25518_, new_n25517_, new_n25126_ );
and  ( new_n25519_, new_n25518_, new_n25516_ );
or   ( new_n25520_, new_n25519_, new_n25512_ );
and  ( new_n25521_, new_n25520_, new_n25511_ );
or   ( new_n25522_, new_n25521_, new_n25297_ );
or   ( new_n25523_, new_n25170_, new_n25128_ );
or   ( new_n25524_, new_n25280_, new_n24903_ );
and  ( new_n25525_, new_n25524_, new_n25523_ );
or   ( new_n25526_, new_n25525_, new_n25285_ );
and  ( new_n25527_, new_n25281_, new_n25130_ );
or   ( new_n25528_, new_n25527_, new_n25137_ );
and  ( new_n25529_, new_n25528_, new_n25526_ );
and  ( new_n25530_, new_n25521_, new_n25297_ );
or   ( new_n25531_, new_n25530_, new_n25529_ );
and  ( new_n25532_, new_n25531_, new_n25522_ );
or   ( new_n25533_, new_n25532_, new_n25294_ );
and  ( new_n25534_, new_n25533_, new_n25152_ );
or   ( new_n25535_, new_n25534_, new_n25151_ );
and  ( new_n25536_, new_n25532_, new_n25294_ );
or   ( new_n25537_, new_n25536_, new_n25151_ );
or   ( new_n25538_, new_n25527_, new_n25285_ );
or   ( new_n25539_, new_n25525_, new_n25137_ );
and  ( new_n25540_, new_n25539_, new_n25538_ );
or   ( new_n25541_, new_n25161_, new_n25158_ );
and  ( new_n25542_, new_n25541_, new_n24888_ );
or   ( new_n25543_, new_n25542_, new_n25521_ );
or   ( new_n25544_, new_n25169_, new_n25166_ );
and  ( new_n25545_, new_n25544_, new_n24903_ );
or   ( new_n25546_, new_n25306_, new_n21261_ );
or   ( new_n25547_, new_n25302_, new_n21009_ );
and  ( new_n25548_, new_n25547_, new_n25546_ );
or   ( new_n25549_, new_n25315_, new_n21013_ );
or   ( new_n25550_, new_n25311_, new_n21265_ );
and  ( new_n25551_, new_n25550_, new_n25549_ );
or   ( new_n25552_, new_n25551_, new_n25548_ );
and  ( new_n25553_, new_n25551_, new_n25548_ );
or   ( new_n25554_, new_n25326_, new_n20156_ );
or   ( new_n25555_, new_n25322_, new_n20443_ );
and  ( new_n25556_, new_n25555_, new_n25554_ );
or   ( new_n25557_, new_n25556_, new_n25553_ );
and  ( new_n25558_, new_n25557_, new_n25552_ );
or   ( new_n25559_, new_n25337_, new_n19394_ );
or   ( new_n25560_, new_n25333_, new_n19659_ );
and  ( new_n25561_, new_n25560_, new_n25559_ );
or   ( new_n25562_, new_n25346_, new_n18742_ );
or   ( new_n25563_, new_n25342_, new_n18977_ );
and  ( new_n25564_, new_n25563_, new_n25562_ );
or   ( new_n25565_, new_n25564_, new_n25561_ );
and  ( new_n25566_, new_n25564_, new_n25561_ );
or   ( new_n25567_, new_n25357_, new_n18066_ );
or   ( new_n25568_, new_n25353_, new_n18309_ );
and  ( new_n25569_, new_n25568_, new_n25567_ );
or   ( new_n25570_, new_n25569_, new_n25566_ );
and  ( new_n25571_, new_n25570_, new_n25565_ );
or   ( new_n25572_, new_n25571_, new_n25558_ );
and  ( new_n25573_, new_n25571_, new_n25558_ );
or   ( new_n25574_, new_n25370_, new_n17238_ );
or   ( new_n25575_, new_n25366_, new_n17650_ );
and  ( new_n25576_, new_n25575_, new_n25574_ );
or   ( new_n25577_, new_n25379_, new_n16814_ );
or   ( new_n25578_, new_n25375_, new_n17142_ );
and  ( new_n25579_, new_n25578_, new_n25577_ );
or   ( new_n25580_, new_n25579_, new_n25576_ );
and  ( new_n25581_, new_n25579_, new_n25576_ );
or   ( new_n25582_, new_n25390_, new_n16505_ );
or   ( new_n25583_, new_n25386_, new_n16438_ );
and  ( new_n25584_, new_n25583_, new_n25582_ );
or   ( new_n25585_, new_n25584_, new_n25581_ );
and  ( new_n25586_, new_n25585_, new_n25580_ );
or   ( new_n25587_, new_n25586_, new_n25573_ );
and  ( new_n25588_, new_n25587_, new_n25572_ );
or   ( new_n25589_, new_n25401_, new_n25207_ );
or   ( new_n25590_, new_n25399_, new_n24984_ );
and  ( new_n25591_, new_n25590_, new_n25589_ );
or   ( new_n25592_, new_n25410_, new_n16085_ );
or   ( new_n25593_, new_n25406_, new_n16048_ );
and  ( new_n25594_, new_n25593_, new_n25592_ );
or   ( new_n25595_, new_n25419_, new_n16052_ );
or   ( new_n25596_, new_n25415_, new_n16071_ );
and  ( new_n25597_, new_n25596_, new_n25595_ );
or   ( new_n25598_, new_n25597_, new_n25594_ );
and  ( new_n25599_, new_n25597_, new_n25594_ );
or   ( new_n25600_, new_n25430_, new_n16009_ );
or   ( new_n25601_, new_n25426_, new_n16029_ );
and  ( new_n25602_, new_n25601_, new_n25600_ );
or   ( new_n25603_, new_n25602_, new_n25599_ );
and  ( new_n25604_, new_n25603_, new_n25598_ );
or   ( new_n25605_, new_n25604_, new_n25591_ );
and  ( new_n25606_, new_n25604_, new_n25591_ );
or   ( new_n25607_, new_n25441_, new_n25194_ );
or   ( new_n25608_, new_n25439_, new_n24957_ );
and  ( new_n25609_, new_n25608_, new_n25607_ );
or   ( new_n25610_, new_n25609_, new_n25606_ );
and  ( new_n25611_, new_n25610_, new_n25605_ );
or   ( new_n25612_, new_n25611_, new_n25588_ );
and  ( new_n25613_, new_n25611_, new_n25588_ );
or   ( new_n25614_, new_n25452_, new_n25252_ );
or   ( new_n25615_, new_n25450_, new_n25082_ );
and  ( new_n25616_, new_n25615_, new_n25614_ );
or   ( new_n25617_, new_n25459_, new_n25227_ );
or   ( new_n25618_, new_n25457_, new_n25028_ );
and  ( new_n25619_, new_n25618_, new_n25617_ );
or   ( new_n25620_, new_n25619_, new_n25616_ );
and  ( new_n25621_, new_n25619_, new_n25616_ );
or   ( new_n25622_, new_n25468_, new_n25237_ );
or   ( new_n25623_, new_n25466_, new_n25049_ );
and  ( new_n25624_, new_n25623_, new_n25622_ );
or   ( new_n25625_, new_n25624_, new_n25621_ );
and  ( new_n25626_, new_n25625_, new_n25620_ );
or   ( new_n25627_, new_n25626_, new_n25613_ );
and  ( new_n25628_, new_n25627_, new_n25612_ );
or   ( new_n25629_, new_n25479_, new_n24816_ );
or   ( new_n25630_, new_n25477_, new_n24568_ );
and  ( new_n25631_, new_n25630_, new_n25629_ );
or   ( new_n25632_, new_n25486_, new_n24803_ );
or   ( new_n25633_, new_n25484_, new_n24537_ );
and  ( new_n25634_, new_n25633_, new_n25632_ );
or   ( new_n25635_, new_n25634_, new_n25631_ );
and  ( new_n25636_, new_n25634_, new_n25631_ );
or   ( new_n25637_, new_n25495_, new_n25269_ );
or   ( new_n25638_, new_n25493_, new_n25113_ );
and  ( new_n25639_, new_n25638_, new_n25637_ );
or   ( new_n25640_, new_n25639_, new_n25636_ );
and  ( new_n25641_, new_n25640_, new_n25635_ );
or   ( new_n25642_, new_n25641_, new_n25628_ );
and  ( new_n25643_, new_n25641_, new_n25628_ );
or   ( new_n25644_, new_n25506_, new_n24833_ );
or   ( new_n25645_, new_n25504_, new_n24603_ );
and  ( new_n25646_, new_n25645_, new_n25644_ );
or   ( new_n25647_, new_n25646_, new_n25643_ );
and  ( new_n25648_, new_n25647_, new_n25642_ );
or   ( new_n25649_, new_n25648_, new_n25545_ );
and  ( new_n25650_, new_n25648_, new_n25545_ );
or   ( new_n25651_, new_n25517_, new_n25278_ );
or   ( new_n25652_, new_n25515_, new_n25126_ );
and  ( new_n25653_, new_n25652_, new_n25651_ );
or   ( new_n25654_, new_n25653_, new_n25650_ );
and  ( new_n25655_, new_n25654_, new_n25649_ );
or   ( new_n25656_, new_n25655_, new_n25297_ );
and  ( new_n25657_, new_n25656_, new_n25543_ );
or   ( new_n25658_, new_n25657_, new_n25540_ );
or   ( new_n25659_, new_n25655_, new_n25542_ );
and  ( new_n25660_, new_n25659_, new_n25522_ );
or   ( new_n25661_, new_n25660_, new_n25529_ );
and  ( new_n25662_, new_n25661_, new_n25658_ );
or   ( new_n25663_, new_n25216_, new_n25086_ );
or   ( new_n25664_, new_n25256_, new_n24999_ );
and  ( new_n25665_, new_n25664_, new_n25663_ );
or   ( new_n25666_, new_n25665_, new_n25271_ );
and  ( new_n25667_, new_n25257_, new_n25088_ );
or   ( new_n25668_, new_n25667_, new_n25115_ );
and  ( new_n25669_, new_n25668_, new_n25666_ );
or   ( new_n25670_, new_n25641_, new_n25474_ );
or   ( new_n25671_, new_n25628_, new_n25499_ );
and  ( new_n25672_, new_n25671_, new_n25670_ );
or   ( new_n25673_, new_n25672_, new_n25646_ );
and  ( new_n25674_, new_n25642_, new_n25500_ );
or   ( new_n25675_, new_n25674_, new_n25508_ );
and  ( new_n25676_, new_n25675_, new_n25673_ );
or   ( new_n25677_, new_n25676_, new_n25669_ );
or   ( new_n25678_, new_n25229_, new_n25051_ );
or   ( new_n25679_, new_n25239_, new_n25030_ );
and  ( new_n25680_, new_n25679_, new_n25678_ );
or   ( new_n25681_, new_n25680_, new_n25254_ );
and  ( new_n25682_, new_n25240_, new_n25053_ );
or   ( new_n25683_, new_n25682_, new_n25084_ );
and  ( new_n25684_, new_n25683_, new_n25681_ );
or   ( new_n25685_, new_n25634_, new_n25481_ );
or   ( new_n25686_, new_n25631_, new_n25488_ );
and  ( new_n25687_, new_n25686_, new_n25685_ );
or   ( new_n25688_, new_n25687_, new_n25639_ );
and  ( new_n25689_, new_n25635_, new_n25489_ );
or   ( new_n25690_, new_n25689_, new_n25497_ );
and  ( new_n25691_, new_n25690_, new_n25688_ );
or   ( new_n25692_, new_n25691_, new_n25684_ );
and  ( new_n25693_, new_n25691_, new_n25684_ );
or   ( new_n25694_, new_n25611_, new_n25396_ );
or   ( new_n25695_, new_n25588_, new_n25445_ );
and  ( new_n25696_, new_n25695_, new_n25694_ );
or   ( new_n25697_, new_n25696_, new_n25626_ );
and  ( new_n25698_, new_n25612_, new_n25446_ );
or   ( new_n25699_, new_n25698_, new_n25472_ );
and  ( new_n25700_, new_n25699_, new_n25697_ );
or   ( new_n25701_, new_n25700_, new_n25693_ );
and  ( new_n25702_, new_n25701_, new_n25692_ );
or   ( new_n25703_, new_n25619_, new_n25454_ );
or   ( new_n25704_, new_n25616_, new_n25461_ );
and  ( new_n25705_, new_n25704_, new_n25703_ );
or   ( new_n25706_, new_n25705_, new_n25624_ );
and  ( new_n25707_, new_n25620_, new_n25462_ );
or   ( new_n25708_, new_n25707_, new_n25470_ );
and  ( new_n25709_, new_n25708_, new_n25706_ );
or   ( new_n25710_, new_n25591_, new_n25434_ );
or   ( new_n25711_, new_n25604_, new_n25403_ );
and  ( new_n25712_, new_n25711_, new_n25710_ );
or   ( new_n25713_, new_n25712_, new_n25609_ );
and  ( new_n25714_, new_n25605_, new_n25435_ );
or   ( new_n25715_, new_n25714_, new_n25443_ );
and  ( new_n25716_, new_n25715_, new_n25713_ );
or   ( new_n25717_, new_n25716_, new_n25709_ );
and  ( new_n25718_, new_n25716_, new_n25709_ );
or   ( new_n25719_, new_n25571_, new_n25330_ );
or   ( new_n25720_, new_n25558_, new_n25361_ );
and  ( new_n25721_, new_n25720_, new_n25719_ );
or   ( new_n25722_, new_n25721_, new_n25586_ );
and  ( new_n25723_, new_n25572_, new_n25362_ );
or   ( new_n25724_, new_n25723_, new_n25394_ );
and  ( new_n25725_, new_n25724_, new_n25722_ );
or   ( new_n25726_, new_n25725_, new_n25718_ );
and  ( new_n25727_, new_n25726_, new_n25717_ );
or   ( new_n25728_, new_n16033_, new_n124_ );
or   ( new_n25729_, new_n16017_, new_n6321_ );
and  ( new_n25730_, new_n25729_, new_n25728_ );
or   ( new_n25731_, new_n25730_, new_n16009_ );
and  ( new_n25732_, new_n16021_, RI2b1c4342e2f0_95 );
and  ( new_n25733_, new_n16024_, RI2b1c4342e278_94 );
or   ( new_n25734_, new_n25733_, new_n25732_ );
or   ( new_n25735_, new_n25734_, new_n16029_ );
and  ( new_n25736_, new_n25735_, new_n25731_ );
or   ( new_n25737_, new_n16194_, new_n7274_ );
or   ( new_n25738_, new_n25737_, new_n16186_ );
and  ( new_n25739_, new_n16199_, RI2b1c4342e368_96 );
or   ( new_n25740_, new_n25739_, new_n16204_ );
and  ( new_n25741_, new_n25740_, new_n25738_ );
or   ( new_n25742_, new_n25741_, new_n25736_ );
or   ( new_n25743_, new_n16607_, new_n132_ );
or   ( new_n25744_, new_n16613_, new_n3902_ );
and  ( new_n25745_, new_n25744_, new_n25743_ );
or   ( new_n25746_, new_n25745_, new_n16505_ );
and  ( new_n25747_, new_n16616_, RI2b1c4342e020_89 );
and  ( new_n25748_, new_n16603_, RI2b1c4342dfa8_88 );
or   ( new_n25749_, new_n25748_, new_n25747_ );
or   ( new_n25750_, new_n25749_, new_n16438_ );
and  ( new_n25751_, new_n25750_, new_n25746_ );
or   ( new_n25752_, new_n16366_, new_n117_ );
or   ( new_n25753_, new_n16355_, new_n4635_ );
and  ( new_n25754_, new_n25753_, new_n25752_ );
or   ( new_n25755_, new_n25754_, new_n16085_ );
and  ( new_n25756_, new_n16358_, RI2b1c4342e110_91 );
and  ( new_n25757_, new_n16362_, RI2b1c4342e098_90 );
or   ( new_n25758_, new_n25757_, new_n25756_ );
or   ( new_n25759_, new_n25758_, new_n16048_ );
and  ( new_n25760_, new_n25759_, new_n25755_ );
or   ( new_n25761_, new_n25760_, new_n25751_ );
and  ( new_n25762_, new_n25760_, new_n25751_ );
or   ( new_n25763_, new_n16075_, new_n6307_ );
or   ( new_n25764_, new_n16060_, new_n5459_ );
and  ( new_n25765_, new_n25764_, new_n25763_ );
or   ( new_n25766_, new_n25765_, new_n16052_ );
and  ( new_n25767_, new_n16063_, RI2b1c4342e200_93 );
and  ( new_n25768_, new_n16066_, RI2b1c4342e188_92 );
or   ( new_n25769_, new_n25768_, new_n25767_ );
or   ( new_n25770_, new_n25769_, new_n16071_ );
and  ( new_n25771_, new_n25770_, new_n25766_ );
or   ( new_n25772_, new_n25771_, new_n25762_ );
and  ( new_n25773_, new_n25772_, new_n25761_ );
or   ( new_n25774_, new_n25773_, new_n25742_ );
and  ( new_n25775_, new_n25773_, new_n25742_ );
or   ( new_n25776_, new_n16208_, new_n7274_ );
or   ( new_n25777_, new_n16194_, new_n124_ );
and  ( new_n25778_, new_n25777_, new_n25776_ );
or   ( new_n25779_, new_n25778_, new_n16186_ );
and  ( new_n25780_, new_n16196_, RI2b1c4342e368_96 );
and  ( new_n25781_, new_n16199_, RI2b1c4342e2f0_95 );
or   ( new_n25782_, new_n25781_, new_n25780_ );
or   ( new_n25783_, new_n25782_, new_n16204_ );
and  ( new_n25784_, new_n25783_, new_n25779_ );
or   ( new_n25785_, new_n25784_, new_n25775_ );
and  ( new_n25786_, new_n25785_, new_n25774_ );
or   ( new_n25787_, new_n20557_, new_n1004_ );
or   ( new_n25788_, new_n20562_, new_n886_ );
and  ( new_n25789_, new_n25788_, new_n25787_ );
or   ( new_n25790_, new_n25789_, new_n20156_ );
and  ( new_n25791_, new_n20566_, RI2b1c4342da80_77 );
and  ( new_n25792_, new_n20553_, RI2b1c4342da08_76 );
or   ( new_n25793_, new_n25792_, new_n25791_ );
or   ( new_n25794_, new_n25793_, new_n20443_ );
and  ( new_n25795_, new_n25794_, new_n25790_ );
or   ( new_n25796_, new_n19758_, new_n1310_ );
or   ( new_n25797_, new_n19763_, new_n1002_ );
and  ( new_n25798_, new_n25797_, new_n25796_ );
or   ( new_n25799_, new_n25798_, new_n19394_ );
and  ( new_n25800_, new_n19767_, RI2b1c4342db70_79 );
and  ( new_n25801_, new_n19754_, RI2b1c4342daf8_78 );
or   ( new_n25802_, new_n25801_, new_n25800_ );
or   ( new_n25803_, new_n25802_, new_n19659_ );
and  ( new_n25804_, new_n25803_, new_n25799_ );
or   ( new_n25805_, new_n25804_, new_n25795_ );
and  ( new_n25806_, new_n25804_, new_n25795_ );
or   ( new_n25807_, new_n19048_, new_n126_ );
or   ( new_n25808_, new_n19055_, new_n1511_ );
and  ( new_n25809_, new_n25808_, new_n25807_ );
or   ( new_n25810_, new_n25809_, new_n18742_ );
and  ( new_n25811_, new_n19057_, RI2b1c4342dc60_81 );
and  ( new_n25812_, new_n19044_, RI2b1c4342dbe8_80 );
or   ( new_n25813_, new_n25812_, new_n25811_ );
or   ( new_n25814_, new_n25813_, new_n18977_ );
and  ( new_n25815_, new_n25814_, new_n25810_ );
or   ( new_n25816_, new_n25815_, new_n25806_ );
and  ( new_n25817_, new_n25816_, new_n25805_ );
nor  ( new_n25818_, new_n22333_, new_n105_ );
nor  ( new_n25819_, new_n25818_, new_n10670_ );
or   ( new_n25820_, new_n25819_, new_n21261_ );
and  ( new_n25821_, new_n22337_, RI2b1c4342d8a0_73 );
and  ( new_n25822_, new_n22330_, RI2b1c4342d828_72 );
or   ( new_n25823_, new_n25822_, new_n25821_ );
or   ( new_n25824_, new_n25823_, new_n21009_ );
and  ( new_n25825_, new_n25824_, new_n25820_ );
and  ( new_n25826_, new_n25825_, new_n16204_ );
or   ( new_n25827_, new_n25825_, new_n16204_ );
or   ( new_n25828_, new_n21419_, new_n843_ );
or   ( new_n25829_, new_n21424_, new_n859_ );
and  ( new_n25830_, new_n25829_, new_n25828_ );
or   ( new_n25831_, new_n25830_, new_n21013_ );
and  ( new_n25832_, new_n21428_, RI2b1c4342d990_75 );
and  ( new_n25833_, new_n21415_, RI2b1c4342d918_74 );
or   ( new_n25834_, new_n25833_, new_n25832_ );
or   ( new_n25835_, new_n25834_, new_n21265_ );
and  ( new_n25836_, new_n25835_, new_n25831_ );
and  ( new_n25837_, new_n25836_, new_n25827_ );
or   ( new_n25838_, new_n25837_, new_n25826_ );
and  ( new_n25839_, new_n25838_, new_n25817_ );
or   ( new_n25840_, new_n25838_, new_n25817_ );
or   ( new_n25841_, new_n18388_, new_n121_ );
or   ( new_n25842_, new_n18395_, new_n2119_ );
and  ( new_n25843_, new_n25842_, new_n25841_ );
or   ( new_n25844_, new_n25843_, new_n18066_ );
and  ( new_n25845_, new_n18397_, RI2b1c4342dd50_83 );
and  ( new_n25846_, new_n18384_, RI2b1c4342dcd8_82 );
or   ( new_n25847_, new_n25846_, new_n25845_ );
or   ( new_n25848_, new_n25847_, new_n18309_ );
and  ( new_n25849_, new_n25848_, new_n25844_ );
or   ( new_n25850_, new_n17727_, new_n2806_ );
or   ( new_n25851_, new_n17734_, new_n2541_ );
and  ( new_n25852_, new_n25851_, new_n25850_ );
or   ( new_n25853_, new_n25852_, new_n17238_ );
and  ( new_n25854_, new_n17736_, RI2b1c4342de40_85 );
and  ( new_n25855_, new_n17723_, RI2b1c4342ddc8_84 );
or   ( new_n25856_, new_n25855_, new_n25854_ );
or   ( new_n25857_, new_n25856_, new_n17650_ );
and  ( new_n25858_, new_n25857_, new_n25853_ );
or   ( new_n25859_, new_n25858_, new_n25849_ );
and  ( new_n25860_, new_n25858_, new_n25849_ );
or   ( new_n25861_, new_n17244_, new_n3924_ );
or   ( new_n25862_, new_n17248_, new_n3239_ );
and  ( new_n25863_, new_n25862_, new_n25861_ );
or   ( new_n25864_, new_n25863_, new_n16814_ );
and  ( new_n25865_, new_n17255_, RI2b1c4342df30_87 );
and  ( new_n25866_, new_n17240_, RI2b1c4342deb8_86 );
or   ( new_n25867_, new_n25866_, new_n25865_ );
or   ( new_n25868_, new_n25867_, new_n17142_ );
and  ( new_n25869_, new_n25868_, new_n25864_ );
or   ( new_n25870_, new_n25869_, new_n25860_ );
and  ( new_n25871_, new_n25870_, new_n25859_ );
and  ( new_n25872_, new_n25871_, new_n25840_ );
or   ( new_n25873_, new_n25872_, new_n25839_ );
and  ( new_n25874_, new_n25873_, new_n25786_ );
or   ( new_n25875_, new_n25873_, new_n25786_ );
or   ( new_n25876_, new_n25597_, new_n25412_ );
or   ( new_n25877_, new_n25594_, new_n25421_ );
and  ( new_n25878_, new_n25877_, new_n25876_ );
or   ( new_n25879_, new_n25878_, new_n25602_ );
and  ( new_n25880_, new_n25598_, new_n25422_ );
or   ( new_n25881_, new_n25880_, new_n25432_ );
and  ( new_n25882_, new_n25881_, new_n25879_ );
or   ( new_n25883_, new_n25579_, new_n25372_ );
or   ( new_n25884_, new_n25576_, new_n25381_ );
and  ( new_n25885_, new_n25884_, new_n25883_ );
or   ( new_n25886_, new_n25885_, new_n25584_ );
and  ( new_n25887_, new_n25580_, new_n25382_ );
or   ( new_n25888_, new_n25887_, new_n25392_ );
and  ( new_n25889_, new_n25888_, new_n25886_ );
or   ( new_n25890_, new_n25889_, new_n25882_ );
and  ( new_n25891_, new_n25889_, new_n25882_ );
or   ( new_n25892_, new_n25564_, new_n25339_ );
or   ( new_n25893_, new_n25561_, new_n25348_ );
and  ( new_n25894_, new_n25893_, new_n25892_ );
or   ( new_n25895_, new_n25894_, new_n25569_ );
and  ( new_n25896_, new_n25565_, new_n25349_ );
or   ( new_n25897_, new_n25896_, new_n25359_ );
and  ( new_n25898_, new_n25897_, new_n25895_ );
or   ( new_n25899_, new_n25898_, new_n25891_ );
and  ( new_n25900_, new_n25899_, new_n25890_ );
and  ( new_n25901_, new_n25900_, new_n25875_ );
or   ( new_n25902_, new_n25901_, new_n25874_ );
and  ( new_n25903_, new_n25902_, new_n25727_ );
or   ( new_n25904_, new_n25902_, new_n25727_ );
or   ( new_n25905_, new_n25209_, new_n24959_ );
or   ( new_n25906_, new_n25196_, new_n24986_ );
and  ( new_n25907_, new_n25906_, new_n25905_ );
or   ( new_n25908_, new_n25907_, new_n25214_ );
and  ( new_n25909_, new_n25210_, new_n24987_ );
or   ( new_n25910_, new_n25909_, new_n24997_ );
and  ( new_n25911_, new_n25910_, new_n25908_ );
and  ( new_n25912_, new_n25911_, new_n25904_ );
or   ( new_n25913_, new_n25912_, new_n25903_ );
and  ( new_n25914_, new_n25913_, new_n25702_ );
or   ( new_n25915_, new_n25913_, new_n25702_ );
or   ( new_n25916_, new_n25176_, new_n24910_ );
or   ( new_n25917_, new_n25173_, new_n24917_ );
and  ( new_n25918_, new_n25917_, new_n25916_ );
or   ( new_n25919_, new_n25918_, new_n25181_ );
and  ( new_n25920_, new_n25177_, new_n24918_ );
or   ( new_n25921_, new_n25920_, new_n24926_ );
and  ( new_n25922_, new_n25921_, new_n25919_ );
and  ( new_n25923_, new_n25922_, new_n25915_ );
or   ( new_n25924_, new_n25923_, new_n25914_ );
and  ( new_n25925_, new_n25924_, new_n25677_ );
or   ( new_n25926_, new_n25924_, new_n25677_ );
or   ( new_n25927_, new_n25545_, new_n25510_ );
or   ( new_n25928_, new_n25648_, new_n25300_ );
and  ( new_n25929_, new_n25928_, new_n25927_ );
or   ( new_n25930_, new_n25929_, new_n25653_ );
and  ( new_n25931_, new_n25649_, new_n25511_ );
or   ( new_n25932_, new_n25931_, new_n25519_ );
and  ( new_n25933_, new_n25932_, new_n25930_ );
and  ( new_n25934_, new_n25933_, new_n25926_ );
or   ( new_n25935_, new_n25934_, new_n25925_ );
and  ( new_n25936_, new_n25935_, new_n25662_ );
or   ( new_n25937_, new_n25935_, new_n25662_ );
or   ( new_n25938_, new_n25931_, new_n25653_ );
or   ( new_n25939_, new_n25929_, new_n25519_ );
and  ( new_n25940_, new_n25939_, new_n25938_ );
or   ( new_n25941_, new_n25667_, new_n25271_ );
or   ( new_n25942_, new_n25665_, new_n25115_ );
and  ( new_n25943_, new_n25942_, new_n25941_ );
or   ( new_n25944_, new_n25674_, new_n25646_ );
or   ( new_n25945_, new_n25672_, new_n25508_ );
and  ( new_n25946_, new_n25945_, new_n25944_ );
and  ( new_n25947_, new_n25946_, new_n25943_ );
or   ( new_n25948_, new_n25947_, new_n25924_ );
or   ( new_n25949_, new_n25682_, new_n25254_ );
or   ( new_n25950_, new_n25680_, new_n25084_ );
and  ( new_n25951_, new_n25950_, new_n25949_ );
or   ( new_n25952_, new_n25689_, new_n25639_ );
or   ( new_n25953_, new_n25687_, new_n25497_ );
and  ( new_n25954_, new_n25953_, new_n25952_ );
or   ( new_n25955_, new_n25954_, new_n25951_ );
and  ( new_n25956_, new_n25954_, new_n25951_ );
or   ( new_n25957_, new_n25698_, new_n25626_ );
or   ( new_n25958_, new_n25696_, new_n25472_ );
and  ( new_n25959_, new_n25958_, new_n25957_ );
or   ( new_n25960_, new_n25959_, new_n25956_ );
and  ( new_n25961_, new_n25960_, new_n25955_ );
or   ( new_n25962_, new_n25707_, new_n25624_ );
or   ( new_n25963_, new_n25705_, new_n25470_ );
and  ( new_n25964_, new_n25963_, new_n25962_ );
or   ( new_n25965_, new_n25714_, new_n25609_ );
or   ( new_n25966_, new_n25712_, new_n25443_ );
and  ( new_n25967_, new_n25966_, new_n25965_ );
or   ( new_n25968_, new_n25967_, new_n25964_ );
and  ( new_n25969_, new_n25967_, new_n25964_ );
or   ( new_n25970_, new_n25723_, new_n25586_ );
or   ( new_n25971_, new_n25721_, new_n25394_ );
and  ( new_n25972_, new_n25971_, new_n25970_ );
or   ( new_n25973_, new_n25972_, new_n25969_ );
and  ( new_n25974_, new_n25973_, new_n25968_ );
or   ( new_n25975_, new_n25734_, new_n16009_ );
or   ( new_n25976_, new_n25730_, new_n16029_ );
and  ( new_n25977_, new_n25976_, new_n25975_ );
or   ( new_n25978_, new_n25739_, new_n16186_ );
or   ( new_n25979_, new_n25737_, new_n16204_ );
and  ( new_n25980_, new_n25979_, new_n25978_ );
and  ( new_n25981_, new_n25980_, new_n25977_ );
or   ( new_n25982_, new_n25749_, new_n16505_ );
or   ( new_n25983_, new_n25745_, new_n16438_ );
and  ( new_n25984_, new_n25983_, new_n25982_ );
or   ( new_n25985_, new_n25758_, new_n16085_ );
or   ( new_n25986_, new_n25754_, new_n16048_ );
and  ( new_n25987_, new_n25986_, new_n25985_ );
or   ( new_n25988_, new_n25987_, new_n25984_ );
and  ( new_n25989_, new_n25987_, new_n25984_ );
or   ( new_n25990_, new_n25769_, new_n16052_ );
or   ( new_n25991_, new_n25765_, new_n16071_ );
and  ( new_n25992_, new_n25991_, new_n25990_ );
or   ( new_n25993_, new_n25992_, new_n25989_ );
and  ( new_n25994_, new_n25993_, new_n25988_ );
or   ( new_n25995_, new_n25994_, new_n25981_ );
and  ( new_n25996_, new_n25994_, new_n25981_ );
or   ( new_n25997_, new_n25782_, new_n16186_ );
or   ( new_n25998_, new_n25778_, new_n16204_ );
and  ( new_n25999_, new_n25998_, new_n25997_ );
or   ( new_n26000_, new_n25999_, new_n25996_ );
and  ( new_n26001_, new_n26000_, new_n25995_ );
or   ( new_n26002_, new_n25793_, new_n20156_ );
or   ( new_n26003_, new_n25789_, new_n20443_ );
and  ( new_n26004_, new_n26003_, new_n26002_ );
or   ( new_n26005_, new_n25802_, new_n19394_ );
or   ( new_n26006_, new_n25798_, new_n19659_ );
and  ( new_n26007_, new_n26006_, new_n26005_ );
or   ( new_n26008_, new_n26007_, new_n26004_ );
and  ( new_n26009_, new_n26007_, new_n26004_ );
or   ( new_n26010_, new_n25813_, new_n18742_ );
or   ( new_n26011_, new_n25809_, new_n18977_ );
and  ( new_n26012_, new_n26011_, new_n26010_ );
or   ( new_n26013_, new_n26012_, new_n26009_ );
and  ( new_n26014_, new_n26013_, new_n26008_ );
or   ( new_n26015_, new_n25823_, new_n21261_ );
or   ( new_n26016_, new_n25819_, new_n21009_ );
and  ( new_n26017_, new_n26016_, new_n26015_ );
or   ( new_n26018_, new_n26017_, new_n16186_ );
and  ( new_n26019_, new_n26017_, new_n16186_ );
or   ( new_n26020_, new_n25834_, new_n21013_ );
or   ( new_n26021_, new_n25830_, new_n21265_ );
and  ( new_n26022_, new_n26021_, new_n26020_ );
or   ( new_n26023_, new_n26022_, new_n26019_ );
and  ( new_n26024_, new_n26023_, new_n26018_ );
or   ( new_n26025_, new_n26024_, new_n26014_ );
and  ( new_n26026_, new_n26024_, new_n26014_ );
or   ( new_n26027_, new_n25847_, new_n18066_ );
or   ( new_n26028_, new_n25843_, new_n18309_ );
and  ( new_n26029_, new_n26028_, new_n26027_ );
or   ( new_n26030_, new_n25856_, new_n17238_ );
or   ( new_n26031_, new_n25852_, new_n17650_ );
and  ( new_n26032_, new_n26031_, new_n26030_ );
or   ( new_n26033_, new_n26032_, new_n26029_ );
and  ( new_n26034_, new_n26032_, new_n26029_ );
or   ( new_n26035_, new_n25867_, new_n16814_ );
or   ( new_n26036_, new_n25863_, new_n17142_ );
and  ( new_n26037_, new_n26036_, new_n26035_ );
or   ( new_n26038_, new_n26037_, new_n26034_ );
and  ( new_n26039_, new_n26038_, new_n26033_ );
or   ( new_n26040_, new_n26039_, new_n26026_ );
and  ( new_n26041_, new_n26040_, new_n26025_ );
or   ( new_n26042_, new_n26041_, new_n26001_ );
and  ( new_n26043_, new_n26041_, new_n26001_ );
or   ( new_n26044_, new_n25880_, new_n25602_ );
or   ( new_n26045_, new_n25878_, new_n25432_ );
and  ( new_n26046_, new_n26045_, new_n26044_ );
or   ( new_n26047_, new_n25887_, new_n25584_ );
or   ( new_n26048_, new_n25885_, new_n25392_ );
and  ( new_n26049_, new_n26048_, new_n26047_ );
or   ( new_n26050_, new_n26049_, new_n26046_ );
and  ( new_n26051_, new_n26049_, new_n26046_ );
or   ( new_n26052_, new_n25896_, new_n25569_ );
or   ( new_n26053_, new_n25894_, new_n25359_ );
and  ( new_n26054_, new_n26053_, new_n26052_ );
or   ( new_n26055_, new_n26054_, new_n26051_ );
and  ( new_n26056_, new_n26055_, new_n26050_ );
or   ( new_n26057_, new_n26056_, new_n26043_ );
and  ( new_n26058_, new_n26057_, new_n26042_ );
or   ( new_n26059_, new_n26058_, new_n25974_ );
and  ( new_n26060_, new_n26058_, new_n25974_ );
or   ( new_n26061_, new_n25909_, new_n25214_ );
or   ( new_n26062_, new_n25907_, new_n24997_ );
and  ( new_n26063_, new_n26062_, new_n26061_ );
or   ( new_n26064_, new_n26063_, new_n26060_ );
and  ( new_n26065_, new_n26064_, new_n26059_ );
or   ( new_n26066_, new_n26065_, new_n25961_ );
and  ( new_n26067_, new_n26065_, new_n25961_ );
or   ( new_n26068_, new_n25920_, new_n25181_ );
or   ( new_n26069_, new_n25918_, new_n24926_ );
and  ( new_n26070_, new_n26069_, new_n26068_ );
or   ( new_n26071_, new_n26070_, new_n26067_ );
and  ( new_n26072_, new_n26071_, new_n26066_ );
or   ( new_n26073_, new_n26072_, new_n25677_ );
and  ( new_n26074_, new_n26073_, new_n25948_ );
or   ( new_n26075_, new_n26074_, new_n25940_ );
or   ( new_n26076_, new_n26072_, new_n25947_ );
and  ( new_n26077_, new_n26076_, new_n25926_ );
or   ( new_n26078_, new_n26077_, new_n25933_ );
and  ( new_n26079_, new_n26078_, new_n26075_ );
or   ( new_n26080_, new_n25946_, new_n25669_ );
or   ( new_n26081_, new_n25943_, new_n25676_ );
and  ( new_n26082_, new_n26081_, new_n26080_ );
or   ( new_n26083_, new_n25954_, new_n25684_ );
or   ( new_n26084_, new_n25951_, new_n25691_ );
and  ( new_n26085_, new_n26084_, new_n26083_ );
or   ( new_n26086_, new_n26085_, new_n25959_ );
and  ( new_n26087_, new_n25955_, new_n25692_ );
or   ( new_n26088_, new_n26087_, new_n25700_ );
and  ( new_n26089_, new_n26088_, new_n26086_ );
nor  ( new_n26090_, new_n22333_, new_n859_ );
nor  ( new_n26091_, new_n26090_, new_n10942_ );
or   ( new_n26092_, new_n26091_, new_n21261_ );
and  ( new_n26093_, new_n22337_, RI2b1c4342d918_74 );
and  ( new_n26094_, new_n22330_, RI2b1c4342d8a0_73 );
or   ( new_n26095_, new_n26094_, new_n26093_ );
or   ( new_n26096_, new_n26095_, new_n21009_ );
and  ( new_n26097_, new_n26096_, new_n26092_ );
or   ( new_n26098_, new_n21419_, new_n886_ );
or   ( new_n26099_, new_n21424_, new_n843_ );
and  ( new_n26100_, new_n26099_, new_n26098_ );
or   ( new_n26101_, new_n26100_, new_n21013_ );
and  ( new_n26102_, new_n21428_, RI2b1c4342da08_76 );
and  ( new_n26103_, new_n21415_, RI2b1c4342d990_75 );
or   ( new_n26104_, new_n26103_, new_n26102_ );
or   ( new_n26105_, new_n26104_, new_n21265_ );
and  ( new_n26106_, new_n26105_, new_n26101_ );
or   ( new_n26107_, new_n26106_, new_n26097_ );
and  ( new_n26108_, new_n26106_, new_n26097_ );
or   ( new_n26109_, new_n20557_, new_n1002_ );
or   ( new_n26110_, new_n20562_, new_n1004_ );
and  ( new_n26111_, new_n26110_, new_n26109_ );
or   ( new_n26112_, new_n26111_, new_n20156_ );
and  ( new_n26113_, new_n20566_, RI2b1c4342daf8_78 );
and  ( new_n26114_, new_n20553_, RI2b1c4342da80_77 );
or   ( new_n26115_, new_n26114_, new_n26113_ );
or   ( new_n26116_, new_n26115_, new_n20443_ );
and  ( new_n26117_, new_n26116_, new_n26112_ );
or   ( new_n26118_, new_n26117_, new_n26108_ );
and  ( new_n26119_, new_n26118_, new_n26107_ );
or   ( new_n26120_, new_n19758_, new_n1511_ );
or   ( new_n26121_, new_n19763_, new_n1310_ );
and  ( new_n26122_, new_n26121_, new_n26120_ );
or   ( new_n26123_, new_n26122_, new_n19394_ );
and  ( new_n26124_, new_n19767_, RI2b1c4342dbe8_80 );
and  ( new_n26125_, new_n19754_, RI2b1c4342db70_79 );
or   ( new_n26126_, new_n26125_, new_n26124_ );
or   ( new_n26127_, new_n26126_, new_n19659_ );
and  ( new_n26128_, new_n26127_, new_n26123_ );
or   ( new_n26129_, new_n19048_, new_n2119_ );
or   ( new_n26130_, new_n19055_, new_n126_ );
and  ( new_n26131_, new_n26130_, new_n26129_ );
or   ( new_n26132_, new_n26131_, new_n18742_ );
and  ( new_n26133_, new_n19057_, RI2b1c4342dcd8_82 );
and  ( new_n26134_, new_n19044_, RI2b1c4342dc60_81 );
or   ( new_n26135_, new_n26134_, new_n26133_ );
or   ( new_n26136_, new_n26135_, new_n18977_ );
and  ( new_n26137_, new_n26136_, new_n26132_ );
or   ( new_n26138_, new_n26137_, new_n26128_ );
and  ( new_n26139_, new_n26137_, new_n26128_ );
or   ( new_n26140_, new_n18388_, new_n2541_ );
or   ( new_n26141_, new_n18395_, new_n121_ );
and  ( new_n26142_, new_n26141_, new_n26140_ );
or   ( new_n26143_, new_n26142_, new_n18066_ );
and  ( new_n26144_, new_n18397_, RI2b1c4342ddc8_84 );
and  ( new_n26145_, new_n18384_, RI2b1c4342dd50_83 );
or   ( new_n26146_, new_n26145_, new_n26144_ );
or   ( new_n26147_, new_n26146_, new_n18309_ );
and  ( new_n26148_, new_n26147_, new_n26143_ );
or   ( new_n26149_, new_n26148_, new_n26139_ );
and  ( new_n26150_, new_n26149_, new_n26138_ );
or   ( new_n26151_, new_n26150_, new_n26119_ );
and  ( new_n26152_, new_n26150_, new_n26119_ );
or   ( new_n26153_, new_n17727_, new_n3239_ );
or   ( new_n26154_, new_n17734_, new_n2806_ );
and  ( new_n26155_, new_n26154_, new_n26153_ );
or   ( new_n26156_, new_n26155_, new_n17238_ );
and  ( new_n26157_, new_n17736_, RI2b1c4342deb8_86 );
and  ( new_n26158_, new_n17723_, RI2b1c4342de40_85 );
or   ( new_n26159_, new_n26158_, new_n26157_ );
or   ( new_n26160_, new_n26159_, new_n17650_ );
and  ( new_n26161_, new_n26160_, new_n26156_ );
or   ( new_n26162_, new_n17244_, new_n3902_ );
or   ( new_n26163_, new_n17248_, new_n3924_ );
and  ( new_n26164_, new_n26163_, new_n26162_ );
or   ( new_n26165_, new_n26164_, new_n16814_ );
and  ( new_n26166_, new_n17255_, RI2b1c4342dfa8_88 );
and  ( new_n26167_, new_n17240_, RI2b1c4342df30_87 );
or   ( new_n26168_, new_n26167_, new_n26166_ );
or   ( new_n26169_, new_n26168_, new_n17142_ );
and  ( new_n26170_, new_n26169_, new_n26165_ );
or   ( new_n26171_, new_n26170_, new_n26161_ );
and  ( new_n26172_, new_n26170_, new_n26161_ );
or   ( new_n26173_, new_n16607_, new_n4635_ );
or   ( new_n26174_, new_n16613_, new_n132_ );
and  ( new_n26175_, new_n26174_, new_n26173_ );
or   ( new_n26176_, new_n26175_, new_n16505_ );
and  ( new_n26177_, new_n16616_, RI2b1c4342e098_90 );
and  ( new_n26178_, new_n16603_, RI2b1c4342e020_89 );
or   ( new_n26179_, new_n26178_, new_n26177_ );
or   ( new_n26180_, new_n26179_, new_n16438_ );
and  ( new_n26181_, new_n26180_, new_n26176_ );
or   ( new_n26182_, new_n26181_, new_n26172_ );
and  ( new_n26183_, new_n26182_, new_n26171_ );
or   ( new_n26184_, new_n26183_, new_n26152_ );
and  ( new_n26185_, new_n26184_, new_n26151_ );
or   ( new_n26186_, new_n25980_, new_n25736_ );
or   ( new_n26187_, new_n25977_, new_n25741_ );
and  ( new_n26188_, new_n26187_, new_n26186_ );
or   ( new_n26189_, new_n16366_, new_n5459_ );
or   ( new_n26190_, new_n16355_, new_n117_ );
and  ( new_n26191_, new_n26190_, new_n26189_ );
or   ( new_n26192_, new_n26191_, new_n16085_ );
and  ( new_n26193_, new_n16358_, RI2b1c4342e188_92 );
and  ( new_n26194_, new_n16362_, RI2b1c4342e110_91 );
or   ( new_n26195_, new_n26194_, new_n26193_ );
or   ( new_n26196_, new_n26195_, new_n16048_ );
and  ( new_n26197_, new_n26196_, new_n26192_ );
or   ( new_n26198_, new_n16075_, new_n6321_ );
or   ( new_n26199_, new_n16060_, new_n6307_ );
and  ( new_n26200_, new_n26199_, new_n26198_ );
or   ( new_n26201_, new_n26200_, new_n16052_ );
and  ( new_n26202_, new_n16063_, RI2b1c4342e278_94 );
and  ( new_n26203_, new_n16066_, RI2b1c4342e200_93 );
or   ( new_n26204_, new_n26203_, new_n26202_ );
or   ( new_n26205_, new_n26204_, new_n16071_ );
and  ( new_n26206_, new_n26205_, new_n26201_ );
or   ( new_n26207_, new_n26206_, new_n26197_ );
and  ( new_n26208_, new_n26206_, new_n26197_ );
or   ( new_n26209_, new_n16033_, new_n7274_ );
or   ( new_n26210_, new_n16017_, new_n124_ );
and  ( new_n26211_, new_n26210_, new_n26209_ );
or   ( new_n26212_, new_n26211_, new_n16009_ );
and  ( new_n26213_, new_n16021_, RI2b1c4342e368_96 );
and  ( new_n26214_, new_n16024_, RI2b1c4342e2f0_95 );
or   ( new_n26215_, new_n26214_, new_n26213_ );
or   ( new_n26216_, new_n26215_, new_n16029_ );
and  ( new_n26217_, new_n26216_, new_n26212_ );
or   ( new_n26218_, new_n26217_, new_n26208_ );
and  ( new_n26219_, new_n26218_, new_n26207_ );
or   ( new_n26220_, new_n26219_, new_n26188_ );
and  ( new_n26221_, new_n26219_, new_n26188_ );
or   ( new_n26222_, new_n25987_, new_n25751_ );
or   ( new_n26223_, new_n25984_, new_n25760_ );
and  ( new_n26224_, new_n26223_, new_n26222_ );
or   ( new_n26225_, new_n26224_, new_n25992_ );
and  ( new_n26226_, new_n25988_, new_n25761_ );
or   ( new_n26227_, new_n26226_, new_n25771_ );
and  ( new_n26228_, new_n26227_, new_n26225_ );
or   ( new_n26229_, new_n26228_, new_n26221_ );
and  ( new_n26230_, new_n26229_, new_n26220_ );
or   ( new_n26231_, new_n26230_, new_n26185_ );
and  ( new_n26232_, new_n26230_, new_n26185_ );
or   ( new_n26233_, new_n26032_, new_n25849_ );
or   ( new_n26234_, new_n26029_, new_n25858_ );
and  ( new_n26235_, new_n26234_, new_n26233_ );
or   ( new_n26236_, new_n26235_, new_n26037_ );
and  ( new_n26237_, new_n26033_, new_n25859_ );
or   ( new_n26238_, new_n26237_, new_n25869_ );
and  ( new_n26239_, new_n26238_, new_n26236_ );
or   ( new_n26240_, new_n26007_, new_n25795_ );
or   ( new_n26241_, new_n26004_, new_n25804_ );
and  ( new_n26242_, new_n26241_, new_n26240_ );
or   ( new_n26243_, new_n26242_, new_n26012_ );
and  ( new_n26244_, new_n26008_, new_n25805_ );
or   ( new_n26245_, new_n26244_, new_n25815_ );
and  ( new_n26246_, new_n26245_, new_n26243_ );
or   ( new_n26247_, new_n26246_, new_n26239_ );
and  ( new_n26248_, new_n26246_, new_n26239_ );
or   ( new_n26249_, new_n26017_, new_n16204_ );
or   ( new_n26250_, new_n25825_, new_n16186_ );
and  ( new_n26251_, new_n26250_, new_n26249_ );
or   ( new_n26252_, new_n26251_, new_n26022_ );
and  ( new_n26253_, new_n26018_, new_n25827_ );
or   ( new_n26254_, new_n26253_, new_n25836_ );
and  ( new_n26255_, new_n26254_, new_n26252_ );
or   ( new_n26256_, new_n26255_, new_n26248_ );
and  ( new_n26257_, new_n26256_, new_n26247_ );
or   ( new_n26258_, new_n26257_, new_n26232_ );
and  ( new_n26259_, new_n26258_, new_n26231_ );
or   ( new_n26260_, new_n25551_, new_n25308_ );
or   ( new_n26261_, new_n25548_, new_n25317_ );
and  ( new_n26262_, new_n26261_, new_n26260_ );
or   ( new_n26263_, new_n26262_, new_n25556_ );
and  ( new_n26264_, new_n25552_, new_n25318_ );
or   ( new_n26265_, new_n26264_, new_n25328_ );
and  ( new_n26266_, new_n26265_, new_n26263_ );
or   ( new_n26267_, new_n26049_, new_n25882_ );
or   ( new_n26268_, new_n26046_, new_n25889_ );
and  ( new_n26269_, new_n26268_, new_n26267_ );
or   ( new_n26270_, new_n26269_, new_n26054_ );
and  ( new_n26271_, new_n26050_, new_n25890_ );
or   ( new_n26272_, new_n26271_, new_n25898_ );
and  ( new_n26273_, new_n26272_, new_n26270_ );
or   ( new_n26274_, new_n26273_, new_n26266_ );
and  ( new_n26275_, new_n26273_, new_n26266_ );
or   ( new_n26276_, new_n25981_, new_n25773_ );
or   ( new_n26277_, new_n25994_, new_n25742_ );
and  ( new_n26278_, new_n26277_, new_n26276_ );
or   ( new_n26279_, new_n26278_, new_n25999_ );
and  ( new_n26280_, new_n25995_, new_n25774_ );
or   ( new_n26281_, new_n26280_, new_n25784_ );
and  ( new_n26282_, new_n26281_, new_n26279_ );
or   ( new_n26283_, new_n26282_, new_n26275_ );
and  ( new_n26284_, new_n26283_, new_n26274_ );
or   ( new_n26285_, new_n26284_, new_n26259_ );
and  ( new_n26286_, new_n26284_, new_n26259_ );
or   ( new_n26287_, new_n25967_, new_n25709_ );
or   ( new_n26288_, new_n25964_, new_n25716_ );
and  ( new_n26289_, new_n26288_, new_n26287_ );
or   ( new_n26290_, new_n26289_, new_n25972_ );
and  ( new_n26291_, new_n25968_, new_n25717_ );
or   ( new_n26292_, new_n26291_, new_n25725_ );
and  ( new_n26293_, new_n26292_, new_n26290_ );
or   ( new_n26294_, new_n26293_, new_n26286_ );
and  ( new_n26295_, new_n26294_, new_n26285_ );
or   ( new_n26296_, new_n26295_, new_n26089_ );
and  ( new_n26297_, new_n26295_, new_n26089_ );
or   ( new_n26298_, new_n25974_, new_n25902_ );
or   ( new_n26299_, new_n26058_, new_n25727_ );
and  ( new_n26300_, new_n26299_, new_n26298_ );
or   ( new_n26301_, new_n26300_, new_n26063_ );
and  ( new_n26302_, new_n26059_, new_n25904_ );
or   ( new_n26303_, new_n26302_, new_n25911_ );
and  ( new_n26304_, new_n26303_, new_n26301_ );
or   ( new_n26305_, new_n26304_, new_n26297_ );
and  ( new_n26306_, new_n26305_, new_n26296_ );
or   ( new_n26307_, new_n26306_, new_n26082_ );
or   ( new_n26308_, new_n25961_, new_n25913_ );
or   ( new_n26309_, new_n26065_, new_n25702_ );
and  ( new_n26310_, new_n26309_, new_n26308_ );
or   ( new_n26311_, new_n26310_, new_n26070_ );
and  ( new_n26312_, new_n26066_, new_n25915_ );
or   ( new_n26313_, new_n26312_, new_n25922_ );
and  ( new_n26314_, new_n26313_, new_n26311_ );
and  ( new_n26315_, new_n26306_, new_n26082_ );
or   ( new_n26316_, new_n26315_, new_n26314_ );
and  ( new_n26317_, new_n26316_, new_n26307_ );
or   ( new_n26318_, new_n26317_, new_n26079_ );
and  ( new_n26319_, new_n26318_, new_n25937_ );
or   ( new_n26320_, new_n26319_, new_n25936_ );
or   ( new_n26321_, new_n26320_, new_n25537_ );
and  ( new_n26322_, new_n26321_, new_n25535_ );
or   ( new_n26323_, new_n26322_, new_n24747_ );
and  ( new_n26324_, new_n26317_, new_n26079_ );
or   ( new_n26325_, new_n26324_, new_n25936_ );
or   ( new_n26326_, new_n26325_, new_n25537_ );
or   ( new_n26327_, new_n26302_, new_n26063_ );
or   ( new_n26328_, new_n26300_, new_n25911_ );
and  ( new_n26329_, new_n26328_, new_n26327_ );
or   ( new_n26330_, new_n26087_, new_n25959_ );
or   ( new_n26331_, new_n26085_, new_n25700_ );
and  ( new_n26332_, new_n26331_, new_n26330_ );
or   ( new_n26333_, new_n26332_, new_n26295_ );
or   ( new_n26334_, new_n26095_, new_n21261_ );
or   ( new_n26335_, new_n26091_, new_n21009_ );
and  ( new_n26336_, new_n26335_, new_n26334_ );
or   ( new_n26337_, new_n26104_, new_n21013_ );
or   ( new_n26338_, new_n26100_, new_n21265_ );
and  ( new_n26339_, new_n26338_, new_n26337_ );
or   ( new_n26340_, new_n26339_, new_n26336_ );
and  ( new_n26341_, new_n26339_, new_n26336_ );
or   ( new_n26342_, new_n26115_, new_n20156_ );
or   ( new_n26343_, new_n26111_, new_n20443_ );
and  ( new_n26344_, new_n26343_, new_n26342_ );
or   ( new_n26345_, new_n26344_, new_n26341_ );
and  ( new_n26346_, new_n26345_, new_n26340_ );
or   ( new_n26347_, new_n26126_, new_n19394_ );
or   ( new_n26348_, new_n26122_, new_n19659_ );
and  ( new_n26349_, new_n26348_, new_n26347_ );
or   ( new_n26350_, new_n26135_, new_n18742_ );
or   ( new_n26351_, new_n26131_, new_n18977_ );
and  ( new_n26352_, new_n26351_, new_n26350_ );
or   ( new_n26353_, new_n26352_, new_n26349_ );
and  ( new_n26354_, new_n26352_, new_n26349_ );
or   ( new_n26355_, new_n26146_, new_n18066_ );
or   ( new_n26356_, new_n26142_, new_n18309_ );
and  ( new_n26357_, new_n26356_, new_n26355_ );
or   ( new_n26358_, new_n26357_, new_n26354_ );
and  ( new_n26359_, new_n26358_, new_n26353_ );
or   ( new_n26360_, new_n26359_, new_n26346_ );
and  ( new_n26361_, new_n26359_, new_n26346_ );
or   ( new_n26362_, new_n26159_, new_n17238_ );
or   ( new_n26363_, new_n26155_, new_n17650_ );
and  ( new_n26364_, new_n26363_, new_n26362_ );
or   ( new_n26365_, new_n26168_, new_n16814_ );
or   ( new_n26366_, new_n26164_, new_n17142_ );
and  ( new_n26367_, new_n26366_, new_n26365_ );
or   ( new_n26368_, new_n26367_, new_n26364_ );
and  ( new_n26369_, new_n26367_, new_n26364_ );
or   ( new_n26370_, new_n26179_, new_n16505_ );
or   ( new_n26371_, new_n26175_, new_n16438_ );
and  ( new_n26372_, new_n26371_, new_n26370_ );
or   ( new_n26373_, new_n26372_, new_n26369_ );
and  ( new_n26374_, new_n26373_, new_n26368_ );
or   ( new_n26375_, new_n26374_, new_n26361_ );
and  ( new_n26376_, new_n26375_, new_n26360_ );
or   ( new_n26377_, new_n25980_, new_n25977_ );
and  ( new_n26378_, new_n26377_, new_n25742_ );
or   ( new_n26379_, new_n26195_, new_n16085_ );
or   ( new_n26380_, new_n26191_, new_n16048_ );
and  ( new_n26381_, new_n26380_, new_n26379_ );
or   ( new_n26382_, new_n26204_, new_n16052_ );
or   ( new_n26383_, new_n26200_, new_n16071_ );
and  ( new_n26384_, new_n26383_, new_n26382_ );
or   ( new_n26385_, new_n26384_, new_n26381_ );
and  ( new_n26386_, new_n26384_, new_n26381_ );
or   ( new_n26387_, new_n26215_, new_n16009_ );
or   ( new_n26388_, new_n26211_, new_n16029_ );
and  ( new_n26389_, new_n26388_, new_n26387_ );
or   ( new_n26390_, new_n26389_, new_n26386_ );
and  ( new_n26391_, new_n26390_, new_n26385_ );
or   ( new_n26392_, new_n26391_, new_n26378_ );
and  ( new_n26393_, new_n26391_, new_n26378_ );
or   ( new_n26394_, new_n26226_, new_n25992_ );
or   ( new_n26395_, new_n26224_, new_n25771_ );
and  ( new_n26396_, new_n26395_, new_n26394_ );
or   ( new_n26397_, new_n26396_, new_n26393_ );
and  ( new_n26398_, new_n26397_, new_n26392_ );
or   ( new_n26399_, new_n26398_, new_n26376_ );
and  ( new_n26400_, new_n26398_, new_n26376_ );
or   ( new_n26401_, new_n26237_, new_n26037_ );
or   ( new_n26402_, new_n26235_, new_n25869_ );
and  ( new_n26403_, new_n26402_, new_n26401_ );
or   ( new_n26404_, new_n26244_, new_n26012_ );
or   ( new_n26405_, new_n26242_, new_n25815_ );
and  ( new_n26406_, new_n26405_, new_n26404_ );
or   ( new_n26407_, new_n26406_, new_n26403_ );
and  ( new_n26408_, new_n26406_, new_n26403_ );
or   ( new_n26409_, new_n26253_, new_n26022_ );
or   ( new_n26410_, new_n26251_, new_n25836_ );
and  ( new_n26411_, new_n26410_, new_n26409_ );
or   ( new_n26412_, new_n26411_, new_n26408_ );
and  ( new_n26413_, new_n26412_, new_n26407_ );
or   ( new_n26414_, new_n26413_, new_n26400_ );
and  ( new_n26415_, new_n26414_, new_n26399_ );
or   ( new_n26416_, new_n26264_, new_n25556_ );
or   ( new_n26417_, new_n26262_, new_n25328_ );
and  ( new_n26418_, new_n26417_, new_n26416_ );
or   ( new_n26419_, new_n26271_, new_n26054_ );
or   ( new_n26420_, new_n26269_, new_n25898_ );
and  ( new_n26421_, new_n26420_, new_n26419_ );
or   ( new_n26422_, new_n26421_, new_n26418_ );
and  ( new_n26423_, new_n26421_, new_n26418_ );
or   ( new_n26424_, new_n26280_, new_n25999_ );
or   ( new_n26425_, new_n26278_, new_n25784_ );
and  ( new_n26426_, new_n26425_, new_n26424_ );
or   ( new_n26427_, new_n26426_, new_n26423_ );
and  ( new_n26428_, new_n26427_, new_n26422_ );
or   ( new_n26429_, new_n26428_, new_n26415_ );
and  ( new_n26430_, new_n26428_, new_n26415_ );
or   ( new_n26431_, new_n26291_, new_n25972_ );
or   ( new_n26432_, new_n26289_, new_n25725_ );
and  ( new_n26433_, new_n26432_, new_n26431_ );
or   ( new_n26434_, new_n26433_, new_n26430_ );
and  ( new_n26435_, new_n26434_, new_n26429_ );
or   ( new_n26436_, new_n26435_, new_n26089_ );
and  ( new_n26437_, new_n26436_, new_n26333_ );
or   ( new_n26438_, new_n26437_, new_n26329_ );
or   ( new_n26439_, new_n26435_, new_n26332_ );
and  ( new_n26440_, new_n26439_, new_n26296_ );
or   ( new_n26441_, new_n26440_, new_n26304_ );
and  ( new_n26442_, new_n26441_, new_n26438_ );
or   ( new_n26443_, new_n26421_, new_n26266_ );
or   ( new_n26444_, new_n26418_, new_n26273_ );
and  ( new_n26445_, new_n26444_, new_n26443_ );
or   ( new_n26446_, new_n26445_, new_n26426_ );
and  ( new_n26447_, new_n26422_, new_n26274_ );
or   ( new_n26448_, new_n26447_, new_n26282_ );
and  ( new_n26449_, new_n26448_, new_n26446_ );
or   ( new_n26450_, new_n26398_, new_n26185_ );
or   ( new_n26451_, new_n26376_, new_n26230_ );
and  ( new_n26452_, new_n26451_, new_n26450_ );
or   ( new_n26453_, new_n26452_, new_n26413_ );
and  ( new_n26454_, new_n26399_, new_n26231_ );
or   ( new_n26455_, new_n26454_, new_n26257_ );
and  ( new_n26456_, new_n26455_, new_n26453_ );
or   ( new_n26457_, new_n26456_, new_n26449_ );
or   ( new_n26458_, new_n26406_, new_n26239_ );
or   ( new_n26459_, new_n26403_, new_n26246_ );
and  ( new_n26460_, new_n26459_, new_n26458_ );
or   ( new_n26461_, new_n26460_, new_n26411_ );
and  ( new_n26462_, new_n26407_, new_n26247_ );
or   ( new_n26463_, new_n26462_, new_n26255_ );
and  ( new_n26464_, new_n26463_, new_n26461_ );
or   ( new_n26465_, new_n26378_, new_n26219_ );
or   ( new_n26466_, new_n26391_, new_n26188_ );
and  ( new_n26467_, new_n26466_, new_n26465_ );
or   ( new_n26468_, new_n26467_, new_n26396_ );
and  ( new_n26469_, new_n26392_, new_n26220_ );
or   ( new_n26470_, new_n26469_, new_n26228_ );
and  ( new_n26471_, new_n26470_, new_n26468_ );
or   ( new_n26472_, new_n26471_, new_n26464_ );
and  ( new_n26473_, new_n26471_, new_n26464_ );
or   ( new_n26474_, new_n26359_, new_n26119_ );
or   ( new_n26475_, new_n26346_, new_n26150_ );
and  ( new_n26476_, new_n26475_, new_n26474_ );
or   ( new_n26477_, new_n26476_, new_n26374_ );
and  ( new_n26478_, new_n26360_, new_n26151_ );
or   ( new_n26479_, new_n26478_, new_n26183_ );
and  ( new_n26480_, new_n26479_, new_n26477_ );
or   ( new_n26481_, new_n26480_, new_n26473_ );
and  ( new_n26482_, new_n26481_, new_n26472_ );
or   ( new_n26483_, new_n26384_, new_n26197_ );
or   ( new_n26484_, new_n26381_, new_n26206_ );
and  ( new_n26485_, new_n26484_, new_n26483_ );
or   ( new_n26486_, new_n26485_, new_n26389_ );
and  ( new_n26487_, new_n26385_, new_n26207_ );
or   ( new_n26488_, new_n26487_, new_n26217_ );
and  ( new_n26489_, new_n26488_, new_n26486_ );
or   ( new_n26490_, new_n16607_, new_n117_ );
or   ( new_n26491_, new_n16613_, new_n4635_ );
and  ( new_n26492_, new_n26491_, new_n26490_ );
or   ( new_n26493_, new_n26492_, new_n16505_ );
and  ( new_n26494_, new_n16616_, RI2b1c4342e110_91 );
and  ( new_n26495_, new_n16603_, RI2b1c4342e098_90 );
or   ( new_n26496_, new_n26495_, new_n26494_ );
or   ( new_n26497_, new_n26496_, new_n16438_ );
and  ( new_n26498_, new_n26497_, new_n26493_ );
or   ( new_n26499_, new_n16366_, new_n6307_ );
or   ( new_n26500_, new_n16355_, new_n5459_ );
and  ( new_n26501_, new_n26500_, new_n26499_ );
or   ( new_n26502_, new_n26501_, new_n16085_ );
and  ( new_n26503_, new_n16358_, RI2b1c4342e200_93 );
and  ( new_n26504_, new_n16362_, RI2b1c4342e188_92 );
or   ( new_n26505_, new_n26504_, new_n26503_ );
or   ( new_n26506_, new_n26505_, new_n16048_ );
and  ( new_n26507_, new_n26506_, new_n26502_ );
or   ( new_n26508_, new_n26507_, new_n26498_ );
and  ( new_n26509_, new_n26507_, new_n26498_ );
or   ( new_n26510_, new_n16075_, new_n124_ );
or   ( new_n26511_, new_n16060_, new_n6321_ );
and  ( new_n26512_, new_n26511_, new_n26510_ );
or   ( new_n26513_, new_n26512_, new_n16052_ );
and  ( new_n26514_, new_n16063_, RI2b1c4342e2f0_95 );
and  ( new_n26515_, new_n16066_, RI2b1c4342e278_94 );
or   ( new_n26516_, new_n26515_, new_n26514_ );
or   ( new_n26517_, new_n26516_, new_n16071_ );
and  ( new_n26518_, new_n26517_, new_n26513_ );
or   ( new_n26519_, new_n26518_, new_n26509_ );
and  ( new_n26520_, new_n26519_, new_n26508_ );
or   ( new_n26521_, new_n26520_, new_n26489_ );
and  ( new_n26522_, new_n26520_, new_n26489_ );
or   ( new_n26523_, new_n26367_, new_n26161_ );
or   ( new_n26524_, new_n26364_, new_n26170_ );
and  ( new_n26525_, new_n26524_, new_n26523_ );
or   ( new_n26526_, new_n26525_, new_n26372_ );
and  ( new_n26527_, new_n26368_, new_n26171_ );
or   ( new_n26528_, new_n26527_, new_n26181_ );
and  ( new_n26529_, new_n26528_, new_n26526_ );
or   ( new_n26530_, new_n26529_, new_n26522_ );
and  ( new_n26531_, new_n26530_, new_n26521_ );
or   ( new_n26532_, new_n20557_, new_n1310_ );
or   ( new_n26533_, new_n20562_, new_n1002_ );
and  ( new_n26534_, new_n26533_, new_n26532_ );
or   ( new_n26535_, new_n26534_, new_n20156_ );
and  ( new_n26536_, new_n20566_, RI2b1c4342db70_79 );
and  ( new_n26537_, new_n20553_, RI2b1c4342daf8_78 );
or   ( new_n26538_, new_n26537_, new_n26536_ );
or   ( new_n26539_, new_n26538_, new_n20443_ );
and  ( new_n26540_, new_n26539_, new_n26535_ );
or   ( new_n26541_, new_n19758_, new_n126_ );
or   ( new_n26542_, new_n19763_, new_n1511_ );
and  ( new_n26543_, new_n26542_, new_n26541_ );
or   ( new_n26544_, new_n26543_, new_n19394_ );
and  ( new_n26545_, new_n19767_, RI2b1c4342dc60_81 );
and  ( new_n26546_, new_n19754_, RI2b1c4342dbe8_80 );
or   ( new_n26547_, new_n26546_, new_n26545_ );
or   ( new_n26548_, new_n26547_, new_n19659_ );
and  ( new_n26549_, new_n26548_, new_n26544_ );
or   ( new_n26550_, new_n26549_, new_n26540_ );
and  ( new_n26551_, new_n26549_, new_n26540_ );
or   ( new_n26552_, new_n19048_, new_n121_ );
or   ( new_n26553_, new_n19055_, new_n2119_ );
and  ( new_n26554_, new_n26553_, new_n26552_ );
or   ( new_n26555_, new_n26554_, new_n18742_ );
and  ( new_n26556_, new_n19057_, RI2b1c4342dd50_83 );
and  ( new_n26557_, new_n19044_, RI2b1c4342dcd8_82 );
or   ( new_n26558_, new_n26557_, new_n26556_ );
or   ( new_n26559_, new_n26558_, new_n18977_ );
and  ( new_n26560_, new_n26559_, new_n26555_ );
or   ( new_n26561_, new_n26560_, new_n26551_ );
and  ( new_n26562_, new_n26561_, new_n26550_ );
nor  ( new_n26563_, new_n22333_, new_n843_ );
nor  ( new_n26564_, new_n26563_, new_n11434_ );
or   ( new_n26565_, new_n26564_, new_n21261_ );
and  ( new_n26566_, new_n22337_, RI2b1c4342d990_75 );
and  ( new_n26567_, new_n22330_, RI2b1c4342d918_74 );
or   ( new_n26568_, new_n26567_, new_n26566_ );
or   ( new_n26569_, new_n26568_, new_n21009_ );
and  ( new_n26570_, new_n26569_, new_n26565_ );
and  ( new_n26571_, new_n26570_, new_n16029_ );
or   ( new_n26572_, new_n26570_, new_n16029_ );
or   ( new_n26573_, new_n21419_, new_n1004_ );
or   ( new_n26574_, new_n21424_, new_n886_ );
and  ( new_n26575_, new_n26574_, new_n26573_ );
or   ( new_n26576_, new_n26575_, new_n21013_ );
and  ( new_n26577_, new_n21428_, RI2b1c4342da80_77 );
and  ( new_n26578_, new_n21415_, RI2b1c4342da08_76 );
or   ( new_n26579_, new_n26578_, new_n26577_ );
or   ( new_n26580_, new_n26579_, new_n21265_ );
and  ( new_n26581_, new_n26580_, new_n26576_ );
and  ( new_n26582_, new_n26581_, new_n26572_ );
or   ( new_n26583_, new_n26582_, new_n26571_ );
and  ( new_n26584_, new_n26583_, new_n26562_ );
or   ( new_n26585_, new_n26583_, new_n26562_ );
or   ( new_n26586_, new_n18388_, new_n2806_ );
or   ( new_n26587_, new_n18395_, new_n2541_ );
and  ( new_n26588_, new_n26587_, new_n26586_ );
or   ( new_n26589_, new_n26588_, new_n18066_ );
and  ( new_n26590_, new_n18397_, RI2b1c4342de40_85 );
and  ( new_n26591_, new_n18384_, RI2b1c4342ddc8_84 );
or   ( new_n26592_, new_n26591_, new_n26590_ );
or   ( new_n26593_, new_n26592_, new_n18309_ );
and  ( new_n26594_, new_n26593_, new_n26589_ );
or   ( new_n26595_, new_n17727_, new_n3924_ );
or   ( new_n26596_, new_n17734_, new_n3239_ );
and  ( new_n26597_, new_n26596_, new_n26595_ );
or   ( new_n26598_, new_n26597_, new_n17238_ );
and  ( new_n26599_, new_n17736_, RI2b1c4342df30_87 );
and  ( new_n26600_, new_n17723_, RI2b1c4342deb8_86 );
or   ( new_n26601_, new_n26600_, new_n26599_ );
or   ( new_n26602_, new_n26601_, new_n17650_ );
and  ( new_n26603_, new_n26602_, new_n26598_ );
or   ( new_n26604_, new_n26603_, new_n26594_ );
and  ( new_n26605_, new_n26603_, new_n26594_ );
or   ( new_n26606_, new_n17244_, new_n132_ );
or   ( new_n26607_, new_n17248_, new_n3902_ );
and  ( new_n26608_, new_n26607_, new_n26606_ );
or   ( new_n26609_, new_n26608_, new_n16814_ );
and  ( new_n26610_, new_n17255_, RI2b1c4342e020_89 );
and  ( new_n26611_, new_n17240_, RI2b1c4342dfa8_88 );
or   ( new_n26612_, new_n26611_, new_n26610_ );
or   ( new_n26613_, new_n26612_, new_n17142_ );
and  ( new_n26614_, new_n26613_, new_n26609_ );
or   ( new_n26615_, new_n26614_, new_n26605_ );
and  ( new_n26616_, new_n26615_, new_n26604_ );
and  ( new_n26617_, new_n26616_, new_n26585_ );
or   ( new_n26618_, new_n26617_, new_n26584_ );
and  ( new_n26619_, new_n26618_, new_n26531_ );
or   ( new_n26620_, new_n26618_, new_n26531_ );
or   ( new_n26621_, new_n26352_, new_n26128_ );
or   ( new_n26622_, new_n26349_, new_n26137_ );
and  ( new_n26623_, new_n26622_, new_n26621_ );
or   ( new_n26624_, new_n26623_, new_n26357_ );
and  ( new_n26625_, new_n26353_, new_n26138_ );
or   ( new_n26626_, new_n26625_, new_n26148_ );
and  ( new_n26627_, new_n26626_, new_n26624_ );
or   ( new_n26628_, new_n26339_, new_n26097_ );
or   ( new_n26629_, new_n26336_, new_n26106_ );
and  ( new_n26630_, new_n26629_, new_n26628_ );
or   ( new_n26631_, new_n26630_, new_n26344_ );
and  ( new_n26632_, new_n26340_, new_n26107_ );
or   ( new_n26633_, new_n26632_, new_n26117_ );
and  ( new_n26634_, new_n26633_, new_n26631_ );
or   ( new_n26635_, new_n26634_, new_n26627_ );
and  ( new_n26636_, new_n26635_, new_n26620_ );
or   ( new_n26637_, new_n26636_, new_n26619_ );
and  ( new_n26638_, new_n26637_, new_n26482_ );
or   ( new_n26639_, new_n26637_, new_n26482_ );
or   ( new_n26640_, new_n26014_, new_n25838_ );
or   ( new_n26641_, new_n26024_, new_n25817_ );
and  ( new_n26642_, new_n26641_, new_n26640_ );
or   ( new_n26643_, new_n26642_, new_n26039_ );
and  ( new_n26644_, new_n26025_, new_n25840_ );
or   ( new_n26645_, new_n26644_, new_n25871_ );
and  ( new_n26646_, new_n26645_, new_n26643_ );
and  ( new_n26647_, new_n26646_, new_n26639_ );
or   ( new_n26648_, new_n26647_, new_n26638_ );
and  ( new_n26649_, new_n26648_, new_n26457_ );
or   ( new_n26650_, new_n26648_, new_n26457_ );
or   ( new_n26651_, new_n26001_, new_n25873_ );
or   ( new_n26652_, new_n26041_, new_n25786_ );
and  ( new_n26653_, new_n26652_, new_n26651_ );
or   ( new_n26654_, new_n26653_, new_n26056_ );
and  ( new_n26655_, new_n26042_, new_n25875_ );
or   ( new_n26656_, new_n26655_, new_n25900_ );
and  ( new_n26657_, new_n26656_, new_n26654_ );
and  ( new_n26658_, new_n26657_, new_n26650_ );
or   ( new_n26659_, new_n26658_, new_n26649_ );
or   ( new_n26660_, new_n26659_, new_n26442_ );
or   ( new_n26661_, new_n26312_, new_n26070_ );
or   ( new_n26662_, new_n26310_, new_n25922_ );
and  ( new_n26663_, new_n26662_, new_n26661_ );
or   ( new_n26664_, new_n25946_, new_n25943_ );
and  ( new_n26665_, new_n26664_, new_n25677_ );
or   ( new_n26666_, new_n26665_, new_n26306_ );
and  ( new_n26667_, new_n26435_, new_n26332_ );
or   ( new_n26668_, new_n26667_, new_n26329_ );
and  ( new_n26669_, new_n26668_, new_n26439_ );
or   ( new_n26670_, new_n26669_, new_n26082_ );
and  ( new_n26671_, new_n26670_, new_n26666_ );
or   ( new_n26672_, new_n26671_, new_n26663_ );
or   ( new_n26673_, new_n26669_, new_n26665_ );
and  ( new_n26674_, new_n26673_, new_n26307_ );
or   ( new_n26675_, new_n26674_, new_n26314_ );
and  ( new_n26676_, new_n26675_, new_n26672_ );
or   ( new_n26677_, new_n26676_, new_n26660_ );
and  ( new_n26678_, new_n26676_, new_n26660_ );
or   ( new_n26679_, new_n26428_, new_n26259_ );
or   ( new_n26680_, new_n26415_, new_n26284_ );
and  ( new_n26681_, new_n26680_, new_n26679_ );
or   ( new_n26682_, new_n26681_, new_n26433_ );
and  ( new_n26683_, new_n26429_, new_n26285_ );
or   ( new_n26684_, new_n26683_, new_n26293_ );
and  ( new_n26685_, new_n26684_, new_n26682_ );
or   ( new_n26686_, new_n26655_, new_n26056_ );
or   ( new_n26687_, new_n26653_, new_n25900_ );
and  ( new_n26688_, new_n26687_, new_n26686_ );
or   ( new_n26689_, new_n26447_, new_n26426_ );
or   ( new_n26690_, new_n26445_, new_n26282_ );
and  ( new_n26691_, new_n26690_, new_n26689_ );
or   ( new_n26692_, new_n26454_, new_n26413_ );
or   ( new_n26693_, new_n26452_, new_n26257_ );
and  ( new_n26694_, new_n26693_, new_n26692_ );
and  ( new_n26695_, new_n26694_, new_n26691_ );
or   ( new_n26696_, new_n26695_, new_n26648_ );
or   ( new_n26697_, new_n26462_, new_n26411_ );
or   ( new_n26698_, new_n26460_, new_n26255_ );
and  ( new_n26699_, new_n26698_, new_n26697_ );
or   ( new_n26700_, new_n26469_, new_n26396_ );
or   ( new_n26701_, new_n26467_, new_n26228_ );
and  ( new_n26702_, new_n26701_, new_n26700_ );
or   ( new_n26703_, new_n26702_, new_n26699_ );
and  ( new_n26704_, new_n26702_, new_n26699_ );
or   ( new_n26705_, new_n26478_, new_n26374_ );
or   ( new_n26706_, new_n26476_, new_n26183_ );
and  ( new_n26707_, new_n26706_, new_n26705_ );
or   ( new_n26708_, new_n26707_, new_n26704_ );
and  ( new_n26709_, new_n26708_, new_n26703_ );
or   ( new_n26710_, new_n26487_, new_n26389_ );
or   ( new_n26711_, new_n26485_, new_n26217_ );
and  ( new_n26712_, new_n26711_, new_n26710_ );
or   ( new_n26713_, new_n26496_, new_n16505_ );
or   ( new_n26714_, new_n26492_, new_n16438_ );
and  ( new_n26715_, new_n26714_, new_n26713_ );
or   ( new_n26716_, new_n26505_, new_n16085_ );
or   ( new_n26717_, new_n26501_, new_n16048_ );
and  ( new_n26718_, new_n26717_, new_n26716_ );
or   ( new_n26719_, new_n26718_, new_n26715_ );
and  ( new_n26720_, new_n26718_, new_n26715_ );
or   ( new_n26721_, new_n26516_, new_n16052_ );
or   ( new_n26722_, new_n26512_, new_n16071_ );
and  ( new_n26723_, new_n26722_, new_n26721_ );
or   ( new_n26724_, new_n26723_, new_n26720_ );
and  ( new_n26725_, new_n26724_, new_n26719_ );
or   ( new_n26726_, new_n26725_, new_n26712_ );
and  ( new_n26727_, new_n26725_, new_n26712_ );
or   ( new_n26728_, new_n26527_, new_n26372_ );
or   ( new_n26729_, new_n26525_, new_n26181_ );
and  ( new_n26730_, new_n26729_, new_n26728_ );
or   ( new_n26731_, new_n26730_, new_n26727_ );
and  ( new_n26732_, new_n26731_, new_n26726_ );
or   ( new_n26733_, new_n26538_, new_n20156_ );
or   ( new_n26734_, new_n26534_, new_n20443_ );
and  ( new_n26735_, new_n26734_, new_n26733_ );
or   ( new_n26736_, new_n26547_, new_n19394_ );
or   ( new_n26737_, new_n26543_, new_n19659_ );
and  ( new_n26738_, new_n26737_, new_n26736_ );
or   ( new_n26739_, new_n26738_, new_n26735_ );
and  ( new_n26740_, new_n26738_, new_n26735_ );
or   ( new_n26741_, new_n26558_, new_n18742_ );
or   ( new_n26742_, new_n26554_, new_n18977_ );
and  ( new_n26743_, new_n26742_, new_n26741_ );
or   ( new_n26744_, new_n26743_, new_n26740_ );
and  ( new_n26745_, new_n26744_, new_n26739_ );
or   ( new_n26746_, new_n26568_, new_n21261_ );
or   ( new_n26747_, new_n26564_, new_n21009_ );
and  ( new_n26748_, new_n26747_, new_n26746_ );
or   ( new_n26749_, new_n26748_, new_n16009_ );
and  ( new_n26750_, new_n26748_, new_n16009_ );
or   ( new_n26751_, new_n26579_, new_n21013_ );
or   ( new_n26752_, new_n26575_, new_n21265_ );
and  ( new_n26753_, new_n26752_, new_n26751_ );
or   ( new_n26754_, new_n26753_, new_n26750_ );
and  ( new_n26755_, new_n26754_, new_n26749_ );
or   ( new_n26756_, new_n26755_, new_n26745_ );
and  ( new_n26757_, new_n26755_, new_n26745_ );
or   ( new_n26758_, new_n26592_, new_n18066_ );
or   ( new_n26759_, new_n26588_, new_n18309_ );
and  ( new_n26760_, new_n26759_, new_n26758_ );
or   ( new_n26761_, new_n26601_, new_n17238_ );
or   ( new_n26762_, new_n26597_, new_n17650_ );
and  ( new_n26763_, new_n26762_, new_n26761_ );
or   ( new_n26764_, new_n26763_, new_n26760_ );
and  ( new_n26765_, new_n26763_, new_n26760_ );
or   ( new_n26766_, new_n26612_, new_n16814_ );
or   ( new_n26767_, new_n26608_, new_n17142_ );
and  ( new_n26768_, new_n26767_, new_n26766_ );
or   ( new_n26769_, new_n26768_, new_n26765_ );
and  ( new_n26770_, new_n26769_, new_n26764_ );
or   ( new_n26771_, new_n26770_, new_n26757_ );
and  ( new_n26772_, new_n26771_, new_n26756_ );
or   ( new_n26773_, new_n26772_, new_n26732_ );
and  ( new_n26774_, new_n26772_, new_n26732_ );
or   ( new_n26775_, new_n26625_, new_n26357_ );
or   ( new_n26776_, new_n26623_, new_n26148_ );
and  ( new_n26777_, new_n26776_, new_n26775_ );
or   ( new_n26778_, new_n26632_, new_n26344_ );
or   ( new_n26779_, new_n26630_, new_n26117_ );
and  ( new_n26780_, new_n26779_, new_n26778_ );
and  ( new_n26781_, new_n26780_, new_n26777_ );
or   ( new_n26782_, new_n26781_, new_n26774_ );
and  ( new_n26783_, new_n26782_, new_n26773_ );
or   ( new_n26784_, new_n26783_, new_n26709_ );
and  ( new_n26785_, new_n26783_, new_n26709_ );
or   ( new_n26786_, new_n26644_, new_n26039_ );
or   ( new_n26787_, new_n26642_, new_n25871_ );
and  ( new_n26788_, new_n26787_, new_n26786_ );
or   ( new_n26789_, new_n26788_, new_n26785_ );
and  ( new_n26790_, new_n26789_, new_n26784_ );
or   ( new_n26791_, new_n26790_, new_n26457_ );
and  ( new_n26792_, new_n26791_, new_n26696_ );
or   ( new_n26793_, new_n26792_, new_n26688_ );
or   ( new_n26794_, new_n26790_, new_n26695_ );
and  ( new_n26795_, new_n26794_, new_n26650_ );
or   ( new_n26796_, new_n26795_, new_n26657_ );
and  ( new_n26797_, new_n26796_, new_n26793_ );
or   ( new_n26798_, new_n26797_, new_n26685_ );
or   ( new_n26799_, new_n26440_, new_n26329_ );
or   ( new_n26800_, new_n26437_, new_n26304_ );
and  ( new_n26801_, new_n26800_, new_n26799_ );
or   ( new_n26802_, new_n26801_, new_n26659_ );
and  ( new_n26803_, new_n26790_, new_n26695_ );
or   ( new_n26804_, new_n26803_, new_n26688_ );
and  ( new_n26805_, new_n26804_, new_n26794_ );
or   ( new_n26806_, new_n26805_, new_n26442_ );
and  ( new_n26807_, new_n26806_, new_n26802_ );
or   ( new_n26808_, new_n26807_, new_n26798_ );
or   ( new_n26809_, new_n26808_, new_n26678_ );
and  ( new_n26810_, new_n26809_, new_n26677_ );
and  ( new_n26811_, new_n26807_, new_n26798_ );
or   ( new_n26812_, new_n26811_, new_n26678_ );
or   ( new_n26813_, new_n26795_, new_n26688_ );
or   ( new_n26814_, new_n26792_, new_n26657_ );
and  ( new_n26815_, new_n26814_, new_n26813_ );
or   ( new_n26816_, new_n26815_, new_n26685_ );
or   ( new_n26817_, new_n26683_, new_n26433_ );
or   ( new_n26818_, new_n26681_, new_n26293_ );
and  ( new_n26819_, new_n26818_, new_n26817_ );
or   ( new_n26820_, new_n26819_, new_n26797_ );
and  ( new_n26821_, new_n26820_, new_n26816_ );
or   ( new_n26822_, new_n26694_, new_n26449_ );
or   ( new_n26823_, new_n26691_, new_n26456_ );
and  ( new_n26824_, new_n26823_, new_n26822_ );
nor  ( new_n26825_, new_n22333_, new_n886_ );
nor  ( new_n26826_, new_n26825_, new_n11680_ );
or   ( new_n26827_, new_n26826_, new_n21261_ );
and  ( new_n26828_, new_n22337_, RI2b1c4342da08_76 );
and  ( new_n26829_, new_n22330_, RI2b1c4342d990_75 );
or   ( new_n26830_, new_n26829_, new_n26828_ );
or   ( new_n26831_, new_n26830_, new_n21009_ );
and  ( new_n26832_, new_n26831_, new_n26827_ );
or   ( new_n26833_, new_n21419_, new_n1002_ );
or   ( new_n26834_, new_n21424_, new_n1004_ );
and  ( new_n26835_, new_n26834_, new_n26833_ );
or   ( new_n26836_, new_n26835_, new_n21013_ );
and  ( new_n26837_, new_n21428_, RI2b1c4342daf8_78 );
and  ( new_n26838_, new_n21415_, RI2b1c4342da80_77 );
or   ( new_n26839_, new_n26838_, new_n26837_ );
or   ( new_n26840_, new_n26839_, new_n21265_ );
and  ( new_n26841_, new_n26840_, new_n26836_ );
or   ( new_n26842_, new_n26841_, new_n26832_ );
and  ( new_n26843_, new_n26841_, new_n26832_ );
or   ( new_n26844_, new_n20557_, new_n1511_ );
or   ( new_n26845_, new_n20562_, new_n1310_ );
and  ( new_n26846_, new_n26845_, new_n26844_ );
or   ( new_n26847_, new_n26846_, new_n20156_ );
and  ( new_n26848_, new_n20566_, RI2b1c4342dbe8_80 );
and  ( new_n26849_, new_n20553_, RI2b1c4342db70_79 );
or   ( new_n26850_, new_n26849_, new_n26848_ );
or   ( new_n26851_, new_n26850_, new_n20443_ );
and  ( new_n26852_, new_n26851_, new_n26847_ );
or   ( new_n26853_, new_n26852_, new_n26843_ );
and  ( new_n26854_, new_n26853_, new_n26842_ );
or   ( new_n26855_, new_n19758_, new_n2119_ );
or   ( new_n26856_, new_n19763_, new_n126_ );
and  ( new_n26857_, new_n26856_, new_n26855_ );
or   ( new_n26858_, new_n26857_, new_n19394_ );
and  ( new_n26859_, new_n19767_, RI2b1c4342dcd8_82 );
and  ( new_n26860_, new_n19754_, RI2b1c4342dc60_81 );
or   ( new_n26861_, new_n26860_, new_n26859_ );
or   ( new_n26862_, new_n26861_, new_n19659_ );
and  ( new_n26863_, new_n26862_, new_n26858_ );
or   ( new_n26864_, new_n19048_, new_n2541_ );
or   ( new_n26865_, new_n19055_, new_n121_ );
and  ( new_n26866_, new_n26865_, new_n26864_ );
or   ( new_n26867_, new_n26866_, new_n18742_ );
and  ( new_n26868_, new_n19057_, RI2b1c4342ddc8_84 );
and  ( new_n26869_, new_n19044_, RI2b1c4342dd50_83 );
or   ( new_n26870_, new_n26869_, new_n26868_ );
or   ( new_n26871_, new_n26870_, new_n18977_ );
and  ( new_n26872_, new_n26871_, new_n26867_ );
or   ( new_n26873_, new_n26872_, new_n26863_ );
and  ( new_n26874_, new_n26872_, new_n26863_ );
or   ( new_n26875_, new_n18388_, new_n3239_ );
or   ( new_n26876_, new_n18395_, new_n2806_ );
and  ( new_n26877_, new_n26876_, new_n26875_ );
or   ( new_n26878_, new_n26877_, new_n18066_ );
and  ( new_n26879_, new_n18397_, RI2b1c4342deb8_86 );
and  ( new_n26880_, new_n18384_, RI2b1c4342de40_85 );
or   ( new_n26881_, new_n26880_, new_n26879_ );
or   ( new_n26882_, new_n26881_, new_n18309_ );
and  ( new_n26883_, new_n26882_, new_n26878_ );
or   ( new_n26884_, new_n26883_, new_n26874_ );
and  ( new_n26885_, new_n26884_, new_n26873_ );
or   ( new_n26886_, new_n26885_, new_n26854_ );
and  ( new_n26887_, new_n26885_, new_n26854_ );
or   ( new_n26888_, new_n17727_, new_n3902_ );
or   ( new_n26889_, new_n17734_, new_n3924_ );
and  ( new_n26890_, new_n26889_, new_n26888_ );
or   ( new_n26891_, new_n26890_, new_n17238_ );
and  ( new_n26892_, new_n17736_, RI2b1c4342dfa8_88 );
and  ( new_n26893_, new_n17723_, RI2b1c4342df30_87 );
or   ( new_n26894_, new_n26893_, new_n26892_ );
or   ( new_n26895_, new_n26894_, new_n17650_ );
and  ( new_n26896_, new_n26895_, new_n26891_ );
or   ( new_n26897_, new_n17244_, new_n4635_ );
or   ( new_n26898_, new_n17248_, new_n132_ );
and  ( new_n26899_, new_n26898_, new_n26897_ );
or   ( new_n26900_, new_n26899_, new_n16814_ );
and  ( new_n26901_, new_n17255_, RI2b1c4342e098_90 );
and  ( new_n26902_, new_n17240_, RI2b1c4342e020_89 );
or   ( new_n26903_, new_n26902_, new_n26901_ );
or   ( new_n26904_, new_n26903_, new_n17142_ );
and  ( new_n26905_, new_n26904_, new_n26900_ );
or   ( new_n26906_, new_n26905_, new_n26896_ );
and  ( new_n26907_, new_n26905_, new_n26896_ );
or   ( new_n26908_, new_n16607_, new_n5459_ );
or   ( new_n26909_, new_n16613_, new_n117_ );
and  ( new_n26910_, new_n26909_, new_n26908_ );
or   ( new_n26911_, new_n26910_, new_n16505_ );
and  ( new_n26912_, new_n16616_, RI2b1c4342e188_92 );
and  ( new_n26913_, new_n16603_, RI2b1c4342e110_91 );
or   ( new_n26914_, new_n26913_, new_n26912_ );
or   ( new_n26915_, new_n26914_, new_n16438_ );
and  ( new_n26916_, new_n26915_, new_n26911_ );
or   ( new_n26917_, new_n26916_, new_n26907_ );
and  ( new_n26918_, new_n26917_, new_n26906_ );
or   ( new_n26919_, new_n26918_, new_n26887_ );
and  ( new_n26920_, new_n26919_, new_n26886_ );
or   ( new_n26921_, new_n16017_, new_n7274_ );
or   ( new_n26922_, new_n26921_, new_n16009_ );
and  ( new_n26923_, new_n16024_, RI2b1c4342e368_96 );
or   ( new_n26924_, new_n26923_, new_n16029_ );
and  ( new_n26925_, new_n26924_, new_n26922_ );
or   ( new_n26926_, new_n26718_, new_n26498_ );
or   ( new_n26927_, new_n26715_, new_n26507_ );
and  ( new_n26928_, new_n26927_, new_n26926_ );
or   ( new_n26929_, new_n26928_, new_n26723_ );
and  ( new_n26930_, new_n26719_, new_n26508_ );
or   ( new_n26931_, new_n26930_, new_n26518_ );
and  ( new_n26932_, new_n26931_, new_n26929_ );
or   ( new_n26933_, new_n26932_, new_n26925_ );
and  ( new_n26934_, new_n26932_, new_n26925_ );
or   ( new_n26935_, new_n26763_, new_n26594_ );
or   ( new_n26936_, new_n26760_, new_n26603_ );
and  ( new_n26937_, new_n26936_, new_n26935_ );
or   ( new_n26938_, new_n26937_, new_n26768_ );
and  ( new_n26939_, new_n26764_, new_n26604_ );
or   ( new_n26940_, new_n26939_, new_n26614_ );
and  ( new_n26941_, new_n26940_, new_n26938_ );
or   ( new_n26942_, new_n26941_, new_n26934_ );
and  ( new_n26943_, new_n26942_, new_n26933_ );
or   ( new_n26944_, new_n26943_, new_n26920_ );
and  ( new_n26945_, new_n26943_, new_n26920_ );
or   ( new_n26946_, new_n26738_, new_n26540_ );
or   ( new_n26947_, new_n26735_, new_n26549_ );
and  ( new_n26948_, new_n26947_, new_n26946_ );
or   ( new_n26949_, new_n26948_, new_n26743_ );
and  ( new_n26950_, new_n26739_, new_n26550_ );
or   ( new_n26951_, new_n26950_, new_n26560_ );
and  ( new_n26952_, new_n26951_, new_n26949_ );
or   ( new_n26953_, new_n26748_, new_n16029_ );
or   ( new_n26954_, new_n26570_, new_n16009_ );
and  ( new_n26955_, new_n26954_, new_n26953_ );
or   ( new_n26956_, new_n26955_, new_n26753_ );
and  ( new_n26957_, new_n26749_, new_n26572_ );
or   ( new_n26958_, new_n26957_, new_n26581_ );
and  ( new_n26959_, new_n26958_, new_n26956_ );
or   ( new_n26960_, new_n26959_, new_n26952_ );
or   ( new_n26961_, new_n26960_, new_n26945_ );
and  ( new_n26962_, new_n26961_, new_n26944_ );
or   ( new_n26963_, new_n26780_, new_n26627_ );
or   ( new_n26964_, new_n26777_, new_n26634_ );
and  ( new_n26965_, new_n26964_, new_n26963_ );
or   ( new_n26966_, new_n26712_, new_n26520_ );
or   ( new_n26967_, new_n26725_, new_n26489_ );
and  ( new_n26968_, new_n26967_, new_n26966_ );
or   ( new_n26969_, new_n26968_, new_n26730_ );
and  ( new_n26970_, new_n26726_, new_n26521_ );
or   ( new_n26971_, new_n26970_, new_n26529_ );
and  ( new_n26972_, new_n26971_, new_n26969_ );
or   ( new_n26973_, new_n26972_, new_n26965_ );
and  ( new_n26974_, new_n26972_, new_n26965_ );
or   ( new_n26975_, new_n26745_, new_n26583_ );
or   ( new_n26976_, new_n26755_, new_n26562_ );
and  ( new_n26977_, new_n26976_, new_n26975_ );
or   ( new_n26978_, new_n26977_, new_n26770_ );
and  ( new_n26979_, new_n26756_, new_n26585_ );
or   ( new_n26980_, new_n26979_, new_n26616_ );
and  ( new_n26981_, new_n26980_, new_n26978_ );
or   ( new_n26982_, new_n26981_, new_n26974_ );
and  ( new_n26983_, new_n26982_, new_n26973_ );
or   ( new_n26984_, new_n26983_, new_n26962_ );
and  ( new_n26985_, new_n26983_, new_n26962_ );
or   ( new_n26986_, new_n26702_, new_n26464_ );
or   ( new_n26987_, new_n26699_, new_n26471_ );
and  ( new_n26988_, new_n26987_, new_n26986_ );
or   ( new_n26989_, new_n26988_, new_n26707_ );
and  ( new_n26990_, new_n26703_, new_n26472_ );
or   ( new_n26991_, new_n26990_, new_n26480_ );
and  ( new_n26992_, new_n26991_, new_n26989_ );
or   ( new_n26993_, new_n26992_, new_n26985_ );
and  ( new_n26994_, new_n26993_, new_n26984_ );
or   ( new_n26995_, new_n26994_, new_n26824_ );
or   ( new_n26996_, new_n26709_, new_n26637_ );
or   ( new_n26997_, new_n26783_, new_n26482_ );
and  ( new_n26998_, new_n26997_, new_n26996_ );
or   ( new_n26999_, new_n26998_, new_n26788_ );
and  ( new_n27000_, new_n26784_, new_n26639_ );
or   ( new_n27001_, new_n27000_, new_n26646_ );
and  ( new_n27002_, new_n27001_, new_n26999_ );
and  ( new_n27003_, new_n26994_, new_n26824_ );
or   ( new_n27004_, new_n27003_, new_n27002_ );
and  ( new_n27005_, new_n27004_, new_n26995_ );
or   ( new_n27006_, new_n27005_, new_n26821_ );
and  ( new_n27007_, new_n27005_, new_n26821_ );
or   ( new_n27008_, new_n27000_, new_n26788_ );
or   ( new_n27009_, new_n26998_, new_n26646_ );
and  ( new_n27010_, new_n27009_, new_n27008_ );
or   ( new_n27011_, new_n26694_, new_n26691_ );
and  ( new_n27012_, new_n27011_, new_n26457_ );
or   ( new_n27013_, new_n27012_, new_n26994_ );
or   ( new_n27014_, new_n26830_, new_n21261_ );
or   ( new_n27015_, new_n26826_, new_n21009_ );
and  ( new_n27016_, new_n27015_, new_n27014_ );
or   ( new_n27017_, new_n26839_, new_n21013_ );
or   ( new_n27018_, new_n26835_, new_n21265_ );
and  ( new_n27019_, new_n27018_, new_n27017_ );
or   ( new_n27020_, new_n27019_, new_n27016_ );
and  ( new_n27021_, new_n27019_, new_n27016_ );
or   ( new_n27022_, new_n26850_, new_n20156_ );
or   ( new_n27023_, new_n26846_, new_n20443_ );
and  ( new_n27024_, new_n27023_, new_n27022_ );
or   ( new_n27025_, new_n27024_, new_n27021_ );
and  ( new_n27026_, new_n27025_, new_n27020_ );
or   ( new_n27027_, new_n26861_, new_n19394_ );
or   ( new_n27028_, new_n26857_, new_n19659_ );
and  ( new_n27029_, new_n27028_, new_n27027_ );
or   ( new_n27030_, new_n26870_, new_n18742_ );
or   ( new_n27031_, new_n26866_, new_n18977_ );
and  ( new_n27032_, new_n27031_, new_n27030_ );
or   ( new_n27033_, new_n27032_, new_n27029_ );
and  ( new_n27034_, new_n27032_, new_n27029_ );
or   ( new_n27035_, new_n26881_, new_n18066_ );
or   ( new_n27036_, new_n26877_, new_n18309_ );
and  ( new_n27037_, new_n27036_, new_n27035_ );
or   ( new_n27038_, new_n27037_, new_n27034_ );
and  ( new_n27039_, new_n27038_, new_n27033_ );
or   ( new_n27040_, new_n27039_, new_n27026_ );
and  ( new_n27041_, new_n27039_, new_n27026_ );
or   ( new_n27042_, new_n26894_, new_n17238_ );
or   ( new_n27043_, new_n26890_, new_n17650_ );
and  ( new_n27044_, new_n27043_, new_n27042_ );
or   ( new_n27045_, new_n26903_, new_n16814_ );
or   ( new_n27046_, new_n26899_, new_n17142_ );
and  ( new_n27047_, new_n27046_, new_n27045_ );
or   ( new_n27048_, new_n27047_, new_n27044_ );
and  ( new_n27049_, new_n27047_, new_n27044_ );
or   ( new_n27050_, new_n26914_, new_n16505_ );
or   ( new_n27051_, new_n26910_, new_n16438_ );
and  ( new_n27052_, new_n27051_, new_n27050_ );
or   ( new_n27053_, new_n27052_, new_n27049_ );
and  ( new_n27054_, new_n27053_, new_n27048_ );
or   ( new_n27055_, new_n27054_, new_n27041_ );
and  ( new_n27056_, new_n27055_, new_n27040_ );
or   ( new_n27057_, new_n26923_, new_n16009_ );
or   ( new_n27058_, new_n26921_, new_n16029_ );
and  ( new_n27059_, new_n27058_, new_n27057_ );
or   ( new_n27060_, new_n26930_, new_n26723_ );
or   ( new_n27061_, new_n26928_, new_n26518_ );
and  ( new_n27062_, new_n27061_, new_n27060_ );
or   ( new_n27063_, new_n27062_, new_n27059_ );
and  ( new_n27064_, new_n27062_, new_n27059_ );
or   ( new_n27065_, new_n26939_, new_n26768_ );
or   ( new_n27066_, new_n26937_, new_n26614_ );
and  ( new_n27067_, new_n27066_, new_n27065_ );
or   ( new_n27068_, new_n27067_, new_n27064_ );
and  ( new_n27069_, new_n27068_, new_n27063_ );
or   ( new_n27070_, new_n27069_, new_n27056_ );
and  ( new_n27071_, new_n27069_, new_n27056_ );
or   ( new_n27072_, new_n26950_, new_n26743_ );
or   ( new_n27073_, new_n26948_, new_n26560_ );
and  ( new_n27074_, new_n27073_, new_n27072_ );
or   ( new_n27075_, new_n26957_, new_n26753_ );
or   ( new_n27076_, new_n26955_, new_n26581_ );
and  ( new_n27077_, new_n27076_, new_n27075_ );
and  ( new_n27078_, new_n27077_, new_n27074_ );
or   ( new_n27079_, new_n27078_, new_n27071_ );
and  ( new_n27080_, new_n27079_, new_n27070_ );
or   ( new_n27081_, new_n26780_, new_n26777_ );
and  ( new_n27082_, new_n27081_, new_n26635_ );
or   ( new_n27083_, new_n26970_, new_n26730_ );
or   ( new_n27084_, new_n26968_, new_n26529_ );
and  ( new_n27085_, new_n27084_, new_n27083_ );
or   ( new_n27086_, new_n27085_, new_n27082_ );
and  ( new_n27087_, new_n27085_, new_n27082_ );
or   ( new_n27088_, new_n26979_, new_n26770_ );
or   ( new_n27089_, new_n26977_, new_n26616_ );
and  ( new_n27090_, new_n27089_, new_n27088_ );
or   ( new_n27091_, new_n27090_, new_n27087_ );
and  ( new_n27092_, new_n27091_, new_n27086_ );
or   ( new_n27093_, new_n27092_, new_n27080_ );
and  ( new_n27094_, new_n27092_, new_n27080_ );
or   ( new_n27095_, new_n26990_, new_n26707_ );
or   ( new_n27096_, new_n26988_, new_n26480_ );
and  ( new_n27097_, new_n27096_, new_n27095_ );
or   ( new_n27098_, new_n27097_, new_n27094_ );
and  ( new_n27099_, new_n27098_, new_n27093_ );
or   ( new_n27100_, new_n27099_, new_n26824_ );
and  ( new_n27101_, new_n27100_, new_n27013_ );
or   ( new_n27102_, new_n27101_, new_n27010_ );
or   ( new_n27103_, new_n27099_, new_n27012_ );
and  ( new_n27104_, new_n27103_, new_n26995_ );
or   ( new_n27105_, new_n27104_, new_n27002_ );
and  ( new_n27106_, new_n27105_, new_n27102_ );
or   ( new_n27107_, new_n26732_, new_n26618_ );
or   ( new_n27108_, new_n26772_, new_n26531_ );
and  ( new_n27109_, new_n27108_, new_n27107_ );
or   ( new_n27110_, new_n27109_, new_n26781_ );
and  ( new_n27111_, new_n26773_, new_n26620_ );
or   ( new_n27112_, new_n27111_, new_n26635_ );
and  ( new_n27113_, new_n27112_, new_n27110_ );
or   ( new_n27114_, new_n27077_, new_n26952_ );
or   ( new_n27115_, new_n27074_, new_n26959_ );
and  ( new_n27116_, new_n27115_, new_n27114_ );
or   ( new_n27117_, new_n27062_, new_n26925_ );
or   ( new_n27118_, new_n27059_, new_n26932_ );
and  ( new_n27119_, new_n27118_, new_n27117_ );
or   ( new_n27120_, new_n27119_, new_n27067_ );
and  ( new_n27121_, new_n27063_, new_n26933_ );
or   ( new_n27122_, new_n27121_, new_n26941_ );
and  ( new_n27123_, new_n27122_, new_n27120_ );
or   ( new_n27124_, new_n27123_, new_n27116_ );
and  ( new_n27125_, new_n27123_, new_n27116_ );
or   ( new_n27126_, new_n27039_, new_n26854_ );
or   ( new_n27127_, new_n27026_, new_n26885_ );
and  ( new_n27128_, new_n27127_, new_n27126_ );
or   ( new_n27129_, new_n27128_, new_n27054_ );
and  ( new_n27130_, new_n27040_, new_n26886_ );
or   ( new_n27131_, new_n27130_, new_n26918_ );
and  ( new_n27132_, new_n27131_, new_n27129_ );
or   ( new_n27133_, new_n27132_, new_n27125_ );
and  ( new_n27134_, new_n27133_, new_n27124_ );
or   ( new_n27135_, new_n16366_, new_n6321_ );
or   ( new_n27136_, new_n16355_, new_n6307_ );
and  ( new_n27137_, new_n27136_, new_n27135_ );
or   ( new_n27138_, new_n27137_, new_n16085_ );
and  ( new_n27139_, new_n16358_, RI2b1c4342e278_94 );
and  ( new_n27140_, new_n16362_, RI2b1c4342e200_93 );
or   ( new_n27141_, new_n27140_, new_n27139_ );
or   ( new_n27142_, new_n27141_, new_n16048_ );
and  ( new_n27143_, new_n27142_, new_n27138_ );
or   ( new_n27144_, new_n16607_, new_n6307_ );
or   ( new_n27145_, new_n16613_, new_n5459_ );
and  ( new_n27146_, new_n27145_, new_n27144_ );
or   ( new_n27147_, new_n27146_, new_n16505_ );
and  ( new_n27148_, new_n16616_, RI2b1c4342e200_93 );
and  ( new_n27149_, new_n16603_, RI2b1c4342e188_92 );
or   ( new_n27150_, new_n27149_, new_n27148_ );
or   ( new_n27151_, new_n27150_, new_n16438_ );
and  ( new_n27152_, new_n27151_, new_n27147_ );
or   ( new_n27153_, new_n16366_, new_n124_ );
or   ( new_n27154_, new_n16355_, new_n6321_ );
and  ( new_n27155_, new_n27154_, new_n27153_ );
or   ( new_n27156_, new_n27155_, new_n16085_ );
and  ( new_n27157_, new_n16358_, RI2b1c4342e2f0_95 );
and  ( new_n27158_, new_n16362_, RI2b1c4342e278_94 );
or   ( new_n27159_, new_n27158_, new_n27157_ );
or   ( new_n27160_, new_n27159_, new_n16048_ );
and  ( new_n27161_, new_n27160_, new_n27156_ );
or   ( new_n27162_, new_n27161_, new_n27152_ );
and  ( new_n27163_, new_n27161_, new_n27152_ );
or   ( new_n27164_, new_n16060_, new_n7274_ );
or   ( new_n27165_, new_n27164_, new_n16052_ );
and  ( new_n27166_, new_n16066_, RI2b1c4342e368_96 );
or   ( new_n27167_, new_n27166_, new_n16071_ );
and  ( new_n27168_, new_n27167_, new_n27165_ );
or   ( new_n27169_, new_n27168_, new_n27163_ );
and  ( new_n27170_, new_n27169_, new_n27162_ );
or   ( new_n27171_, new_n27170_, new_n27143_ );
and  ( new_n27172_, new_n27170_, new_n27143_ );
or   ( new_n27173_, new_n16075_, new_n7274_ );
or   ( new_n27174_, new_n16060_, new_n124_ );
and  ( new_n27175_, new_n27174_, new_n27173_ );
or   ( new_n27176_, new_n27175_, new_n16052_ );
and  ( new_n27177_, new_n16063_, RI2b1c4342e368_96 );
and  ( new_n27178_, new_n16066_, RI2b1c4342e2f0_95 );
or   ( new_n27179_, new_n27178_, new_n27177_ );
or   ( new_n27180_, new_n27179_, new_n16071_ );
and  ( new_n27181_, new_n27180_, new_n27176_ );
or   ( new_n27182_, new_n27181_, new_n27172_ );
and  ( new_n27183_, new_n27182_, new_n27171_ );
or   ( new_n27184_, new_n20557_, new_n126_ );
or   ( new_n27185_, new_n20562_, new_n1511_ );
and  ( new_n27186_, new_n27185_, new_n27184_ );
or   ( new_n27187_, new_n27186_, new_n20156_ );
and  ( new_n27188_, new_n20566_, RI2b1c4342dc60_81 );
and  ( new_n27189_, new_n20553_, RI2b1c4342dbe8_80 );
or   ( new_n27190_, new_n27189_, new_n27188_ );
or   ( new_n27191_, new_n27190_, new_n20443_ );
and  ( new_n27192_, new_n27191_, new_n27187_ );
or   ( new_n27193_, new_n19758_, new_n121_ );
or   ( new_n27194_, new_n19763_, new_n2119_ );
and  ( new_n27195_, new_n27194_, new_n27193_ );
or   ( new_n27196_, new_n27195_, new_n19394_ );
and  ( new_n27197_, new_n19767_, RI2b1c4342dd50_83 );
and  ( new_n27198_, new_n19754_, RI2b1c4342dcd8_82 );
or   ( new_n27199_, new_n27198_, new_n27197_ );
or   ( new_n27200_, new_n27199_, new_n19659_ );
and  ( new_n27201_, new_n27200_, new_n27196_ );
or   ( new_n27202_, new_n27201_, new_n27192_ );
and  ( new_n27203_, new_n27201_, new_n27192_ );
or   ( new_n27204_, new_n19048_, new_n2806_ );
or   ( new_n27205_, new_n19055_, new_n2541_ );
and  ( new_n27206_, new_n27205_, new_n27204_ );
or   ( new_n27207_, new_n27206_, new_n18742_ );
and  ( new_n27208_, new_n19057_, RI2b1c4342de40_85 );
and  ( new_n27209_, new_n19044_, RI2b1c4342ddc8_84 );
or   ( new_n27210_, new_n27209_, new_n27208_ );
or   ( new_n27211_, new_n27210_, new_n18977_ );
and  ( new_n27212_, new_n27211_, new_n27207_ );
or   ( new_n27213_, new_n27212_, new_n27203_ );
and  ( new_n27214_, new_n27213_, new_n27202_ );
nor  ( new_n27215_, new_n22333_, new_n1004_ );
nor  ( new_n27216_, new_n27215_, new_n12071_ );
or   ( new_n27217_, new_n27216_, new_n21261_ );
and  ( new_n27218_, new_n22337_, RI2b1c4342da80_77 );
and  ( new_n27219_, new_n22330_, RI2b1c4342da08_76 );
or   ( new_n27220_, new_n27219_, new_n27218_ );
or   ( new_n27221_, new_n27220_, new_n21009_ );
and  ( new_n27222_, new_n27221_, new_n27217_ );
and  ( new_n27223_, new_n27222_, new_n16071_ );
or   ( new_n27224_, new_n27222_, new_n16071_ );
or   ( new_n27225_, new_n21419_, new_n1310_ );
or   ( new_n27226_, new_n21424_, new_n1002_ );
and  ( new_n27227_, new_n27226_, new_n27225_ );
or   ( new_n27228_, new_n27227_, new_n21013_ );
and  ( new_n27229_, new_n21428_, RI2b1c4342db70_79 );
and  ( new_n27230_, new_n21415_, RI2b1c4342daf8_78 );
or   ( new_n27231_, new_n27230_, new_n27229_ );
or   ( new_n27232_, new_n27231_, new_n21265_ );
and  ( new_n27233_, new_n27232_, new_n27228_ );
and  ( new_n27234_, new_n27233_, new_n27224_ );
or   ( new_n27235_, new_n27234_, new_n27223_ );
and  ( new_n27236_, new_n27235_, new_n27214_ );
or   ( new_n27237_, new_n27235_, new_n27214_ );
or   ( new_n27238_, new_n18388_, new_n3924_ );
or   ( new_n27239_, new_n18395_, new_n3239_ );
and  ( new_n27240_, new_n27239_, new_n27238_ );
or   ( new_n27241_, new_n27240_, new_n18066_ );
and  ( new_n27242_, new_n18397_, RI2b1c4342df30_87 );
and  ( new_n27243_, new_n18384_, RI2b1c4342deb8_86 );
or   ( new_n27244_, new_n27243_, new_n27242_ );
or   ( new_n27245_, new_n27244_, new_n18309_ );
and  ( new_n27246_, new_n27245_, new_n27241_ );
or   ( new_n27247_, new_n17727_, new_n132_ );
or   ( new_n27248_, new_n17734_, new_n3902_ );
and  ( new_n27249_, new_n27248_, new_n27247_ );
or   ( new_n27250_, new_n27249_, new_n17238_ );
and  ( new_n27251_, new_n17736_, RI2b1c4342e020_89 );
and  ( new_n27252_, new_n17723_, RI2b1c4342dfa8_88 );
or   ( new_n27253_, new_n27252_, new_n27251_ );
or   ( new_n27254_, new_n27253_, new_n17650_ );
and  ( new_n27255_, new_n27254_, new_n27250_ );
or   ( new_n27256_, new_n27255_, new_n27246_ );
and  ( new_n27257_, new_n27255_, new_n27246_ );
or   ( new_n27258_, new_n17244_, new_n117_ );
or   ( new_n27259_, new_n17248_, new_n4635_ );
and  ( new_n27260_, new_n27259_, new_n27258_ );
or   ( new_n27261_, new_n27260_, new_n16814_ );
and  ( new_n27262_, new_n17255_, RI2b1c4342e110_91 );
and  ( new_n27263_, new_n17240_, RI2b1c4342e098_90 );
or   ( new_n27264_, new_n27263_, new_n27262_ );
or   ( new_n27265_, new_n27264_, new_n17142_ );
and  ( new_n27266_, new_n27265_, new_n27261_ );
or   ( new_n27267_, new_n27266_, new_n27257_ );
and  ( new_n27268_, new_n27267_, new_n27256_ );
and  ( new_n27269_, new_n27268_, new_n27237_ );
or   ( new_n27270_, new_n27269_, new_n27236_ );
and  ( new_n27271_, new_n27270_, new_n27183_ );
or   ( new_n27272_, new_n27270_, new_n27183_ );
or   ( new_n27273_, new_n27047_, new_n26896_ );
or   ( new_n27274_, new_n27044_, new_n26905_ );
and  ( new_n27275_, new_n27274_, new_n27273_ );
or   ( new_n27276_, new_n27275_, new_n27052_ );
and  ( new_n27277_, new_n27048_, new_n26906_ );
or   ( new_n27278_, new_n27277_, new_n26916_ );
and  ( new_n27279_, new_n27278_, new_n27276_ );
or   ( new_n27280_, new_n27032_, new_n26863_ );
or   ( new_n27281_, new_n27029_, new_n26872_ );
and  ( new_n27282_, new_n27281_, new_n27280_ );
or   ( new_n27283_, new_n27282_, new_n27037_ );
and  ( new_n27284_, new_n27033_, new_n26873_ );
or   ( new_n27285_, new_n27284_, new_n26883_ );
and  ( new_n27286_, new_n27285_, new_n27283_ );
or   ( new_n27287_, new_n27286_, new_n27279_ );
and  ( new_n27288_, new_n27286_, new_n27279_ );
or   ( new_n27289_, new_n27019_, new_n26832_ );
or   ( new_n27290_, new_n27016_, new_n26841_ );
and  ( new_n27291_, new_n27290_, new_n27289_ );
or   ( new_n27292_, new_n27291_, new_n27024_ );
and  ( new_n27293_, new_n27020_, new_n26842_ );
or   ( new_n27294_, new_n27293_, new_n26852_ );
and  ( new_n27295_, new_n27294_, new_n27292_ );
or   ( new_n27296_, new_n27295_, new_n27288_ );
and  ( new_n27297_, new_n27296_, new_n27287_ );
and  ( new_n27298_, new_n27297_, new_n27272_ );
or   ( new_n27299_, new_n27298_, new_n27271_ );
and  ( new_n27300_, new_n27299_, new_n27134_ );
or   ( new_n27301_, new_n27299_, new_n27134_ );
or   ( new_n27302_, new_n27085_, new_n26965_ );
or   ( new_n27303_, new_n27082_, new_n26972_ );
and  ( new_n27304_, new_n27303_, new_n27302_ );
or   ( new_n27305_, new_n27304_, new_n27090_ );
and  ( new_n27306_, new_n27086_, new_n26973_ );
or   ( new_n27307_, new_n27306_, new_n26981_ );
and  ( new_n27308_, new_n27307_, new_n27305_ );
and  ( new_n27309_, new_n27308_, new_n27301_ );
or   ( new_n27310_, new_n27309_, new_n27300_ );
and  ( new_n27311_, new_n27310_, new_n27113_ );
or   ( new_n27312_, new_n27310_, new_n27113_ );
or   ( new_n27313_, new_n27092_, new_n26962_ );
or   ( new_n27314_, new_n27080_, new_n26983_ );
and  ( new_n27315_, new_n27314_, new_n27313_ );
or   ( new_n27316_, new_n27315_, new_n27097_ );
and  ( new_n27317_, new_n27093_, new_n26984_ );
or   ( new_n27318_, new_n27317_, new_n26992_ );
and  ( new_n27319_, new_n27318_, new_n27316_ );
and  ( new_n27320_, new_n27319_, new_n27312_ );
or   ( new_n27321_, new_n27320_, new_n27311_ );
or   ( new_n27322_, new_n27321_, new_n27106_ );
or   ( new_n27323_, new_n27322_, new_n27007_ );
and  ( new_n27324_, new_n27323_, new_n27006_ );
or   ( new_n27325_, new_n27324_, new_n26812_ );
and  ( new_n27326_, new_n27325_, new_n26810_ );
and  ( new_n27327_, new_n27321_, new_n27106_ );
or   ( new_n27328_, new_n27327_, new_n27007_ );
or   ( new_n27329_, new_n27328_, new_n26812_ );
or   ( new_n27330_, new_n27317_, new_n27097_ );
or   ( new_n27331_, new_n27315_, new_n26992_ );
and  ( new_n27332_, new_n27331_, new_n27330_ );
or   ( new_n27333_, new_n27111_, new_n26781_ );
or   ( new_n27334_, new_n27109_, new_n26635_ );
and  ( new_n27335_, new_n27334_, new_n27333_ );
or   ( new_n27336_, new_n27335_, new_n27310_ );
or   ( new_n27337_, new_n27077_, new_n27074_ );
and  ( new_n27338_, new_n27337_, new_n26960_ );
or   ( new_n27339_, new_n27121_, new_n27067_ );
or   ( new_n27340_, new_n27119_, new_n26941_ );
and  ( new_n27341_, new_n27340_, new_n27339_ );
or   ( new_n27342_, new_n27341_, new_n27338_ );
and  ( new_n27343_, new_n27341_, new_n27338_ );
or   ( new_n27344_, new_n27130_, new_n27054_ );
or   ( new_n27345_, new_n27128_, new_n26918_ );
and  ( new_n27346_, new_n27345_, new_n27344_ );
or   ( new_n27347_, new_n27346_, new_n27343_ );
and  ( new_n27348_, new_n27347_, new_n27342_ );
or   ( new_n27349_, new_n27141_, new_n16085_ );
or   ( new_n27350_, new_n27137_, new_n16048_ );
and  ( new_n27351_, new_n27350_, new_n27349_ );
or   ( new_n27352_, new_n27150_, new_n16505_ );
or   ( new_n27353_, new_n27146_, new_n16438_ );
and  ( new_n27354_, new_n27353_, new_n27352_ );
or   ( new_n27355_, new_n27159_, new_n16085_ );
or   ( new_n27356_, new_n27155_, new_n16048_ );
and  ( new_n27357_, new_n27356_, new_n27355_ );
or   ( new_n27358_, new_n27357_, new_n27354_ );
and  ( new_n27359_, new_n27357_, new_n27354_ );
or   ( new_n27360_, new_n27166_, new_n16052_ );
or   ( new_n27361_, new_n27164_, new_n16071_ );
and  ( new_n27362_, new_n27361_, new_n27360_ );
or   ( new_n27363_, new_n27362_, new_n27359_ );
and  ( new_n27364_, new_n27363_, new_n27358_ );
or   ( new_n27365_, new_n27364_, new_n27351_ );
and  ( new_n27366_, new_n27364_, new_n27351_ );
or   ( new_n27367_, new_n27179_, new_n16052_ );
or   ( new_n27368_, new_n27175_, new_n16071_ );
and  ( new_n27369_, new_n27368_, new_n27367_ );
or   ( new_n27370_, new_n27369_, new_n27366_ );
and  ( new_n27371_, new_n27370_, new_n27365_ );
or   ( new_n27372_, new_n27190_, new_n20156_ );
or   ( new_n27373_, new_n27186_, new_n20443_ );
and  ( new_n27374_, new_n27373_, new_n27372_ );
or   ( new_n27375_, new_n27199_, new_n19394_ );
or   ( new_n27376_, new_n27195_, new_n19659_ );
and  ( new_n27377_, new_n27376_, new_n27375_ );
or   ( new_n27378_, new_n27377_, new_n27374_ );
and  ( new_n27379_, new_n27377_, new_n27374_ );
or   ( new_n27380_, new_n27210_, new_n18742_ );
or   ( new_n27381_, new_n27206_, new_n18977_ );
and  ( new_n27382_, new_n27381_, new_n27380_ );
or   ( new_n27383_, new_n27382_, new_n27379_ );
and  ( new_n27384_, new_n27383_, new_n27378_ );
or   ( new_n27385_, new_n27220_, new_n21261_ );
or   ( new_n27386_, new_n27216_, new_n21009_ );
and  ( new_n27387_, new_n27386_, new_n27385_ );
or   ( new_n27388_, new_n27387_, new_n16052_ );
and  ( new_n27389_, new_n27387_, new_n16052_ );
or   ( new_n27390_, new_n27231_, new_n21013_ );
or   ( new_n27391_, new_n27227_, new_n21265_ );
and  ( new_n27392_, new_n27391_, new_n27390_ );
or   ( new_n27393_, new_n27392_, new_n27389_ );
and  ( new_n27394_, new_n27393_, new_n27388_ );
or   ( new_n27395_, new_n27394_, new_n27384_ );
and  ( new_n27396_, new_n27394_, new_n27384_ );
or   ( new_n27397_, new_n27244_, new_n18066_ );
or   ( new_n27398_, new_n27240_, new_n18309_ );
and  ( new_n27399_, new_n27398_, new_n27397_ );
or   ( new_n27400_, new_n27253_, new_n17238_ );
or   ( new_n27401_, new_n27249_, new_n17650_ );
and  ( new_n27402_, new_n27401_, new_n27400_ );
or   ( new_n27403_, new_n27402_, new_n27399_ );
and  ( new_n27404_, new_n27402_, new_n27399_ );
or   ( new_n27405_, new_n27264_, new_n16814_ );
or   ( new_n27406_, new_n27260_, new_n17142_ );
and  ( new_n27407_, new_n27406_, new_n27405_ );
or   ( new_n27408_, new_n27407_, new_n27404_ );
and  ( new_n27409_, new_n27408_, new_n27403_ );
or   ( new_n27410_, new_n27409_, new_n27396_ );
and  ( new_n27411_, new_n27410_, new_n27395_ );
or   ( new_n27412_, new_n27411_, new_n27371_ );
and  ( new_n27413_, new_n27411_, new_n27371_ );
or   ( new_n27414_, new_n27277_, new_n27052_ );
or   ( new_n27415_, new_n27275_, new_n26916_ );
and  ( new_n27416_, new_n27415_, new_n27414_ );
or   ( new_n27417_, new_n27284_, new_n27037_ );
or   ( new_n27418_, new_n27282_, new_n26883_ );
and  ( new_n27419_, new_n27418_, new_n27417_ );
or   ( new_n27420_, new_n27419_, new_n27416_ );
and  ( new_n27421_, new_n27419_, new_n27416_ );
or   ( new_n27422_, new_n27293_, new_n27024_ );
or   ( new_n27423_, new_n27291_, new_n26852_ );
and  ( new_n27424_, new_n27423_, new_n27422_ );
or   ( new_n27425_, new_n27424_, new_n27421_ );
and  ( new_n27426_, new_n27425_, new_n27420_ );
or   ( new_n27427_, new_n27426_, new_n27413_ );
and  ( new_n27428_, new_n27427_, new_n27412_ );
or   ( new_n27429_, new_n27428_, new_n27348_ );
and  ( new_n27430_, new_n27428_, new_n27348_ );
or   ( new_n27431_, new_n27306_, new_n27090_ );
or   ( new_n27432_, new_n27304_, new_n26981_ );
and  ( new_n27433_, new_n27432_, new_n27431_ );
or   ( new_n27434_, new_n27433_, new_n27430_ );
and  ( new_n27435_, new_n27434_, new_n27429_ );
or   ( new_n27436_, new_n27435_, new_n27113_ );
and  ( new_n27437_, new_n27436_, new_n27336_ );
or   ( new_n27438_, new_n27437_, new_n27332_ );
or   ( new_n27439_, new_n27435_, new_n27335_ );
and  ( new_n27440_, new_n27439_, new_n27312_ );
or   ( new_n27441_, new_n27440_, new_n27319_ );
and  ( new_n27442_, new_n27441_, new_n27438_ );
or   ( new_n27443_, new_n27069_, new_n26920_ );
or   ( new_n27444_, new_n27056_, new_n26943_ );
and  ( new_n27445_, new_n27444_, new_n27443_ );
or   ( new_n27446_, new_n27445_, new_n27078_ );
and  ( new_n27447_, new_n27070_, new_n26944_ );
or   ( new_n27448_, new_n27447_, new_n26960_ );
and  ( new_n27449_, new_n27448_, new_n27446_ );
or   ( new_n27450_, new_n27341_, new_n27116_ );
or   ( new_n27451_, new_n27338_, new_n27123_ );
and  ( new_n27452_, new_n27451_, new_n27450_ );
or   ( new_n27453_, new_n27452_, new_n27346_ );
and  ( new_n27454_, new_n27342_, new_n27124_ );
or   ( new_n27455_, new_n27454_, new_n27132_ );
and  ( new_n27456_, new_n27455_, new_n27453_ );
nor  ( new_n27457_, new_n22333_, new_n1002_ );
nor  ( new_n27458_, new_n27457_, new_n12315_ );
or   ( new_n27459_, new_n27458_, new_n21261_ );
and  ( new_n27460_, new_n22337_, RI2b1c4342daf8_78 );
and  ( new_n27461_, new_n22330_, RI2b1c4342da80_77 );
or   ( new_n27462_, new_n27461_, new_n27460_ );
or   ( new_n27463_, new_n27462_, new_n21009_ );
and  ( new_n27464_, new_n27463_, new_n27459_ );
or   ( new_n27465_, new_n21419_, new_n1511_ );
or   ( new_n27466_, new_n21424_, new_n1310_ );
and  ( new_n27467_, new_n27466_, new_n27465_ );
or   ( new_n27468_, new_n27467_, new_n21013_ );
and  ( new_n27469_, new_n21428_, RI2b1c4342dbe8_80 );
and  ( new_n27470_, new_n21415_, RI2b1c4342db70_79 );
or   ( new_n27471_, new_n27470_, new_n27469_ );
or   ( new_n27472_, new_n27471_, new_n21265_ );
and  ( new_n27473_, new_n27472_, new_n27468_ );
or   ( new_n27474_, new_n27473_, new_n27464_ );
and  ( new_n27475_, new_n27473_, new_n27464_ );
or   ( new_n27476_, new_n20557_, new_n2119_ );
or   ( new_n27477_, new_n20562_, new_n126_ );
and  ( new_n27478_, new_n27477_, new_n27476_ );
or   ( new_n27479_, new_n27478_, new_n20156_ );
and  ( new_n27480_, new_n20566_, RI2b1c4342dcd8_82 );
and  ( new_n27481_, new_n20553_, RI2b1c4342dc60_81 );
or   ( new_n27482_, new_n27481_, new_n27480_ );
or   ( new_n27483_, new_n27482_, new_n20443_ );
and  ( new_n27484_, new_n27483_, new_n27479_ );
or   ( new_n27485_, new_n27484_, new_n27475_ );
and  ( new_n27486_, new_n27485_, new_n27474_ );
or   ( new_n27487_, new_n19758_, new_n2541_ );
or   ( new_n27488_, new_n19763_, new_n121_ );
and  ( new_n27489_, new_n27488_, new_n27487_ );
or   ( new_n27490_, new_n27489_, new_n19394_ );
and  ( new_n27491_, new_n19767_, RI2b1c4342ddc8_84 );
and  ( new_n27492_, new_n19754_, RI2b1c4342dd50_83 );
or   ( new_n27493_, new_n27492_, new_n27491_ );
or   ( new_n27494_, new_n27493_, new_n19659_ );
and  ( new_n27495_, new_n27494_, new_n27490_ );
or   ( new_n27496_, new_n19048_, new_n3239_ );
or   ( new_n27497_, new_n19055_, new_n2806_ );
and  ( new_n27498_, new_n27497_, new_n27496_ );
or   ( new_n27499_, new_n27498_, new_n18742_ );
and  ( new_n27500_, new_n19057_, RI2b1c4342deb8_86 );
and  ( new_n27501_, new_n19044_, RI2b1c4342de40_85 );
or   ( new_n27502_, new_n27501_, new_n27500_ );
or   ( new_n27503_, new_n27502_, new_n18977_ );
and  ( new_n27504_, new_n27503_, new_n27499_ );
or   ( new_n27505_, new_n27504_, new_n27495_ );
and  ( new_n27506_, new_n27504_, new_n27495_ );
or   ( new_n27507_, new_n18388_, new_n3902_ );
or   ( new_n27508_, new_n18395_, new_n3924_ );
and  ( new_n27509_, new_n27508_, new_n27507_ );
or   ( new_n27510_, new_n27509_, new_n18066_ );
and  ( new_n27511_, new_n18397_, RI2b1c4342dfa8_88 );
and  ( new_n27512_, new_n18384_, RI2b1c4342df30_87 );
or   ( new_n27513_, new_n27512_, new_n27511_ );
or   ( new_n27514_, new_n27513_, new_n18309_ );
and  ( new_n27515_, new_n27514_, new_n27510_ );
or   ( new_n27516_, new_n27515_, new_n27506_ );
and  ( new_n27517_, new_n27516_, new_n27505_ );
or   ( new_n27518_, new_n27517_, new_n27486_ );
and  ( new_n27519_, new_n27517_, new_n27486_ );
or   ( new_n27520_, new_n17727_, new_n4635_ );
or   ( new_n27521_, new_n17734_, new_n132_ );
and  ( new_n27522_, new_n27521_, new_n27520_ );
or   ( new_n27523_, new_n27522_, new_n17238_ );
and  ( new_n27524_, new_n17736_, RI2b1c4342e098_90 );
and  ( new_n27525_, new_n17723_, RI2b1c4342e020_89 );
or   ( new_n27526_, new_n27525_, new_n27524_ );
or   ( new_n27527_, new_n27526_, new_n17650_ );
and  ( new_n27528_, new_n27527_, new_n27523_ );
or   ( new_n27529_, new_n17244_, new_n5459_ );
or   ( new_n27530_, new_n17248_, new_n117_ );
and  ( new_n27531_, new_n27530_, new_n27529_ );
or   ( new_n27532_, new_n27531_, new_n16814_ );
and  ( new_n27533_, new_n17255_, RI2b1c4342e188_92 );
and  ( new_n27534_, new_n17240_, RI2b1c4342e110_91 );
or   ( new_n27535_, new_n27534_, new_n27533_ );
or   ( new_n27536_, new_n27535_, new_n17142_ );
and  ( new_n27537_, new_n27536_, new_n27532_ );
or   ( new_n27538_, new_n27537_, new_n27528_ );
and  ( new_n27539_, new_n27537_, new_n27528_ );
or   ( new_n27540_, new_n16607_, new_n6321_ );
or   ( new_n27541_, new_n16613_, new_n6307_ );
and  ( new_n27542_, new_n27541_, new_n27540_ );
or   ( new_n27543_, new_n27542_, new_n16505_ );
and  ( new_n27544_, new_n16616_, RI2b1c4342e278_94 );
and  ( new_n27545_, new_n16603_, RI2b1c4342e200_93 );
or   ( new_n27546_, new_n27545_, new_n27544_ );
or   ( new_n27547_, new_n27546_, new_n16438_ );
and  ( new_n27548_, new_n27547_, new_n27543_ );
or   ( new_n27549_, new_n27548_, new_n27539_ );
and  ( new_n27550_, new_n27549_, new_n27538_ );
or   ( new_n27551_, new_n27550_, new_n27519_ );
and  ( new_n27552_, new_n27551_, new_n27518_ );
or   ( new_n27553_, new_n27357_, new_n27152_ );
or   ( new_n27554_, new_n27354_, new_n27161_ );
and  ( new_n27555_, new_n27554_, new_n27553_ );
or   ( new_n27556_, new_n27555_, new_n27362_ );
and  ( new_n27557_, new_n27358_, new_n27162_ );
or   ( new_n27558_, new_n27557_, new_n27168_ );
and  ( new_n27559_, new_n27558_, new_n27556_ );
or   ( new_n27560_, new_n27402_, new_n27246_ );
or   ( new_n27561_, new_n27399_, new_n27255_ );
and  ( new_n27562_, new_n27561_, new_n27560_ );
or   ( new_n27563_, new_n27562_, new_n27407_ );
and  ( new_n27564_, new_n27403_, new_n27256_ );
or   ( new_n27565_, new_n27564_, new_n27266_ );
and  ( new_n27566_, new_n27565_, new_n27563_ );
or   ( new_n27567_, new_n27566_, new_n27559_ );
and  ( new_n27568_, new_n27566_, new_n27559_ );
or   ( new_n27569_, new_n27377_, new_n27192_ );
or   ( new_n27570_, new_n27374_, new_n27201_ );
and  ( new_n27571_, new_n27570_, new_n27569_ );
or   ( new_n27572_, new_n27571_, new_n27382_ );
and  ( new_n27573_, new_n27378_, new_n27202_ );
or   ( new_n27574_, new_n27573_, new_n27212_ );
and  ( new_n27575_, new_n27574_, new_n27572_ );
or   ( new_n27576_, new_n27575_, new_n27568_ );
and  ( new_n27577_, new_n27576_, new_n27567_ );
or   ( new_n27578_, new_n27577_, new_n27552_ );
and  ( new_n27579_, new_n27577_, new_n27552_ );
or   ( new_n27580_, new_n27419_, new_n27279_ );
or   ( new_n27581_, new_n27416_, new_n27286_ );
and  ( new_n27582_, new_n27581_, new_n27580_ );
or   ( new_n27583_, new_n27582_, new_n27424_ );
and  ( new_n27584_, new_n27420_, new_n27287_ );
or   ( new_n27585_, new_n27584_, new_n27295_ );
and  ( new_n27586_, new_n27585_, new_n27583_ );
or   ( new_n27587_, new_n27586_, new_n27579_ );
and  ( new_n27588_, new_n27587_, new_n27578_ );
or   ( new_n27589_, new_n27588_, new_n27456_ );
and  ( new_n27590_, new_n27588_, new_n27456_ );
or   ( new_n27591_, new_n27371_, new_n27270_ );
or   ( new_n27592_, new_n27411_, new_n27183_ );
and  ( new_n27593_, new_n27592_, new_n27591_ );
or   ( new_n27594_, new_n27593_, new_n27426_ );
and  ( new_n27595_, new_n27412_, new_n27272_ );
or   ( new_n27596_, new_n27595_, new_n27297_ );
and  ( new_n27597_, new_n27596_, new_n27594_ );
or   ( new_n27598_, new_n27597_, new_n27590_ );
and  ( new_n27599_, new_n27598_, new_n27589_ );
or   ( new_n27600_, new_n27599_, new_n27449_ );
or   ( new_n27601_, new_n27348_, new_n27299_ );
or   ( new_n27602_, new_n27428_, new_n27134_ );
and  ( new_n27603_, new_n27602_, new_n27601_ );
or   ( new_n27604_, new_n27603_, new_n27433_ );
and  ( new_n27605_, new_n27429_, new_n27301_ );
or   ( new_n27606_, new_n27605_, new_n27308_ );
and  ( new_n27607_, new_n27606_, new_n27604_ );
and  ( new_n27608_, new_n27599_, new_n27449_ );
or   ( new_n27609_, new_n27608_, new_n27607_ );
and  ( new_n27610_, new_n27609_, new_n27600_ );
and  ( new_n27611_, new_n27610_, new_n27442_ );
or   ( new_n27612_, new_n27605_, new_n27433_ );
or   ( new_n27613_, new_n27603_, new_n27308_ );
and  ( new_n27614_, new_n27613_, new_n27612_ );
or   ( new_n27615_, new_n27447_, new_n27078_ );
or   ( new_n27616_, new_n27445_, new_n26960_ );
and  ( new_n27617_, new_n27616_, new_n27615_ );
or   ( new_n27618_, new_n27617_, new_n27599_ );
or   ( new_n27619_, new_n27454_, new_n27346_ );
or   ( new_n27620_, new_n27452_, new_n27132_ );
and  ( new_n27621_, new_n27620_, new_n27619_ );
or   ( new_n27622_, new_n27462_, new_n21261_ );
or   ( new_n27623_, new_n27458_, new_n21009_ );
and  ( new_n27624_, new_n27623_, new_n27622_ );
or   ( new_n27625_, new_n27471_, new_n21013_ );
or   ( new_n27626_, new_n27467_, new_n21265_ );
and  ( new_n27627_, new_n27626_, new_n27625_ );
or   ( new_n27628_, new_n27627_, new_n27624_ );
and  ( new_n27629_, new_n27627_, new_n27624_ );
or   ( new_n27630_, new_n27482_, new_n20156_ );
or   ( new_n27631_, new_n27478_, new_n20443_ );
and  ( new_n27632_, new_n27631_, new_n27630_ );
or   ( new_n27633_, new_n27632_, new_n27629_ );
and  ( new_n27634_, new_n27633_, new_n27628_ );
or   ( new_n27635_, new_n27493_, new_n19394_ );
or   ( new_n27636_, new_n27489_, new_n19659_ );
and  ( new_n27637_, new_n27636_, new_n27635_ );
or   ( new_n27638_, new_n27502_, new_n18742_ );
or   ( new_n27639_, new_n27498_, new_n18977_ );
and  ( new_n27640_, new_n27639_, new_n27638_ );
or   ( new_n27641_, new_n27640_, new_n27637_ );
and  ( new_n27642_, new_n27640_, new_n27637_ );
or   ( new_n27643_, new_n27513_, new_n18066_ );
or   ( new_n27644_, new_n27509_, new_n18309_ );
and  ( new_n27645_, new_n27644_, new_n27643_ );
or   ( new_n27646_, new_n27645_, new_n27642_ );
and  ( new_n27647_, new_n27646_, new_n27641_ );
or   ( new_n27648_, new_n27647_, new_n27634_ );
and  ( new_n27649_, new_n27647_, new_n27634_ );
or   ( new_n27650_, new_n27526_, new_n17238_ );
or   ( new_n27651_, new_n27522_, new_n17650_ );
and  ( new_n27652_, new_n27651_, new_n27650_ );
or   ( new_n27653_, new_n27535_, new_n16814_ );
or   ( new_n27654_, new_n27531_, new_n17142_ );
and  ( new_n27655_, new_n27654_, new_n27653_ );
or   ( new_n27656_, new_n27655_, new_n27652_ );
and  ( new_n27657_, new_n27655_, new_n27652_ );
or   ( new_n27658_, new_n27546_, new_n16505_ );
or   ( new_n27659_, new_n27542_, new_n16438_ );
and  ( new_n27660_, new_n27659_, new_n27658_ );
or   ( new_n27661_, new_n27660_, new_n27657_ );
and  ( new_n27662_, new_n27661_, new_n27656_ );
or   ( new_n27663_, new_n27662_, new_n27649_ );
and  ( new_n27664_, new_n27663_, new_n27648_ );
or   ( new_n27665_, new_n27557_, new_n27362_ );
or   ( new_n27666_, new_n27555_, new_n27168_ );
and  ( new_n27667_, new_n27666_, new_n27665_ );
or   ( new_n27668_, new_n27564_, new_n27407_ );
or   ( new_n27669_, new_n27562_, new_n27266_ );
and  ( new_n27670_, new_n27669_, new_n27668_ );
or   ( new_n27671_, new_n27670_, new_n27667_ );
and  ( new_n27672_, new_n27670_, new_n27667_ );
or   ( new_n27673_, new_n27573_, new_n27382_ );
or   ( new_n27674_, new_n27571_, new_n27212_ );
and  ( new_n27675_, new_n27674_, new_n27673_ );
or   ( new_n27676_, new_n27675_, new_n27672_ );
and  ( new_n27677_, new_n27676_, new_n27671_ );
or   ( new_n27678_, new_n27677_, new_n27664_ );
and  ( new_n27679_, new_n27677_, new_n27664_ );
or   ( new_n27680_, new_n27584_, new_n27424_ );
or   ( new_n27681_, new_n27582_, new_n27295_ );
and  ( new_n27682_, new_n27681_, new_n27680_ );
or   ( new_n27683_, new_n27682_, new_n27679_ );
and  ( new_n27684_, new_n27683_, new_n27678_ );
or   ( new_n27685_, new_n27684_, new_n27621_ );
and  ( new_n27686_, new_n27684_, new_n27621_ );
or   ( new_n27687_, new_n27595_, new_n27426_ );
or   ( new_n27688_, new_n27593_, new_n27297_ );
and  ( new_n27689_, new_n27688_, new_n27687_ );
or   ( new_n27690_, new_n27689_, new_n27686_ );
and  ( new_n27691_, new_n27690_, new_n27685_ );
or   ( new_n27692_, new_n27691_, new_n27449_ );
and  ( new_n27693_, new_n27692_, new_n27618_ );
or   ( new_n27694_, new_n27693_, new_n27614_ );
or   ( new_n27695_, new_n27691_, new_n27617_ );
and  ( new_n27696_, new_n27695_, new_n27600_ );
or   ( new_n27697_, new_n27696_, new_n27607_ );
and  ( new_n27698_, new_n27697_, new_n27694_ );
or   ( new_n27699_, new_n27384_, new_n27235_ );
or   ( new_n27700_, new_n27394_, new_n27214_ );
and  ( new_n27701_, new_n27700_, new_n27699_ );
or   ( new_n27702_, new_n27701_, new_n27409_ );
and  ( new_n27703_, new_n27395_, new_n27237_ );
or   ( new_n27704_, new_n27703_, new_n27268_ );
and  ( new_n27705_, new_n27704_, new_n27702_ );
or   ( new_n27706_, new_n27677_, new_n27552_ );
or   ( new_n27707_, new_n27664_, new_n27577_ );
and  ( new_n27708_, new_n27707_, new_n27706_ );
or   ( new_n27709_, new_n27708_, new_n27682_ );
and  ( new_n27710_, new_n27678_, new_n27578_ );
or   ( new_n27711_, new_n27710_, new_n27586_ );
and  ( new_n27712_, new_n27711_, new_n27709_ );
or   ( new_n27713_, new_n27712_, new_n27705_ );
or   ( new_n27714_, new_n27670_, new_n27559_ );
or   ( new_n27715_, new_n27667_, new_n27566_ );
and  ( new_n27716_, new_n27715_, new_n27714_ );
or   ( new_n27717_, new_n27716_, new_n27675_ );
and  ( new_n27718_, new_n27671_, new_n27567_ );
or   ( new_n27719_, new_n27718_, new_n27575_ );
and  ( new_n27720_, new_n27719_, new_n27717_ );
or   ( new_n27721_, new_n27647_, new_n27486_ );
or   ( new_n27722_, new_n27634_, new_n27517_ );
and  ( new_n27723_, new_n27722_, new_n27721_ );
or   ( new_n27724_, new_n27723_, new_n27662_ );
and  ( new_n27725_, new_n27648_, new_n27518_ );
or   ( new_n27726_, new_n27725_, new_n27550_ );
and  ( new_n27727_, new_n27726_, new_n27724_ );
or   ( new_n27728_, new_n27727_, new_n27720_ );
or   ( new_n27729_, new_n16366_, new_n7274_ );
or   ( new_n27730_, new_n16355_, new_n124_ );
and  ( new_n27731_, new_n27730_, new_n27729_ );
or   ( new_n27732_, new_n27731_, new_n16085_ );
and  ( new_n27733_, new_n16358_, RI2b1c4342e368_96 );
and  ( new_n27734_, new_n16362_, RI2b1c4342e2f0_95 );
or   ( new_n27735_, new_n27734_, new_n27733_ );
or   ( new_n27736_, new_n27735_, new_n16048_ );
and  ( new_n27737_, new_n27736_, new_n27732_ );
or   ( new_n27738_, new_n27655_, new_n27528_ );
or   ( new_n27739_, new_n27652_, new_n27537_ );
and  ( new_n27740_, new_n27739_, new_n27738_ );
or   ( new_n27741_, new_n27740_, new_n27660_ );
and  ( new_n27742_, new_n27656_, new_n27538_ );
or   ( new_n27743_, new_n27742_, new_n27548_ );
and  ( new_n27744_, new_n27743_, new_n27741_ );
or   ( new_n27745_, new_n27744_, new_n27737_ );
and  ( new_n27746_, new_n27744_, new_n27737_ );
or   ( new_n27747_, new_n27640_, new_n27495_ );
or   ( new_n27748_, new_n27637_, new_n27504_ );
and  ( new_n27749_, new_n27748_, new_n27747_ );
or   ( new_n27750_, new_n27749_, new_n27645_ );
and  ( new_n27751_, new_n27641_, new_n27505_ );
or   ( new_n27752_, new_n27751_, new_n27515_ );
and  ( new_n27753_, new_n27752_, new_n27750_ );
or   ( new_n27754_, new_n27753_, new_n27746_ );
and  ( new_n27755_, new_n27754_, new_n27745_ );
or   ( new_n27756_, new_n20557_, new_n121_ );
or   ( new_n27757_, new_n20562_, new_n2119_ );
and  ( new_n27758_, new_n27757_, new_n27756_ );
or   ( new_n27759_, new_n27758_, new_n20156_ );
and  ( new_n27760_, new_n20566_, RI2b1c4342dd50_83 );
and  ( new_n27761_, new_n20553_, RI2b1c4342dcd8_82 );
or   ( new_n27762_, new_n27761_, new_n27760_ );
or   ( new_n27763_, new_n27762_, new_n20443_ );
and  ( new_n27764_, new_n27763_, new_n27759_ );
or   ( new_n27765_, new_n19758_, new_n2806_ );
or   ( new_n27766_, new_n19763_, new_n2541_ );
and  ( new_n27767_, new_n27766_, new_n27765_ );
or   ( new_n27768_, new_n27767_, new_n19394_ );
and  ( new_n27769_, new_n19767_, RI2b1c4342de40_85 );
and  ( new_n27770_, new_n19754_, RI2b1c4342ddc8_84 );
or   ( new_n27771_, new_n27770_, new_n27769_ );
or   ( new_n27772_, new_n27771_, new_n19659_ );
and  ( new_n27773_, new_n27772_, new_n27768_ );
or   ( new_n27774_, new_n27773_, new_n27764_ );
and  ( new_n27775_, new_n27773_, new_n27764_ );
or   ( new_n27776_, new_n19048_, new_n3924_ );
or   ( new_n27777_, new_n19055_, new_n3239_ );
and  ( new_n27778_, new_n27777_, new_n27776_ );
or   ( new_n27779_, new_n27778_, new_n18742_ );
and  ( new_n27780_, new_n19057_, RI2b1c4342df30_87 );
and  ( new_n27781_, new_n19044_, RI2b1c4342deb8_86 );
or   ( new_n27782_, new_n27781_, new_n27780_ );
or   ( new_n27783_, new_n27782_, new_n18977_ );
and  ( new_n27784_, new_n27783_, new_n27779_ );
or   ( new_n27785_, new_n27784_, new_n27775_ );
and  ( new_n27786_, new_n27785_, new_n27774_ );
nor  ( new_n27787_, new_n22333_, new_n1310_ );
nor  ( new_n27788_, new_n27787_, new_n12619_ );
or   ( new_n27789_, new_n27788_, new_n21261_ );
and  ( new_n27790_, new_n22337_, RI2b1c4342db70_79 );
and  ( new_n27791_, new_n22330_, RI2b1c4342daf8_78 );
or   ( new_n27792_, new_n27791_, new_n27790_ );
or   ( new_n27793_, new_n27792_, new_n21009_ );
and  ( new_n27794_, new_n27793_, new_n27789_ );
and  ( new_n27795_, new_n27794_, new_n16048_ );
or   ( new_n27796_, new_n27794_, new_n16048_ );
or   ( new_n27797_, new_n21419_, new_n126_ );
or   ( new_n27798_, new_n21424_, new_n1511_ );
and  ( new_n27799_, new_n27798_, new_n27797_ );
or   ( new_n27800_, new_n27799_, new_n21013_ );
and  ( new_n27801_, new_n21428_, RI2b1c4342dc60_81 );
and  ( new_n27802_, new_n21415_, RI2b1c4342dbe8_80 );
or   ( new_n27803_, new_n27802_, new_n27801_ );
or   ( new_n27804_, new_n27803_, new_n21265_ );
and  ( new_n27805_, new_n27804_, new_n27800_ );
and  ( new_n27806_, new_n27805_, new_n27796_ );
or   ( new_n27807_, new_n27806_, new_n27795_ );
and  ( new_n27808_, new_n27807_, new_n27786_ );
or   ( new_n27809_, new_n27807_, new_n27786_ );
or   ( new_n27810_, new_n18388_, new_n132_ );
or   ( new_n27811_, new_n18395_, new_n3902_ );
and  ( new_n27812_, new_n27811_, new_n27810_ );
or   ( new_n27813_, new_n27812_, new_n18066_ );
and  ( new_n27814_, new_n18397_, RI2b1c4342e020_89 );
and  ( new_n27815_, new_n18384_, RI2b1c4342dfa8_88 );
or   ( new_n27816_, new_n27815_, new_n27814_ );
or   ( new_n27817_, new_n27816_, new_n18309_ );
and  ( new_n27818_, new_n27817_, new_n27813_ );
or   ( new_n27819_, new_n17727_, new_n117_ );
or   ( new_n27820_, new_n17734_, new_n4635_ );
and  ( new_n27821_, new_n27820_, new_n27819_ );
or   ( new_n27822_, new_n27821_, new_n17238_ );
and  ( new_n27823_, new_n17736_, RI2b1c4342e110_91 );
and  ( new_n27824_, new_n17723_, RI2b1c4342e098_90 );
or   ( new_n27825_, new_n27824_, new_n27823_ );
or   ( new_n27826_, new_n27825_, new_n17650_ );
and  ( new_n27827_, new_n27826_, new_n27822_ );
or   ( new_n27828_, new_n27827_, new_n27818_ );
and  ( new_n27829_, new_n27827_, new_n27818_ );
or   ( new_n27830_, new_n17244_, new_n6307_ );
or   ( new_n27831_, new_n17248_, new_n5459_ );
and  ( new_n27832_, new_n27831_, new_n27830_ );
or   ( new_n27833_, new_n27832_, new_n16814_ );
and  ( new_n27834_, new_n17255_, RI2b1c4342e200_93 );
and  ( new_n27835_, new_n17240_, RI2b1c4342e188_92 );
or   ( new_n27836_, new_n27835_, new_n27834_ );
or   ( new_n27837_, new_n27836_, new_n17142_ );
and  ( new_n27838_, new_n27837_, new_n27833_ );
or   ( new_n27839_, new_n27838_, new_n27829_ );
and  ( new_n27840_, new_n27839_, new_n27828_ );
and  ( new_n27841_, new_n27840_, new_n27809_ );
or   ( new_n27842_, new_n27841_, new_n27808_ );
and  ( new_n27843_, new_n27842_, new_n27755_ );
or   ( new_n27844_, new_n27842_, new_n27755_ );
or   ( new_n27845_, new_n27387_, new_n16071_ );
or   ( new_n27846_, new_n27222_, new_n16052_ );
and  ( new_n27847_, new_n27846_, new_n27845_ );
or   ( new_n27848_, new_n27847_, new_n27392_ );
and  ( new_n27849_, new_n27388_, new_n27224_ );
or   ( new_n27850_, new_n27849_, new_n27233_ );
and  ( new_n27851_, new_n27850_, new_n27848_ );
and  ( new_n27852_, new_n27851_, new_n27844_ );
or   ( new_n27853_, new_n27852_, new_n27843_ );
and  ( new_n27854_, new_n27853_, new_n27728_ );
or   ( new_n27855_, new_n27853_, new_n27728_ );
or   ( new_n27856_, new_n27351_, new_n27170_ );
or   ( new_n27857_, new_n27364_, new_n27143_ );
and  ( new_n27858_, new_n27857_, new_n27856_ );
or   ( new_n27859_, new_n27858_, new_n27369_ );
and  ( new_n27860_, new_n27365_, new_n27171_ );
or   ( new_n27861_, new_n27860_, new_n27181_ );
and  ( new_n27862_, new_n27861_, new_n27859_ );
and  ( new_n27863_, new_n27862_, new_n27855_ );
or   ( new_n27864_, new_n27863_, new_n27854_ );
and  ( new_n27865_, new_n27864_, new_n27713_ );
or   ( new_n27866_, new_n27864_, new_n27713_ );
or   ( new_n27867_, new_n27621_, new_n27588_ );
or   ( new_n27868_, new_n27684_, new_n27456_ );
and  ( new_n27869_, new_n27868_, new_n27867_ );
or   ( new_n27870_, new_n27869_, new_n27689_ );
and  ( new_n27871_, new_n27685_, new_n27589_ );
or   ( new_n27872_, new_n27871_, new_n27597_ );
and  ( new_n27873_, new_n27872_, new_n27870_ );
and  ( new_n27874_, new_n27873_, new_n27866_ );
or   ( new_n27875_, new_n27874_, new_n27865_ );
and  ( new_n27876_, new_n27875_, new_n27698_ );
or   ( new_n27877_, new_n27876_, new_n27611_ );
or   ( new_n27878_, new_n27871_, new_n27689_ );
or   ( new_n27879_, new_n27869_, new_n27597_ );
and  ( new_n27880_, new_n27879_, new_n27878_ );
or   ( new_n27881_, new_n27703_, new_n27409_ );
or   ( new_n27882_, new_n27701_, new_n27268_ );
and  ( new_n27883_, new_n27882_, new_n27881_ );
or   ( new_n27884_, new_n27710_, new_n27682_ );
or   ( new_n27885_, new_n27708_, new_n27586_ );
and  ( new_n27886_, new_n27885_, new_n27884_ );
and  ( new_n27887_, new_n27886_, new_n27883_ );
or   ( new_n27888_, new_n27887_, new_n27864_ );
or   ( new_n27889_, new_n27718_, new_n27675_ );
or   ( new_n27890_, new_n27716_, new_n27575_ );
and  ( new_n27891_, new_n27890_, new_n27889_ );
or   ( new_n27892_, new_n27725_, new_n27662_ );
or   ( new_n27893_, new_n27723_, new_n27550_ );
and  ( new_n27894_, new_n27893_, new_n27892_ );
and  ( new_n27895_, new_n27894_, new_n27891_ );
or   ( new_n27896_, new_n27762_, new_n20156_ );
or   ( new_n27897_, new_n27758_, new_n20443_ );
and  ( new_n27898_, new_n27897_, new_n27896_ );
or   ( new_n27899_, new_n27771_, new_n19394_ );
or   ( new_n27900_, new_n27767_, new_n19659_ );
and  ( new_n27901_, new_n27900_, new_n27899_ );
or   ( new_n27902_, new_n27901_, new_n27898_ );
and  ( new_n27903_, new_n27901_, new_n27898_ );
or   ( new_n27904_, new_n27782_, new_n18742_ );
or   ( new_n27905_, new_n27778_, new_n18977_ );
and  ( new_n27906_, new_n27905_, new_n27904_ );
or   ( new_n27907_, new_n27906_, new_n27903_ );
and  ( new_n27908_, new_n27907_, new_n27902_ );
or   ( new_n27909_, new_n27792_, new_n21261_ );
or   ( new_n27910_, new_n27788_, new_n21009_ );
and  ( new_n27911_, new_n27910_, new_n27909_ );
or   ( new_n27912_, new_n27911_, new_n16085_ );
and  ( new_n27913_, new_n27911_, new_n16085_ );
or   ( new_n27914_, new_n27803_, new_n21013_ );
or   ( new_n27915_, new_n27799_, new_n21265_ );
and  ( new_n27916_, new_n27915_, new_n27914_ );
or   ( new_n27917_, new_n27916_, new_n27913_ );
and  ( new_n27918_, new_n27917_, new_n27912_ );
or   ( new_n27919_, new_n27918_, new_n27908_ );
and  ( new_n27920_, new_n27918_, new_n27908_ );
or   ( new_n27921_, new_n27816_, new_n18066_ );
or   ( new_n27922_, new_n27812_, new_n18309_ );
and  ( new_n27923_, new_n27922_, new_n27921_ );
or   ( new_n27924_, new_n27825_, new_n17238_ );
or   ( new_n27925_, new_n27821_, new_n17650_ );
and  ( new_n27926_, new_n27925_, new_n27924_ );
or   ( new_n27927_, new_n27926_, new_n27923_ );
and  ( new_n27928_, new_n27926_, new_n27923_ );
or   ( new_n27929_, new_n27836_, new_n16814_ );
or   ( new_n27930_, new_n27832_, new_n17142_ );
and  ( new_n27931_, new_n27930_, new_n27929_ );
or   ( new_n27932_, new_n27931_, new_n27928_ );
and  ( new_n27933_, new_n27932_, new_n27927_ );
or   ( new_n27934_, new_n27933_, new_n27920_ );
and  ( new_n27935_, new_n27934_, new_n27919_ );
or   ( new_n27936_, new_n27735_, new_n16085_ );
or   ( new_n27937_, new_n27731_, new_n16048_ );
and  ( new_n27938_, new_n27937_, new_n27936_ );
or   ( new_n27939_, new_n27742_, new_n27660_ );
or   ( new_n27940_, new_n27740_, new_n27548_ );
and  ( new_n27941_, new_n27940_, new_n27939_ );
or   ( new_n27942_, new_n27941_, new_n27938_ );
and  ( new_n27943_, new_n27941_, new_n27938_ );
or   ( new_n27944_, new_n27751_, new_n27645_ );
or   ( new_n27945_, new_n27749_, new_n27515_ );
and  ( new_n27946_, new_n27945_, new_n27944_ );
or   ( new_n27947_, new_n27946_, new_n27943_ );
and  ( new_n27948_, new_n27947_, new_n27942_ );
or   ( new_n27949_, new_n27948_, new_n27935_ );
and  ( new_n27950_, new_n27948_, new_n27935_ );
or   ( new_n27951_, new_n27849_, new_n27392_ );
or   ( new_n27952_, new_n27847_, new_n27233_ );
and  ( new_n27953_, new_n27952_, new_n27951_ );
or   ( new_n27954_, new_n27953_, new_n27950_ );
and  ( new_n27955_, new_n27954_, new_n27949_ );
or   ( new_n27956_, new_n27955_, new_n27895_ );
and  ( new_n27957_, new_n27955_, new_n27895_ );
or   ( new_n27958_, new_n27860_, new_n27369_ );
or   ( new_n27959_, new_n27858_, new_n27181_ );
and  ( new_n27960_, new_n27959_, new_n27958_ );
or   ( new_n27961_, new_n27960_, new_n27957_ );
and  ( new_n27962_, new_n27961_, new_n27956_ );
or   ( new_n27963_, new_n27962_, new_n27713_ );
and  ( new_n27964_, new_n27963_, new_n27888_ );
or   ( new_n27965_, new_n27964_, new_n27880_ );
or   ( new_n27966_, new_n27962_, new_n27887_ );
and  ( new_n27967_, new_n27966_, new_n27866_ );
or   ( new_n27968_, new_n27967_, new_n27873_ );
and  ( new_n27969_, new_n27968_, new_n27965_ );
or   ( new_n27970_, new_n27886_, new_n27705_ );
or   ( new_n27971_, new_n27883_, new_n27712_ );
and  ( new_n27972_, new_n27971_, new_n27970_ );
or   ( new_n27973_, new_n27894_, new_n27720_ );
or   ( new_n27974_, new_n27891_, new_n27727_ );
and  ( new_n27975_, new_n27974_, new_n27973_ );
nor  ( new_n27976_, new_n22333_, new_n1511_ );
nor  ( new_n27977_, new_n27976_, new_n12834_ );
or   ( new_n27978_, new_n27977_, new_n21261_ );
and  ( new_n27979_, new_n22337_, RI2b1c4342dbe8_80 );
and  ( new_n27980_, new_n22330_, RI2b1c4342db70_79 );
or   ( new_n27981_, new_n27980_, new_n27979_ );
or   ( new_n27982_, new_n27981_, new_n21009_ );
and  ( new_n27983_, new_n27982_, new_n27978_ );
or   ( new_n27984_, new_n21419_, new_n2119_ );
or   ( new_n27985_, new_n21424_, new_n126_ );
and  ( new_n27986_, new_n27985_, new_n27984_ );
or   ( new_n27987_, new_n27986_, new_n21013_ );
and  ( new_n27988_, new_n21428_, RI2b1c4342dcd8_82 );
and  ( new_n27989_, new_n21415_, RI2b1c4342dc60_81 );
or   ( new_n27990_, new_n27989_, new_n27988_ );
or   ( new_n27991_, new_n27990_, new_n21265_ );
and  ( new_n27992_, new_n27991_, new_n27987_ );
or   ( new_n27993_, new_n27992_, new_n27983_ );
and  ( new_n27994_, new_n27992_, new_n27983_ );
or   ( new_n27995_, new_n20557_, new_n2541_ );
or   ( new_n27996_, new_n20562_, new_n121_ );
and  ( new_n27997_, new_n27996_, new_n27995_ );
or   ( new_n27998_, new_n27997_, new_n20156_ );
and  ( new_n27999_, new_n20566_, RI2b1c4342ddc8_84 );
and  ( new_n28000_, new_n20553_, RI2b1c4342dd50_83 );
or   ( new_n28001_, new_n28000_, new_n27999_ );
or   ( new_n28002_, new_n28001_, new_n20443_ );
and  ( new_n28003_, new_n28002_, new_n27998_ );
or   ( new_n28004_, new_n28003_, new_n27994_ );
and  ( new_n28005_, new_n28004_, new_n27993_ );
or   ( new_n28006_, new_n19758_, new_n3239_ );
or   ( new_n28007_, new_n19763_, new_n2806_ );
and  ( new_n28008_, new_n28007_, new_n28006_ );
or   ( new_n28009_, new_n28008_, new_n19394_ );
and  ( new_n28010_, new_n19767_, RI2b1c4342deb8_86 );
and  ( new_n28011_, new_n19754_, RI2b1c4342de40_85 );
or   ( new_n28012_, new_n28011_, new_n28010_ );
or   ( new_n28013_, new_n28012_, new_n19659_ );
and  ( new_n28014_, new_n28013_, new_n28009_ );
or   ( new_n28015_, new_n19048_, new_n3902_ );
or   ( new_n28016_, new_n19055_, new_n3924_ );
and  ( new_n28017_, new_n28016_, new_n28015_ );
or   ( new_n28018_, new_n28017_, new_n18742_ );
and  ( new_n28019_, new_n19057_, RI2b1c4342dfa8_88 );
and  ( new_n28020_, new_n19044_, RI2b1c4342df30_87 );
or   ( new_n28021_, new_n28020_, new_n28019_ );
or   ( new_n28022_, new_n28021_, new_n18977_ );
and  ( new_n28023_, new_n28022_, new_n28018_ );
or   ( new_n28024_, new_n28023_, new_n28014_ );
and  ( new_n28025_, new_n28023_, new_n28014_ );
or   ( new_n28026_, new_n18388_, new_n4635_ );
or   ( new_n28027_, new_n18395_, new_n132_ );
and  ( new_n28028_, new_n28027_, new_n28026_ );
or   ( new_n28029_, new_n28028_, new_n18066_ );
and  ( new_n28030_, new_n18397_, RI2b1c4342e098_90 );
and  ( new_n28031_, new_n18384_, RI2b1c4342e020_89 );
or   ( new_n28032_, new_n28031_, new_n28030_ );
or   ( new_n28033_, new_n28032_, new_n18309_ );
and  ( new_n28034_, new_n28033_, new_n28029_ );
or   ( new_n28035_, new_n28034_, new_n28025_ );
and  ( new_n28036_, new_n28035_, new_n28024_ );
or   ( new_n28037_, new_n28036_, new_n28005_ );
and  ( new_n28038_, new_n28036_, new_n28005_ );
or   ( new_n28039_, new_n17727_, new_n5459_ );
or   ( new_n28040_, new_n17734_, new_n117_ );
and  ( new_n28041_, new_n28040_, new_n28039_ );
or   ( new_n28042_, new_n28041_, new_n17238_ );
and  ( new_n28043_, new_n17736_, RI2b1c4342e188_92 );
and  ( new_n28044_, new_n17723_, RI2b1c4342e110_91 );
or   ( new_n28045_, new_n28044_, new_n28043_ );
or   ( new_n28046_, new_n28045_, new_n17650_ );
and  ( new_n28047_, new_n28046_, new_n28042_ );
or   ( new_n28048_, new_n17244_, new_n6321_ );
or   ( new_n28049_, new_n17248_, new_n6307_ );
and  ( new_n28050_, new_n28049_, new_n28048_ );
or   ( new_n28051_, new_n28050_, new_n16814_ );
and  ( new_n28052_, new_n17255_, RI2b1c4342e278_94 );
and  ( new_n28053_, new_n17240_, RI2b1c4342e200_93 );
or   ( new_n28054_, new_n28053_, new_n28052_ );
or   ( new_n28055_, new_n28054_, new_n17142_ );
and  ( new_n28056_, new_n28055_, new_n28051_ );
or   ( new_n28057_, new_n28056_, new_n28047_ );
and  ( new_n28058_, new_n28056_, new_n28047_ );
or   ( new_n28059_, new_n16607_, new_n7274_ );
or   ( new_n28060_, new_n16613_, new_n124_ );
and  ( new_n28061_, new_n28060_, new_n28059_ );
or   ( new_n28062_, new_n28061_, new_n16505_ );
and  ( new_n28063_, new_n16616_, RI2b1c4342e368_96 );
and  ( new_n28064_, new_n16603_, RI2b1c4342e2f0_95 );
or   ( new_n28065_, new_n28064_, new_n28063_ );
or   ( new_n28066_, new_n28065_, new_n16438_ );
and  ( new_n28067_, new_n28066_, new_n28062_ );
or   ( new_n28068_, new_n28067_, new_n28058_ );
and  ( new_n28069_, new_n28068_, new_n28057_ );
or   ( new_n28070_, new_n28069_, new_n28038_ );
and  ( new_n28071_, new_n28070_, new_n28037_ );
or   ( new_n28072_, new_n16607_, new_n124_ );
or   ( new_n28073_, new_n16613_, new_n6321_ );
and  ( new_n28074_, new_n28073_, new_n28072_ );
or   ( new_n28075_, new_n28074_, new_n16505_ );
and  ( new_n28076_, new_n16616_, RI2b1c4342e2f0_95 );
and  ( new_n28077_, new_n16603_, RI2b1c4342e278_94 );
or   ( new_n28078_, new_n28077_, new_n28076_ );
or   ( new_n28079_, new_n28078_, new_n16438_ );
and  ( new_n28080_, new_n28079_, new_n28075_ );
or   ( new_n28081_, new_n16355_, new_n7274_ );
or   ( new_n28082_, new_n28081_, new_n16085_ );
and  ( new_n28083_, new_n16362_, RI2b1c4342e368_96 );
or   ( new_n28084_, new_n28083_, new_n16048_ );
and  ( new_n28085_, new_n28084_, new_n28082_ );
or   ( new_n28086_, new_n28085_, new_n28080_ );
and  ( new_n28087_, new_n28085_, new_n28080_ );
or   ( new_n28088_, new_n27926_, new_n27818_ );
or   ( new_n28089_, new_n27923_, new_n27827_ );
and  ( new_n28090_, new_n28089_, new_n28088_ );
or   ( new_n28091_, new_n28090_, new_n27931_ );
and  ( new_n28092_, new_n27927_, new_n27828_ );
or   ( new_n28093_, new_n28092_, new_n27838_ );
and  ( new_n28094_, new_n28093_, new_n28091_ );
or   ( new_n28095_, new_n28094_, new_n28087_ );
and  ( new_n28096_, new_n28095_, new_n28086_ );
or   ( new_n28097_, new_n28096_, new_n28071_ );
and  ( new_n28098_, new_n28096_, new_n28071_ );
or   ( new_n28099_, new_n27627_, new_n27464_ );
or   ( new_n28100_, new_n27624_, new_n27473_ );
and  ( new_n28101_, new_n28100_, new_n28099_ );
or   ( new_n28102_, new_n28101_, new_n27632_ );
and  ( new_n28103_, new_n27628_, new_n27474_ );
or   ( new_n28104_, new_n28103_, new_n27484_ );
and  ( new_n28105_, new_n28104_, new_n28102_ );
or   ( new_n28106_, new_n28105_, new_n28098_ );
and  ( new_n28107_, new_n28106_, new_n28097_ );
or   ( new_n28108_, new_n28107_, new_n27975_ );
and  ( new_n28109_, new_n28107_, new_n27975_ );
or   ( new_n28110_, new_n27948_, new_n27842_ );
or   ( new_n28111_, new_n27935_, new_n27755_ );
and  ( new_n28112_, new_n28111_, new_n28110_ );
or   ( new_n28113_, new_n28112_, new_n27953_ );
and  ( new_n28114_, new_n27949_, new_n27844_ );
or   ( new_n28115_, new_n28114_, new_n27851_ );
and  ( new_n28116_, new_n28115_, new_n28113_ );
or   ( new_n28117_, new_n28116_, new_n28109_ );
and  ( new_n28118_, new_n28117_, new_n28108_ );
or   ( new_n28119_, new_n28118_, new_n27972_ );
or   ( new_n28120_, new_n27895_, new_n27853_ );
or   ( new_n28121_, new_n27955_, new_n27728_ );
and  ( new_n28122_, new_n28121_, new_n28120_ );
or   ( new_n28123_, new_n28122_, new_n27960_ );
and  ( new_n28124_, new_n27956_, new_n27855_ );
or   ( new_n28125_, new_n28124_, new_n27862_ );
and  ( new_n28126_, new_n28125_, new_n28123_ );
and  ( new_n28127_, new_n28118_, new_n27972_ );
or   ( new_n28128_, new_n28127_, new_n28126_ );
and  ( new_n28129_, new_n28128_, new_n28119_ );
and  ( new_n28130_, new_n28129_, new_n27969_ );
or   ( new_n28131_, new_n28124_, new_n27960_ );
or   ( new_n28132_, new_n28122_, new_n27862_ );
and  ( new_n28133_, new_n28132_, new_n28131_ );
or   ( new_n28134_, new_n27886_, new_n27883_ );
and  ( new_n28135_, new_n28134_, new_n27713_ );
or   ( new_n28136_, new_n28135_, new_n28118_ );
or   ( new_n28137_, new_n27894_, new_n27891_ );
and  ( new_n28138_, new_n28137_, new_n27728_ );
or   ( new_n28139_, new_n27981_, new_n21261_ );
or   ( new_n28140_, new_n27977_, new_n21009_ );
and  ( new_n28141_, new_n28140_, new_n28139_ );
or   ( new_n28142_, new_n27990_, new_n21013_ );
or   ( new_n28143_, new_n27986_, new_n21265_ );
and  ( new_n28144_, new_n28143_, new_n28142_ );
or   ( new_n28145_, new_n28144_, new_n28141_ );
and  ( new_n28146_, new_n28144_, new_n28141_ );
or   ( new_n28147_, new_n28001_, new_n20156_ );
or   ( new_n28148_, new_n27997_, new_n20443_ );
and  ( new_n28149_, new_n28148_, new_n28147_ );
or   ( new_n28150_, new_n28149_, new_n28146_ );
and  ( new_n28151_, new_n28150_, new_n28145_ );
or   ( new_n28152_, new_n28012_, new_n19394_ );
or   ( new_n28153_, new_n28008_, new_n19659_ );
and  ( new_n28154_, new_n28153_, new_n28152_ );
or   ( new_n28155_, new_n28021_, new_n18742_ );
or   ( new_n28156_, new_n28017_, new_n18977_ );
and  ( new_n28157_, new_n28156_, new_n28155_ );
or   ( new_n28158_, new_n28157_, new_n28154_ );
and  ( new_n28159_, new_n28157_, new_n28154_ );
or   ( new_n28160_, new_n28032_, new_n18066_ );
or   ( new_n28161_, new_n28028_, new_n18309_ );
and  ( new_n28162_, new_n28161_, new_n28160_ );
or   ( new_n28163_, new_n28162_, new_n28159_ );
and  ( new_n28164_, new_n28163_, new_n28158_ );
or   ( new_n28165_, new_n28164_, new_n28151_ );
and  ( new_n28166_, new_n28164_, new_n28151_ );
or   ( new_n28167_, new_n28045_, new_n17238_ );
or   ( new_n28168_, new_n28041_, new_n17650_ );
and  ( new_n28169_, new_n28168_, new_n28167_ );
or   ( new_n28170_, new_n28054_, new_n16814_ );
or   ( new_n28171_, new_n28050_, new_n17142_ );
and  ( new_n28172_, new_n28171_, new_n28170_ );
or   ( new_n28173_, new_n28172_, new_n28169_ );
and  ( new_n28174_, new_n28172_, new_n28169_ );
or   ( new_n28175_, new_n28065_, new_n16505_ );
or   ( new_n28176_, new_n28061_, new_n16438_ );
and  ( new_n28177_, new_n28176_, new_n28175_ );
or   ( new_n28178_, new_n28177_, new_n28174_ );
and  ( new_n28179_, new_n28178_, new_n28173_ );
or   ( new_n28180_, new_n28179_, new_n28166_ );
and  ( new_n28181_, new_n28180_, new_n28165_ );
or   ( new_n28182_, new_n28078_, new_n16505_ );
or   ( new_n28183_, new_n28074_, new_n16438_ );
and  ( new_n28184_, new_n28183_, new_n28182_ );
or   ( new_n28185_, new_n28083_, new_n16085_ );
or   ( new_n28186_, new_n28081_, new_n16048_ );
and  ( new_n28187_, new_n28186_, new_n28185_ );
or   ( new_n28188_, new_n28187_, new_n28184_ );
and  ( new_n28189_, new_n28187_, new_n28184_ );
or   ( new_n28190_, new_n28092_, new_n27931_ );
or   ( new_n28191_, new_n28090_, new_n27838_ );
and  ( new_n28192_, new_n28191_, new_n28190_ );
or   ( new_n28193_, new_n28192_, new_n28189_ );
and  ( new_n28194_, new_n28193_, new_n28188_ );
or   ( new_n28195_, new_n28194_, new_n28181_ );
and  ( new_n28196_, new_n28194_, new_n28181_ );
or   ( new_n28197_, new_n28103_, new_n27632_ );
or   ( new_n28198_, new_n28101_, new_n27484_ );
and  ( new_n28199_, new_n28198_, new_n28197_ );
or   ( new_n28200_, new_n28199_, new_n28196_ );
and  ( new_n28201_, new_n28200_, new_n28195_ );
or   ( new_n28202_, new_n28201_, new_n28138_ );
and  ( new_n28203_, new_n28201_, new_n28138_ );
or   ( new_n28204_, new_n28114_, new_n27953_ );
or   ( new_n28205_, new_n28112_, new_n27851_ );
and  ( new_n28206_, new_n28205_, new_n28204_ );
or   ( new_n28207_, new_n28206_, new_n28203_ );
and  ( new_n28208_, new_n28207_, new_n28202_ );
or   ( new_n28209_, new_n28208_, new_n27972_ );
and  ( new_n28210_, new_n28209_, new_n28136_ );
or   ( new_n28211_, new_n28210_, new_n28133_ );
or   ( new_n28212_, new_n28208_, new_n28135_ );
and  ( new_n28213_, new_n28212_, new_n28119_ );
or   ( new_n28214_, new_n28213_, new_n28126_ );
and  ( new_n28215_, new_n28214_, new_n28211_ );
or   ( new_n28216_, new_n27908_, new_n27807_ );
or   ( new_n28217_, new_n27918_, new_n27786_ );
and  ( new_n28218_, new_n28217_, new_n28216_ );
or   ( new_n28219_, new_n28218_, new_n27933_ );
and  ( new_n28220_, new_n27919_, new_n27809_ );
or   ( new_n28221_, new_n28220_, new_n27840_ );
and  ( new_n28222_, new_n28221_, new_n28219_ );
or   ( new_n28223_, new_n28194_, new_n28071_ );
or   ( new_n28224_, new_n28181_, new_n28096_ );
and  ( new_n28225_, new_n28224_, new_n28223_ );
or   ( new_n28226_, new_n28225_, new_n28199_ );
and  ( new_n28227_, new_n28195_, new_n28097_ );
or   ( new_n28228_, new_n28227_, new_n28105_ );
and  ( new_n28229_, new_n28228_, new_n28226_ );
or   ( new_n28230_, new_n28229_, new_n28222_ );
or   ( new_n28231_, new_n27911_, new_n16048_ );
or   ( new_n28232_, new_n27794_, new_n16085_ );
and  ( new_n28233_, new_n28232_, new_n28231_ );
or   ( new_n28234_, new_n28233_, new_n27916_ );
and  ( new_n28235_, new_n27912_, new_n27796_ );
or   ( new_n28236_, new_n28235_, new_n27805_ );
and  ( new_n28237_, new_n28236_, new_n28234_ );
or   ( new_n28238_, new_n28187_, new_n28080_ );
or   ( new_n28239_, new_n28184_, new_n28085_ );
and  ( new_n28240_, new_n28239_, new_n28238_ );
or   ( new_n28241_, new_n28240_, new_n28192_ );
and  ( new_n28242_, new_n28188_, new_n28086_ );
or   ( new_n28243_, new_n28242_, new_n28094_ );
and  ( new_n28244_, new_n28243_, new_n28241_ );
or   ( new_n28245_, new_n28244_, new_n28237_ );
and  ( new_n28246_, new_n28244_, new_n28237_ );
or   ( new_n28247_, new_n28164_, new_n28005_ );
or   ( new_n28248_, new_n28151_, new_n28036_ );
and  ( new_n28249_, new_n28248_, new_n28247_ );
or   ( new_n28250_, new_n28249_, new_n28179_ );
and  ( new_n28251_, new_n28165_, new_n28037_ );
or   ( new_n28252_, new_n28251_, new_n28069_ );
and  ( new_n28253_, new_n28252_, new_n28250_ );
or   ( new_n28254_, new_n28253_, new_n28246_ );
and  ( new_n28255_, new_n28254_, new_n28245_ );
or   ( new_n28256_, new_n28172_, new_n28047_ );
or   ( new_n28257_, new_n28169_, new_n28056_ );
and  ( new_n28258_, new_n28257_, new_n28256_ );
or   ( new_n28259_, new_n28258_, new_n28177_ );
and  ( new_n28260_, new_n28173_, new_n28057_ );
or   ( new_n28261_, new_n28260_, new_n28067_ );
and  ( new_n28262_, new_n28261_, new_n28259_ );
or   ( new_n28263_, new_n28157_, new_n28014_ );
or   ( new_n28264_, new_n28154_, new_n28023_ );
and  ( new_n28265_, new_n28264_, new_n28263_ );
or   ( new_n28266_, new_n28265_, new_n28162_ );
and  ( new_n28267_, new_n28158_, new_n28024_ );
or   ( new_n28268_, new_n28267_, new_n28034_ );
and  ( new_n28269_, new_n28268_, new_n28266_ );
or   ( new_n28270_, new_n28269_, new_n28262_ );
and  ( new_n28271_, new_n28269_, new_n28262_ );
or   ( new_n28272_, new_n28144_, new_n27983_ );
or   ( new_n28273_, new_n28141_, new_n27992_ );
and  ( new_n28274_, new_n28273_, new_n28272_ );
or   ( new_n28275_, new_n28274_, new_n28149_ );
and  ( new_n28276_, new_n28145_, new_n27993_ );
or   ( new_n28277_, new_n28276_, new_n28003_ );
and  ( new_n28278_, new_n28277_, new_n28275_ );
or   ( new_n28279_, new_n28278_, new_n28271_ );
and  ( new_n28280_, new_n28279_, new_n28270_ );
or   ( new_n28281_, new_n20557_, new_n2806_ );
or   ( new_n28282_, new_n20562_, new_n2541_ );
and  ( new_n28283_, new_n28282_, new_n28281_ );
or   ( new_n28284_, new_n28283_, new_n20156_ );
and  ( new_n28285_, new_n20566_, RI2b1c4342de40_85 );
and  ( new_n28286_, new_n20553_, RI2b1c4342ddc8_84 );
or   ( new_n28287_, new_n28286_, new_n28285_ );
or   ( new_n28288_, new_n28287_, new_n20443_ );
and  ( new_n28289_, new_n28288_, new_n28284_ );
or   ( new_n28290_, new_n19758_, new_n3924_ );
or   ( new_n28291_, new_n19763_, new_n3239_ );
and  ( new_n28292_, new_n28291_, new_n28290_ );
or   ( new_n28293_, new_n28292_, new_n19394_ );
and  ( new_n28294_, new_n19767_, RI2b1c4342df30_87 );
and  ( new_n28295_, new_n19754_, RI2b1c4342deb8_86 );
or   ( new_n28296_, new_n28295_, new_n28294_ );
or   ( new_n28297_, new_n28296_, new_n19659_ );
and  ( new_n28298_, new_n28297_, new_n28293_ );
or   ( new_n28299_, new_n28298_, new_n28289_ );
and  ( new_n28300_, new_n28298_, new_n28289_ );
or   ( new_n28301_, new_n19048_, new_n132_ );
or   ( new_n28302_, new_n19055_, new_n3902_ );
and  ( new_n28303_, new_n28302_, new_n28301_ );
or   ( new_n28304_, new_n28303_, new_n18742_ );
and  ( new_n28305_, new_n19057_, RI2b1c4342e020_89 );
and  ( new_n28306_, new_n19044_, RI2b1c4342dfa8_88 );
or   ( new_n28307_, new_n28306_, new_n28305_ );
or   ( new_n28308_, new_n28307_, new_n18977_ );
and  ( new_n28309_, new_n28308_, new_n28304_ );
or   ( new_n28310_, new_n28309_, new_n28300_ );
and  ( new_n28311_, new_n28310_, new_n28299_ );
nor  ( new_n28312_, new_n22333_, new_n126_ );
nor  ( new_n28313_, new_n28312_, new_n13173_ );
or   ( new_n28314_, new_n28313_, new_n21261_ );
and  ( new_n28315_, new_n22337_, RI2b1c4342dc60_81 );
and  ( new_n28316_, new_n22330_, RI2b1c4342dbe8_80 );
or   ( new_n28317_, new_n28316_, new_n28315_ );
or   ( new_n28318_, new_n28317_, new_n21009_ );
and  ( new_n28319_, new_n28318_, new_n28314_ );
and  ( new_n28320_, new_n28319_, new_n16438_ );
or   ( new_n28321_, new_n28319_, new_n16438_ );
or   ( new_n28322_, new_n21419_, new_n121_ );
or   ( new_n28323_, new_n21424_, new_n2119_ );
and  ( new_n28324_, new_n28323_, new_n28322_ );
or   ( new_n28325_, new_n28324_, new_n21013_ );
and  ( new_n28326_, new_n21428_, RI2b1c4342dd50_83 );
and  ( new_n28327_, new_n21415_, RI2b1c4342dcd8_82 );
or   ( new_n28328_, new_n28327_, new_n28326_ );
or   ( new_n28329_, new_n28328_, new_n21265_ );
and  ( new_n28330_, new_n28329_, new_n28325_ );
and  ( new_n28331_, new_n28330_, new_n28321_ );
or   ( new_n28332_, new_n28331_, new_n28320_ );
and  ( new_n28333_, new_n28332_, new_n28311_ );
or   ( new_n28334_, new_n28332_, new_n28311_ );
or   ( new_n28335_, new_n18388_, new_n117_ );
or   ( new_n28336_, new_n18395_, new_n4635_ );
and  ( new_n28337_, new_n28336_, new_n28335_ );
or   ( new_n28338_, new_n28337_, new_n18066_ );
and  ( new_n28339_, new_n18397_, RI2b1c4342e110_91 );
and  ( new_n28340_, new_n18384_, RI2b1c4342e098_90 );
or   ( new_n28341_, new_n28340_, new_n28339_ );
or   ( new_n28342_, new_n28341_, new_n18309_ );
and  ( new_n28343_, new_n28342_, new_n28338_ );
or   ( new_n28344_, new_n17727_, new_n6307_ );
or   ( new_n28345_, new_n17734_, new_n5459_ );
and  ( new_n28346_, new_n28345_, new_n28344_ );
or   ( new_n28347_, new_n28346_, new_n17238_ );
and  ( new_n28348_, new_n17736_, RI2b1c4342e200_93 );
and  ( new_n28349_, new_n17723_, RI2b1c4342e188_92 );
or   ( new_n28350_, new_n28349_, new_n28348_ );
or   ( new_n28351_, new_n28350_, new_n17650_ );
and  ( new_n28352_, new_n28351_, new_n28347_ );
or   ( new_n28353_, new_n28352_, new_n28343_ );
and  ( new_n28354_, new_n28352_, new_n28343_ );
or   ( new_n28355_, new_n17244_, new_n124_ );
or   ( new_n28356_, new_n17248_, new_n6321_ );
and  ( new_n28357_, new_n28356_, new_n28355_ );
or   ( new_n28358_, new_n28357_, new_n16814_ );
and  ( new_n28359_, new_n17255_, RI2b1c4342e2f0_95 );
and  ( new_n28360_, new_n17240_, RI2b1c4342e278_94 );
or   ( new_n28361_, new_n28360_, new_n28359_ );
or   ( new_n28362_, new_n28361_, new_n17142_ );
and  ( new_n28363_, new_n28362_, new_n28358_ );
or   ( new_n28364_, new_n28363_, new_n28354_ );
and  ( new_n28365_, new_n28364_, new_n28353_ );
and  ( new_n28366_, new_n28365_, new_n28334_ );
or   ( new_n28367_, new_n28366_, new_n28333_ );
and  ( new_n28368_, new_n28367_, new_n28280_ );
or   ( new_n28369_, new_n28367_, new_n28280_ );
or   ( new_n28370_, new_n27901_, new_n27764_ );
or   ( new_n28371_, new_n27898_, new_n27773_ );
and  ( new_n28372_, new_n28371_, new_n28370_ );
or   ( new_n28373_, new_n28372_, new_n27906_ );
and  ( new_n28374_, new_n27902_, new_n27774_ );
or   ( new_n28375_, new_n28374_, new_n27784_ );
and  ( new_n28376_, new_n28375_, new_n28373_ );
and  ( new_n28377_, new_n28376_, new_n28369_ );
or   ( new_n28378_, new_n28377_, new_n28368_ );
and  ( new_n28379_, new_n28378_, new_n28255_ );
or   ( new_n28380_, new_n28378_, new_n28255_ );
or   ( new_n28381_, new_n27941_, new_n27737_ );
or   ( new_n28382_, new_n27938_, new_n27744_ );
and  ( new_n28383_, new_n28382_, new_n28381_ );
or   ( new_n28384_, new_n28383_, new_n27946_ );
and  ( new_n28385_, new_n27942_, new_n27745_ );
or   ( new_n28386_, new_n28385_, new_n27753_ );
and  ( new_n28387_, new_n28386_, new_n28384_ );
and  ( new_n28388_, new_n28387_, new_n28380_ );
or   ( new_n28389_, new_n28388_, new_n28379_ );
and  ( new_n28390_, new_n28389_, new_n28230_ );
or   ( new_n28391_, new_n28389_, new_n28230_ );
or   ( new_n28392_, new_n28138_, new_n28107_ );
or   ( new_n28393_, new_n28201_, new_n27975_ );
and  ( new_n28394_, new_n28393_, new_n28392_ );
or   ( new_n28395_, new_n28394_, new_n28206_ );
and  ( new_n28396_, new_n28202_, new_n28108_ );
or   ( new_n28397_, new_n28396_, new_n28116_ );
and  ( new_n28398_, new_n28397_, new_n28395_ );
and  ( new_n28399_, new_n28398_, new_n28391_ );
or   ( new_n28400_, new_n28399_, new_n28390_ );
and  ( new_n28401_, new_n28400_, new_n28215_ );
or   ( new_n28402_, new_n28401_, new_n28130_ );
or   ( new_n28403_, new_n28396_, new_n28206_ );
or   ( new_n28404_, new_n28394_, new_n28116_ );
and  ( new_n28405_, new_n28404_, new_n28403_ );
or   ( new_n28406_, new_n28220_, new_n27933_ );
or   ( new_n28407_, new_n28218_, new_n27840_ );
and  ( new_n28408_, new_n28407_, new_n28406_ );
or   ( new_n28409_, new_n28227_, new_n28199_ );
or   ( new_n28410_, new_n28225_, new_n28105_ );
and  ( new_n28411_, new_n28410_, new_n28409_ );
and  ( new_n28412_, new_n28411_, new_n28408_ );
or   ( new_n28413_, new_n28412_, new_n28389_ );
or   ( new_n28414_, new_n28235_, new_n27916_ );
or   ( new_n28415_, new_n28233_, new_n27805_ );
and  ( new_n28416_, new_n28415_, new_n28414_ );
or   ( new_n28417_, new_n28242_, new_n28192_ );
or   ( new_n28418_, new_n28240_, new_n28094_ );
and  ( new_n28419_, new_n28418_, new_n28417_ );
or   ( new_n28420_, new_n28419_, new_n28416_ );
and  ( new_n28421_, new_n28419_, new_n28416_ );
or   ( new_n28422_, new_n28251_, new_n28179_ );
or   ( new_n28423_, new_n28249_, new_n28069_ );
and  ( new_n28424_, new_n28423_, new_n28422_ );
or   ( new_n28425_, new_n28424_, new_n28421_ );
and  ( new_n28426_, new_n28425_, new_n28420_ );
or   ( new_n28427_, new_n28260_, new_n28177_ );
or   ( new_n28428_, new_n28258_, new_n28067_ );
and  ( new_n28429_, new_n28428_, new_n28427_ );
or   ( new_n28430_, new_n28267_, new_n28162_ );
or   ( new_n28431_, new_n28265_, new_n28034_ );
and  ( new_n28432_, new_n28431_, new_n28430_ );
or   ( new_n28433_, new_n28432_, new_n28429_ );
and  ( new_n28434_, new_n28432_, new_n28429_ );
or   ( new_n28435_, new_n28276_, new_n28149_ );
or   ( new_n28436_, new_n28274_, new_n28003_ );
and  ( new_n28437_, new_n28436_, new_n28435_ );
or   ( new_n28438_, new_n28437_, new_n28434_ );
and  ( new_n28439_, new_n28438_, new_n28433_ );
or   ( new_n28440_, new_n28287_, new_n20156_ );
or   ( new_n28441_, new_n28283_, new_n20443_ );
and  ( new_n28442_, new_n28441_, new_n28440_ );
or   ( new_n28443_, new_n28296_, new_n19394_ );
or   ( new_n28444_, new_n28292_, new_n19659_ );
and  ( new_n28445_, new_n28444_, new_n28443_ );
or   ( new_n28446_, new_n28445_, new_n28442_ );
and  ( new_n28447_, new_n28445_, new_n28442_ );
or   ( new_n28448_, new_n28307_, new_n18742_ );
or   ( new_n28449_, new_n28303_, new_n18977_ );
and  ( new_n28450_, new_n28449_, new_n28448_ );
or   ( new_n28451_, new_n28450_, new_n28447_ );
and  ( new_n28452_, new_n28451_, new_n28446_ );
or   ( new_n28453_, new_n28317_, new_n21261_ );
or   ( new_n28454_, new_n28313_, new_n21009_ );
and  ( new_n28455_, new_n28454_, new_n28453_ );
or   ( new_n28456_, new_n28455_, new_n16505_ );
and  ( new_n28457_, new_n28455_, new_n16505_ );
or   ( new_n28458_, new_n28328_, new_n21013_ );
or   ( new_n28459_, new_n28324_, new_n21265_ );
and  ( new_n28460_, new_n28459_, new_n28458_ );
or   ( new_n28461_, new_n28460_, new_n28457_ );
and  ( new_n28462_, new_n28461_, new_n28456_ );
or   ( new_n28463_, new_n28462_, new_n28452_ );
and  ( new_n28464_, new_n28462_, new_n28452_ );
or   ( new_n28465_, new_n28341_, new_n18066_ );
or   ( new_n28466_, new_n28337_, new_n18309_ );
and  ( new_n28467_, new_n28466_, new_n28465_ );
or   ( new_n28468_, new_n28350_, new_n17238_ );
or   ( new_n28469_, new_n28346_, new_n17650_ );
and  ( new_n28470_, new_n28469_, new_n28468_ );
or   ( new_n28471_, new_n28470_, new_n28467_ );
and  ( new_n28472_, new_n28470_, new_n28467_ );
or   ( new_n28473_, new_n28361_, new_n16814_ );
or   ( new_n28474_, new_n28357_, new_n17142_ );
and  ( new_n28475_, new_n28474_, new_n28473_ );
or   ( new_n28476_, new_n28475_, new_n28472_ );
and  ( new_n28477_, new_n28476_, new_n28471_ );
or   ( new_n28478_, new_n28477_, new_n28464_ );
and  ( new_n28479_, new_n28478_, new_n28463_ );
or   ( new_n28480_, new_n28479_, new_n28439_ );
and  ( new_n28481_, new_n28479_, new_n28439_ );
or   ( new_n28482_, new_n28374_, new_n27906_ );
or   ( new_n28483_, new_n28372_, new_n27784_ );
and  ( new_n28484_, new_n28483_, new_n28482_ );
or   ( new_n28485_, new_n28484_, new_n28481_ );
and  ( new_n28486_, new_n28485_, new_n28480_ );
or   ( new_n28487_, new_n28486_, new_n28426_ );
and  ( new_n28488_, new_n28486_, new_n28426_ );
or   ( new_n28489_, new_n28385_, new_n27946_ );
or   ( new_n28490_, new_n28383_, new_n27753_ );
and  ( new_n28491_, new_n28490_, new_n28489_ );
or   ( new_n28492_, new_n28491_, new_n28488_ );
and  ( new_n28493_, new_n28492_, new_n28487_ );
or   ( new_n28494_, new_n28493_, new_n28230_ );
and  ( new_n28495_, new_n28494_, new_n28413_ );
or   ( new_n28496_, new_n28495_, new_n28405_ );
or   ( new_n28497_, new_n28493_, new_n28412_ );
and  ( new_n28498_, new_n28497_, new_n28391_ );
or   ( new_n28499_, new_n28498_, new_n28398_ );
and  ( new_n28500_, new_n28499_, new_n28496_ );
or   ( new_n28501_, new_n28411_, new_n28222_ );
or   ( new_n28502_, new_n28408_, new_n28229_ );
and  ( new_n28503_, new_n28502_, new_n28501_ );
or   ( new_n28504_, new_n28419_, new_n28237_ );
or   ( new_n28505_, new_n28416_, new_n28244_ );
and  ( new_n28506_, new_n28505_, new_n28504_ );
or   ( new_n28507_, new_n28506_, new_n28424_ );
and  ( new_n28508_, new_n28420_, new_n28245_ );
or   ( new_n28509_, new_n28508_, new_n28253_ );
and  ( new_n28510_, new_n28509_, new_n28507_ );
nor  ( new_n28511_, new_n22333_, new_n2119_ );
nor  ( new_n28512_, new_n28511_, new_n13372_ );
or   ( new_n28513_, new_n28512_, new_n21261_ );
and  ( new_n28514_, new_n22337_, RI2b1c4342dcd8_82 );
and  ( new_n28515_, new_n22330_, RI2b1c4342dc60_81 );
or   ( new_n28516_, new_n28515_, new_n28514_ );
or   ( new_n28517_, new_n28516_, new_n21009_ );
and  ( new_n28518_, new_n28517_, new_n28513_ );
or   ( new_n28519_, new_n21419_, new_n2541_ );
or   ( new_n28520_, new_n21424_, new_n121_ );
and  ( new_n28521_, new_n28520_, new_n28519_ );
or   ( new_n28522_, new_n28521_, new_n21013_ );
and  ( new_n28523_, new_n21428_, RI2b1c4342ddc8_84 );
and  ( new_n28524_, new_n21415_, RI2b1c4342dd50_83 );
or   ( new_n28525_, new_n28524_, new_n28523_ );
or   ( new_n28526_, new_n28525_, new_n21265_ );
and  ( new_n28527_, new_n28526_, new_n28522_ );
or   ( new_n28528_, new_n28527_, new_n28518_ );
and  ( new_n28529_, new_n28527_, new_n28518_ );
or   ( new_n28530_, new_n20557_, new_n3239_ );
or   ( new_n28531_, new_n20562_, new_n2806_ );
and  ( new_n28532_, new_n28531_, new_n28530_ );
or   ( new_n28533_, new_n28532_, new_n20156_ );
and  ( new_n28534_, new_n20566_, RI2b1c4342deb8_86 );
and  ( new_n28535_, new_n20553_, RI2b1c4342de40_85 );
or   ( new_n28536_, new_n28535_, new_n28534_ );
or   ( new_n28537_, new_n28536_, new_n20443_ );
and  ( new_n28538_, new_n28537_, new_n28533_ );
or   ( new_n28539_, new_n28538_, new_n28529_ );
and  ( new_n28540_, new_n28539_, new_n28528_ );
or   ( new_n28541_, new_n19758_, new_n3902_ );
or   ( new_n28542_, new_n19763_, new_n3924_ );
and  ( new_n28543_, new_n28542_, new_n28541_ );
or   ( new_n28544_, new_n28543_, new_n19394_ );
and  ( new_n28545_, new_n19767_, RI2b1c4342dfa8_88 );
and  ( new_n28546_, new_n19754_, RI2b1c4342df30_87 );
or   ( new_n28547_, new_n28546_, new_n28545_ );
or   ( new_n28548_, new_n28547_, new_n19659_ );
and  ( new_n28549_, new_n28548_, new_n28544_ );
or   ( new_n28550_, new_n19048_, new_n4635_ );
or   ( new_n28551_, new_n19055_, new_n132_ );
and  ( new_n28552_, new_n28551_, new_n28550_ );
or   ( new_n28553_, new_n28552_, new_n18742_ );
and  ( new_n28554_, new_n19057_, RI2b1c4342e098_90 );
and  ( new_n28555_, new_n19044_, RI2b1c4342e020_89 );
or   ( new_n28556_, new_n28555_, new_n28554_ );
or   ( new_n28557_, new_n28556_, new_n18977_ );
and  ( new_n28558_, new_n28557_, new_n28553_ );
or   ( new_n28559_, new_n28558_, new_n28549_ );
and  ( new_n28560_, new_n28558_, new_n28549_ );
or   ( new_n28561_, new_n18388_, new_n5459_ );
or   ( new_n28562_, new_n18395_, new_n117_ );
and  ( new_n28563_, new_n28562_, new_n28561_ );
or   ( new_n28564_, new_n28563_, new_n18066_ );
and  ( new_n28565_, new_n18397_, RI2b1c4342e188_92 );
and  ( new_n28566_, new_n18384_, RI2b1c4342e110_91 );
or   ( new_n28567_, new_n28566_, new_n28565_ );
or   ( new_n28568_, new_n28567_, new_n18309_ );
and  ( new_n28569_, new_n28568_, new_n28564_ );
or   ( new_n28570_, new_n28569_, new_n28560_ );
and  ( new_n28571_, new_n28570_, new_n28559_ );
or   ( new_n28572_, new_n28571_, new_n28540_ );
and  ( new_n28573_, new_n28571_, new_n28540_ );
or   ( new_n28574_, new_n17727_, new_n6321_ );
or   ( new_n28575_, new_n17734_, new_n6307_ );
and  ( new_n28576_, new_n28575_, new_n28574_ );
or   ( new_n28577_, new_n28576_, new_n17238_ );
and  ( new_n28578_, new_n17736_, RI2b1c4342e278_94 );
and  ( new_n28579_, new_n17723_, RI2b1c4342e200_93 );
or   ( new_n28580_, new_n28579_, new_n28578_ );
or   ( new_n28581_, new_n28580_, new_n17650_ );
and  ( new_n28582_, new_n28581_, new_n28577_ );
or   ( new_n28583_, new_n17244_, new_n7274_ );
or   ( new_n28584_, new_n17248_, new_n124_ );
and  ( new_n28585_, new_n28584_, new_n28583_ );
or   ( new_n28586_, new_n28585_, new_n16814_ );
and  ( new_n28587_, new_n17255_, RI2b1c4342e368_96 );
and  ( new_n28588_, new_n17240_, RI2b1c4342e2f0_95 );
or   ( new_n28589_, new_n28588_, new_n28587_ );
or   ( new_n28590_, new_n28589_, new_n17142_ );
and  ( new_n28591_, new_n28590_, new_n28586_ );
or   ( new_n28592_, new_n28591_, new_n28582_ );
or   ( new_n28593_, new_n28592_, new_n28573_ );
and  ( new_n28594_, new_n28593_, new_n28572_ );
or   ( new_n28595_, new_n16613_, new_n7274_ );
or   ( new_n28596_, new_n28595_, new_n16505_ );
and  ( new_n28597_, new_n16603_, RI2b1c4342e368_96 );
or   ( new_n28598_, new_n28597_, new_n16438_ );
and  ( new_n28599_, new_n28598_, new_n28596_ );
or   ( new_n28600_, new_n28470_, new_n28343_ );
or   ( new_n28601_, new_n28467_, new_n28352_ );
and  ( new_n28602_, new_n28601_, new_n28600_ );
or   ( new_n28603_, new_n28602_, new_n28475_ );
and  ( new_n28604_, new_n28471_, new_n28353_ );
or   ( new_n28605_, new_n28604_, new_n28363_ );
and  ( new_n28606_, new_n28605_, new_n28603_ );
or   ( new_n28607_, new_n28606_, new_n28599_ );
and  ( new_n28608_, new_n28606_, new_n28599_ );
or   ( new_n28609_, new_n28445_, new_n28289_ );
or   ( new_n28610_, new_n28442_, new_n28298_ );
and  ( new_n28611_, new_n28610_, new_n28609_ );
or   ( new_n28612_, new_n28611_, new_n28450_ );
and  ( new_n28613_, new_n28446_, new_n28299_ );
or   ( new_n28614_, new_n28613_, new_n28309_ );
and  ( new_n28615_, new_n28614_, new_n28612_ );
or   ( new_n28616_, new_n28615_, new_n28608_ );
and  ( new_n28617_, new_n28616_, new_n28607_ );
or   ( new_n28618_, new_n28617_, new_n28594_ );
and  ( new_n28619_, new_n28617_, new_n28594_ );
or   ( new_n28620_, new_n28432_, new_n28262_ );
or   ( new_n28621_, new_n28429_, new_n28269_ );
and  ( new_n28622_, new_n28621_, new_n28620_ );
or   ( new_n28623_, new_n28622_, new_n28437_ );
and  ( new_n28624_, new_n28433_, new_n28270_ );
or   ( new_n28625_, new_n28624_, new_n28278_ );
and  ( new_n28626_, new_n28625_, new_n28623_ );
or   ( new_n28627_, new_n28626_, new_n28619_ );
and  ( new_n28628_, new_n28627_, new_n28618_ );
or   ( new_n28629_, new_n28628_, new_n28510_ );
and  ( new_n28630_, new_n28628_, new_n28510_ );
or   ( new_n28631_, new_n28439_, new_n28367_ );
or   ( new_n28632_, new_n28479_, new_n28280_ );
and  ( new_n28633_, new_n28632_, new_n28631_ );
or   ( new_n28634_, new_n28633_, new_n28484_ );
and  ( new_n28635_, new_n28480_, new_n28369_ );
or   ( new_n28636_, new_n28635_, new_n28376_ );
and  ( new_n28637_, new_n28636_, new_n28634_ );
or   ( new_n28638_, new_n28637_, new_n28630_ );
and  ( new_n28639_, new_n28638_, new_n28629_ );
or   ( new_n28640_, new_n28639_, new_n28503_ );
or   ( new_n28641_, new_n28426_, new_n28378_ );
or   ( new_n28642_, new_n28486_, new_n28255_ );
and  ( new_n28643_, new_n28642_, new_n28641_ );
or   ( new_n28644_, new_n28643_, new_n28491_ );
and  ( new_n28645_, new_n28487_, new_n28380_ );
or   ( new_n28646_, new_n28645_, new_n28387_ );
and  ( new_n28647_, new_n28646_, new_n28644_ );
and  ( new_n28648_, new_n28639_, new_n28503_ );
or   ( new_n28649_, new_n28648_, new_n28647_ );
and  ( new_n28650_, new_n28649_, new_n28640_ );
and  ( new_n28651_, new_n28650_, new_n28500_ );
or   ( new_n28652_, new_n28635_, new_n28484_ );
or   ( new_n28653_, new_n28633_, new_n28376_ );
and  ( new_n28654_, new_n28653_, new_n28652_ );
or   ( new_n28655_, new_n28508_, new_n28424_ );
or   ( new_n28656_, new_n28506_, new_n28253_ );
and  ( new_n28657_, new_n28656_, new_n28655_ );
or   ( new_n28658_, new_n28657_, new_n28628_ );
or   ( new_n28659_, new_n28516_, new_n21261_ );
or   ( new_n28660_, new_n28512_, new_n21009_ );
and  ( new_n28661_, new_n28660_, new_n28659_ );
or   ( new_n28662_, new_n28525_, new_n21013_ );
or   ( new_n28663_, new_n28521_, new_n21265_ );
and  ( new_n28664_, new_n28663_, new_n28662_ );
or   ( new_n28665_, new_n28664_, new_n28661_ );
and  ( new_n28666_, new_n28664_, new_n28661_ );
or   ( new_n28667_, new_n28536_, new_n20156_ );
or   ( new_n28668_, new_n28532_, new_n20443_ );
and  ( new_n28669_, new_n28668_, new_n28667_ );
or   ( new_n28670_, new_n28669_, new_n28666_ );
and  ( new_n28671_, new_n28670_, new_n28665_ );
or   ( new_n28672_, new_n28547_, new_n19394_ );
or   ( new_n28673_, new_n28543_, new_n19659_ );
and  ( new_n28674_, new_n28673_, new_n28672_ );
or   ( new_n28675_, new_n28556_, new_n18742_ );
or   ( new_n28676_, new_n28552_, new_n18977_ );
and  ( new_n28677_, new_n28676_, new_n28675_ );
or   ( new_n28678_, new_n28677_, new_n28674_ );
and  ( new_n28679_, new_n28677_, new_n28674_ );
or   ( new_n28680_, new_n28567_, new_n18066_ );
or   ( new_n28681_, new_n28563_, new_n18309_ );
and  ( new_n28682_, new_n28681_, new_n28680_ );
or   ( new_n28683_, new_n28682_, new_n28679_ );
and  ( new_n28684_, new_n28683_, new_n28678_ );
or   ( new_n28685_, new_n28684_, new_n28671_ );
and  ( new_n28686_, new_n28684_, new_n28671_ );
or   ( new_n28687_, new_n28580_, new_n17238_ );
or   ( new_n28688_, new_n28576_, new_n17650_ );
and  ( new_n28689_, new_n28688_, new_n28687_ );
or   ( new_n28690_, new_n28589_, new_n16814_ );
or   ( new_n28691_, new_n28585_, new_n17142_ );
and  ( new_n28692_, new_n28691_, new_n28690_ );
and  ( new_n28693_, new_n28692_, new_n28689_ );
or   ( new_n28694_, new_n28693_, new_n28686_ );
and  ( new_n28695_, new_n28694_, new_n28685_ );
or   ( new_n28696_, new_n28597_, new_n16505_ );
or   ( new_n28697_, new_n28595_, new_n16438_ );
and  ( new_n28698_, new_n28697_, new_n28696_ );
or   ( new_n28699_, new_n28604_, new_n28475_ );
or   ( new_n28700_, new_n28602_, new_n28363_ );
and  ( new_n28701_, new_n28700_, new_n28699_ );
or   ( new_n28702_, new_n28701_, new_n28698_ );
and  ( new_n28703_, new_n28701_, new_n28698_ );
or   ( new_n28704_, new_n28613_, new_n28450_ );
or   ( new_n28705_, new_n28611_, new_n28309_ );
and  ( new_n28706_, new_n28705_, new_n28704_ );
or   ( new_n28707_, new_n28706_, new_n28703_ );
and  ( new_n28708_, new_n28707_, new_n28702_ );
or   ( new_n28709_, new_n28708_, new_n28695_ );
and  ( new_n28710_, new_n28708_, new_n28695_ );
or   ( new_n28711_, new_n28624_, new_n28437_ );
or   ( new_n28712_, new_n28622_, new_n28278_ );
and  ( new_n28713_, new_n28712_, new_n28711_ );
or   ( new_n28714_, new_n28713_, new_n28710_ );
and  ( new_n28715_, new_n28714_, new_n28709_ );
or   ( new_n28716_, new_n28715_, new_n28510_ );
and  ( new_n28717_, new_n28716_, new_n28658_ );
or   ( new_n28718_, new_n28717_, new_n28654_ );
or   ( new_n28719_, new_n28715_, new_n28657_ );
and  ( new_n28720_, new_n28719_, new_n28629_ );
or   ( new_n28721_, new_n28720_, new_n28637_ );
and  ( new_n28722_, new_n28721_, new_n28718_ );
or   ( new_n28723_, new_n28692_, new_n28582_ );
or   ( new_n28724_, new_n28689_, new_n28591_ );
and  ( new_n28725_, new_n28724_, new_n28723_ );
or   ( new_n28726_, new_n28677_, new_n28549_ );
or   ( new_n28727_, new_n28674_, new_n28558_ );
and  ( new_n28728_, new_n28727_, new_n28726_ );
or   ( new_n28729_, new_n28728_, new_n28682_ );
and  ( new_n28730_, new_n28678_, new_n28559_ );
or   ( new_n28731_, new_n28730_, new_n28569_ );
and  ( new_n28732_, new_n28731_, new_n28729_ );
or   ( new_n28733_, new_n28732_, new_n28725_ );
and  ( new_n28734_, new_n28732_, new_n28725_ );
or   ( new_n28735_, new_n28664_, new_n28518_ );
or   ( new_n28736_, new_n28661_, new_n28527_ );
and  ( new_n28737_, new_n28736_, new_n28735_ );
or   ( new_n28738_, new_n28737_, new_n28669_ );
and  ( new_n28739_, new_n28665_, new_n28528_ );
or   ( new_n28740_, new_n28739_, new_n28538_ );
and  ( new_n28741_, new_n28740_, new_n28738_ );
or   ( new_n28742_, new_n28741_, new_n28734_ );
and  ( new_n28743_, new_n28742_, new_n28733_ );
or   ( new_n28744_, new_n20557_, new_n3924_ );
or   ( new_n28745_, new_n20562_, new_n3239_ );
and  ( new_n28746_, new_n28745_, new_n28744_ );
or   ( new_n28747_, new_n28746_, new_n20156_ );
and  ( new_n28748_, new_n20566_, RI2b1c4342df30_87 );
and  ( new_n28749_, new_n20553_, RI2b1c4342deb8_86 );
or   ( new_n28750_, new_n28749_, new_n28748_ );
or   ( new_n28751_, new_n28750_, new_n20443_ );
and  ( new_n28752_, new_n28751_, new_n28747_ );
or   ( new_n28753_, new_n19758_, new_n132_ );
or   ( new_n28754_, new_n19763_, new_n3902_ );
and  ( new_n28755_, new_n28754_, new_n28753_ );
or   ( new_n28756_, new_n28755_, new_n19394_ );
and  ( new_n28757_, new_n19767_, RI2b1c4342e020_89 );
and  ( new_n28758_, new_n19754_, RI2b1c4342dfa8_88 );
or   ( new_n28759_, new_n28758_, new_n28757_ );
or   ( new_n28760_, new_n28759_, new_n19659_ );
and  ( new_n28761_, new_n28760_, new_n28756_ );
or   ( new_n28762_, new_n28761_, new_n28752_ );
and  ( new_n28763_, new_n28761_, new_n28752_ );
or   ( new_n28764_, new_n19048_, new_n117_ );
or   ( new_n28765_, new_n19055_, new_n4635_ );
and  ( new_n28766_, new_n28765_, new_n28764_ );
or   ( new_n28767_, new_n28766_, new_n18742_ );
and  ( new_n28768_, new_n19057_, RI2b1c4342e110_91 );
and  ( new_n28769_, new_n19044_, RI2b1c4342e098_90 );
or   ( new_n28770_, new_n28769_, new_n28768_ );
or   ( new_n28771_, new_n28770_, new_n18977_ );
and  ( new_n28772_, new_n28771_, new_n28767_ );
or   ( new_n28773_, new_n28772_, new_n28763_ );
and  ( new_n28774_, new_n28773_, new_n28762_ );
nor  ( new_n28775_, new_n22333_, new_n121_ );
nor  ( new_n28776_, new_n28775_, new_n13668_ );
or   ( new_n28777_, new_n28776_, new_n21261_ );
and  ( new_n28778_, new_n22337_, RI2b1c4342dd50_83 );
and  ( new_n28779_, new_n22330_, RI2b1c4342dcd8_82 );
or   ( new_n28780_, new_n28779_, new_n28778_ );
or   ( new_n28781_, new_n28780_, new_n21009_ );
and  ( new_n28782_, new_n28781_, new_n28777_ );
and  ( new_n28783_, new_n28782_, new_n17142_ );
or   ( new_n28784_, new_n28782_, new_n17142_ );
or   ( new_n28785_, new_n21419_, new_n2806_ );
or   ( new_n28786_, new_n21424_, new_n2541_ );
and  ( new_n28787_, new_n28786_, new_n28785_ );
or   ( new_n28788_, new_n28787_, new_n21013_ );
and  ( new_n28789_, new_n21428_, RI2b1c4342de40_85 );
and  ( new_n28790_, new_n21415_, RI2b1c4342ddc8_84 );
or   ( new_n28791_, new_n28790_, new_n28789_ );
or   ( new_n28792_, new_n28791_, new_n21265_ );
and  ( new_n28793_, new_n28792_, new_n28788_ );
and  ( new_n28794_, new_n28793_, new_n28784_ );
or   ( new_n28795_, new_n28794_, new_n28783_ );
and  ( new_n28796_, new_n28795_, new_n28774_ );
or   ( new_n28797_, new_n28795_, new_n28774_ );
or   ( new_n28798_, new_n18388_, new_n6307_ );
or   ( new_n28799_, new_n18395_, new_n5459_ );
and  ( new_n28800_, new_n28799_, new_n28798_ );
or   ( new_n28801_, new_n28800_, new_n18066_ );
and  ( new_n28802_, new_n18397_, RI2b1c4342e200_93 );
and  ( new_n28803_, new_n18384_, RI2b1c4342e188_92 );
or   ( new_n28804_, new_n28803_, new_n28802_ );
or   ( new_n28805_, new_n28804_, new_n18309_ );
and  ( new_n28806_, new_n28805_, new_n28801_ );
or   ( new_n28807_, new_n17727_, new_n124_ );
or   ( new_n28808_, new_n17734_, new_n6321_ );
and  ( new_n28809_, new_n28808_, new_n28807_ );
or   ( new_n28810_, new_n28809_, new_n17238_ );
and  ( new_n28811_, new_n17736_, RI2b1c4342e2f0_95 );
and  ( new_n28812_, new_n17723_, RI2b1c4342e278_94 );
or   ( new_n28813_, new_n28812_, new_n28811_ );
or   ( new_n28814_, new_n28813_, new_n17650_ );
and  ( new_n28815_, new_n28814_, new_n28810_ );
or   ( new_n28816_, new_n28815_, new_n28806_ );
and  ( new_n28817_, new_n28815_, new_n28806_ );
or   ( new_n28818_, new_n17248_, new_n7274_ );
or   ( new_n28819_, new_n28818_, new_n16814_ );
and  ( new_n28820_, new_n17240_, RI2b1c4342e368_96 );
or   ( new_n28821_, new_n28820_, new_n17142_ );
and  ( new_n28822_, new_n28821_, new_n28819_ );
or   ( new_n28823_, new_n28822_, new_n28817_ );
and  ( new_n28824_, new_n28823_, new_n28816_ );
and  ( new_n28825_, new_n28824_, new_n28797_ );
or   ( new_n28826_, new_n28825_, new_n28796_ );
and  ( new_n28827_, new_n28826_, new_n28743_ );
or   ( new_n28828_, new_n28826_, new_n28743_ );
or   ( new_n28829_, new_n28455_, new_n16438_ );
or   ( new_n28830_, new_n28319_, new_n16505_ );
and  ( new_n28831_, new_n28830_, new_n28829_ );
or   ( new_n28832_, new_n28831_, new_n28460_ );
and  ( new_n28833_, new_n28456_, new_n28321_ );
or   ( new_n28834_, new_n28833_, new_n28330_ );
and  ( new_n28835_, new_n28834_, new_n28832_ );
and  ( new_n28836_, new_n28835_, new_n28828_ );
or   ( new_n28837_, new_n28836_, new_n28827_ );
or   ( new_n28838_, new_n28701_, new_n28599_ );
or   ( new_n28839_, new_n28698_, new_n28606_ );
and  ( new_n28840_, new_n28839_, new_n28838_ );
or   ( new_n28841_, new_n28840_, new_n28706_ );
and  ( new_n28842_, new_n28702_, new_n28607_ );
or   ( new_n28843_, new_n28842_, new_n28615_ );
and  ( new_n28844_, new_n28843_, new_n28841_ );
or   ( new_n28845_, new_n28684_, new_n28540_ );
or   ( new_n28846_, new_n28671_, new_n28571_ );
and  ( new_n28847_, new_n28846_, new_n28845_ );
or   ( new_n28848_, new_n28847_, new_n28693_ );
and  ( new_n28849_, new_n28685_, new_n28572_ );
or   ( new_n28850_, new_n28849_, new_n28592_ );
and  ( new_n28851_, new_n28850_, new_n28848_ );
or   ( new_n28852_, new_n28851_, new_n28844_ );
and  ( new_n28853_, new_n28852_, new_n28837_ );
or   ( new_n28854_, new_n28452_, new_n28332_ );
or   ( new_n28855_, new_n28462_, new_n28311_ );
and  ( new_n28856_, new_n28855_, new_n28854_ );
or   ( new_n28857_, new_n28856_, new_n28477_ );
and  ( new_n28858_, new_n28463_, new_n28334_ );
or   ( new_n28859_, new_n28858_, new_n28365_ );
and  ( new_n28860_, new_n28859_, new_n28857_ );
or   ( new_n28861_, new_n28852_, new_n28837_ );
and  ( new_n28862_, new_n28861_, new_n28860_ );
or   ( new_n28863_, new_n28862_, new_n28853_ );
or   ( new_n28864_, new_n28863_, new_n28722_ );
or   ( new_n28865_, new_n28645_, new_n28491_ );
or   ( new_n28866_, new_n28643_, new_n28387_ );
and  ( new_n28867_, new_n28866_, new_n28865_ );
or   ( new_n28868_, new_n28411_, new_n28408_ );
and  ( new_n28869_, new_n28868_, new_n28230_ );
or   ( new_n28870_, new_n28869_, new_n28639_ );
and  ( new_n28871_, new_n28715_, new_n28657_ );
or   ( new_n28872_, new_n28871_, new_n28654_ );
and  ( new_n28873_, new_n28872_, new_n28719_ );
or   ( new_n28874_, new_n28873_, new_n28503_ );
and  ( new_n28875_, new_n28874_, new_n28870_ );
or   ( new_n28876_, new_n28875_, new_n28867_ );
or   ( new_n28877_, new_n28873_, new_n28869_ );
and  ( new_n28878_, new_n28877_, new_n28640_ );
or   ( new_n28879_, new_n28878_, new_n28647_ );
and  ( new_n28880_, new_n28879_, new_n28876_ );
and  ( new_n28881_, new_n28880_, new_n28864_ );
or   ( new_n28882_, new_n28881_, new_n28651_ );
or   ( new_n28883_, new_n28708_, new_n28594_ );
or   ( new_n28884_, new_n28695_, new_n28617_ );
and  ( new_n28885_, new_n28884_, new_n28883_ );
or   ( new_n28886_, new_n28885_, new_n28713_ );
and  ( new_n28887_, new_n28709_, new_n28618_ );
or   ( new_n28888_, new_n28887_, new_n28626_ );
and  ( new_n28889_, new_n28888_, new_n28886_ );
or   ( new_n28890_, new_n28858_, new_n28477_ );
or   ( new_n28891_, new_n28856_, new_n28365_ );
and  ( new_n28892_, new_n28891_, new_n28890_ );
or   ( new_n28893_, new_n28842_, new_n28706_ );
or   ( new_n28894_, new_n28840_, new_n28615_ );
and  ( new_n28895_, new_n28894_, new_n28893_ );
or   ( new_n28896_, new_n28849_, new_n28693_ );
or   ( new_n28897_, new_n28847_, new_n28592_ );
and  ( new_n28898_, new_n28897_, new_n28896_ );
and  ( new_n28899_, new_n28898_, new_n28895_ );
or   ( new_n28900_, new_n28692_, new_n28689_ );
and  ( new_n28901_, new_n28900_, new_n28592_ );
or   ( new_n28902_, new_n28730_, new_n28682_ );
or   ( new_n28903_, new_n28728_, new_n28569_ );
and  ( new_n28904_, new_n28903_, new_n28902_ );
or   ( new_n28905_, new_n28904_, new_n28901_ );
and  ( new_n28906_, new_n28904_, new_n28901_ );
or   ( new_n28907_, new_n28739_, new_n28669_ );
or   ( new_n28908_, new_n28737_, new_n28538_ );
and  ( new_n28909_, new_n28908_, new_n28907_ );
or   ( new_n28910_, new_n28909_, new_n28906_ );
and  ( new_n28911_, new_n28910_, new_n28905_ );
or   ( new_n28912_, new_n28759_, new_n19394_ );
or   ( new_n28913_, new_n28755_, new_n19659_ );
and  ( new_n28914_, new_n28913_, new_n28912_ );
or   ( new_n28915_, new_n28750_, new_n20156_ );
or   ( new_n28916_, new_n28746_, new_n20443_ );
and  ( new_n28917_, new_n28916_, new_n28915_ );
or   ( new_n28918_, new_n28917_, new_n28914_ );
and  ( new_n28919_, new_n28917_, new_n28914_ );
or   ( new_n28920_, new_n28770_, new_n18742_ );
or   ( new_n28921_, new_n28766_, new_n18977_ );
and  ( new_n28922_, new_n28921_, new_n28920_ );
or   ( new_n28923_, new_n28922_, new_n28919_ );
and  ( new_n28924_, new_n28923_, new_n28918_ );
or   ( new_n28925_, new_n28780_, new_n21261_ );
or   ( new_n28926_, new_n28776_, new_n21009_ );
and  ( new_n28927_, new_n28926_, new_n28925_ );
or   ( new_n28928_, new_n28927_, new_n16814_ );
and  ( new_n28929_, new_n28927_, new_n16814_ );
or   ( new_n28930_, new_n28791_, new_n21013_ );
or   ( new_n28931_, new_n28787_, new_n21265_ );
and  ( new_n28932_, new_n28931_, new_n28930_ );
or   ( new_n28933_, new_n28932_, new_n28929_ );
and  ( new_n28934_, new_n28933_, new_n28928_ );
or   ( new_n28935_, new_n28934_, new_n28924_ );
and  ( new_n28936_, new_n28934_, new_n28924_ );
or   ( new_n28937_, new_n28804_, new_n18066_ );
or   ( new_n28938_, new_n28800_, new_n18309_ );
and  ( new_n28939_, new_n28938_, new_n28937_ );
or   ( new_n28940_, new_n28813_, new_n17238_ );
or   ( new_n28941_, new_n28809_, new_n17650_ );
and  ( new_n28942_, new_n28941_, new_n28940_ );
or   ( new_n28943_, new_n28942_, new_n28939_ );
and  ( new_n28944_, new_n28942_, new_n28939_ );
or   ( new_n28945_, new_n28820_, new_n16814_ );
or   ( new_n28946_, new_n28818_, new_n17142_ );
and  ( new_n28947_, new_n28946_, new_n28945_ );
or   ( new_n28948_, new_n28947_, new_n28944_ );
and  ( new_n28949_, new_n28948_, new_n28943_ );
or   ( new_n28950_, new_n28949_, new_n28936_ );
and  ( new_n28951_, new_n28950_, new_n28935_ );
or   ( new_n28952_, new_n28951_, new_n28911_ );
and  ( new_n28953_, new_n28951_, new_n28911_ );
or   ( new_n28954_, new_n28833_, new_n28460_ );
or   ( new_n28955_, new_n28831_, new_n28330_ );
and  ( new_n28956_, new_n28955_, new_n28954_ );
or   ( new_n28957_, new_n28956_, new_n28953_ );
and  ( new_n28958_, new_n28957_, new_n28952_ );
or   ( new_n28959_, new_n28958_, new_n28899_ );
and  ( new_n28960_, new_n28959_, new_n28861_ );
or   ( new_n28961_, new_n28960_, new_n28892_ );
or   ( new_n28962_, new_n28899_, new_n28837_ );
or   ( new_n28963_, new_n28958_, new_n28852_ );
and  ( new_n28964_, new_n28963_, new_n28962_ );
or   ( new_n28965_, new_n28964_, new_n28860_ );
and  ( new_n28966_, new_n28965_, new_n28961_ );
or   ( new_n28967_, new_n28966_, new_n28889_ );
or   ( new_n28968_, new_n28964_, new_n28892_ );
or   ( new_n28969_, new_n28960_, new_n28860_ );
and  ( new_n28970_, new_n28969_, new_n28968_ );
or   ( new_n28971_, new_n28887_, new_n28713_ );
or   ( new_n28972_, new_n28885_, new_n28626_ );
and  ( new_n28973_, new_n28972_, new_n28971_ );
or   ( new_n28974_, new_n28973_, new_n28970_ );
and  ( new_n28975_, new_n28974_, new_n28967_ );
or   ( new_n28976_, new_n28898_, new_n28844_ );
or   ( new_n28977_, new_n28895_, new_n28851_ );
and  ( new_n28978_, new_n28977_, new_n28976_ );
or   ( new_n28979_, new_n28914_, new_n28752_ );
or   ( new_n28980_, new_n28917_, new_n28761_ );
and  ( new_n28981_, new_n28980_, new_n28979_ );
or   ( new_n28982_, new_n28981_, new_n28922_ );
and  ( new_n28983_, new_n28918_, new_n28762_ );
or   ( new_n28984_, new_n28983_, new_n28772_ );
and  ( new_n28985_, new_n28984_, new_n28982_ );
or   ( new_n28986_, new_n28927_, new_n17142_ );
or   ( new_n28987_, new_n28782_, new_n16814_ );
and  ( new_n28988_, new_n28987_, new_n28986_ );
or   ( new_n28989_, new_n28988_, new_n28932_ );
and  ( new_n28990_, new_n28928_, new_n28784_ );
or   ( new_n28991_, new_n28990_, new_n28793_ );
and  ( new_n28992_, new_n28991_, new_n28989_ );
or   ( new_n28993_, new_n28992_, new_n28985_ );
nor  ( new_n28994_, new_n22333_, new_n2541_ );
nor  ( new_n28995_, new_n28994_, new_n13857_ );
or   ( new_n28996_, new_n28995_, new_n21261_ );
and  ( new_n28997_, new_n22337_, RI2b1c4342ddc8_84 );
and  ( new_n28998_, new_n22330_, RI2b1c4342dd50_83 );
or   ( new_n28999_, new_n28998_, new_n28997_ );
or   ( new_n29000_, new_n28999_, new_n21009_ );
and  ( new_n29001_, new_n29000_, new_n28996_ );
or   ( new_n29002_, new_n21419_, new_n3239_ );
or   ( new_n29003_, new_n21424_, new_n2806_ );
and  ( new_n29004_, new_n29003_, new_n29002_ );
or   ( new_n29005_, new_n29004_, new_n21013_ );
and  ( new_n29006_, new_n21428_, RI2b1c4342deb8_86 );
and  ( new_n29007_, new_n21415_, RI2b1c4342de40_85 );
or   ( new_n29008_, new_n29007_, new_n29006_ );
or   ( new_n29009_, new_n29008_, new_n21265_ );
and  ( new_n29010_, new_n29009_, new_n29005_ );
or   ( new_n29011_, new_n29010_, new_n29001_ );
and  ( new_n29012_, new_n29010_, new_n29001_ );
or   ( new_n29013_, new_n20557_, new_n3902_ );
or   ( new_n29014_, new_n20562_, new_n3924_ );
and  ( new_n29015_, new_n29014_, new_n29013_ );
or   ( new_n29016_, new_n29015_, new_n20156_ );
and  ( new_n29017_, new_n20566_, RI2b1c4342dfa8_88 );
and  ( new_n29018_, new_n20553_, RI2b1c4342df30_87 );
or   ( new_n29019_, new_n29018_, new_n29017_ );
or   ( new_n29020_, new_n29019_, new_n20443_ );
and  ( new_n29021_, new_n29020_, new_n29016_ );
or   ( new_n29022_, new_n29021_, new_n29012_ );
and  ( new_n29023_, new_n29022_, new_n29011_ );
or   ( new_n29024_, new_n19758_, new_n4635_ );
or   ( new_n29025_, new_n19763_, new_n132_ );
and  ( new_n29026_, new_n29025_, new_n29024_ );
or   ( new_n29027_, new_n29026_, new_n19394_ );
and  ( new_n29028_, new_n19767_, RI2b1c4342e098_90 );
and  ( new_n29029_, new_n19754_, RI2b1c4342e020_89 );
or   ( new_n29030_, new_n29029_, new_n29028_ );
or   ( new_n29031_, new_n29030_, new_n19659_ );
and  ( new_n29032_, new_n29031_, new_n29027_ );
or   ( new_n29033_, new_n19048_, new_n5459_ );
or   ( new_n29034_, new_n19055_, new_n117_ );
and  ( new_n29035_, new_n29034_, new_n29033_ );
or   ( new_n29036_, new_n29035_, new_n18742_ );
and  ( new_n29037_, new_n19057_, RI2b1c4342e188_92 );
and  ( new_n29038_, new_n19044_, RI2b1c4342e110_91 );
or   ( new_n29039_, new_n29038_, new_n29037_ );
or   ( new_n29040_, new_n29039_, new_n18977_ );
and  ( new_n29041_, new_n29040_, new_n29036_ );
or   ( new_n29042_, new_n29041_, new_n29032_ );
and  ( new_n29043_, new_n29041_, new_n29032_ );
or   ( new_n29044_, new_n18388_, new_n6321_ );
or   ( new_n29045_, new_n18395_, new_n6307_ );
and  ( new_n29046_, new_n29045_, new_n29044_ );
or   ( new_n29047_, new_n29046_, new_n18066_ );
and  ( new_n29048_, new_n18397_, RI2b1c4342e278_94 );
and  ( new_n29049_, new_n18384_, RI2b1c4342e200_93 );
or   ( new_n29050_, new_n29049_, new_n29048_ );
or   ( new_n29051_, new_n29050_, new_n18309_ );
and  ( new_n29052_, new_n29051_, new_n29047_ );
or   ( new_n29053_, new_n29052_, new_n29043_ );
and  ( new_n29054_, new_n29053_, new_n29042_ );
or   ( new_n29055_, new_n29054_, new_n29023_ );
and  ( new_n29056_, new_n29054_, new_n29023_ );
or   ( new_n29057_, new_n28942_, new_n28806_ );
or   ( new_n29058_, new_n28939_, new_n28815_ );
and  ( new_n29059_, new_n29058_, new_n29057_ );
or   ( new_n29060_, new_n29059_, new_n28947_ );
and  ( new_n29061_, new_n28943_, new_n28816_ );
or   ( new_n29062_, new_n29061_, new_n28822_ );
and  ( new_n29063_, new_n29062_, new_n29060_ );
or   ( new_n29064_, new_n29063_, new_n29056_ );
and  ( new_n29065_, new_n29064_, new_n29055_ );
or   ( new_n29066_, new_n29065_, new_n28993_ );
and  ( new_n29067_, new_n29065_, new_n28993_ );
or   ( new_n29068_, new_n28904_, new_n28725_ );
or   ( new_n29069_, new_n28901_, new_n28732_ );
and  ( new_n29070_, new_n29069_, new_n29068_ );
or   ( new_n29071_, new_n29070_, new_n28909_ );
and  ( new_n29072_, new_n28905_, new_n28733_ );
or   ( new_n29073_, new_n29072_, new_n28741_ );
and  ( new_n29074_, new_n29073_, new_n29071_ );
or   ( new_n29075_, new_n29074_, new_n29067_ );
and  ( new_n29076_, new_n29075_, new_n29066_ );
or   ( new_n29077_, new_n29076_, new_n28978_ );
or   ( new_n29078_, new_n28911_, new_n28826_ );
or   ( new_n29079_, new_n28951_, new_n28743_ );
and  ( new_n29080_, new_n29079_, new_n29078_ );
or   ( new_n29081_, new_n29080_, new_n28956_ );
and  ( new_n29082_, new_n28952_, new_n28828_ );
or   ( new_n29083_, new_n29082_, new_n28835_ );
and  ( new_n29084_, new_n29083_, new_n29081_ );
and  ( new_n29085_, new_n29076_, new_n28978_ );
or   ( new_n29086_, new_n29085_, new_n29084_ );
and  ( new_n29087_, new_n29086_, new_n29077_ );
and  ( new_n29088_, new_n29087_, new_n28975_ );
or   ( new_n29089_, new_n28970_, new_n28889_ );
or   ( new_n29090_, new_n28720_, new_n28654_ );
or   ( new_n29091_, new_n28717_, new_n28637_ );
and  ( new_n29092_, new_n29091_, new_n29090_ );
or   ( new_n29093_, new_n29092_, new_n28863_ );
and  ( new_n29094_, new_n28958_, new_n28899_ );
or   ( new_n29095_, new_n29094_, new_n28892_ );
and  ( new_n29096_, new_n29095_, new_n28959_ );
or   ( new_n29097_, new_n29096_, new_n28722_ );
and  ( new_n29098_, new_n29097_, new_n29093_ );
and  ( new_n29099_, new_n29098_, new_n29089_ );
or   ( new_n29100_, new_n29099_, new_n29088_ );
or   ( new_n29101_, new_n29082_, new_n28956_ );
or   ( new_n29102_, new_n29080_, new_n28835_ );
and  ( new_n29103_, new_n29102_, new_n29101_ );
or   ( new_n29104_, new_n28898_, new_n28895_ );
and  ( new_n29105_, new_n29104_, new_n28852_ );
or   ( new_n29106_, new_n29105_, new_n29076_ );
or   ( new_n29107_, new_n28990_, new_n28932_ );
or   ( new_n29108_, new_n28988_, new_n28793_ );
and  ( new_n29109_, new_n29108_, new_n29107_ );
or   ( new_n29110_, new_n28983_, new_n28922_ );
or   ( new_n29111_, new_n28981_, new_n28772_ );
and  ( new_n29112_, new_n29111_, new_n29110_ );
and  ( new_n29113_, new_n29112_, new_n29109_ );
or   ( new_n29114_, new_n28999_, new_n21261_ );
or   ( new_n29115_, new_n28995_, new_n21009_ );
and  ( new_n29116_, new_n29115_, new_n29114_ );
or   ( new_n29117_, new_n29008_, new_n21013_ );
or   ( new_n29118_, new_n29004_, new_n21265_ );
and  ( new_n29119_, new_n29118_, new_n29117_ );
or   ( new_n29120_, new_n29119_, new_n29116_ );
and  ( new_n29121_, new_n29119_, new_n29116_ );
or   ( new_n29122_, new_n29019_, new_n20156_ );
or   ( new_n29123_, new_n29015_, new_n20443_ );
and  ( new_n29124_, new_n29123_, new_n29122_ );
or   ( new_n29125_, new_n29124_, new_n29121_ );
and  ( new_n29126_, new_n29125_, new_n29120_ );
or   ( new_n29127_, new_n29030_, new_n19394_ );
or   ( new_n29128_, new_n29026_, new_n19659_ );
and  ( new_n29129_, new_n29128_, new_n29127_ );
or   ( new_n29130_, new_n29039_, new_n18742_ );
or   ( new_n29131_, new_n29035_, new_n18977_ );
and  ( new_n29132_, new_n29131_, new_n29130_ );
or   ( new_n29133_, new_n29132_, new_n29129_ );
and  ( new_n29134_, new_n29132_, new_n29129_ );
or   ( new_n29135_, new_n29050_, new_n18066_ );
or   ( new_n29136_, new_n29046_, new_n18309_ );
and  ( new_n29137_, new_n29136_, new_n29135_ );
or   ( new_n29138_, new_n29137_, new_n29134_ );
and  ( new_n29139_, new_n29138_, new_n29133_ );
or   ( new_n29140_, new_n29139_, new_n29126_ );
and  ( new_n29141_, new_n29139_, new_n29126_ );
or   ( new_n29142_, new_n29061_, new_n28947_ );
or   ( new_n29143_, new_n29059_, new_n28822_ );
and  ( new_n29144_, new_n29143_, new_n29142_ );
or   ( new_n29145_, new_n29144_, new_n29141_ );
and  ( new_n29146_, new_n29145_, new_n29140_ );
or   ( new_n29147_, new_n29146_, new_n29113_ );
and  ( new_n29148_, new_n29146_, new_n29113_ );
or   ( new_n29149_, new_n29072_, new_n28909_ );
or   ( new_n29150_, new_n29070_, new_n28741_ );
and  ( new_n29151_, new_n29150_, new_n29149_ );
or   ( new_n29152_, new_n29151_, new_n29148_ );
and  ( new_n29153_, new_n29152_, new_n29147_ );
or   ( new_n29154_, new_n29153_, new_n28978_ );
and  ( new_n29155_, new_n29154_, new_n29106_ );
or   ( new_n29156_, new_n29155_, new_n29103_ );
or   ( new_n29157_, new_n29153_, new_n29105_ );
and  ( new_n29158_, new_n29157_, new_n29077_ );
or   ( new_n29159_, new_n29158_, new_n29084_ );
and  ( new_n29160_, new_n29159_, new_n29156_ );
or   ( new_n29161_, new_n28924_, new_n28795_ );
or   ( new_n29162_, new_n28934_, new_n28774_ );
and  ( new_n29163_, new_n29162_, new_n29161_ );
or   ( new_n29164_, new_n29163_, new_n28949_ );
and  ( new_n29165_, new_n28935_, new_n28797_ );
or   ( new_n29166_, new_n29165_, new_n28824_ );
and  ( new_n29167_, new_n29166_, new_n29164_ );
or   ( new_n29168_, new_n29109_, new_n28985_ );
or   ( new_n29169_, new_n29112_, new_n28992_ );
and  ( new_n29170_, new_n29169_, new_n29168_ );
or   ( new_n29171_, new_n20557_, new_n132_ );
or   ( new_n29172_, new_n20562_, new_n3902_ );
and  ( new_n29173_, new_n29172_, new_n29171_ );
or   ( new_n29174_, new_n29173_, new_n20156_ );
and  ( new_n29175_, new_n20566_, RI2b1c4342e020_89 );
and  ( new_n29176_, new_n20553_, RI2b1c4342dfa8_88 );
or   ( new_n29177_, new_n29176_, new_n29175_ );
or   ( new_n29178_, new_n29177_, new_n20443_ );
and  ( new_n29179_, new_n29178_, new_n29174_ );
or   ( new_n29180_, new_n19758_, new_n117_ );
or   ( new_n29181_, new_n19763_, new_n4635_ );
and  ( new_n29182_, new_n29181_, new_n29180_ );
or   ( new_n29183_, new_n29182_, new_n19394_ );
and  ( new_n29184_, new_n19767_, RI2b1c4342e110_91 );
and  ( new_n29185_, new_n19754_, RI2b1c4342e098_90 );
or   ( new_n29186_, new_n29185_, new_n29184_ );
or   ( new_n29187_, new_n29186_, new_n19659_ );
and  ( new_n29188_, new_n29187_, new_n29183_ );
or   ( new_n29189_, new_n29188_, new_n29179_ );
and  ( new_n29190_, new_n29188_, new_n29179_ );
or   ( new_n29191_, new_n19048_, new_n6307_ );
or   ( new_n29192_, new_n19055_, new_n5459_ );
and  ( new_n29193_, new_n29192_, new_n29191_ );
or   ( new_n29194_, new_n29193_, new_n18742_ );
and  ( new_n29195_, new_n19057_, RI2b1c4342e200_93 );
and  ( new_n29196_, new_n19044_, RI2b1c4342e188_92 );
or   ( new_n29197_, new_n29196_, new_n29195_ );
or   ( new_n29198_, new_n29197_, new_n18977_ );
and  ( new_n29199_, new_n29198_, new_n29194_ );
or   ( new_n29200_, new_n29199_, new_n29190_ );
and  ( new_n29201_, new_n29200_, new_n29189_ );
nor  ( new_n29202_, new_n22333_, new_n2806_ );
nor  ( new_n29203_, new_n29202_, new_n14066_ );
or   ( new_n29204_, new_n29203_, new_n21261_ );
and  ( new_n29205_, new_n22337_, RI2b1c4342de40_85 );
and  ( new_n29206_, new_n22330_, RI2b1c4342ddc8_84 );
or   ( new_n29207_, new_n29206_, new_n29205_ );
or   ( new_n29208_, new_n29207_, new_n21009_ );
and  ( new_n29209_, new_n29208_, new_n29204_ );
and  ( new_n29210_, new_n29209_, new_n17650_ );
or   ( new_n29211_, new_n29209_, new_n17650_ );
or   ( new_n29212_, new_n21419_, new_n3924_ );
or   ( new_n29213_, new_n21424_, new_n3239_ );
and  ( new_n29214_, new_n29213_, new_n29212_ );
or   ( new_n29215_, new_n29214_, new_n21013_ );
and  ( new_n29216_, new_n21428_, RI2b1c4342df30_87 );
and  ( new_n29217_, new_n21415_, RI2b1c4342deb8_86 );
or   ( new_n29218_, new_n29217_, new_n29216_ );
or   ( new_n29219_, new_n29218_, new_n21265_ );
and  ( new_n29220_, new_n29219_, new_n29215_ );
and  ( new_n29221_, new_n29220_, new_n29211_ );
or   ( new_n29222_, new_n29221_, new_n29210_ );
and  ( new_n29223_, new_n29222_, new_n29201_ );
or   ( new_n29224_, new_n29222_, new_n29201_ );
or   ( new_n29225_, new_n17727_, new_n7274_ );
or   ( new_n29226_, new_n17734_, new_n124_ );
and  ( new_n29227_, new_n29226_, new_n29225_ );
or   ( new_n29228_, new_n29227_, new_n17238_ );
and  ( new_n29229_, new_n17736_, RI2b1c4342e368_96 );
and  ( new_n29230_, new_n17723_, RI2b1c4342e2f0_95 );
or   ( new_n29231_, new_n29230_, new_n29229_ );
or   ( new_n29232_, new_n29231_, new_n17650_ );
and  ( new_n29233_, new_n29232_, new_n29228_ );
and  ( new_n29234_, new_n29233_, new_n29224_ );
or   ( new_n29235_, new_n29234_, new_n29223_ );
and  ( new_n29236_, new_n29235_, new_n29170_ );
or   ( new_n29237_, new_n29235_, new_n29170_ );
or   ( new_n29238_, new_n29139_, new_n29023_ );
or   ( new_n29239_, new_n29126_, new_n29054_ );
and  ( new_n29240_, new_n29239_, new_n29238_ );
or   ( new_n29241_, new_n29240_, new_n29144_ );
and  ( new_n29242_, new_n29140_, new_n29055_ );
or   ( new_n29243_, new_n29242_, new_n29063_ );
and  ( new_n29244_, new_n29243_, new_n29241_ );
and  ( new_n29245_, new_n29244_, new_n29237_ );
or   ( new_n29246_, new_n29245_, new_n29236_ );
and  ( new_n29247_, new_n29246_, new_n29167_ );
or   ( new_n29248_, new_n29246_, new_n29167_ );
or   ( new_n29249_, new_n29113_, new_n29065_ );
or   ( new_n29250_, new_n29146_, new_n28993_ );
and  ( new_n29251_, new_n29250_, new_n29249_ );
or   ( new_n29252_, new_n29251_, new_n29151_ );
and  ( new_n29253_, new_n29147_, new_n29066_ );
or   ( new_n29254_, new_n29253_, new_n29074_ );
and  ( new_n29255_, new_n29254_, new_n29252_ );
and  ( new_n29256_, new_n29255_, new_n29248_ );
or   ( new_n29257_, new_n29256_, new_n29247_ );
and  ( new_n29258_, new_n29257_, new_n29160_ );
or   ( new_n29259_, new_n29253_, new_n29151_ );
or   ( new_n29260_, new_n29251_, new_n29074_ );
and  ( new_n29261_, new_n29260_, new_n29259_ );
or   ( new_n29262_, new_n29165_, new_n28949_ );
or   ( new_n29263_, new_n29163_, new_n28824_ );
and  ( new_n29264_, new_n29263_, new_n29262_ );
or   ( new_n29265_, new_n29264_, new_n29246_ );
or   ( new_n29266_, new_n29112_, new_n29109_ );
and  ( new_n29267_, new_n29266_, new_n28993_ );
or   ( new_n29268_, new_n29177_, new_n20156_ );
or   ( new_n29269_, new_n29173_, new_n20443_ );
and  ( new_n29270_, new_n29269_, new_n29268_ );
or   ( new_n29271_, new_n29186_, new_n19394_ );
or   ( new_n29272_, new_n29182_, new_n19659_ );
and  ( new_n29273_, new_n29272_, new_n29271_ );
or   ( new_n29274_, new_n29273_, new_n29270_ );
and  ( new_n29275_, new_n29273_, new_n29270_ );
or   ( new_n29276_, new_n29197_, new_n18742_ );
or   ( new_n29277_, new_n29193_, new_n18977_ );
and  ( new_n29278_, new_n29277_, new_n29276_ );
or   ( new_n29279_, new_n29278_, new_n29275_ );
and  ( new_n29280_, new_n29279_, new_n29274_ );
or   ( new_n29281_, new_n29207_, new_n21261_ );
or   ( new_n29282_, new_n29203_, new_n21009_ );
and  ( new_n29283_, new_n29282_, new_n29281_ );
or   ( new_n29284_, new_n29283_, new_n17238_ );
and  ( new_n29285_, new_n29283_, new_n17238_ );
or   ( new_n29286_, new_n29218_, new_n21013_ );
or   ( new_n29287_, new_n29214_, new_n21265_ );
and  ( new_n29288_, new_n29287_, new_n29286_ );
or   ( new_n29289_, new_n29288_, new_n29285_ );
and  ( new_n29290_, new_n29289_, new_n29284_ );
or   ( new_n29291_, new_n29290_, new_n29280_ );
and  ( new_n29292_, new_n29290_, new_n29280_ );
or   ( new_n29293_, new_n29231_, new_n17238_ );
or   ( new_n29294_, new_n29227_, new_n17650_ );
and  ( new_n29295_, new_n29294_, new_n29293_ );
or   ( new_n29296_, new_n29295_, new_n29292_ );
and  ( new_n29297_, new_n29296_, new_n29291_ );
or   ( new_n29298_, new_n29297_, new_n29267_ );
and  ( new_n29299_, new_n29297_, new_n29267_ );
or   ( new_n29300_, new_n29242_, new_n29144_ );
or   ( new_n29301_, new_n29240_, new_n29063_ );
and  ( new_n29302_, new_n29301_, new_n29300_ );
or   ( new_n29303_, new_n29302_, new_n29299_ );
and  ( new_n29304_, new_n29303_, new_n29298_ );
or   ( new_n29305_, new_n29304_, new_n29167_ );
and  ( new_n29306_, new_n29305_, new_n29265_ );
or   ( new_n29307_, new_n29306_, new_n29261_ );
or   ( new_n29308_, new_n29304_, new_n29264_ );
and  ( new_n29309_, new_n29308_, new_n29248_ );
or   ( new_n29310_, new_n29309_, new_n29255_ );
and  ( new_n29311_, new_n29310_, new_n29307_ );
or   ( new_n29312_, new_n29119_, new_n29001_ );
or   ( new_n29313_, new_n29116_, new_n29010_ );
and  ( new_n29314_, new_n29313_, new_n29312_ );
or   ( new_n29315_, new_n29314_, new_n29124_ );
and  ( new_n29316_, new_n29120_, new_n29011_ );
or   ( new_n29317_, new_n29316_, new_n29021_ );
and  ( new_n29318_, new_n29317_, new_n29315_ );
or   ( new_n29319_, new_n29280_, new_n29222_ );
or   ( new_n29320_, new_n29290_, new_n29201_ );
and  ( new_n29321_, new_n29320_, new_n29319_ );
or   ( new_n29322_, new_n29321_, new_n29295_ );
and  ( new_n29323_, new_n29291_, new_n29224_ );
or   ( new_n29324_, new_n29323_, new_n29233_ );
and  ( new_n29325_, new_n29324_, new_n29322_ );
or   ( new_n29326_, new_n29325_, new_n29318_ );
nor  ( new_n29327_, new_n22333_, new_n3239_ );
nor  ( new_n29328_, new_n29327_, new_n14193_ );
or   ( new_n29329_, new_n29328_, new_n21261_ );
and  ( new_n29330_, new_n22337_, RI2b1c4342deb8_86 );
and  ( new_n29331_, new_n22330_, RI2b1c4342de40_85 );
or   ( new_n29332_, new_n29331_, new_n29330_ );
or   ( new_n29333_, new_n29332_, new_n21009_ );
and  ( new_n29334_, new_n29333_, new_n29329_ );
or   ( new_n29335_, new_n21419_, new_n3902_ );
or   ( new_n29336_, new_n21424_, new_n3924_ );
and  ( new_n29337_, new_n29336_, new_n29335_ );
or   ( new_n29338_, new_n29337_, new_n21013_ );
and  ( new_n29339_, new_n21428_, RI2b1c4342dfa8_88 );
and  ( new_n29340_, new_n21415_, RI2b1c4342df30_87 );
or   ( new_n29341_, new_n29340_, new_n29339_ );
or   ( new_n29342_, new_n29341_, new_n21265_ );
and  ( new_n29343_, new_n29342_, new_n29338_ );
or   ( new_n29344_, new_n29343_, new_n29334_ );
and  ( new_n29345_, new_n29343_, new_n29334_ );
or   ( new_n29346_, new_n20557_, new_n4635_ );
or   ( new_n29347_, new_n20562_, new_n132_ );
and  ( new_n29348_, new_n29347_, new_n29346_ );
or   ( new_n29349_, new_n29348_, new_n20156_ );
and  ( new_n29350_, new_n20566_, RI2b1c4342e098_90 );
and  ( new_n29351_, new_n20553_, RI2b1c4342e020_89 );
or   ( new_n29352_, new_n29351_, new_n29350_ );
or   ( new_n29353_, new_n29352_, new_n20443_ );
and  ( new_n29354_, new_n29353_, new_n29349_ );
or   ( new_n29355_, new_n29354_, new_n29345_ );
and  ( new_n29356_, new_n29355_, new_n29344_ );
or   ( new_n29357_, new_n19758_, new_n5459_ );
or   ( new_n29358_, new_n19763_, new_n117_ );
and  ( new_n29359_, new_n29358_, new_n29357_ );
or   ( new_n29360_, new_n29359_, new_n19394_ );
and  ( new_n29361_, new_n19767_, RI2b1c4342e188_92 );
and  ( new_n29362_, new_n19754_, RI2b1c4342e110_91 );
or   ( new_n29363_, new_n29362_, new_n29361_ );
or   ( new_n29364_, new_n29363_, new_n19659_ );
and  ( new_n29365_, new_n29364_, new_n29360_ );
or   ( new_n29366_, new_n19048_, new_n6321_ );
or   ( new_n29367_, new_n19055_, new_n6307_ );
and  ( new_n29368_, new_n29367_, new_n29366_ );
or   ( new_n29369_, new_n29368_, new_n18742_ );
and  ( new_n29370_, new_n19057_, RI2b1c4342e278_94 );
and  ( new_n29371_, new_n19044_, RI2b1c4342e200_93 );
or   ( new_n29372_, new_n29371_, new_n29370_ );
or   ( new_n29373_, new_n29372_, new_n18977_ );
and  ( new_n29374_, new_n29373_, new_n29369_ );
or   ( new_n29375_, new_n29374_, new_n29365_ );
and  ( new_n29376_, new_n29374_, new_n29365_ );
or   ( new_n29377_, new_n18388_, new_n7274_ );
or   ( new_n29378_, new_n18395_, new_n124_ );
and  ( new_n29379_, new_n29378_, new_n29377_ );
or   ( new_n29380_, new_n29379_, new_n18066_ );
and  ( new_n29381_, new_n18397_, RI2b1c4342e368_96 );
and  ( new_n29382_, new_n18384_, RI2b1c4342e2f0_95 );
or   ( new_n29383_, new_n29382_, new_n29381_ );
or   ( new_n29384_, new_n29383_, new_n18309_ );
and  ( new_n29385_, new_n29384_, new_n29380_ );
or   ( new_n29386_, new_n29385_, new_n29376_ );
and  ( new_n29387_, new_n29386_, new_n29375_ );
or   ( new_n29388_, new_n29387_, new_n29356_ );
and  ( new_n29389_, new_n29387_, new_n29356_ );
or   ( new_n29390_, new_n18388_, new_n124_ );
or   ( new_n29391_, new_n18395_, new_n6321_ );
and  ( new_n29392_, new_n29391_, new_n29390_ );
or   ( new_n29393_, new_n29392_, new_n18066_ );
and  ( new_n29394_, new_n18397_, RI2b1c4342e2f0_95 );
and  ( new_n29395_, new_n18384_, RI2b1c4342e278_94 );
or   ( new_n29396_, new_n29395_, new_n29394_ );
or   ( new_n29397_, new_n29396_, new_n18309_ );
and  ( new_n29398_, new_n29397_, new_n29393_ );
or   ( new_n29399_, new_n29398_, new_n29389_ );
and  ( new_n29400_, new_n29399_, new_n29388_ );
or   ( new_n29401_, new_n17734_, new_n7274_ );
or   ( new_n29402_, new_n29401_, new_n17238_ );
and  ( new_n29403_, new_n17723_, RI2b1c4342e368_96 );
or   ( new_n29404_, new_n29403_, new_n17650_ );
and  ( new_n29405_, new_n29404_, new_n29402_ );
or   ( new_n29406_, new_n29273_, new_n29179_ );
or   ( new_n29407_, new_n29270_, new_n29188_ );
and  ( new_n29408_, new_n29407_, new_n29406_ );
or   ( new_n29409_, new_n29408_, new_n29278_ );
and  ( new_n29410_, new_n29274_, new_n29189_ );
or   ( new_n29411_, new_n29410_, new_n29199_ );
and  ( new_n29412_, new_n29411_, new_n29409_ );
or   ( new_n29413_, new_n29412_, new_n29405_ );
and  ( new_n29414_, new_n29412_, new_n29405_ );
or   ( new_n29415_, new_n29283_, new_n17650_ );
or   ( new_n29416_, new_n29209_, new_n17238_ );
and  ( new_n29417_, new_n29416_, new_n29415_ );
or   ( new_n29418_, new_n29417_, new_n29288_ );
and  ( new_n29419_, new_n29284_, new_n29211_ );
or   ( new_n29420_, new_n29419_, new_n29220_ );
and  ( new_n29421_, new_n29420_, new_n29418_ );
or   ( new_n29422_, new_n29421_, new_n29414_ );
and  ( new_n29423_, new_n29422_, new_n29413_ );
or   ( new_n29424_, new_n29423_, new_n29400_ );
or   ( new_n29425_, new_n29132_, new_n29032_ );
or   ( new_n29426_, new_n29129_, new_n29041_ );
and  ( new_n29427_, new_n29426_, new_n29425_ );
or   ( new_n29428_, new_n29427_, new_n29137_ );
and  ( new_n29429_, new_n29133_, new_n29042_ );
or   ( new_n29430_, new_n29429_, new_n29052_ );
and  ( new_n29431_, new_n29430_, new_n29428_ );
and  ( new_n29432_, new_n29423_, new_n29400_ );
or   ( new_n29433_, new_n29432_, new_n29431_ );
and  ( new_n29434_, new_n29433_, new_n29424_ );
or   ( new_n29435_, new_n29434_, new_n29326_ );
or   ( new_n29436_, new_n29267_, new_n29235_ );
or   ( new_n29437_, new_n29297_, new_n29170_ );
and  ( new_n29438_, new_n29437_, new_n29436_ );
or   ( new_n29439_, new_n29438_, new_n29302_ );
and  ( new_n29440_, new_n29298_, new_n29237_ );
or   ( new_n29441_, new_n29440_, new_n29244_ );
and  ( new_n29442_, new_n29441_, new_n29439_ );
and  ( new_n29443_, new_n29434_, new_n29326_ );
or   ( new_n29444_, new_n29443_, new_n29442_ );
and  ( new_n29445_, new_n29444_, new_n29435_ );
and  ( new_n29446_, new_n29445_, new_n29311_ );
or   ( new_n29447_, new_n29446_, new_n29258_ );
or   ( new_n29448_, new_n29396_, new_n18066_ );
or   ( new_n29449_, new_n29392_, new_n18309_ );
and  ( new_n29450_, new_n29449_, new_n29448_ );
or   ( new_n29451_, new_n29332_, new_n21261_ );
or   ( new_n29452_, new_n29328_, new_n21009_ );
and  ( new_n29453_, new_n29452_, new_n29451_ );
or   ( new_n29454_, new_n29341_, new_n21013_ );
or   ( new_n29455_, new_n29337_, new_n21265_ );
and  ( new_n29456_, new_n29455_, new_n29454_ );
or   ( new_n29457_, new_n29456_, new_n29453_ );
and  ( new_n29458_, new_n29456_, new_n29453_ );
or   ( new_n29459_, new_n29352_, new_n20156_ );
or   ( new_n29460_, new_n29348_, new_n20443_ );
and  ( new_n29461_, new_n29460_, new_n29459_ );
or   ( new_n29462_, new_n29461_, new_n29458_ );
and  ( new_n29463_, new_n29462_, new_n29457_ );
or   ( new_n29464_, new_n29363_, new_n19394_ );
or   ( new_n29465_, new_n29359_, new_n19659_ );
and  ( new_n29466_, new_n29465_, new_n29464_ );
or   ( new_n29467_, new_n29372_, new_n18742_ );
or   ( new_n29468_, new_n29368_, new_n18977_ );
and  ( new_n29469_, new_n29468_, new_n29467_ );
or   ( new_n29470_, new_n29469_, new_n29466_ );
and  ( new_n29471_, new_n29469_, new_n29466_ );
or   ( new_n29472_, new_n29383_, new_n18066_ );
or   ( new_n29473_, new_n29379_, new_n18309_ );
and  ( new_n29474_, new_n29473_, new_n29472_ );
or   ( new_n29475_, new_n29474_, new_n29471_ );
and  ( new_n29476_, new_n29475_, new_n29470_ );
or   ( new_n29477_, new_n29476_, new_n29463_ );
and  ( new_n29478_, new_n29477_, new_n29388_ );
or   ( new_n29479_, new_n29478_, new_n29450_ );
or   ( new_n29480_, new_n29476_, new_n29356_ );
or   ( new_n29481_, new_n29463_, new_n29387_ );
and  ( new_n29482_, new_n29481_, new_n29480_ );
or   ( new_n29483_, new_n29482_, new_n29398_ );
and  ( new_n29484_, new_n29483_, new_n29479_ );
or   ( new_n29485_, new_n29419_, new_n29288_ );
or   ( new_n29486_, new_n29417_, new_n29220_ );
and  ( new_n29487_, new_n29486_, new_n29485_ );
or   ( new_n29488_, new_n29403_, new_n17238_ );
or   ( new_n29489_, new_n29401_, new_n17650_ );
and  ( new_n29490_, new_n29489_, new_n29488_ );
or   ( new_n29491_, new_n29410_, new_n29278_ );
or   ( new_n29492_, new_n29408_, new_n29199_ );
and  ( new_n29493_, new_n29492_, new_n29491_ );
or   ( new_n29494_, new_n29493_, new_n29490_ );
and  ( new_n29495_, new_n29494_, new_n29413_ );
or   ( new_n29496_, new_n29495_, new_n29487_ );
or   ( new_n29497_, new_n29493_, new_n29405_ );
or   ( new_n29498_, new_n29490_, new_n29412_ );
and  ( new_n29499_, new_n29498_, new_n29497_ );
or   ( new_n29500_, new_n29499_, new_n29421_ );
and  ( new_n29501_, new_n29500_, new_n29496_ );
or   ( new_n29502_, new_n20557_, new_n117_ );
or   ( new_n29503_, new_n20562_, new_n4635_ );
and  ( new_n29504_, new_n29503_, new_n29502_ );
or   ( new_n29505_, new_n29504_, new_n20156_ );
and  ( new_n29506_, new_n20566_, RI2b1c4342e110_91 );
and  ( new_n29507_, new_n20553_, RI2b1c4342e098_90 );
or   ( new_n29508_, new_n29507_, new_n29506_ );
or   ( new_n29509_, new_n29508_, new_n20443_ );
and  ( new_n29510_, new_n29509_, new_n29505_ );
or   ( new_n29511_, new_n19758_, new_n6307_ );
or   ( new_n29512_, new_n19763_, new_n5459_ );
and  ( new_n29513_, new_n29512_, new_n29511_ );
or   ( new_n29514_, new_n29513_, new_n19394_ );
and  ( new_n29515_, new_n19767_, RI2b1c4342e200_93 );
and  ( new_n29516_, new_n19754_, RI2b1c4342e188_92 );
or   ( new_n29517_, new_n29516_, new_n29515_ );
or   ( new_n29518_, new_n29517_, new_n19659_ );
and  ( new_n29519_, new_n29518_, new_n29514_ );
or   ( new_n29520_, new_n29519_, new_n29510_ );
and  ( new_n29521_, new_n29519_, new_n29510_ );
or   ( new_n29522_, new_n19048_, new_n124_ );
or   ( new_n29523_, new_n19055_, new_n6321_ );
and  ( new_n29524_, new_n29523_, new_n29522_ );
or   ( new_n29525_, new_n29524_, new_n18742_ );
and  ( new_n29526_, new_n19057_, RI2b1c4342e2f0_95 );
and  ( new_n29527_, new_n19044_, RI2b1c4342e278_94 );
or   ( new_n29528_, new_n29527_, new_n29526_ );
or   ( new_n29529_, new_n29528_, new_n18977_ );
and  ( new_n29530_, new_n29529_, new_n29525_ );
or   ( new_n29531_, new_n29530_, new_n29521_ );
and  ( new_n29532_, new_n29531_, new_n29520_ );
nor  ( new_n29533_, new_n22333_, new_n3924_ );
nor  ( new_n29534_, new_n29533_, new_n14372_ );
or   ( new_n29535_, new_n29534_, new_n21261_ );
and  ( new_n29536_, new_n22337_, RI2b1c4342df30_87 );
and  ( new_n29537_, new_n22330_, RI2b1c4342deb8_86 );
or   ( new_n29538_, new_n29537_, new_n29536_ );
or   ( new_n29539_, new_n29538_, new_n21009_ );
and  ( new_n29540_, new_n29539_, new_n29535_ );
and  ( new_n29541_, new_n29540_, new_n18309_ );
or   ( new_n29542_, new_n29540_, new_n18309_ );
or   ( new_n29543_, new_n21419_, new_n132_ );
or   ( new_n29544_, new_n21424_, new_n3902_ );
and  ( new_n29545_, new_n29544_, new_n29543_ );
or   ( new_n29546_, new_n29545_, new_n21013_ );
and  ( new_n29547_, new_n21428_, RI2b1c4342e020_89 );
and  ( new_n29548_, new_n21415_, RI2b1c4342dfa8_88 );
or   ( new_n29549_, new_n29548_, new_n29547_ );
or   ( new_n29550_, new_n29549_, new_n21265_ );
and  ( new_n29551_, new_n29550_, new_n29546_ );
and  ( new_n29552_, new_n29551_, new_n29542_ );
or   ( new_n29553_, new_n29552_, new_n29541_ );
and  ( new_n29554_, new_n29553_, new_n29532_ );
or   ( new_n29555_, new_n29553_, new_n29532_ );
or   ( new_n29556_, new_n29469_, new_n29365_ );
or   ( new_n29557_, new_n29466_, new_n29374_ );
and  ( new_n29558_, new_n29557_, new_n29556_ );
or   ( new_n29559_, new_n29558_, new_n29474_ );
and  ( new_n29560_, new_n29470_, new_n29375_ );
or   ( new_n29561_, new_n29560_, new_n29385_ );
and  ( new_n29562_, new_n29561_, new_n29559_ );
and  ( new_n29563_, new_n29562_, new_n29555_ );
or   ( new_n29564_, new_n29563_, new_n29554_ );
or   ( new_n29565_, new_n29564_, new_n29501_ );
or   ( new_n29566_, new_n29508_, new_n20156_ );
or   ( new_n29567_, new_n29504_, new_n20443_ );
and  ( new_n29568_, new_n29567_, new_n29566_ );
or   ( new_n29569_, new_n29517_, new_n19394_ );
or   ( new_n29570_, new_n29513_, new_n19659_ );
and  ( new_n29571_, new_n29570_, new_n29569_ );
or   ( new_n29572_, new_n29571_, new_n29568_ );
and  ( new_n29573_, new_n29571_, new_n29568_ );
or   ( new_n29574_, new_n29528_, new_n18742_ );
or   ( new_n29575_, new_n29524_, new_n18977_ );
and  ( new_n29576_, new_n29575_, new_n29574_ );
or   ( new_n29577_, new_n29576_, new_n29573_ );
and  ( new_n29578_, new_n29577_, new_n29572_ );
or   ( new_n29579_, new_n29538_, new_n21261_ );
or   ( new_n29580_, new_n29534_, new_n21009_ );
and  ( new_n29581_, new_n29580_, new_n29579_ );
or   ( new_n29582_, new_n29581_, new_n18066_ );
and  ( new_n29583_, new_n29581_, new_n18066_ );
or   ( new_n29584_, new_n29549_, new_n21013_ );
or   ( new_n29585_, new_n29545_, new_n21265_ );
and  ( new_n29586_, new_n29585_, new_n29584_ );
or   ( new_n29587_, new_n29586_, new_n29583_ );
and  ( new_n29588_, new_n29587_, new_n29582_ );
or   ( new_n29589_, new_n29588_, new_n29578_ );
and  ( new_n29590_, new_n29588_, new_n29578_ );
or   ( new_n29591_, new_n29560_, new_n29474_ );
or   ( new_n29592_, new_n29558_, new_n29385_ );
and  ( new_n29593_, new_n29592_, new_n29591_ );
or   ( new_n29594_, new_n29593_, new_n29590_ );
and  ( new_n29595_, new_n29594_, new_n29589_ );
or   ( new_n29596_, new_n29499_, new_n29487_ );
or   ( new_n29597_, new_n29495_, new_n29421_ );
and  ( new_n29598_, new_n29597_, new_n29596_ );
or   ( new_n29599_, new_n29598_, new_n29595_ );
and  ( new_n29600_, new_n29599_, new_n29565_ );
or   ( new_n29601_, new_n29600_, new_n29484_ );
or   ( new_n29602_, new_n29482_, new_n29450_ );
or   ( new_n29603_, new_n29478_, new_n29398_ );
and  ( new_n29604_, new_n29603_, new_n29602_ );
or   ( new_n29605_, new_n29595_, new_n29501_ );
or   ( new_n29606_, new_n29598_, new_n29564_ );
and  ( new_n29607_, new_n29606_, new_n29605_ );
or   ( new_n29608_, new_n29607_, new_n29604_ );
and  ( new_n29609_, new_n29608_, new_n29601_ );
or   ( new_n29610_, new_n29456_, new_n29334_ );
or   ( new_n29611_, new_n29453_, new_n29343_ );
and  ( new_n29612_, new_n29611_, new_n29610_ );
or   ( new_n29613_, new_n29612_, new_n29461_ );
and  ( new_n29614_, new_n29457_, new_n29344_ );
or   ( new_n29615_, new_n29614_, new_n29354_ );
and  ( new_n29616_, new_n29615_, new_n29613_ );
or   ( new_n29617_, new_n18395_, new_n7274_ );
or   ( new_n29618_, new_n29617_, new_n18066_ );
and  ( new_n29619_, new_n18384_, RI2b1c4342e368_96 );
or   ( new_n29620_, new_n29619_, new_n18309_ );
and  ( new_n29621_, new_n29620_, new_n29618_ );
nor  ( new_n29622_, new_n22333_, new_n3902_ );
nor  ( new_n29623_, new_n29622_, new_n14537_ );
or   ( new_n29624_, new_n29623_, new_n21261_ );
and  ( new_n29625_, new_n22337_, RI2b1c4342dfa8_88 );
and  ( new_n29626_, new_n22330_, RI2b1c4342df30_87 );
or   ( new_n29627_, new_n29626_, new_n29625_ );
or   ( new_n29628_, new_n29627_, new_n21009_ );
and  ( new_n29629_, new_n29628_, new_n29624_ );
or   ( new_n29630_, new_n21419_, new_n4635_ );
or   ( new_n29631_, new_n21424_, new_n132_ );
and  ( new_n29632_, new_n29631_, new_n29630_ );
or   ( new_n29633_, new_n29632_, new_n21013_ );
and  ( new_n29634_, new_n21428_, RI2b1c4342e098_90 );
and  ( new_n29635_, new_n21415_, RI2b1c4342e020_89 );
or   ( new_n29636_, new_n29635_, new_n29634_ );
or   ( new_n29637_, new_n29636_, new_n21265_ );
and  ( new_n29638_, new_n29637_, new_n29633_ );
or   ( new_n29639_, new_n29638_, new_n29629_ );
and  ( new_n29640_, new_n29638_, new_n29629_ );
or   ( new_n29641_, new_n20557_, new_n5459_ );
or   ( new_n29642_, new_n20562_, new_n117_ );
and  ( new_n29643_, new_n29642_, new_n29641_ );
or   ( new_n29644_, new_n29643_, new_n20156_ );
and  ( new_n29645_, new_n20566_, RI2b1c4342e188_92 );
and  ( new_n29646_, new_n20553_, RI2b1c4342e110_91 );
or   ( new_n29647_, new_n29646_, new_n29645_ );
or   ( new_n29648_, new_n29647_, new_n20443_ );
and  ( new_n29649_, new_n29648_, new_n29644_ );
or   ( new_n29650_, new_n29649_, new_n29640_ );
and  ( new_n29651_, new_n29650_, new_n29639_ );
or   ( new_n29652_, new_n29651_, new_n29621_ );
and  ( new_n29653_, new_n29651_, new_n29621_ );
or   ( new_n29654_, new_n29571_, new_n29510_ );
or   ( new_n29655_, new_n29568_, new_n29519_ );
and  ( new_n29656_, new_n29655_, new_n29654_ );
or   ( new_n29657_, new_n29656_, new_n29576_ );
and  ( new_n29658_, new_n29572_, new_n29520_ );
or   ( new_n29659_, new_n29658_, new_n29530_ );
and  ( new_n29660_, new_n29659_, new_n29657_ );
or   ( new_n29661_, new_n29660_, new_n29653_ );
and  ( new_n29662_, new_n29661_, new_n29652_ );
or   ( new_n29663_, new_n29662_, new_n29616_ );
and  ( new_n29664_, new_n29662_, new_n29616_ );
or   ( new_n29665_, new_n29578_, new_n29553_ );
or   ( new_n29666_, new_n29588_, new_n29532_ );
and  ( new_n29667_, new_n29666_, new_n29665_ );
or   ( new_n29668_, new_n29667_, new_n29593_ );
and  ( new_n29669_, new_n29589_, new_n29555_ );
or   ( new_n29670_, new_n29669_, new_n29562_ );
and  ( new_n29671_, new_n29670_, new_n29668_ );
or   ( new_n29672_, new_n29671_, new_n29664_ );
and  ( new_n29673_, new_n29672_, new_n29663_ );
or   ( new_n29674_, new_n29673_, new_n29609_ );
or   ( new_n29675_, new_n29429_, new_n29137_ );
or   ( new_n29676_, new_n29427_, new_n29052_ );
and  ( new_n29677_, new_n29676_, new_n29675_ );
and  ( new_n29678_, new_n29476_, new_n29463_ );
or   ( new_n29679_, new_n29678_, new_n29450_ );
and  ( new_n29680_, new_n29679_, new_n29477_ );
and  ( new_n29681_, new_n29493_, new_n29490_ );
or   ( new_n29682_, new_n29681_, new_n29487_ );
and  ( new_n29683_, new_n29682_, new_n29494_ );
or   ( new_n29684_, new_n29683_, new_n29680_ );
and  ( new_n29685_, new_n29684_, new_n29424_ );
or   ( new_n29686_, new_n29685_, new_n29677_ );
or   ( new_n29687_, new_n29683_, new_n29400_ );
or   ( new_n29688_, new_n29680_, new_n29423_ );
and  ( new_n29689_, new_n29688_, new_n29687_ );
or   ( new_n29690_, new_n29689_, new_n29431_ );
and  ( new_n29691_, new_n29690_, new_n29686_ );
or   ( new_n29692_, new_n29316_, new_n29124_ );
or   ( new_n29693_, new_n29314_, new_n29021_ );
and  ( new_n29694_, new_n29693_, new_n29692_ );
or   ( new_n29695_, new_n29323_, new_n29295_ );
or   ( new_n29696_, new_n29321_, new_n29233_ );
and  ( new_n29697_, new_n29696_, new_n29695_ );
or   ( new_n29698_, new_n29697_, new_n29694_ );
and  ( new_n29699_, new_n29698_, new_n29326_ );
and  ( new_n29700_, new_n29598_, new_n29564_ );
and  ( new_n29701_, new_n29606_, new_n29604_ );
or   ( new_n29702_, new_n29701_, new_n29700_ );
or   ( new_n29703_, new_n29702_, new_n29699_ );
and  ( new_n29704_, new_n29595_, new_n29501_ );
or   ( new_n29705_, new_n29704_, new_n29484_ );
and  ( new_n29706_, new_n29705_, new_n29605_ );
or   ( new_n29707_, new_n29697_, new_n29318_ );
or   ( new_n29708_, new_n29694_, new_n29325_ );
and  ( new_n29709_, new_n29708_, new_n29707_ );
or   ( new_n29710_, new_n29709_, new_n29706_ );
and  ( new_n29711_, new_n29710_, new_n29703_ );
or   ( new_n29712_, new_n29711_, new_n29691_ );
or   ( new_n29713_, new_n29706_, new_n29699_ );
or   ( new_n29714_, new_n29709_, new_n29702_ );
and  ( new_n29715_, new_n29714_, new_n29713_ );
or   ( new_n29716_, new_n29689_, new_n29677_ );
or   ( new_n29717_, new_n29685_, new_n29431_ );
and  ( new_n29718_, new_n29717_, new_n29716_ );
or   ( new_n29719_, new_n29718_, new_n29715_ );
and  ( new_n29720_, new_n29719_, new_n29712_ );
and  ( new_n29721_, new_n29720_, new_n29674_ );
or   ( new_n29722_, new_n29440_, new_n29302_ );
or   ( new_n29723_, new_n29438_, new_n29244_ );
and  ( new_n29724_, new_n29723_, new_n29722_ );
and  ( new_n29725_, new_n29697_, new_n29694_ );
or   ( new_n29726_, new_n29725_, new_n29434_ );
and  ( new_n29727_, new_n29683_, new_n29680_ );
or   ( new_n29728_, new_n29727_, new_n29677_ );
and  ( new_n29729_, new_n29728_, new_n29684_ );
or   ( new_n29730_, new_n29729_, new_n29326_ );
and  ( new_n29731_, new_n29730_, new_n29726_ );
or   ( new_n29732_, new_n29731_, new_n29724_ );
or   ( new_n29733_, new_n29729_, new_n29725_ );
and  ( new_n29734_, new_n29733_, new_n29435_ );
or   ( new_n29735_, new_n29734_, new_n29442_ );
and  ( new_n29736_, new_n29735_, new_n29732_ );
and  ( new_n29737_, new_n29709_, new_n29702_ );
and  ( new_n29738_, new_n29718_, new_n29714_ );
or   ( new_n29739_, new_n29738_, new_n29737_ );
and  ( new_n29740_, new_n29739_, new_n29736_ );
or   ( new_n29741_, new_n29740_, new_n29721_ );
or   ( new_n29742_, new_n29669_, new_n29593_ );
or   ( new_n29743_, new_n29667_, new_n29562_ );
and  ( new_n29744_, new_n29743_, new_n29742_ );
or   ( new_n29745_, new_n29614_, new_n29461_ );
or   ( new_n29746_, new_n29612_, new_n29354_ );
and  ( new_n29747_, new_n29746_, new_n29745_ );
or   ( new_n29748_, new_n29747_, new_n29662_ );
or   ( new_n29749_, new_n29619_, new_n18066_ );
or   ( new_n29750_, new_n29617_, new_n18309_ );
and  ( new_n29751_, new_n29750_, new_n29749_ );
or   ( new_n29752_, new_n29627_, new_n21261_ );
or   ( new_n29753_, new_n29623_, new_n21009_ );
and  ( new_n29754_, new_n29753_, new_n29752_ );
or   ( new_n29755_, new_n29636_, new_n21013_ );
or   ( new_n29756_, new_n29632_, new_n21265_ );
and  ( new_n29757_, new_n29756_, new_n29755_ );
or   ( new_n29758_, new_n29757_, new_n29754_ );
and  ( new_n29759_, new_n29757_, new_n29754_ );
or   ( new_n29760_, new_n29647_, new_n20156_ );
or   ( new_n29761_, new_n29643_, new_n20443_ );
and  ( new_n29762_, new_n29761_, new_n29760_ );
or   ( new_n29763_, new_n29762_, new_n29759_ );
and  ( new_n29764_, new_n29763_, new_n29758_ );
or   ( new_n29765_, new_n29764_, new_n29751_ );
and  ( new_n29766_, new_n29764_, new_n29751_ );
or   ( new_n29767_, new_n29658_, new_n29576_ );
or   ( new_n29768_, new_n29656_, new_n29530_ );
and  ( new_n29769_, new_n29768_, new_n29767_ );
or   ( new_n29770_, new_n29769_, new_n29766_ );
and  ( new_n29771_, new_n29770_, new_n29765_ );
or   ( new_n29772_, new_n29771_, new_n29616_ );
and  ( new_n29773_, new_n29772_, new_n29748_ );
or   ( new_n29774_, new_n29773_, new_n29744_ );
or   ( new_n29775_, new_n29771_, new_n29747_ );
and  ( new_n29776_, new_n29775_, new_n29663_ );
or   ( new_n29777_, new_n29776_, new_n29671_ );
and  ( new_n29778_, new_n29777_, new_n29774_ );
or   ( new_n29779_, new_n19048_, new_n7274_ );
or   ( new_n29780_, new_n19055_, new_n124_ );
and  ( new_n29781_, new_n29780_, new_n29779_ );
or   ( new_n29782_, new_n29781_, new_n18742_ );
and  ( new_n29783_, new_n19057_, RI2b1c4342e368_96 );
and  ( new_n29784_, new_n19044_, RI2b1c4342e2f0_95 );
or   ( new_n29785_, new_n29784_, new_n29783_ );
or   ( new_n29786_, new_n29785_, new_n18977_ );
and  ( new_n29787_, new_n29786_, new_n29782_ );
or   ( new_n29788_, new_n29757_, new_n29629_ );
or   ( new_n29789_, new_n29754_, new_n29638_ );
and  ( new_n29790_, new_n29789_, new_n29788_ );
or   ( new_n29791_, new_n29790_, new_n29762_ );
and  ( new_n29792_, new_n29758_, new_n29639_ );
or   ( new_n29793_, new_n29792_, new_n29649_ );
and  ( new_n29794_, new_n29793_, new_n29791_ );
or   ( new_n29795_, new_n29794_, new_n29787_ );
or   ( new_n29796_, new_n20557_, new_n6307_ );
or   ( new_n29797_, new_n20562_, new_n5459_ );
and  ( new_n29798_, new_n29797_, new_n29796_ );
or   ( new_n29799_, new_n29798_, new_n20156_ );
and  ( new_n29800_, new_n20566_, RI2b1c4342e200_93 );
and  ( new_n29801_, new_n20553_, RI2b1c4342e188_92 );
or   ( new_n29802_, new_n29801_, new_n29800_ );
or   ( new_n29803_, new_n29802_, new_n20443_ );
and  ( new_n29804_, new_n29803_, new_n29799_ );
or   ( new_n29805_, new_n19758_, new_n124_ );
or   ( new_n29806_, new_n19763_, new_n6321_ );
and  ( new_n29807_, new_n29806_, new_n29805_ );
or   ( new_n29808_, new_n29807_, new_n19394_ );
and  ( new_n29809_, new_n19767_, RI2b1c4342e2f0_95 );
and  ( new_n29810_, new_n19754_, RI2b1c4342e278_94 );
or   ( new_n29811_, new_n29810_, new_n29809_ );
or   ( new_n29812_, new_n29811_, new_n19659_ );
and  ( new_n29813_, new_n29812_, new_n29808_ );
or   ( new_n29814_, new_n29813_, new_n29804_ );
and  ( new_n29815_, new_n29813_, new_n29804_ );
or   ( new_n29816_, new_n19055_, new_n7274_ );
or   ( new_n29817_, new_n29816_, new_n18742_ );
and  ( new_n29818_, new_n19044_, RI2b1c4342e368_96 );
or   ( new_n29819_, new_n29818_, new_n18977_ );
and  ( new_n29820_, new_n29819_, new_n29817_ );
or   ( new_n29821_, new_n29820_, new_n29815_ );
and  ( new_n29822_, new_n29821_, new_n29814_ );
nor  ( new_n29823_, new_n22333_, new_n132_ );
nor  ( new_n29824_, new_n29823_, new_n14701_ );
or   ( new_n29825_, new_n29824_, new_n21261_ );
and  ( new_n29826_, new_n22337_, RI2b1c4342e020_89 );
and  ( new_n29827_, new_n22330_, RI2b1c4342dfa8_88 );
or   ( new_n29828_, new_n29827_, new_n29826_ );
or   ( new_n29829_, new_n29828_, new_n21009_ );
and  ( new_n29830_, new_n29829_, new_n29825_ );
and  ( new_n29831_, new_n29830_, new_n18977_ );
or   ( new_n29832_, new_n29830_, new_n18977_ );
or   ( new_n29833_, new_n21419_, new_n117_ );
or   ( new_n29834_, new_n21424_, new_n4635_ );
and  ( new_n29835_, new_n29834_, new_n29833_ );
or   ( new_n29836_, new_n29835_, new_n21013_ );
and  ( new_n29837_, new_n21428_, RI2b1c4342e110_91 );
and  ( new_n29838_, new_n21415_, RI2b1c4342e098_90 );
or   ( new_n29839_, new_n29838_, new_n29837_ );
or   ( new_n29840_, new_n29839_, new_n21265_ );
and  ( new_n29841_, new_n29840_, new_n29836_ );
and  ( new_n29842_, new_n29841_, new_n29832_ );
or   ( new_n29843_, new_n29842_, new_n29831_ );
and  ( new_n29844_, new_n29843_, new_n29822_ );
or   ( new_n29845_, new_n29843_, new_n29822_ );
or   ( new_n29846_, new_n19758_, new_n6321_ );
or   ( new_n29847_, new_n19763_, new_n6307_ );
and  ( new_n29848_, new_n29847_, new_n29846_ );
or   ( new_n29849_, new_n29848_, new_n19394_ );
and  ( new_n29850_, new_n19767_, RI2b1c4342e278_94 );
and  ( new_n29851_, new_n19754_, RI2b1c4342e200_93 );
or   ( new_n29852_, new_n29851_, new_n29850_ );
or   ( new_n29853_, new_n29852_, new_n19659_ );
and  ( new_n29854_, new_n29853_, new_n29849_ );
and  ( new_n29855_, new_n29854_, new_n29845_ );
or   ( new_n29856_, new_n29855_, new_n29844_ );
and  ( new_n29857_, new_n29856_, new_n29795_ );
or   ( new_n29858_, new_n29856_, new_n29795_ );
or   ( new_n29859_, new_n29581_, new_n18309_ );
or   ( new_n29860_, new_n29540_, new_n18066_ );
and  ( new_n29861_, new_n29860_, new_n29859_ );
or   ( new_n29862_, new_n29861_, new_n29586_ );
and  ( new_n29863_, new_n29582_, new_n29542_ );
or   ( new_n29864_, new_n29863_, new_n29551_ );
and  ( new_n29865_, new_n29864_, new_n29862_ );
and  ( new_n29866_, new_n29865_, new_n29858_ );
or   ( new_n29867_, new_n29866_, new_n29857_ );
or   ( new_n29868_, new_n29867_, new_n29778_ );
or   ( new_n29869_, new_n29607_, new_n29484_ );
or   ( new_n29870_, new_n29604_, new_n29600_ );
and  ( new_n29871_, new_n29870_, new_n29869_ );
or   ( new_n29872_, new_n29871_, new_n29673_ );
and  ( new_n29873_, new_n29771_, new_n29747_ );
or   ( new_n29874_, new_n29873_, new_n29744_ );
and  ( new_n29875_, new_n29874_, new_n29775_ );
or   ( new_n29876_, new_n29875_, new_n29609_ );
and  ( new_n29877_, new_n29876_, new_n29872_ );
and  ( new_n29878_, new_n29877_, new_n29868_ );
or   ( new_n29879_, new_n29751_, new_n29651_ );
or   ( new_n29880_, new_n29764_, new_n29621_ );
and  ( new_n29881_, new_n29880_, new_n29879_ );
or   ( new_n29882_, new_n29881_, new_n29769_ );
and  ( new_n29883_, new_n29765_, new_n29652_ );
or   ( new_n29884_, new_n29883_, new_n29660_ );
and  ( new_n29885_, new_n29884_, new_n29882_ );
or   ( new_n29886_, new_n29863_, new_n29586_ );
or   ( new_n29887_, new_n29861_, new_n29551_ );
and  ( new_n29888_, new_n29887_, new_n29886_ );
or   ( new_n29889_, new_n29785_, new_n18742_ );
or   ( new_n29890_, new_n29781_, new_n18977_ );
and  ( new_n29891_, new_n29890_, new_n29889_ );
or   ( new_n29892_, new_n29792_, new_n29762_ );
or   ( new_n29893_, new_n29790_, new_n29649_ );
and  ( new_n29894_, new_n29893_, new_n29892_ );
and  ( new_n29895_, new_n29894_, new_n29891_ );
or   ( new_n29896_, new_n29895_, new_n29856_ );
or   ( new_n29897_, new_n29802_, new_n20156_ );
or   ( new_n29898_, new_n29798_, new_n20443_ );
and  ( new_n29899_, new_n29898_, new_n29897_ );
or   ( new_n29900_, new_n29811_, new_n19394_ );
or   ( new_n29901_, new_n29807_, new_n19659_ );
and  ( new_n29902_, new_n29901_, new_n29900_ );
or   ( new_n29903_, new_n29902_, new_n29899_ );
and  ( new_n29904_, new_n29902_, new_n29899_ );
or   ( new_n29905_, new_n29818_, new_n18742_ );
or   ( new_n29906_, new_n29816_, new_n18977_ );
and  ( new_n29907_, new_n29906_, new_n29905_ );
or   ( new_n29908_, new_n29907_, new_n29904_ );
and  ( new_n29909_, new_n29908_, new_n29903_ );
or   ( new_n29910_, new_n29828_, new_n21261_ );
or   ( new_n29911_, new_n29824_, new_n21009_ );
and  ( new_n29912_, new_n29911_, new_n29910_ );
or   ( new_n29913_, new_n29912_, new_n18742_ );
and  ( new_n29914_, new_n29912_, new_n18742_ );
or   ( new_n29915_, new_n29839_, new_n21013_ );
or   ( new_n29916_, new_n29835_, new_n21265_ );
and  ( new_n29917_, new_n29916_, new_n29915_ );
or   ( new_n29918_, new_n29917_, new_n29914_ );
and  ( new_n29919_, new_n29918_, new_n29913_ );
or   ( new_n29920_, new_n29919_, new_n29909_ );
and  ( new_n29921_, new_n29919_, new_n29909_ );
or   ( new_n29922_, new_n29852_, new_n19394_ );
or   ( new_n29923_, new_n29848_, new_n19659_ );
and  ( new_n29924_, new_n29923_, new_n29922_ );
or   ( new_n29925_, new_n29924_, new_n29921_ );
and  ( new_n29926_, new_n29925_, new_n29920_ );
or   ( new_n29927_, new_n29926_, new_n29795_ );
and  ( new_n29928_, new_n29927_, new_n29896_ );
or   ( new_n29929_, new_n29928_, new_n29888_ );
or   ( new_n29930_, new_n29926_, new_n29895_ );
and  ( new_n29931_, new_n29930_, new_n29858_ );
or   ( new_n29932_, new_n29931_, new_n29865_ );
and  ( new_n29933_, new_n29932_, new_n29929_ );
or   ( new_n29934_, new_n29933_, new_n29885_ );
or   ( new_n29935_, new_n29776_, new_n29744_ );
or   ( new_n29936_, new_n29773_, new_n29671_ );
and  ( new_n29937_, new_n29936_, new_n29935_ );
or   ( new_n29938_, new_n29937_, new_n29867_ );
and  ( new_n29939_, new_n29926_, new_n29895_ );
or   ( new_n29940_, new_n29939_, new_n29888_ );
and  ( new_n29941_, new_n29940_, new_n29930_ );
or   ( new_n29942_, new_n29941_, new_n29778_ );
and  ( new_n29943_, new_n29942_, new_n29938_ );
and  ( new_n29944_, new_n29943_, new_n29934_ );
or   ( new_n29945_, new_n29944_, new_n29878_ );
and  ( new_n29946_, new_n29913_, new_n29832_ );
or   ( new_n29947_, new_n29946_, new_n29917_ );
or   ( new_n29948_, new_n29912_, new_n18977_ );
or   ( new_n29949_, new_n29830_, new_n18742_ );
and  ( new_n29950_, new_n29949_, new_n29948_ );
or   ( new_n29951_, new_n29950_, new_n29841_ );
and  ( new_n29952_, new_n29951_, new_n29947_ );
and  ( new_n29953_, new_n29903_, new_n29814_ );
or   ( new_n29954_, new_n29953_, new_n29907_ );
or   ( new_n29955_, new_n29902_, new_n29804_ );
or   ( new_n29956_, new_n29899_, new_n29813_ );
and  ( new_n29957_, new_n29956_, new_n29955_ );
or   ( new_n29958_, new_n29957_, new_n29820_ );
and  ( new_n29959_, new_n29958_, new_n29954_ );
nor  ( new_n29960_, new_n22333_, new_n4635_ );
nor  ( new_n29961_, new_n29960_, new_n14825_ );
or   ( new_n29962_, new_n29961_, new_n21261_ );
and  ( new_n29963_, new_n22337_, RI2b1c4342e098_90 );
and  ( new_n29964_, new_n22330_, RI2b1c4342e020_89 );
or   ( new_n29965_, new_n29964_, new_n29963_ );
or   ( new_n29966_, new_n29965_, new_n21009_ );
and  ( new_n29967_, new_n29966_, new_n29962_ );
or   ( new_n29968_, new_n21419_, new_n5459_ );
or   ( new_n29969_, new_n21424_, new_n117_ );
and  ( new_n29970_, new_n29969_, new_n29968_ );
or   ( new_n29971_, new_n29970_, new_n21013_ );
and  ( new_n29972_, new_n21428_, RI2b1c4342e188_92 );
and  ( new_n29973_, new_n21415_, RI2b1c4342e110_91 );
or   ( new_n29974_, new_n29973_, new_n29972_ );
or   ( new_n29975_, new_n29974_, new_n21265_ );
and  ( new_n29976_, new_n29975_, new_n29971_ );
or   ( new_n29977_, new_n29976_, new_n29967_ );
and  ( new_n29978_, new_n29976_, new_n29967_ );
or   ( new_n29979_, new_n20557_, new_n6321_ );
or   ( new_n29980_, new_n20562_, new_n6307_ );
and  ( new_n29981_, new_n29980_, new_n29979_ );
or   ( new_n29982_, new_n29981_, new_n20156_ );
and  ( new_n29983_, new_n20566_, RI2b1c4342e278_94 );
and  ( new_n29984_, new_n20553_, RI2b1c4342e200_93 );
or   ( new_n29985_, new_n29984_, new_n29983_ );
or   ( new_n29986_, new_n29985_, new_n20443_ );
and  ( new_n29987_, new_n29986_, new_n29982_ );
or   ( new_n29988_, new_n29987_, new_n29978_ );
and  ( new_n29989_, new_n29988_, new_n29977_ );
or   ( new_n29990_, new_n29989_, new_n29959_ );
or   ( new_n29991_, new_n29974_, new_n21013_ );
or   ( new_n29992_, new_n29970_, new_n21265_ );
and  ( new_n29993_, new_n29992_, new_n29991_ );
or   ( new_n29994_, new_n29965_, new_n21261_ );
or   ( new_n29995_, new_n29961_, new_n21009_ );
and  ( new_n29996_, new_n29995_, new_n29994_ );
or   ( new_n29997_, new_n29996_, new_n29993_ );
and  ( new_n29998_, new_n29996_, new_n29993_ );
or   ( new_n29999_, new_n29985_, new_n20156_ );
or   ( new_n30000_, new_n29981_, new_n20443_ );
and  ( new_n30001_, new_n30000_, new_n29999_ );
or   ( new_n30002_, new_n30001_, new_n29998_ );
and  ( new_n30003_, new_n30002_, new_n29997_ );
or   ( new_n30004_, new_n29957_, new_n29907_ );
or   ( new_n30005_, new_n29953_, new_n29820_ );
and  ( new_n30006_, new_n30005_, new_n30004_ );
or   ( new_n30007_, new_n30006_, new_n30003_ );
and  ( new_n30008_, new_n30007_, new_n29990_ );
or   ( new_n30009_, new_n30008_, new_n29952_ );
or   ( new_n30010_, new_n29950_, new_n29917_ );
or   ( new_n30011_, new_n29946_, new_n29841_ );
and  ( new_n30012_, new_n30011_, new_n30010_ );
or   ( new_n30013_, new_n30003_, new_n29959_ );
or   ( new_n30014_, new_n30006_, new_n29989_ );
and  ( new_n30015_, new_n30014_, new_n30013_ );
or   ( new_n30016_, new_n30015_, new_n30012_ );
and  ( new_n30017_, new_n30016_, new_n30009_ );
or   ( new_n30018_, new_n20557_, new_n124_ );
or   ( new_n30019_, new_n20562_, new_n6321_ );
and  ( new_n30020_, new_n30019_, new_n30018_ );
or   ( new_n30021_, new_n30020_, new_n20156_ );
and  ( new_n30022_, new_n20566_, RI2b1c4342e2f0_95 );
and  ( new_n30023_, new_n20553_, RI2b1c4342e278_94 );
or   ( new_n30024_, new_n30023_, new_n30022_ );
or   ( new_n30025_, new_n30024_, new_n20443_ );
and  ( new_n30026_, new_n30025_, new_n30021_ );
or   ( new_n30027_, new_n19763_, new_n7274_ );
or   ( new_n30028_, new_n30027_, new_n19394_ );
and  ( new_n30029_, new_n19754_, RI2b1c4342e368_96 );
or   ( new_n30030_, new_n30029_, new_n19659_ );
and  ( new_n30031_, new_n30030_, new_n30028_ );
or   ( new_n30032_, new_n30031_, new_n30026_ );
nor  ( new_n30033_, new_n22333_, new_n117_ );
nor  ( new_n30034_, new_n30033_, new_n14934_ );
or   ( new_n30035_, new_n30034_, new_n21261_ );
and  ( new_n30036_, new_n22337_, RI2b1c4342e110_91 );
and  ( new_n30037_, new_n22330_, RI2b1c4342e098_90 );
or   ( new_n30038_, new_n30037_, new_n30036_ );
or   ( new_n30039_, new_n30038_, new_n21009_ );
and  ( new_n30040_, new_n30039_, new_n30035_ );
and  ( new_n30041_, new_n30040_, new_n19659_ );
or   ( new_n30042_, new_n30040_, new_n19659_ );
or   ( new_n30043_, new_n21419_, new_n6307_ );
or   ( new_n30044_, new_n21424_, new_n5459_ );
and  ( new_n30045_, new_n30044_, new_n30043_ );
or   ( new_n30046_, new_n30045_, new_n21013_ );
and  ( new_n30047_, new_n21428_, RI2b1c4342e200_93 );
and  ( new_n30048_, new_n21415_, RI2b1c4342e188_92 );
or   ( new_n30049_, new_n30048_, new_n30047_ );
or   ( new_n30050_, new_n30049_, new_n21265_ );
and  ( new_n30051_, new_n30050_, new_n30046_ );
and  ( new_n30052_, new_n30051_, new_n30042_ );
or   ( new_n30053_, new_n30052_, new_n30041_ );
and  ( new_n30054_, new_n30053_, new_n30032_ );
or   ( new_n30055_, new_n30053_, new_n30032_ );
or   ( new_n30056_, new_n19758_, new_n7274_ );
or   ( new_n30057_, new_n19763_, new_n124_ );
and  ( new_n30058_, new_n30057_, new_n30056_ );
or   ( new_n30059_, new_n30058_, new_n19394_ );
and  ( new_n30060_, new_n19767_, RI2b1c4342e368_96 );
and  ( new_n30061_, new_n19754_, RI2b1c4342e2f0_95 );
or   ( new_n30062_, new_n30061_, new_n30060_ );
or   ( new_n30063_, new_n30062_, new_n19659_ );
and  ( new_n30064_, new_n30063_, new_n30059_ );
and  ( new_n30065_, new_n30064_, new_n30055_ );
or   ( new_n30066_, new_n30065_, new_n30054_ );
or   ( new_n30067_, new_n30066_, new_n30017_ );
and  ( new_n30068_, new_n29920_, new_n29845_ );
or   ( new_n30069_, new_n30068_, new_n29924_ );
or   ( new_n30070_, new_n29909_, new_n29843_ );
or   ( new_n30071_, new_n29919_, new_n29822_ );
and  ( new_n30072_, new_n30071_, new_n30070_ );
or   ( new_n30073_, new_n30072_, new_n29854_ );
and  ( new_n30074_, new_n30073_, new_n30069_ );
or   ( new_n30075_, new_n29894_, new_n29891_ );
and  ( new_n30076_, new_n30075_, new_n29795_ );
and  ( new_n30077_, new_n30006_, new_n29989_ );
or   ( new_n30078_, new_n30077_, new_n30012_ );
and  ( new_n30079_, new_n30078_, new_n30014_ );
or   ( new_n30080_, new_n30079_, new_n30076_ );
and  ( new_n30081_, new_n30003_, new_n29959_ );
or   ( new_n30082_, new_n30081_, new_n29952_ );
and  ( new_n30083_, new_n30082_, new_n30013_ );
or   ( new_n30084_, new_n29894_, new_n29787_ );
or   ( new_n30085_, new_n29891_, new_n29794_ );
and  ( new_n30086_, new_n30085_, new_n30084_ );
or   ( new_n30087_, new_n30086_, new_n30083_ );
and  ( new_n30088_, new_n30087_, new_n30080_ );
or   ( new_n30089_, new_n30088_, new_n30074_ );
or   ( new_n30090_, new_n30083_, new_n30076_ );
or   ( new_n30091_, new_n30086_, new_n30079_ );
and  ( new_n30092_, new_n30091_, new_n30090_ );
or   ( new_n30093_, new_n30072_, new_n29924_ );
or   ( new_n30094_, new_n30068_, new_n29854_ );
and  ( new_n30095_, new_n30094_, new_n30093_ );
or   ( new_n30096_, new_n30095_, new_n30092_ );
and  ( new_n30097_, new_n30096_, new_n30089_ );
and  ( new_n30098_, new_n30097_, new_n30067_ );
or   ( new_n30099_, new_n29931_, new_n29888_ );
or   ( new_n30100_, new_n29928_, new_n29865_ );
and  ( new_n30101_, new_n30100_, new_n30099_ );
or   ( new_n30102_, new_n30101_, new_n29885_ );
or   ( new_n30103_, new_n29883_, new_n29769_ );
or   ( new_n30104_, new_n29881_, new_n29660_ );
and  ( new_n30105_, new_n30104_, new_n30103_ );
or   ( new_n30106_, new_n30105_, new_n29933_ );
and  ( new_n30107_, new_n30106_, new_n30102_ );
and  ( new_n30108_, new_n30086_, new_n30079_ );
or   ( new_n30109_, new_n30108_, new_n30095_ );
and  ( new_n30110_, new_n30109_, new_n30091_ );
and  ( new_n30111_, new_n30110_, new_n30107_ );
or   ( new_n30112_, new_n30111_, new_n30098_ );
or   ( new_n30113_, new_n29993_, new_n29967_ );
or   ( new_n30114_, new_n29996_, new_n29976_ );
and  ( new_n30115_, new_n30114_, new_n30113_ );
or   ( new_n30116_, new_n30115_, new_n30001_ );
and  ( new_n30117_, new_n29997_, new_n29977_ );
or   ( new_n30118_, new_n30117_, new_n29987_ );
and  ( new_n30119_, new_n30118_, new_n30116_ );
or   ( new_n30120_, new_n30062_, new_n19394_ );
or   ( new_n30121_, new_n30058_, new_n19659_ );
and  ( new_n30122_, new_n30121_, new_n30120_ );
or   ( new_n30123_, new_n30024_, new_n20156_ );
or   ( new_n30124_, new_n30020_, new_n20443_ );
and  ( new_n30125_, new_n30124_, new_n30123_ );
or   ( new_n30126_, new_n30029_, new_n19394_ );
or   ( new_n30127_, new_n30027_, new_n19659_ );
and  ( new_n30128_, new_n30127_, new_n30126_ );
and  ( new_n30129_, new_n30128_, new_n30125_ );
or   ( new_n30130_, new_n30129_, new_n30053_ );
or   ( new_n30131_, new_n30038_, new_n21261_ );
or   ( new_n30132_, new_n30034_, new_n21009_ );
and  ( new_n30133_, new_n30132_, new_n30131_ );
or   ( new_n30134_, new_n30133_, new_n19394_ );
and  ( new_n30135_, new_n30133_, new_n19394_ );
or   ( new_n30136_, new_n30049_, new_n21013_ );
or   ( new_n30137_, new_n30045_, new_n21265_ );
and  ( new_n30138_, new_n30137_, new_n30136_ );
or   ( new_n30139_, new_n30138_, new_n30135_ );
and  ( new_n30140_, new_n30139_, new_n30134_ );
or   ( new_n30141_, new_n30140_, new_n30032_ );
and  ( new_n30142_, new_n30141_, new_n30130_ );
or   ( new_n30143_, new_n30142_, new_n30122_ );
or   ( new_n30144_, new_n30140_, new_n30129_ );
and  ( new_n30145_, new_n30144_, new_n30055_ );
or   ( new_n30146_, new_n30145_, new_n30064_ );
and  ( new_n30147_, new_n30146_, new_n30143_ );
or   ( new_n30148_, new_n30147_, new_n30119_ );
or   ( new_n30149_, new_n30015_, new_n29952_ );
or   ( new_n30150_, new_n30012_, new_n30008_ );
and  ( new_n30151_, new_n30150_, new_n30149_ );
or   ( new_n30152_, new_n30151_, new_n30066_ );
and  ( new_n30153_, new_n30140_, new_n30129_ );
or   ( new_n30154_, new_n30153_, new_n30122_ );
and  ( new_n30155_, new_n30154_, new_n30144_ );
or   ( new_n30156_, new_n30155_, new_n30017_ );
and  ( new_n30157_, new_n30156_, new_n30152_ );
or   ( new_n30158_, new_n30157_, new_n30148_ );
and  ( new_n30159_, new_n30157_, new_n30148_ );
or   ( new_n30160_, new_n30145_, new_n30122_ );
or   ( new_n30161_, new_n30142_, new_n30064_ );
and  ( new_n30162_, new_n30161_, new_n30160_ );
or   ( new_n30163_, new_n30162_, new_n30119_ );
or   ( new_n30164_, new_n30117_, new_n30001_ );
or   ( new_n30165_, new_n30115_, new_n29987_ );
and  ( new_n30166_, new_n30165_, new_n30164_ );
or   ( new_n30167_, new_n30166_, new_n30147_ );
and  ( new_n30168_, new_n30167_, new_n30163_ );
or   ( new_n30169_, new_n30128_, new_n30026_ );
or   ( new_n30170_, new_n30125_, new_n30031_ );
and  ( new_n30171_, new_n30170_, new_n30169_ );
nor  ( new_n30172_, new_n22333_, new_n5459_ );
nor  ( new_n30173_, new_n30172_, new_n15043_ );
or   ( new_n30174_, new_n30173_, new_n21261_ );
and  ( new_n30175_, new_n22337_, RI2b1c4342e188_92 );
and  ( new_n30176_, new_n22330_, RI2b1c4342e110_91 );
or   ( new_n30177_, new_n30176_, new_n30175_ );
or   ( new_n30178_, new_n30177_, new_n21009_ );
and  ( new_n30179_, new_n30178_, new_n30174_ );
or   ( new_n30180_, new_n21419_, new_n6321_ );
or   ( new_n30181_, new_n21424_, new_n6307_ );
and  ( new_n30182_, new_n30181_, new_n30180_ );
or   ( new_n30183_, new_n30182_, new_n21013_ );
and  ( new_n30184_, new_n21428_, RI2b1c4342e278_94 );
and  ( new_n30185_, new_n21415_, RI2b1c4342e200_93 );
or   ( new_n30186_, new_n30185_, new_n30184_ );
or   ( new_n30187_, new_n30186_, new_n21265_ );
and  ( new_n30188_, new_n30187_, new_n30183_ );
or   ( new_n30189_, new_n30188_, new_n30179_ );
and  ( new_n30190_, new_n30188_, new_n30179_ );
or   ( new_n30191_, new_n20557_, new_n7274_ );
or   ( new_n30192_, new_n20562_, new_n124_ );
and  ( new_n30193_, new_n30192_, new_n30191_ );
or   ( new_n30194_, new_n30193_, new_n20156_ );
and  ( new_n30195_, new_n20566_, RI2b1c4342e368_96 );
and  ( new_n30196_, new_n20553_, RI2b1c4342e2f0_95 );
or   ( new_n30197_, new_n30196_, new_n30195_ );
or   ( new_n30198_, new_n30197_, new_n20443_ );
and  ( new_n30199_, new_n30198_, new_n30194_ );
or   ( new_n30200_, new_n30199_, new_n30190_ );
and  ( new_n30201_, new_n30200_, new_n30189_ );
or   ( new_n30202_, new_n30201_, new_n30171_ );
or   ( new_n30203_, new_n30133_, new_n19659_ );
or   ( new_n30204_, new_n30040_, new_n19394_ );
and  ( new_n30205_, new_n30204_, new_n30203_ );
or   ( new_n30206_, new_n30205_, new_n30138_ );
and  ( new_n30207_, new_n30134_, new_n30042_ );
or   ( new_n30208_, new_n30207_, new_n30051_ );
and  ( new_n30209_, new_n30208_, new_n30206_ );
and  ( new_n30210_, new_n30201_, new_n30171_ );
or   ( new_n30211_, new_n30210_, new_n30209_ );
and  ( new_n30212_, new_n30211_, new_n30202_ );
or   ( new_n30213_, new_n30212_, new_n30168_ );
or   ( new_n30214_, new_n30213_, new_n30159_ );
and  ( new_n30215_, new_n30214_, new_n30158_ );
and  ( new_n30216_, new_n30212_, new_n30168_ );
or   ( new_n30217_, new_n30216_, new_n30159_ );
nor  ( new_n30218_, new_n22333_, new_n6321_ );
nor  ( new_n30219_, new_n30218_, new_n15191_ );
or   ( new_n30220_, new_n30219_, new_n21261_ );
and  ( new_n30221_, new_n22337_, RI2b1c4342e278_94 );
and  ( new_n30222_, new_n22330_, RI2b1c4342e200_93 );
or   ( new_n30223_, new_n30222_, new_n30221_ );
or   ( new_n30224_, new_n30223_, new_n21009_ );
and  ( new_n30225_, new_n30224_, new_n30220_ );
or   ( new_n30226_, new_n21419_, new_n7274_ );
or   ( new_n30227_, new_n21424_, new_n124_ );
and  ( new_n30228_, new_n30227_, new_n30226_ );
or   ( new_n30229_, new_n30228_, new_n21013_ );
and  ( new_n30230_, new_n21428_, RI2b1c4342e368_96 );
and  ( new_n30231_, new_n21415_, RI2b1c4342e2f0_95 );
or   ( new_n30232_, new_n30231_, new_n30230_ );
or   ( new_n30233_, new_n30232_, new_n21265_ );
and  ( new_n30234_, new_n30233_, new_n30229_ );
or   ( new_n30235_, new_n30234_, new_n30225_ );
and  ( new_n30236_, new_n21428_, RI2b1c4342e2f0_95 );
and  ( new_n30237_, new_n21415_, RI2b1c4342e278_94 );
or   ( new_n30238_, new_n30237_, new_n30236_ );
or   ( new_n30239_, new_n30238_, new_n21013_ );
or   ( new_n30240_, new_n21419_, new_n124_ );
or   ( new_n30241_, new_n21424_, new_n6321_ );
and  ( new_n30242_, new_n30241_, new_n30240_ );
or   ( new_n30243_, new_n30242_, new_n21265_ );
and  ( new_n30244_, new_n30243_, new_n30239_ );
and  ( new_n30245_, new_n22337_, RI2b1c4342e200_93 );
and  ( new_n30246_, new_n22330_, RI2b1c4342e188_92 );
or   ( new_n30247_, new_n30246_, new_n30245_ );
or   ( new_n30248_, new_n30247_, new_n21261_ );
nor  ( new_n30249_, new_n22333_, new_n6307_ );
nor  ( new_n30250_, new_n30249_, new_n15124_ );
or   ( new_n30251_, new_n30250_, new_n21009_ );
and  ( new_n30252_, new_n30251_, new_n30248_ );
or   ( new_n30253_, new_n30252_, new_n20156_ );
or   ( new_n30254_, new_n30250_, new_n21261_ );
or   ( new_n30255_, new_n30247_, new_n21009_ );
and  ( new_n30256_, new_n30255_, new_n30254_ );
or   ( new_n30257_, new_n30256_, new_n20443_ );
and  ( new_n30258_, new_n30257_, new_n30253_ );
or   ( new_n30259_, new_n30258_, new_n30244_ );
or   ( new_n30260_, new_n30242_, new_n21013_ );
or   ( new_n30261_, new_n30238_, new_n21265_ );
and  ( new_n30262_, new_n30261_, new_n30260_ );
or   ( new_n30263_, new_n30252_, new_n20443_ );
or   ( new_n30264_, new_n30256_, new_n20156_ );
and  ( new_n30265_, new_n30264_, new_n30263_ );
or   ( new_n30266_, new_n30265_, new_n30262_ );
and  ( new_n30267_, new_n30266_, new_n30259_ );
or   ( new_n30268_, new_n20562_, new_n7274_ );
or   ( new_n30269_, new_n30268_, new_n20156_ );
and  ( new_n30270_, new_n20553_, RI2b1c4342e368_96 );
or   ( new_n30271_, new_n30270_, new_n20443_ );
and  ( new_n30272_, new_n30271_, new_n30269_ );
or   ( new_n30273_, new_n30272_, new_n30267_ );
or   ( new_n30274_, new_n30270_, new_n20156_ );
or   ( new_n30275_, new_n30268_, new_n20443_ );
and  ( new_n30276_, new_n30275_, new_n30274_ );
or   ( new_n30277_, new_n30265_, new_n30244_ );
or   ( new_n30278_, new_n30262_, new_n30258_ );
and  ( new_n30279_, new_n30278_, new_n30277_ );
or   ( new_n30280_, new_n30279_, new_n30276_ );
and  ( new_n30281_, new_n30280_, new_n30273_ );
or   ( new_n30282_, new_n30281_, new_n30235_ );
nor  ( new_n30283_, new_n22333_, new_n124_ );
nor  ( new_n30284_, new_n30283_, new_n15222_ );
or   ( new_n30285_, new_n30284_, new_n21261_ );
and  ( new_n30286_, new_n22337_, RI2b1c4342e2f0_95 );
and  ( new_n30287_, new_n22330_, RI2b1c4342e278_94 );
or   ( new_n30288_, new_n30287_, new_n30286_ );
or   ( new_n30289_, new_n30288_, new_n21009_ );
and  ( new_n30290_, new_n30289_, new_n30285_ );
or   ( new_n30291_, new_n30290_, new_n21265_ );
or   ( new_n30292_, new_n30232_, new_n21013_ );
or   ( new_n30293_, new_n30228_, new_n21265_ );
and  ( new_n30294_, new_n30293_, new_n30292_ );
or   ( new_n30295_, new_n30294_, new_n30225_ );
or   ( new_n30296_, new_n30223_, new_n21261_ );
or   ( new_n30297_, new_n30219_, new_n21009_ );
and  ( new_n30298_, new_n30297_, new_n30296_ );
or   ( new_n30299_, new_n30298_, new_n30234_ );
and  ( new_n30300_, new_n30299_, new_n30295_ );
and  ( new_n30301_, new_n30300_, new_n30291_ );
or   ( new_n30302_, new_n30290_, new_n21013_ );
or   ( new_n30303_, new_n30288_, new_n21261_ );
or   ( new_n30304_, new_n30284_, new_n21009_ );
and  ( new_n30305_, new_n30304_, new_n30303_ );
or   ( new_n30306_, new_n30305_, new_n21265_ );
and  ( new_n30307_, new_n30306_, new_n30302_ );
or   ( new_n30308_, new_n21424_, new_n7274_ );
or   ( new_n30309_, new_n30308_, new_n21013_ );
and  ( new_n30310_, new_n21415_, RI2b1c4342e368_96 );
or   ( new_n30311_, new_n30310_, new_n21265_ );
and  ( new_n30312_, new_n30311_, new_n30309_ );
or   ( new_n30313_, new_n30312_, new_n30307_ );
or   ( new_n30314_, new_n30300_, new_n30291_ );
and  ( new_n30315_, new_n30314_, new_n30313_ );
or   ( new_n30316_, new_n30315_, new_n30301_ );
and  ( new_n30317_, new_n30312_, new_n30307_ );
and  ( new_n30318_, new_n22330_, RI2b1c4342e2f0_95 );
or   ( new_n30319_, new_n30318_, RI2b1c4342e368_96 );
and  ( new_n30320_, new_n7097_, new_n137_ );
or   ( new_n30321_, new_n30320_, new_n21261_ );
and  ( new_n30322_, new_n30321_, new_n30319_ );
or   ( new_n30323_, new_n30322_, new_n21009_ );
or   ( new_n30324_, new_n30323_, new_n30301_ );
or   ( new_n30325_, new_n30324_, new_n30317_ );
and  ( new_n30326_, new_n30325_, new_n30316_ );
and  ( new_n30327_, new_n30281_, new_n30235_ );
or   ( new_n30328_, new_n30327_, new_n30326_ );
and  ( new_n30329_, new_n30328_, new_n30282_ );
or   ( new_n30330_, new_n30197_, new_n20156_ );
or   ( new_n30331_, new_n30193_, new_n20443_ );
and  ( new_n30332_, new_n30331_, new_n30330_ );
or   ( new_n30333_, new_n30186_, new_n21013_ );
or   ( new_n30334_, new_n30182_, new_n21265_ );
and  ( new_n30335_, new_n30334_, new_n30333_ );
or   ( new_n30336_, new_n30335_, new_n30179_ );
or   ( new_n30337_, new_n30177_, new_n21261_ );
or   ( new_n30338_, new_n30173_, new_n21009_ );
and  ( new_n30339_, new_n30338_, new_n30337_ );
or   ( new_n30340_, new_n30339_, new_n30188_ );
and  ( new_n30341_, new_n30340_, new_n30336_ );
or   ( new_n30342_, new_n30341_, new_n30332_ );
or   ( new_n30343_, new_n30339_, new_n30335_ );
and  ( new_n30344_, new_n30343_, new_n30189_ );
or   ( new_n30345_, new_n30344_, new_n30199_ );
and  ( new_n30346_, new_n30345_, new_n30342_ );
and  ( new_n30347_, new_n30256_, new_n20443_ );
or   ( new_n30348_, new_n30347_, new_n30262_ );
and  ( new_n30349_, new_n30348_, new_n30257_ );
or   ( new_n30350_, new_n30349_, new_n30346_ );
or   ( new_n30351_, new_n30207_, new_n30138_ );
or   ( new_n30352_, new_n30205_, new_n30051_ );
and  ( new_n30353_, new_n30352_, new_n30351_ );
or   ( new_n30354_, new_n30128_, new_n30125_ );
and  ( new_n30355_, new_n30354_, new_n30032_ );
or   ( new_n30356_, new_n30355_, new_n30201_ );
and  ( new_n30357_, new_n30339_, new_n30335_ );
or   ( new_n30358_, new_n30357_, new_n30332_ );
and  ( new_n30359_, new_n30358_, new_n30343_ );
or   ( new_n30360_, new_n30359_, new_n30171_ );
and  ( new_n30361_, new_n30360_, new_n30356_ );
or   ( new_n30362_, new_n30361_, new_n30353_ );
or   ( new_n30363_, new_n30359_, new_n30355_ );
and  ( new_n30364_, new_n30363_, new_n30202_ );
or   ( new_n30365_, new_n30364_, new_n30209_ );
and  ( new_n30366_, new_n30365_, new_n30362_ );
and  ( new_n30367_, new_n30366_, new_n30350_ );
or   ( new_n30368_, new_n30279_, new_n30272_ );
or   ( new_n30369_, new_n30344_, new_n30332_ );
or   ( new_n30370_, new_n30341_, new_n30199_ );
and  ( new_n30371_, new_n30370_, new_n30369_ );
or   ( new_n30372_, new_n30371_, new_n30349_ );
and  ( new_n30373_, new_n30252_, new_n20156_ );
or   ( new_n30374_, new_n30373_, new_n30244_ );
and  ( new_n30375_, new_n30374_, new_n30253_ );
or   ( new_n30376_, new_n30375_, new_n30346_ );
and  ( new_n30377_, new_n30376_, new_n30372_ );
and  ( new_n30378_, new_n30377_, new_n30368_ );
or   ( new_n30379_, new_n30378_, new_n30367_ );
or   ( new_n30380_, new_n30379_, new_n30329_ );
or   ( new_n30381_, new_n30366_, new_n30350_ );
or   ( new_n30382_, new_n30377_, new_n30368_ );
or   ( new_n30383_, new_n30382_, new_n30367_ );
and  ( new_n30384_, new_n30383_, new_n30381_ );
and  ( new_n30385_, new_n30384_, new_n30380_ );
or   ( new_n30386_, new_n30385_, new_n30217_ );
and  ( new_n30387_, new_n30386_, new_n30215_ );
or   ( new_n30388_, new_n30387_, new_n30112_ );
or   ( new_n30389_, new_n30388_, new_n29945_ );
or   ( new_n30390_, new_n29877_, new_n29868_ );
or   ( new_n30391_, new_n29943_, new_n29934_ );
or   ( new_n30392_, new_n30391_, new_n29878_ );
and  ( new_n30393_, new_n30392_, new_n30390_ );
or   ( new_n30394_, new_n30110_, new_n30107_ );
or   ( new_n30395_, new_n30097_, new_n30067_ );
or   ( new_n30396_, new_n30395_, new_n30111_ );
and  ( new_n30397_, new_n30396_, new_n30394_ );
or   ( new_n30398_, new_n30397_, new_n29945_ );
and  ( new_n30399_, new_n30398_, new_n30393_ );
and  ( new_n30400_, new_n30399_, new_n30389_ );
or   ( new_n30401_, new_n30400_, new_n29741_ );
or   ( new_n30402_, new_n30401_, new_n29447_ );
or   ( new_n30403_, new_n29257_, new_n29160_ );
or   ( new_n30404_, new_n29445_, new_n29311_ );
and  ( new_n30405_, new_n30404_, new_n30403_ );
or   ( new_n30406_, new_n30405_, new_n29258_ );
or   ( new_n30407_, new_n29739_, new_n29736_ );
or   ( new_n30408_, new_n29720_, new_n29674_ );
and  ( new_n30409_, new_n30408_, new_n30407_ );
or   ( new_n30410_, new_n30409_, new_n29740_ );
or   ( new_n30411_, new_n30410_, new_n29447_ );
and  ( new_n30412_, new_n30411_, new_n30406_ );
and  ( new_n30413_, new_n30412_, new_n30402_ );
or   ( new_n30414_, new_n30413_, new_n29100_ );
or   ( new_n30415_, new_n30414_, new_n28882_ );
or   ( new_n30416_, new_n28650_, new_n28500_ );
or   ( new_n30417_, new_n28880_, new_n28864_ );
or   ( new_n30418_, new_n30417_, new_n28651_ );
and  ( new_n30419_, new_n30418_, new_n30416_ );
or   ( new_n30420_, new_n29098_, new_n29089_ );
or   ( new_n30421_, new_n29087_, new_n28975_ );
or   ( new_n30422_, new_n30421_, new_n29099_ );
and  ( new_n30423_, new_n30422_, new_n30420_ );
or   ( new_n30424_, new_n30423_, new_n28882_ );
and  ( new_n30425_, new_n30424_, new_n30419_ );
and  ( new_n30426_, new_n30425_, new_n30415_ );
or   ( new_n30427_, new_n30426_, new_n28402_ );
or   ( new_n30428_, new_n30427_, new_n27877_ );
or   ( new_n30429_, new_n27610_, new_n27442_ );
or   ( new_n30430_, new_n27875_, new_n27698_ );
or   ( new_n30431_, new_n30430_, new_n27611_ );
and  ( new_n30432_, new_n30431_, new_n30429_ );
or   ( new_n30433_, new_n28129_, new_n27969_ );
or   ( new_n30434_, new_n28400_, new_n28215_ );
or   ( new_n30435_, new_n30434_, new_n28130_ );
and  ( new_n30436_, new_n30435_, new_n30433_ );
or   ( new_n30437_, new_n30436_, new_n27877_ );
and  ( new_n30438_, new_n30437_, new_n30432_ );
and  ( new_n30439_, new_n30438_, new_n30428_ );
or   ( new_n30440_, new_n30439_, new_n27329_ );
and  ( new_n30441_, new_n30440_, new_n27326_ );
or   ( new_n30442_, new_n30441_, new_n26326_ );
or   ( new_n30443_, new_n30442_, new_n24747_ );
and  ( new_n30444_, new_n30443_, new_n26323_ );
and  ( new_n30445_, new_n30444_, new_n24744_ );
or   ( new_n30446_, new_n30445_, new_n23019_ );
and  ( new_n30447_, new_n30446_, new_n23016_ );
or   ( new_n30448_, new_n30447_, new_n21196_ );
and  ( new_n30449_, new_n30448_, new_n21193_ );
or   ( new_n30450_, new_n30449_, new_n19620_ );
and  ( new_n30451_, new_n30450_, new_n19617_ );
or   ( new_n30452_, new_n30451_, new_n18249_ );
and  ( new_n30453_, new_n30452_, new_n18246_ );
and  ( new_n30454_, new_n16196_, RI2b1c4342d648_68 );
and  ( new_n30455_, new_n16199_, RI2b1c4342d5d0_67 );
or   ( new_n30456_, new_n30455_, new_n30454_ );
or   ( new_n30457_, new_n30456_, new_n16186_ );
or   ( new_n30458_, new_n16208_, new_n612_ );
or   ( new_n30459_, new_n16194_, new_n112_ );
and  ( new_n30460_, new_n30459_, new_n30458_ );
or   ( new_n30461_, new_n30460_, new_n16204_ );
and  ( new_n30462_, new_n30461_, new_n30457_ );
or   ( new_n30463_, new_n16033_, new_n526_ );
or   ( new_n30464_, new_n16017_, new_n99_ );
and  ( new_n30465_, new_n30464_, new_n30463_ );
or   ( new_n30466_, new_n30465_, new_n16009_ );
and  ( new_n30467_, new_n16021_, RI2b1c4342d558_66 );
and  ( new_n30468_, new_n16024_, RI2b1c4342d4e0_65 );
or   ( new_n30469_, new_n30468_, new_n30467_ );
or   ( new_n30470_, new_n30469_, new_n16029_ );
and  ( new_n30471_, new_n30470_, new_n30466_ );
or   ( new_n30472_, new_n30471_, new_n16052_ );
or   ( new_n30473_, new_n30469_, new_n16009_ );
or   ( new_n30474_, new_n30465_, new_n16029_ );
and  ( new_n30475_, new_n30474_, new_n30473_ );
or   ( new_n30476_, new_n30475_, new_n16071_ );
and  ( new_n30477_, new_n30476_, new_n30472_ );
or   ( new_n30478_, new_n30477_, new_n30462_ );
or   ( new_n30479_, new_n30460_, new_n16186_ );
or   ( new_n30480_, new_n30456_, new_n16204_ );
and  ( new_n30481_, new_n30480_, new_n30479_ );
or   ( new_n30482_, new_n30475_, new_n16052_ );
or   ( new_n30483_, new_n30471_, new_n16071_ );
and  ( new_n30484_, new_n30483_, new_n30482_ );
or   ( new_n30485_, new_n30484_, new_n30481_ );
and  ( new_n30486_, new_n30485_, new_n30478_ );
and  ( new_n30487_, new_n16102_, RI2b1c4342d990_75 );
and  ( new_n30488_, new_n16132_, RI2b1c4342d918_74 );
and  ( new_n30489_, new_n16114_, RI2b1c4342d8a0_73 );
or   ( new_n30490_, new_n30489_, new_n30488_ );
or   ( new_n30491_, new_n30490_, new_n16108_ );
or   ( new_n30492_, new_n16119_, new_n859_ );
or   ( new_n30493_, new_n16123_, new_n105_ );
and  ( new_n30494_, new_n30493_, new_n30492_ );
or   ( new_n30495_, new_n30494_, new_n16128_ );
and  ( new_n30496_, new_n30495_, new_n30491_ );
and  ( new_n30497_, new_n16226_, RI2b1c4342d738_70 );
and  ( new_n30498_, new_n16229_, RI2b1c4342d6c0_69 );
or   ( new_n30499_, new_n30498_, new_n30497_ );
or   ( new_n30500_, new_n30499_, new_n16217_ );
or   ( new_n30501_, new_n16238_, new_n755_ );
or   ( new_n30502_, new_n16224_, new_n591_ );
and  ( new_n30503_, new_n30502_, new_n30501_ );
or   ( new_n30504_, new_n30503_, new_n16234_ );
and  ( new_n30505_, new_n30504_, new_n30500_ );
and  ( new_n30506_, new_n16162_, RI2b1c4342d828_72 );
and  ( new_n30507_, new_n16165_, RI2b1c4342d7b0_71 );
or   ( new_n30508_, new_n30507_, new_n30506_ );
or   ( new_n30509_, new_n30508_, new_n16151_ );
or   ( new_n30510_, new_n16174_, new_n806_ );
or   ( new_n30511_, new_n16160_, new_n110_ );
and  ( new_n30512_, new_n30511_, new_n30510_ );
or   ( new_n30513_, new_n30512_, new_n16170_ );
and  ( new_n30514_, new_n30513_, new_n30509_ );
or   ( new_n30515_, new_n30514_, new_n30505_ );
or   ( new_n30516_, new_n30503_, new_n16217_ );
or   ( new_n30517_, new_n30499_, new_n16234_ );
and  ( new_n30518_, new_n30517_, new_n30516_ );
or   ( new_n30519_, new_n30512_, new_n16151_ );
or   ( new_n30520_, new_n30508_, new_n16170_ );
and  ( new_n30521_, new_n30520_, new_n30519_ );
or   ( new_n30522_, new_n30521_, new_n30518_ );
and  ( new_n30523_, new_n30522_, new_n30515_ );
or   ( new_n30524_, new_n30523_, new_n30496_ );
or   ( new_n30525_, new_n30494_, new_n16108_ );
or   ( new_n30526_, new_n30490_, new_n16128_ );
and  ( new_n30527_, new_n30526_, new_n30525_ );
or   ( new_n30528_, new_n30518_, new_n30514_ );
or   ( new_n30529_, new_n30521_, new_n30505_ );
and  ( new_n30530_, new_n30529_, new_n30528_ );
or   ( new_n30531_, new_n30530_, new_n30527_ );
and  ( new_n30532_, new_n30531_, new_n30524_ );
or   ( new_n30533_, new_n30532_, new_n30487_ );
or   ( new_n30534_, new_n16115_, new_n843_ );
or   ( new_n30535_, new_n30530_, new_n30496_ );
or   ( new_n30536_, new_n30527_, new_n30523_ );
and  ( new_n30537_, new_n30536_, new_n30535_ );
or   ( new_n30538_, new_n30537_, new_n30534_ );
and  ( new_n30539_, new_n30538_, new_n30533_ );
or   ( new_n30540_, new_n30539_, new_n30486_ );
or   ( new_n30541_, new_n30484_, new_n30462_ );
or   ( new_n30542_, new_n30481_, new_n30477_ );
and  ( new_n30543_, new_n30542_, new_n30541_ );
or   ( new_n30544_, new_n30534_, new_n30532_ );
or   ( new_n30545_, new_n30537_, new_n30487_ );
and  ( new_n30546_, new_n30545_, new_n30544_ );
or   ( new_n30547_, new_n30546_, new_n30543_ );
and  ( new_n30548_, new_n30547_, new_n30540_ );
and  ( new_n30549_, new_n17059_, new_n17056_ );
or   ( new_n30550_, new_n30549_, new_n17053_ );
and  ( new_n30551_, new_n30550_, new_n17060_ );
and  ( new_n30552_, new_n17012_, new_n16967_ );
or   ( new_n30553_, new_n30552_, new_n16966_ );
and  ( new_n30554_, new_n30553_, new_n17013_ );
or   ( new_n30555_, new_n30554_, new_n30551_ );
and  ( new_n30556_, new_n17017_, new_n17014_ );
or   ( new_n30557_, new_n30556_, new_n17023_ );
and  ( new_n30558_, new_n30557_, new_n17018_ );
and  ( new_n30559_, new_n17066_, new_n17063_ );
and  ( new_n30560_, new_n17067_, new_n16139_ );
or   ( new_n30561_, new_n30560_, new_n30559_ );
or   ( new_n30562_, new_n30561_, new_n30558_ );
and  ( new_n30563_, new_n30562_, new_n30555_ );
or   ( new_n30564_, new_n30563_, new_n30548_ );
or   ( new_n30565_, new_n30546_, new_n30486_ );
or   ( new_n30566_, new_n30543_, new_n30539_ );
and  ( new_n30567_, new_n30566_, new_n30565_ );
or   ( new_n30568_, new_n30561_, new_n30554_ );
or   ( new_n30569_, new_n30558_, new_n30551_ );
and  ( new_n30570_, new_n30569_, new_n30568_ );
or   ( new_n30571_, new_n30570_, new_n30567_ );
and  ( new_n30572_, new_n30571_, new_n30564_ );
and  ( new_n30573_, new_n16948_, new_n16939_ );
or   ( new_n30574_, new_n30573_, new_n16934_ );
and  ( new_n30575_, new_n30574_, new_n16949_ );
and  ( new_n30576_, new_n16994_, new_n16985_ );
or   ( new_n30577_, new_n30576_, new_n16976_ );
and  ( new_n30578_, new_n30577_, new_n16995_ );
or   ( new_n30579_, new_n30578_, new_n30575_ );
and  ( new_n30580_, new_n16955_, new_n16952_ );
or   ( new_n30581_, new_n30580_, new_n16961_ );
and  ( new_n30582_, new_n30581_, new_n16956_ );
and  ( new_n30583_, new_n17001_, new_n16998_ );
or   ( new_n30584_, new_n30583_, new_n17007_ );
and  ( new_n30585_, new_n30584_, new_n17002_ );
or   ( new_n30586_, new_n30585_, new_n30582_ );
and  ( new_n30587_, new_n30586_, new_n30579_ );
or   ( new_n30588_, new_n30587_, new_n17014_ );
or   ( new_n30589_, new_n30582_, new_n30578_ );
or   ( new_n30590_, new_n30585_, new_n30575_ );
and  ( new_n30591_, new_n30590_, new_n30589_ );
or   ( new_n30592_, new_n30591_, new_n16967_ );
and  ( new_n30593_, new_n30592_, new_n30588_ );
and  ( new_n30594_, new_n17041_, new_n17038_ );
or   ( new_n30595_, new_n30594_, new_n17047_ );
and  ( new_n30596_, new_n30595_, new_n17042_ );
or   ( new_n30597_, new_n30596_, new_n30593_ );
and  ( new_n30598_, new_n17034_, new_n17031_ );
or   ( new_n30599_, new_n30598_, new_n17028_ );
and  ( new_n30600_, new_n30599_, new_n17035_ );
or   ( new_n30601_, new_n30591_, new_n17014_ );
or   ( new_n30602_, new_n30587_, new_n16967_ );
and  ( new_n30603_, new_n30602_, new_n30601_ );
or   ( new_n30604_, new_n30603_, new_n30600_ );
and  ( new_n30605_, new_n30604_, new_n30597_ );
or   ( new_n30606_, new_n30605_, new_n30572_ );
or   ( new_n30607_, new_n30570_, new_n30548_ );
or   ( new_n30608_, new_n30567_, new_n30563_ );
and  ( new_n30609_, new_n30608_, new_n30607_ );
or   ( new_n30610_, new_n30600_, new_n30593_ );
or   ( new_n30611_, new_n30603_, new_n30596_ );
and  ( new_n30612_, new_n30611_, new_n30610_ );
or   ( new_n30613_, new_n30612_, new_n30609_ );
and  ( new_n30614_, new_n30613_, new_n30606_ );
and  ( new_n30615_, new_n17084_, new_n17081_ );
and  ( new_n30616_, new_n17090_, new_n17085_ );
or   ( new_n30617_, new_n30616_, new_n30615_ );
or   ( new_n30618_, new_n30617_, new_n30614_ );
or   ( new_n30619_, new_n30612_, new_n30572_ );
or   ( new_n30620_, new_n30609_, new_n30605_ );
and  ( new_n30621_, new_n30620_, new_n30619_ );
and  ( new_n30622_, new_n17077_, new_n17074_ );
or   ( new_n30623_, new_n30622_, new_n17052_ );
and  ( new_n30624_, new_n30623_, new_n17078_ );
or   ( new_n30625_, new_n30624_, new_n30621_ );
and  ( new_n30626_, new_n30625_, new_n30618_ );
and  ( new_n30627_, new_n17102_, new_n17095_ );
or   ( new_n30628_, new_n30627_, new_n30626_ );
or   ( new_n30629_, new_n17105_, new_n17098_ );
or   ( new_n30630_, new_n30621_, new_n30617_ );
or   ( new_n30631_, new_n30624_, new_n30614_ );
and  ( new_n30632_, new_n30631_, new_n30630_ );
or   ( new_n30633_, new_n30632_, new_n30629_ );
and  ( new_n30634_, new_n30633_, new_n30628_ );
or   ( new_n30635_, new_n30634_, new_n30453_ );
and  ( new_n30636_, new_n30627_, new_n30626_ );
and  ( new_n30637_, new_n30632_, new_n30629_ );
or   ( new_n30638_, new_n30637_, new_n30636_ );
or   ( new_n30639_, new_n17102_, new_n17095_ );
and  ( new_n30640_, new_n30639_, new_n30629_ );
and  ( new_n30641_, new_n17183_, new_n17112_ );
or   ( new_n30642_, new_n30641_, new_n30640_ );
or   ( new_n30643_, new_n17183_, new_n17112_ );
and  ( new_n30644_, new_n30643_, new_n16925_ );
and  ( new_n30645_, new_n17914_, new_n17910_ );
or   ( new_n30646_, new_n30645_, new_n17907_ );
and  ( new_n30647_, new_n30646_, new_n17918_ );
and  ( new_n30648_, new_n30647_, new_n30644_ );
and  ( new_n30649_, new_n30641_, new_n30640_ );
or   ( new_n30650_, new_n30649_, new_n30648_ );
and  ( new_n30651_, new_n30650_, new_n30642_ );
or   ( new_n30652_, new_n30647_, new_n30644_ );
and  ( new_n30653_, new_n30652_, new_n30642_ );
or   ( new_n30654_, new_n17919_, new_n17907_ );
or   ( new_n30655_, new_n17916_, new_n17594_ );
and  ( new_n30656_, new_n30655_, new_n30654_ );
and  ( new_n30657_, new_n18239_, new_n18235_ );
or   ( new_n30658_, new_n30657_, new_n30656_ );
and  ( new_n30659_, new_n30657_, new_n30656_ );
or   ( new_n30660_, new_n18239_, new_n18235_ );
and  ( new_n30661_, new_n30660_, new_n17904_ );
and  ( new_n30662_, new_n18585_, new_n18581_ );
and  ( new_n30663_, new_n30662_, new_n30661_ );
or   ( new_n30664_, new_n30663_, new_n30659_ );
and  ( new_n30665_, new_n30664_, new_n30658_ );
and  ( new_n30666_, new_n30665_, new_n30653_ );
or   ( new_n30667_, new_n30666_, new_n30651_ );
or   ( new_n30668_, new_n30662_, new_n30661_ );
and  ( new_n30669_, new_n30668_, new_n30658_ );
and  ( new_n30670_, new_n30669_, new_n30653_ );
or   ( new_n30671_, new_n18585_, new_n18581_ );
and  ( new_n30672_, new_n30671_, new_n18232_ );
and  ( new_n30673_, new_n18917_, new_n18913_ );
or   ( new_n30674_, new_n30673_, new_n30672_ );
and  ( new_n30675_, new_n30673_, new_n30672_ );
or   ( new_n30676_, new_n18917_, new_n18913_ );
and  ( new_n30677_, new_n30676_, new_n18578_ );
and  ( new_n30678_, new_n19264_, new_n19260_ );
and  ( new_n30679_, new_n30678_, new_n30677_ );
or   ( new_n30680_, new_n30679_, new_n30675_ );
and  ( new_n30681_, new_n30680_, new_n30674_ );
or   ( new_n30682_, new_n19264_, new_n19260_ );
and  ( new_n30683_, new_n30682_, new_n18910_ );
and  ( new_n30684_, new_n19608_, new_n19604_ );
or   ( new_n30685_, new_n30684_, new_n30683_ );
and  ( new_n30686_, new_n30684_, new_n30683_ );
or   ( new_n30687_, new_n19608_, new_n19604_ );
and  ( new_n30688_, new_n30687_, new_n19257_ );
and  ( new_n30689_, new_n19991_, new_n19987_ );
and  ( new_n30690_, new_n30689_, new_n30688_ );
or   ( new_n30691_, new_n30690_, new_n30686_ );
and  ( new_n30692_, new_n30691_, new_n30685_ );
or   ( new_n30693_, new_n30678_, new_n30677_ );
and  ( new_n30694_, new_n30693_, new_n30674_ );
and  ( new_n30695_, new_n30694_, new_n30692_ );
or   ( new_n30696_, new_n30695_, new_n30681_ );
or   ( new_n30697_, new_n30689_, new_n30688_ );
and  ( new_n30698_, new_n30697_, new_n30685_ );
and  ( new_n30699_, new_n30698_, new_n30694_ );
or   ( new_n30700_, new_n19991_, new_n19987_ );
and  ( new_n30701_, new_n30700_, new_n19601_ );
and  ( new_n30702_, new_n20116_, new_n19998_ );
or   ( new_n30703_, new_n30702_, new_n30701_ );
and  ( new_n30704_, new_n30702_, new_n30701_ );
or   ( new_n30705_, new_n20116_, new_n19998_ );
and  ( new_n30706_, new_n30705_, new_n19984_ );
and  ( new_n30707_, new_n20784_, new_n20780_ );
or   ( new_n30708_, new_n30707_, new_n20777_ );
and  ( new_n30709_, new_n30708_, new_n20788_ );
and  ( new_n30710_, new_n30709_, new_n30706_ );
or   ( new_n30711_, new_n30710_, new_n30704_ );
and  ( new_n30712_, new_n30711_, new_n30703_ );
or   ( new_n30713_, new_n30709_, new_n30706_ );
and  ( new_n30714_, new_n30713_, new_n30703_ );
or   ( new_n30715_, new_n20789_, new_n20777_ );
or   ( new_n30716_, new_n20786_, new_n20367_ );
and  ( new_n30717_, new_n30716_, new_n30715_ );
and  ( new_n30718_, new_n20928_, new_n20796_ );
or   ( new_n30719_, new_n30718_, new_n30717_ );
and  ( new_n30720_, new_n30718_, new_n30717_ );
or   ( new_n30721_, new_n20928_, new_n20796_ );
and  ( new_n30722_, new_n30721_, new_n20774_ );
and  ( new_n30723_, new_n21323_, new_n21202_ );
or   ( new_n30724_, new_n30723_, new_n21199_ );
and  ( new_n30725_, new_n30724_, new_n21327_ );
and  ( new_n30726_, new_n30725_, new_n30722_ );
or   ( new_n30727_, new_n30726_, new_n30720_ );
and  ( new_n30728_, new_n30727_, new_n30719_ );
and  ( new_n30729_, new_n30728_, new_n30714_ );
or   ( new_n30730_, new_n30729_, new_n30712_ );
or   ( new_n30731_, new_n30725_, new_n30722_ );
and  ( new_n30732_, new_n30731_, new_n30719_ );
and  ( new_n30733_, new_n30732_, new_n30714_ );
or   ( new_n30734_, new_n21328_, new_n21199_ );
or   ( new_n30735_, new_n21325_, new_n21185_ );
and  ( new_n30736_, new_n30735_, new_n30734_ );
and  ( new_n30737_, new_n21817_, new_n21667_ );
or   ( new_n30738_, new_n30737_, new_n21660_ );
and  ( new_n30739_, new_n30738_, new_n21821_ );
or   ( new_n30740_, new_n30739_, new_n30736_ );
and  ( new_n30741_, new_n30739_, new_n30736_ );
or   ( new_n30742_, new_n21822_, new_n21660_ );
or   ( new_n30743_, new_n21819_, new_n21653_ );
and  ( new_n30744_, new_n30743_, new_n30742_ );
and  ( new_n30745_, new_n22237_, new_n22107_ );
or   ( new_n30746_, new_n30745_, new_n22105_ );
and  ( new_n30747_, new_n30746_, new_n22241_ );
and  ( new_n30748_, new_n30747_, new_n30744_ );
or   ( new_n30749_, new_n30748_, new_n30741_ );
and  ( new_n30750_, new_n30749_, new_n30740_ );
or   ( new_n30751_, new_n30747_, new_n30744_ );
and  ( new_n30752_, new_n30751_, new_n30740_ );
or   ( new_n30753_, new_n22242_, new_n22105_ );
or   ( new_n30754_, new_n22239_, new_n22094_ );
and  ( new_n30755_, new_n30754_, new_n30753_ );
and  ( new_n30756_, new_n22720_, new_n22574_ );
or   ( new_n30757_, new_n30756_, new_n22567_ );
and  ( new_n30758_, new_n30757_, new_n22724_ );
or   ( new_n30759_, new_n30758_, new_n30755_ );
and  ( new_n30760_, new_n30758_, new_n30755_ );
or   ( new_n30761_, new_n22725_, new_n22567_ );
or   ( new_n30762_, new_n22722_, new_n22560_ );
and  ( new_n30763_, new_n30762_, new_n30761_ );
and  ( new_n30764_, new_n23158_, new_n23024_ );
or   ( new_n30765_, new_n30764_, new_n23022_ );
and  ( new_n30766_, new_n30765_, new_n23162_ );
and  ( new_n30767_, new_n30766_, new_n30763_ );
or   ( new_n30768_, new_n30767_, new_n30760_ );
and  ( new_n30769_, new_n30768_, new_n30759_ );
and  ( new_n30770_, new_n30769_, new_n30752_ );
or   ( new_n30771_, new_n30770_, new_n30750_ );
or   ( new_n30772_, new_n30766_, new_n30763_ );
and  ( new_n30773_, new_n30772_, new_n30759_ );
and  ( new_n30774_, new_n30773_, new_n30752_ );
or   ( new_n30775_, new_n23163_, new_n23022_ );
or   ( new_n30776_, new_n23160_, new_n23008_ );
and  ( new_n30777_, new_n30776_, new_n30775_ );
and  ( new_n30778_, new_n23592_, new_n23458_ );
or   ( new_n30779_, new_n30778_, new_n23455_ );
and  ( new_n30780_, new_n30779_, new_n23596_ );
or   ( new_n30781_, new_n30780_, new_n30777_ );
and  ( new_n30782_, new_n30780_, new_n30777_ );
or   ( new_n30783_, new_n23597_, new_n23455_ );
or   ( new_n30784_, new_n23594_, new_n23448_ );
and  ( new_n30785_, new_n30784_, new_n30783_ );
and  ( new_n30786_, new_n24083_, new_n23930_ );
or   ( new_n30787_, new_n30786_, new_n23927_ );
and  ( new_n30788_, new_n30787_, new_n24087_ );
and  ( new_n30789_, new_n30788_, new_n30785_ );
or   ( new_n30790_, new_n30789_, new_n30782_ );
and  ( new_n30791_, new_n30790_, new_n30781_ );
or   ( new_n30792_, new_n30788_, new_n30785_ );
and  ( new_n30793_, new_n30792_, new_n30781_ );
or   ( new_n30794_, new_n24088_, new_n23927_ );
or   ( new_n30795_, new_n24085_, new_n23916_ );
and  ( new_n30796_, new_n30795_, new_n30794_ );
and  ( new_n30797_, new_n24492_, new_n24367_ );
or   ( new_n30798_, new_n30797_, new_n24364_ );
and  ( new_n30799_, new_n30798_, new_n24496_ );
or   ( new_n30800_, new_n30799_, new_n30796_ );
and  ( new_n30801_, new_n30799_, new_n30796_ );
or   ( new_n30802_, new_n24497_, new_n24364_ );
or   ( new_n30803_, new_n24494_, new_n24357_ );
and  ( new_n30804_, new_n30803_, new_n30802_ );
and  ( new_n30805_, new_n24866_, new_n24753_ );
or   ( new_n30806_, new_n30805_, new_n24750_ );
and  ( new_n30807_, new_n30806_, new_n24870_ );
and  ( new_n30808_, new_n30807_, new_n30804_ );
or   ( new_n30809_, new_n30808_, new_n30801_ );
and  ( new_n30810_, new_n30809_, new_n30800_ );
and  ( new_n30811_, new_n30810_, new_n30793_ );
or   ( new_n30812_, new_n30811_, new_n30791_ );
or   ( new_n30813_, new_n30807_, new_n30804_ );
and  ( new_n30814_, new_n30813_, new_n30800_ );
and  ( new_n30815_, new_n30814_, new_n30793_ );
or   ( new_n30816_, new_n24871_, new_n24750_ );
or   ( new_n30817_, new_n24868_, new_n24736_ );
and  ( new_n30818_, new_n30817_, new_n30816_ );
and  ( new_n30819_, new_n25287_, new_n25162_ );
or   ( new_n30820_, new_n30819_, new_n25155_ );
and  ( new_n30821_, new_n30820_, new_n25291_ );
or   ( new_n30822_, new_n30821_, new_n30818_ );
and  ( new_n30823_, new_n30821_, new_n30818_ );
or   ( new_n30824_, new_n25292_, new_n25155_ );
or   ( new_n30825_, new_n25289_, new_n25148_ );
and  ( new_n30826_, new_n30825_, new_n30824_ );
and  ( new_n30827_, new_n25655_, new_n25542_ );
or   ( new_n30828_, new_n30827_, new_n25540_ );
and  ( new_n30829_, new_n30828_, new_n25659_ );
and  ( new_n30830_, new_n30829_, new_n30826_ );
or   ( new_n30831_, new_n30830_, new_n30823_ );
and  ( new_n30832_, new_n30831_, new_n30822_ );
or   ( new_n30833_, new_n30829_, new_n30826_ );
and  ( new_n30834_, new_n30833_, new_n30822_ );
or   ( new_n30835_, new_n25660_, new_n25540_ );
or   ( new_n30836_, new_n25657_, new_n25529_ );
and  ( new_n30837_, new_n30836_, new_n30835_ );
and  ( new_n30838_, new_n26072_, new_n25947_ );
or   ( new_n30839_, new_n30838_, new_n25940_ );
and  ( new_n30840_, new_n30839_, new_n26076_ );
or   ( new_n30841_, new_n30840_, new_n30837_ );
and  ( new_n30842_, new_n30840_, new_n30837_ );
or   ( new_n30843_, new_n26077_, new_n25940_ );
or   ( new_n30844_, new_n26074_, new_n25933_ );
and  ( new_n30845_, new_n30844_, new_n30843_ );
and  ( new_n30846_, new_n26669_, new_n26665_ );
or   ( new_n30847_, new_n30846_, new_n26663_ );
and  ( new_n30848_, new_n30847_, new_n26673_ );
and  ( new_n30849_, new_n30848_, new_n30845_ );
or   ( new_n30850_, new_n30849_, new_n30842_ );
and  ( new_n30851_, new_n30850_, new_n30841_ );
and  ( new_n30852_, new_n30851_, new_n30834_ );
or   ( new_n30853_, new_n30852_, new_n30832_ );
and  ( new_n30854_, new_n30853_, new_n30815_ );
or   ( new_n30855_, new_n30848_, new_n30845_ );
and  ( new_n30856_, new_n30855_, new_n30841_ );
and  ( new_n30857_, new_n30856_, new_n30834_ );
or   ( new_n30858_, new_n26674_, new_n26663_ );
or   ( new_n30859_, new_n26671_, new_n26314_ );
and  ( new_n30860_, new_n30859_, new_n30858_ );
and  ( new_n30861_, new_n26805_, new_n26801_ );
or   ( new_n30862_, new_n30861_, new_n30860_ );
and  ( new_n30863_, new_n30861_, new_n30860_ );
or   ( new_n30864_, new_n26805_, new_n26801_ );
and  ( new_n30865_, new_n30864_, new_n26660_ );
and  ( new_n30866_, new_n26819_, new_n26815_ );
and  ( new_n30867_, new_n30866_, new_n30865_ );
or   ( new_n30868_, new_n30867_, new_n30863_ );
and  ( new_n30869_, new_n30868_, new_n30862_ );
or   ( new_n30870_, new_n30866_, new_n30865_ );
and  ( new_n30871_, new_n30870_, new_n30862_ );
or   ( new_n30872_, new_n26819_, new_n26815_ );
and  ( new_n30873_, new_n30872_, new_n26798_ );
and  ( new_n30874_, new_n27099_, new_n27012_ );
or   ( new_n30875_, new_n30874_, new_n27010_ );
and  ( new_n30876_, new_n30875_, new_n27103_ );
or   ( new_n30877_, new_n30876_, new_n30873_ );
and  ( new_n30878_, new_n30876_, new_n30873_ );
or   ( new_n30879_, new_n27104_, new_n27010_ );
or   ( new_n30880_, new_n27101_, new_n27002_ );
and  ( new_n30881_, new_n30880_, new_n30879_ );
and  ( new_n30882_, new_n27435_, new_n27335_ );
or   ( new_n30883_, new_n30882_, new_n27332_ );
and  ( new_n30884_, new_n30883_, new_n27439_ );
and  ( new_n30885_, new_n30884_, new_n30881_ );
or   ( new_n30886_, new_n30885_, new_n30878_ );
and  ( new_n30887_, new_n30886_, new_n30877_ );
and  ( new_n30888_, new_n30887_, new_n30871_ );
or   ( new_n30889_, new_n30888_, new_n30869_ );
or   ( new_n30890_, new_n30884_, new_n30881_ );
and  ( new_n30891_, new_n30890_, new_n30877_ );
and  ( new_n30892_, new_n30891_, new_n30871_ );
or   ( new_n30893_, new_n27440_, new_n27332_ );
or   ( new_n30894_, new_n27437_, new_n27319_ );
and  ( new_n30895_, new_n30894_, new_n30893_ );
and  ( new_n30896_, new_n27691_, new_n27617_ );
or   ( new_n30897_, new_n30896_, new_n27614_ );
and  ( new_n30898_, new_n30897_, new_n27695_ );
or   ( new_n30899_, new_n30898_, new_n30895_ );
or   ( new_n30900_, new_n27696_, new_n27614_ );
or   ( new_n30901_, new_n27693_, new_n27607_ );
and  ( new_n30902_, new_n30901_, new_n30900_ );
and  ( new_n30903_, new_n27962_, new_n27887_ );
or   ( new_n30904_, new_n30903_, new_n27880_ );
and  ( new_n30905_, new_n30904_, new_n27966_ );
or   ( new_n30906_, new_n30905_, new_n30902_ );
and  ( new_n30907_, new_n30906_, new_n30899_ );
or   ( new_n30908_, new_n27967_, new_n27880_ );
or   ( new_n30909_, new_n27964_, new_n27873_ );
and  ( new_n30910_, new_n30909_, new_n30908_ );
and  ( new_n30911_, new_n28208_, new_n28135_ );
or   ( new_n30912_, new_n30911_, new_n28133_ );
and  ( new_n30913_, new_n30912_, new_n28212_ );
or   ( new_n30914_, new_n30913_, new_n30910_ );
or   ( new_n30915_, new_n28213_, new_n28133_ );
or   ( new_n30916_, new_n28210_, new_n28126_ );
and  ( new_n30917_, new_n30916_, new_n30915_ );
and  ( new_n30918_, new_n28493_, new_n28412_ );
or   ( new_n30919_, new_n30918_, new_n28405_ );
and  ( new_n30920_, new_n30919_, new_n28497_ );
or   ( new_n30921_, new_n30920_, new_n30917_ );
and  ( new_n30922_, new_n30921_, new_n30914_ );
or   ( new_n30923_, new_n28498_, new_n28405_ );
or   ( new_n30924_, new_n28495_, new_n28398_ );
and  ( new_n30925_, new_n30924_, new_n30923_ );
and  ( new_n30926_, new_n28873_, new_n28869_ );
or   ( new_n30927_, new_n30926_, new_n28867_ );
and  ( new_n30928_, new_n30927_, new_n28877_ );
or   ( new_n30929_, new_n30928_, new_n30925_ );
or   ( new_n30930_, new_n28878_, new_n28867_ );
or   ( new_n30931_, new_n28875_, new_n28647_ );
and  ( new_n30932_, new_n30931_, new_n30930_ );
and  ( new_n30933_, new_n29096_, new_n29092_ );
or   ( new_n30934_, new_n30933_, new_n30932_ );
and  ( new_n30935_, new_n30934_, new_n30929_ );
or   ( new_n30936_, new_n28973_, new_n28966_ );
and  ( new_n30937_, new_n30936_, new_n29089_ );
and  ( new_n30938_, new_n29153_, new_n29105_ );
or   ( new_n30939_, new_n30938_, new_n29103_ );
and  ( new_n30940_, new_n30939_, new_n29157_ );
or   ( new_n30941_, new_n30940_, new_n30937_ );
or   ( new_n30942_, new_n29096_, new_n29092_ );
and  ( new_n30943_, new_n30942_, new_n28864_ );
and  ( new_n30944_, new_n28973_, new_n28966_ );
or   ( new_n30945_, new_n30944_, new_n30943_ );
and  ( new_n30946_, new_n30945_, new_n30941_ );
or   ( new_n30947_, new_n29158_, new_n29103_ );
or   ( new_n30948_, new_n29155_, new_n29084_ );
and  ( new_n30949_, new_n30948_, new_n30947_ );
and  ( new_n30950_, new_n29304_, new_n29264_ );
or   ( new_n30951_, new_n30950_, new_n29261_ );
and  ( new_n30952_, new_n30951_, new_n29308_ );
or   ( new_n30953_, new_n30952_, new_n30949_ );
or   ( new_n30954_, new_n29309_, new_n29261_ );
or   ( new_n30955_, new_n29306_, new_n29255_ );
and  ( new_n30956_, new_n30955_, new_n30954_ );
and  ( new_n30957_, new_n29729_, new_n29725_ );
or   ( new_n30958_, new_n30957_, new_n29724_ );
and  ( new_n30959_, new_n30958_, new_n29733_ );
or   ( new_n30960_, new_n30959_, new_n30956_ );
and  ( new_n30961_, new_n30960_, new_n30953_ );
or   ( new_n30962_, new_n29715_, new_n29691_ );
or   ( new_n30963_, new_n29718_, new_n29711_ );
and  ( new_n30964_, new_n30963_, new_n30962_ );
and  ( new_n30965_, new_n29875_, new_n29871_ );
or   ( new_n30966_, new_n30965_, new_n30964_ );
or   ( new_n30967_, new_n29734_, new_n29724_ );
or   ( new_n30968_, new_n29731_, new_n29442_ );
and  ( new_n30969_, new_n30968_, new_n30967_ );
and  ( new_n30970_, new_n29706_, new_n29699_ );
or   ( new_n30971_, new_n30970_, new_n29691_ );
and  ( new_n30972_, new_n30971_, new_n29713_ );
or   ( new_n30973_, new_n30972_, new_n30969_ );
and  ( new_n30974_, new_n30973_, new_n30966_ );
or   ( new_n30975_, new_n29875_, new_n29871_ );
and  ( new_n30976_, new_n30975_, new_n29674_ );
and  ( new_n30977_, new_n29941_, new_n29937_ );
or   ( new_n30978_, new_n30977_, new_n30976_ );
or   ( new_n30979_, new_n29941_, new_n29937_ );
and  ( new_n30980_, new_n30979_, new_n29868_ );
and  ( new_n30981_, new_n30105_, new_n30101_ );
or   ( new_n30982_, new_n30981_, new_n30980_ );
and  ( new_n30983_, new_n30982_, new_n30978_ );
or   ( new_n30984_, new_n30092_, new_n30074_ );
or   ( new_n30985_, new_n30095_, new_n30088_ );
and  ( new_n30986_, new_n30985_, new_n30984_ );
and  ( new_n30987_, new_n30155_, new_n30151_ );
or   ( new_n30988_, new_n30987_, new_n30986_ );
or   ( new_n30989_, new_n30105_, new_n30101_ );
and  ( new_n30990_, new_n30989_, new_n29934_ );
and  ( new_n30991_, new_n30083_, new_n30076_ );
or   ( new_n30992_, new_n30991_, new_n30074_ );
and  ( new_n30993_, new_n30992_, new_n30090_ );
or   ( new_n30994_, new_n30993_, new_n30990_ );
and  ( new_n30995_, new_n30994_, new_n30988_ );
or   ( new_n30996_, new_n30155_, new_n30151_ );
and  ( new_n30997_, new_n30996_, new_n30067_ );
and  ( new_n30998_, new_n30166_, new_n30162_ );
or   ( new_n30999_, new_n30998_, new_n30997_ );
and  ( new_n31000_, new_n30998_, new_n30997_ );
or   ( new_n31001_, new_n30166_, new_n30162_ );
and  ( new_n31002_, new_n31001_, new_n30148_ );
and  ( new_n31003_, new_n30359_, new_n30355_ );
or   ( new_n31004_, new_n31003_, new_n30353_ );
and  ( new_n31005_, new_n31004_, new_n30363_ );
and  ( new_n31006_, new_n31005_, new_n31002_ );
or   ( new_n31007_, new_n31006_, new_n31000_ );
and  ( new_n31008_, new_n31007_, new_n30999_ );
or   ( new_n31009_, new_n31005_, new_n31002_ );
and  ( new_n31010_, new_n31009_, new_n30999_ );
or   ( new_n31011_, new_n30364_, new_n30353_ );
or   ( new_n31012_, new_n30361_, new_n30209_ );
and  ( new_n31013_, new_n31012_, new_n31011_ );
and  ( new_n31014_, new_n30375_, new_n30371_ );
or   ( new_n31015_, new_n31014_, new_n31013_ );
and  ( new_n31016_, new_n31014_, new_n31013_ );
or   ( new_n31017_, new_n30375_, new_n30371_ );
and  ( new_n31018_, new_n31017_, new_n30350_ );
and  ( new_n31019_, new_n30276_, new_n30267_ );
and  ( new_n31020_, new_n31019_, new_n31018_ );
or   ( new_n31021_, new_n31020_, new_n31016_ );
and  ( new_n31022_, new_n31021_, new_n31015_ );
or   ( new_n31023_, new_n30276_, new_n30267_ );
and  ( new_n31024_, new_n31023_, new_n30368_ );
and  ( new_n31025_, new_n30298_, new_n30294_ );
and  ( new_n31026_, new_n31025_, new_n31024_ );
or   ( new_n31027_, new_n30298_, new_n30294_ );
and  ( new_n31028_, new_n31027_, new_n30235_ );
and  ( new_n31029_, new_n30305_, new_n21013_ );
or   ( new_n31030_, new_n31029_, new_n31028_ );
or   ( new_n31031_, new_n30305_, new_n21013_ );
and  ( new_n31032_, new_n31031_, new_n30291_ );
or   ( new_n31033_, new_n30310_, new_n21013_ );
or   ( new_n31034_, new_n30308_, new_n21265_ );
and  ( new_n31035_, new_n31034_, new_n31033_ );
and  ( new_n31036_, new_n31035_, new_n31032_ );
and  ( new_n31037_, new_n31029_, new_n31028_ );
or   ( new_n31038_, new_n31037_, new_n31036_ );
and  ( new_n31039_, new_n31038_, new_n31030_ );
or   ( new_n31040_, new_n31035_, new_n31032_ );
nor  ( new_n31041_, new_n22333_, new_n7274_ );
nor  ( new_n31042_, new_n31041_, new_n15247_ );
or   ( new_n31043_, new_n31042_, new_n21009_ );
and  ( new_n31044_, new_n31043_, new_n21261_ );
and  ( new_n31045_, new_n31044_, new_n31030_ );
and  ( new_n31046_, new_n31045_, new_n31040_ );
or   ( new_n31047_, new_n31046_, new_n31039_ );
or   ( new_n31048_, new_n31047_, new_n31026_ );
or   ( new_n31049_, new_n31019_, new_n31018_ );
or   ( new_n31050_, new_n31025_, new_n31024_ );
and  ( new_n31051_, new_n31050_, new_n31049_ );
and  ( new_n31052_, new_n31051_, new_n31015_ );
and  ( new_n31053_, new_n31052_, new_n31048_ );
or   ( new_n31054_, new_n31053_, new_n31022_ );
and  ( new_n31055_, new_n31054_, new_n31010_ );
or   ( new_n31056_, new_n31055_, new_n31008_ );
and  ( new_n31057_, new_n31056_, new_n30995_ );
and  ( new_n31058_, new_n31057_, new_n30983_ );
and  ( new_n31059_, new_n30977_, new_n30976_ );
and  ( new_n31060_, new_n30981_, new_n30980_ );
or   ( new_n31061_, new_n31060_, new_n31059_ );
and  ( new_n31062_, new_n31061_, new_n30978_ );
and  ( new_n31063_, new_n30993_, new_n30990_ );
and  ( new_n31064_, new_n30987_, new_n30986_ );
or   ( new_n31065_, new_n31064_, new_n31063_ );
and  ( new_n31066_, new_n31065_, new_n30994_ );
and  ( new_n31067_, new_n31066_, new_n30983_ );
or   ( new_n31068_, new_n31067_, new_n31062_ );
or   ( new_n31069_, new_n31068_, new_n31058_ );
and  ( new_n31070_, new_n31069_, new_n30974_ );
and  ( new_n31071_, new_n31070_, new_n30961_ );
and  ( new_n31072_, new_n30952_, new_n30949_ );
and  ( new_n31073_, new_n30959_, new_n30956_ );
or   ( new_n31074_, new_n31073_, new_n31072_ );
and  ( new_n31075_, new_n31074_, new_n30953_ );
and  ( new_n31076_, new_n30972_, new_n30969_ );
and  ( new_n31077_, new_n30965_, new_n30964_ );
or   ( new_n31078_, new_n31077_, new_n31076_ );
and  ( new_n31079_, new_n31078_, new_n30973_ );
and  ( new_n31080_, new_n31079_, new_n30961_ );
or   ( new_n31081_, new_n31080_, new_n31075_ );
or   ( new_n31082_, new_n31081_, new_n31071_ );
and  ( new_n31083_, new_n31082_, new_n30946_ );
and  ( new_n31084_, new_n31083_, new_n30935_ );
and  ( new_n31085_, new_n30928_, new_n30925_ );
and  ( new_n31086_, new_n30933_, new_n30932_ );
or   ( new_n31087_, new_n31086_, new_n31085_ );
and  ( new_n31088_, new_n31087_, new_n30929_ );
and  ( new_n31089_, new_n30944_, new_n30943_ );
and  ( new_n31090_, new_n30940_, new_n30937_ );
or   ( new_n31091_, new_n31090_, new_n31089_ );
and  ( new_n31092_, new_n31091_, new_n30945_ );
and  ( new_n31093_, new_n31092_, new_n30935_ );
or   ( new_n31094_, new_n31093_, new_n31088_ );
or   ( new_n31095_, new_n31094_, new_n31084_ );
and  ( new_n31096_, new_n31095_, new_n30922_ );
and  ( new_n31097_, new_n31096_, new_n30907_ );
and  ( new_n31098_, new_n30898_, new_n30895_ );
and  ( new_n31099_, new_n30905_, new_n30902_ );
or   ( new_n31100_, new_n31099_, new_n31098_ );
and  ( new_n31101_, new_n31100_, new_n30899_ );
and  ( new_n31102_, new_n30913_, new_n30910_ );
and  ( new_n31103_, new_n30920_, new_n30917_ );
or   ( new_n31104_, new_n31103_, new_n31102_ );
and  ( new_n31105_, new_n31104_, new_n30914_ );
and  ( new_n31106_, new_n31105_, new_n30907_ );
or   ( new_n31107_, new_n31106_, new_n31101_ );
or   ( new_n31108_, new_n31107_, new_n31097_ );
and  ( new_n31109_, new_n31108_, new_n30892_ );
or   ( new_n31110_, new_n31109_, new_n30889_ );
and  ( new_n31111_, new_n31110_, new_n30857_ );
and  ( new_n31112_, new_n31111_, new_n30815_ );
or   ( new_n31113_, new_n31112_, new_n30854_ );
or   ( new_n31114_, new_n31113_, new_n30812_ );
and  ( new_n31115_, new_n31114_, new_n30774_ );
or   ( new_n31116_, new_n31115_, new_n30771_ );
and  ( new_n31117_, new_n31116_, new_n30733_ );
or   ( new_n31118_, new_n31117_, new_n30730_ );
and  ( new_n31119_, new_n31118_, new_n30699_ );
or   ( new_n31120_, new_n31119_, new_n30696_ );
and  ( new_n31121_, new_n31120_, new_n30670_ );
or   ( new_n31122_, new_n31121_, new_n30667_ );
or   ( new_n31123_, new_n31122_, new_n30638_ );
and  ( new_n31124_, new_n31123_, new_n30635_ );
and  ( new_n31125_, new_n31124_, new_n16000_ );
or   ( new_n31126_, new_n841_, new_n112_ );
and  ( new_n31127_, new_n870_, RI2b1c4342d558_66 );
and  ( new_n31128_, new_n855_, RI2b1c4342d4e0_65 );
or   ( new_n31129_, new_n31128_, new_n31127_ );
and  ( new_n31130_, new_n31129_, new_n842_ );
or   ( new_n31131_, new_n857_, new_n526_ );
or   ( new_n31132_, new_n861_, new_n99_ );
and  ( new_n31133_, new_n31132_, new_n31131_ );
and  ( new_n31134_, new_n31133_, new_n866_ );
or   ( new_n31135_, new_n31134_, new_n31130_ );
and  ( new_n31136_, new_n31135_, new_n785_ );
and  ( new_n31137_, new_n31133_, new_n842_ );
and  ( new_n31138_, new_n31129_, new_n866_ );
or   ( new_n31139_, new_n31138_, new_n31137_ );
and  ( new_n31140_, new_n31139_, new_n813_ );
or   ( new_n31141_, new_n31140_, new_n31136_ );
and  ( new_n31142_, new_n31141_, new_n31126_ );
and  ( new_n31143_, new_n720_, RI2b1c4342d5d0_67 );
and  ( new_n31144_, new_n31139_, new_n785_ );
and  ( new_n31145_, new_n31135_, new_n813_ );
or   ( new_n31146_, new_n31145_, new_n31144_ );
and  ( new_n31147_, new_n31146_, new_n31143_ );
or   ( new_n31148_, new_n31147_, new_n31142_ );
or   ( new_n31149_, new_n804_, new_n99_ );
and  ( new_n31150_, new_n31149_, new_n785_ );
and  ( new_n31151_, new_n817_, RI2b1c4342d4e0_65 );
and  ( new_n31152_, new_n31151_, new_n813_ );
or   ( new_n31153_, new_n31152_, new_n31150_ );
or   ( new_n31154_, new_n857_, new_n112_ );
or   ( new_n31155_, new_n861_, new_n526_ );
and  ( new_n31156_, new_n31155_, new_n31154_ );
and  ( new_n31157_, new_n31156_, new_n842_ );
and  ( new_n31158_, new_n870_, RI2b1c4342d5d0_67 );
and  ( new_n31159_, new_n855_, RI2b1c4342d558_66 );
or   ( new_n31160_, new_n31159_, new_n31158_ );
and  ( new_n31161_, new_n31160_, new_n866_ );
or   ( new_n31162_, new_n31161_, new_n31157_ );
and  ( new_n31163_, new_n31162_, new_n31153_ );
and  ( new_n31164_, new_n31151_, new_n785_ );
and  ( new_n31165_, new_n31149_, new_n813_ );
or   ( new_n31166_, new_n31165_, new_n31164_ );
and  ( new_n31167_, new_n31160_, new_n842_ );
and  ( new_n31168_, new_n31156_, new_n866_ );
or   ( new_n31169_, new_n31168_, new_n31167_ );
and  ( new_n31170_, new_n31169_, new_n31166_ );
or   ( new_n31171_, new_n31170_, new_n31163_ );
or   ( new_n31172_, new_n841_, new_n612_ );
and  ( new_n31173_, new_n31172_, new_n31171_ );
and  ( new_n31174_, new_n31166_, new_n31162_ );
and  ( new_n31175_, new_n31169_, new_n31153_ );
or   ( new_n31176_, new_n31175_, new_n31174_ );
and  ( new_n31177_, new_n720_, RI2b1c4342d648_68 );
and  ( new_n31178_, new_n31177_, new_n31176_ );
or   ( new_n31179_, new_n31178_, new_n31173_ );
or   ( new_n31180_, new_n804_, new_n526_ );
or   ( new_n31181_, new_n808_, new_n99_ );
and  ( new_n31182_, new_n31181_, new_n31180_ );
and  ( new_n31183_, new_n31182_, new_n785_ );
and  ( new_n31184_, new_n817_, RI2b1c4342d558_66 );
and  ( new_n31185_, new_n802_, RI2b1c4342d4e0_65 );
or   ( new_n31186_, new_n31185_, new_n31184_ );
and  ( new_n31187_, new_n31186_, new_n813_ );
or   ( new_n31188_, new_n31187_, new_n31183_ );
and  ( new_n31189_, new_n31188_, new_n762_ );
or   ( new_n31190_, new_n857_, new_n612_ );
or   ( new_n31191_, new_n861_, new_n112_ );
and  ( new_n31192_, new_n31191_, new_n31190_ );
and  ( new_n31193_, new_n31192_, new_n842_ );
and  ( new_n31194_, new_n870_, RI2b1c4342d648_68 );
and  ( new_n31195_, new_n855_, RI2b1c4342d5d0_67 );
or   ( new_n31196_, new_n31195_, new_n31194_ );
and  ( new_n31197_, new_n31196_, new_n866_ );
or   ( new_n31198_, new_n31197_, new_n31193_ );
or   ( new_n31199_, new_n31188_, new_n762_ );
and  ( new_n31200_, new_n31199_, new_n31198_ );
or   ( new_n31201_, new_n31200_, new_n31189_ );
and  ( new_n31202_, new_n31201_, new_n31179_ );
or   ( new_n31203_, new_n31162_, new_n31153_ );
and  ( new_n31204_, new_n31203_, new_n31172_ );
or   ( new_n31205_, new_n31204_, new_n31163_ );
and  ( new_n31206_, new_n31205_, new_n31202_ );
and  ( new_n31207_, new_n31176_, new_n31172_ );
and  ( new_n31208_, new_n31177_, new_n31171_ );
or   ( new_n31209_, new_n31208_, new_n31207_ );
and  ( new_n31210_, new_n31186_, new_n785_ );
and  ( new_n31211_, new_n31182_, new_n813_ );
or   ( new_n31212_, new_n31211_, new_n31210_ );
and  ( new_n31213_, new_n31212_, new_n734_ );
and  ( new_n31214_, new_n31196_, new_n842_ );
and  ( new_n31215_, new_n31192_, new_n866_ );
or   ( new_n31216_, new_n31215_, new_n31214_ );
or   ( new_n31217_, new_n31212_, new_n734_ );
and  ( new_n31218_, new_n31217_, new_n31216_ );
or   ( new_n31219_, new_n31218_, new_n31213_ );
or   ( new_n31220_, new_n31219_, new_n31209_ );
or   ( new_n31221_, new_n31169_, new_n31166_ );
or   ( new_n31222_, new_n31177_, new_n31170_ );
and  ( new_n31223_, new_n31222_, new_n31221_ );
and  ( new_n31224_, new_n31223_, new_n31220_ );
or   ( new_n31225_, new_n31224_, new_n31206_ );
and  ( new_n31226_, new_n31225_, new_n31148_ );
and  ( new_n31227_, new_n31146_, new_n31126_ );
and  ( new_n31228_, new_n31143_, new_n31141_ );
or   ( new_n31229_, new_n31228_, new_n31227_ );
and  ( new_n31230_, new_n31220_, new_n31205_ );
and  ( new_n31231_, new_n31223_, new_n31202_ );
or   ( new_n31232_, new_n31231_, new_n31230_ );
and  ( new_n31233_, new_n31232_, new_n31229_ );
or   ( new_n31234_, new_n31233_, new_n31226_ );
or   ( new_n31235_, new_n841_, new_n755_ );
or   ( new_n31236_, new_n753_, new_n99_ );
and  ( new_n31237_, new_n31236_, new_n734_ );
and  ( new_n31238_, new_n766_, RI2b1c4342d4e0_65 );
and  ( new_n31239_, new_n31238_, new_n762_ );
or   ( new_n31240_, new_n31239_, new_n31237_ );
or   ( new_n31241_, new_n804_, new_n112_ );
or   ( new_n31242_, new_n808_, new_n526_ );
and  ( new_n31243_, new_n31242_, new_n31241_ );
and  ( new_n31244_, new_n31243_, new_n785_ );
and  ( new_n31245_, new_n817_, RI2b1c4342d5d0_67 );
and  ( new_n31246_, new_n802_, RI2b1c4342d558_66 );
or   ( new_n31247_, new_n31246_, new_n31245_ );
and  ( new_n31248_, new_n31247_, new_n813_ );
or   ( new_n31249_, new_n31248_, new_n31244_ );
and  ( new_n31250_, new_n31249_, new_n31240_ );
or   ( new_n31251_, new_n857_, new_n591_ );
or   ( new_n31252_, new_n861_, new_n612_ );
and  ( new_n31253_, new_n31252_, new_n31251_ );
and  ( new_n31254_, new_n31253_, new_n842_ );
and  ( new_n31255_, new_n870_, RI2b1c4342d6c0_69 );
and  ( new_n31256_, new_n855_, RI2b1c4342d648_68 );
or   ( new_n31257_, new_n31256_, new_n31255_ );
and  ( new_n31258_, new_n31257_, new_n866_ );
or   ( new_n31259_, new_n31258_, new_n31254_ );
or   ( new_n31260_, new_n31249_, new_n31240_ );
and  ( new_n31261_, new_n31260_, new_n31259_ );
or   ( new_n31262_, new_n31261_, new_n31250_ );
and  ( new_n31263_, new_n31262_, new_n31235_ );
or   ( new_n31264_, new_n841_, new_n591_ );
or   ( new_n31265_, new_n31262_, new_n31235_ );
and  ( new_n31266_, new_n31265_, new_n31264_ );
or   ( new_n31267_, new_n31266_, new_n31263_ );
or   ( new_n31268_, new_n31213_, new_n31189_ );
and  ( new_n31269_, new_n31268_, new_n31198_ );
and  ( new_n31270_, new_n31188_, new_n734_ );
and  ( new_n31271_, new_n31212_, new_n762_ );
or   ( new_n31272_, new_n31271_, new_n31270_ );
and  ( new_n31273_, new_n31272_, new_n31216_ );
or   ( new_n31274_, new_n31273_, new_n31269_ );
and  ( new_n31275_, new_n720_, RI2b1c4342d738_70 );
or   ( new_n31276_, new_n753_, new_n526_ );
or   ( new_n31277_, new_n757_, new_n99_ );
and  ( new_n31278_, new_n31277_, new_n31276_ );
and  ( new_n31279_, new_n31278_, new_n734_ );
and  ( new_n31280_, new_n766_, RI2b1c4342d558_66 );
and  ( new_n31281_, new_n751_, RI2b1c4342d4e0_65 );
or   ( new_n31282_, new_n31281_, new_n31280_ );
and  ( new_n31283_, new_n31282_, new_n762_ );
or   ( new_n31284_, new_n31283_, new_n31279_ );
and  ( new_n31285_, new_n31284_, new_n619_ );
or   ( new_n31286_, new_n804_, new_n612_ );
or   ( new_n31287_, new_n808_, new_n112_ );
and  ( new_n31288_, new_n31287_, new_n31286_ );
and  ( new_n31289_, new_n31288_, new_n785_ );
and  ( new_n31290_, new_n817_, RI2b1c4342d648_68 );
and  ( new_n31291_, new_n802_, RI2b1c4342d5d0_67 );
or   ( new_n31292_, new_n31291_, new_n31290_ );
and  ( new_n31293_, new_n31292_, new_n813_ );
or   ( new_n31294_, new_n31293_, new_n31289_ );
or   ( new_n31295_, new_n31284_, new_n619_ );
and  ( new_n31296_, new_n31295_, new_n31294_ );
or   ( new_n31297_, new_n31296_, new_n31285_ );
and  ( new_n31298_, new_n31297_, new_n31275_ );
and  ( new_n31299_, new_n31238_, new_n734_ );
and  ( new_n31300_, new_n31236_, new_n762_ );
or   ( new_n31301_, new_n31300_, new_n31299_ );
and  ( new_n31302_, new_n31247_, new_n785_ );
and  ( new_n31303_, new_n31243_, new_n813_ );
or   ( new_n31304_, new_n31303_, new_n31302_ );
and  ( new_n31305_, new_n31304_, new_n31301_ );
or   ( new_n31306_, new_n31305_, new_n31250_ );
and  ( new_n31307_, new_n31306_, new_n31259_ );
and  ( new_n31308_, new_n31301_, new_n31249_ );
and  ( new_n31309_, new_n31304_, new_n31240_ );
or   ( new_n31310_, new_n31309_, new_n31308_ );
and  ( new_n31311_, new_n31257_, new_n842_ );
and  ( new_n31312_, new_n31253_, new_n866_ );
or   ( new_n31313_, new_n31312_, new_n31311_ );
and  ( new_n31314_, new_n31313_, new_n31310_ );
or   ( new_n31315_, new_n31314_, new_n31307_ );
or   ( new_n31316_, new_n31297_, new_n31275_ );
and  ( new_n31317_, new_n31316_, new_n31315_ );
or   ( new_n31318_, new_n31317_, new_n31298_ );
and  ( new_n31319_, new_n31318_, new_n31274_ );
or   ( new_n31320_, new_n31304_, new_n31301_ );
and  ( new_n31321_, new_n31320_, new_n31313_ );
or   ( new_n31322_, new_n31321_, new_n31305_ );
and  ( new_n31323_, new_n31322_, new_n31275_ );
or   ( new_n31324_, new_n31323_, new_n31263_ );
and  ( new_n31325_, new_n31324_, new_n31264_ );
and  ( new_n31326_, new_n31322_, new_n31235_ );
and  ( new_n31327_, new_n31275_, new_n31262_ );
or   ( new_n31328_, new_n31327_, new_n31326_ );
and  ( new_n31329_, new_n720_, RI2b1c4342d6c0_69 );
and  ( new_n31330_, new_n31329_, new_n31328_ );
or   ( new_n31331_, new_n31330_, new_n31325_ );
or   ( new_n31332_, new_n31318_, new_n31274_ );
and  ( new_n31333_, new_n31332_, new_n31331_ );
or   ( new_n31334_, new_n31333_, new_n31319_ );
and  ( new_n31335_, new_n31334_, new_n31267_ );
and  ( new_n31336_, new_n31219_, new_n31179_ );
and  ( new_n31337_, new_n31209_, new_n31201_ );
or   ( new_n31338_, new_n31337_, new_n31336_ );
or   ( new_n31339_, new_n31334_, new_n31267_ );
and  ( new_n31340_, new_n31339_, new_n31338_ );
or   ( new_n31341_, new_n31340_, new_n31335_ );
or   ( new_n31342_, new_n31341_, new_n31234_ );
and  ( new_n31343_, new_n31232_, new_n31148_ );
and  ( new_n31344_, new_n31229_, new_n31225_ );
or   ( new_n31345_, new_n31344_, new_n31343_ );
and  ( new_n31346_, new_n31272_, new_n31198_ );
and  ( new_n31347_, new_n31268_, new_n31216_ );
or   ( new_n31348_, new_n31347_, new_n31346_ );
and  ( new_n31349_, new_n31282_, new_n734_ );
and  ( new_n31350_, new_n31278_, new_n762_ );
or   ( new_n31351_, new_n31350_, new_n31349_ );
and  ( new_n31352_, new_n31351_, new_n590_ );
and  ( new_n31353_, new_n31292_, new_n785_ );
and  ( new_n31354_, new_n31288_, new_n813_ );
or   ( new_n31355_, new_n31354_, new_n31353_ );
or   ( new_n31356_, new_n31351_, new_n590_ );
and  ( new_n31357_, new_n31356_, new_n31355_ );
or   ( new_n31358_, new_n31357_, new_n31352_ );
and  ( new_n31359_, new_n31358_, new_n31235_ );
and  ( new_n31360_, new_n31310_, new_n31259_ );
and  ( new_n31361_, new_n31313_, new_n31306_ );
or   ( new_n31362_, new_n31361_, new_n31360_ );
or   ( new_n31363_, new_n31358_, new_n31235_ );
and  ( new_n31364_, new_n31363_, new_n31362_ );
or   ( new_n31365_, new_n31364_, new_n31359_ );
and  ( new_n31366_, new_n31365_, new_n31348_ );
and  ( new_n31367_, new_n31328_, new_n31264_ );
and  ( new_n31368_, new_n31329_, new_n31324_ );
or   ( new_n31369_, new_n31368_, new_n31367_ );
or   ( new_n31370_, new_n31365_, new_n31348_ );
and  ( new_n31371_, new_n31370_, new_n31369_ );
or   ( new_n31372_, new_n31371_, new_n31366_ );
or   ( new_n31373_, new_n31322_, new_n31275_ );
and  ( new_n31374_, new_n31373_, new_n31329_ );
or   ( new_n31375_, new_n31374_, new_n31323_ );
and  ( new_n31376_, new_n31375_, new_n31372_ );
and  ( new_n31377_, new_n31219_, new_n31209_ );
or   ( new_n31378_, new_n31377_, new_n31202_ );
or   ( new_n31379_, new_n31375_, new_n31372_ );
and  ( new_n31380_, new_n31379_, new_n31378_ );
or   ( new_n31381_, new_n31380_, new_n31376_ );
or   ( new_n31382_, new_n31381_, new_n31345_ );
and  ( new_n31383_, new_n31382_, new_n31342_ );
or   ( new_n31384_, new_n15321_, new_n11172_ );
and  ( new_n31385_, new_n31384_, new_n7860_ );
or   ( new_n31386_, new_n524_, new_n99_ );
and  ( new_n31387_, new_n31386_, new_n505_ );
and  ( new_n31388_, new_n537_, RI2b1c4342d4e0_65 );
and  ( new_n31389_, new_n31388_, new_n533_ );
or   ( new_n31390_, new_n31389_, new_n31387_ );
or   ( new_n31391_, new_n610_, new_n112_ );
or   ( new_n31392_, new_n614_, new_n526_ );
and  ( new_n31393_, new_n31392_, new_n31391_ );
and  ( new_n31394_, new_n31393_, new_n590_ );
and  ( new_n31395_, new_n623_, RI2b1c4342d5d0_67 );
and  ( new_n31396_, new_n608_, RI2b1c4342d558_66 );
or   ( new_n31397_, new_n31396_, new_n31395_ );
and  ( new_n31398_, new_n31397_, new_n619_ );
or   ( new_n31399_, new_n31398_, new_n31394_ );
and  ( new_n31400_, new_n31399_, new_n31390_ );
and  ( new_n31401_, new_n31388_, new_n505_ );
and  ( new_n31402_, new_n31386_, new_n533_ );
or   ( new_n31403_, new_n31402_, new_n31401_ );
and  ( new_n31404_, new_n31397_, new_n590_ );
and  ( new_n31405_, new_n31393_, new_n619_ );
or   ( new_n31406_, new_n31405_, new_n31404_ );
and  ( new_n31407_, new_n31406_, new_n31403_ );
or   ( new_n31408_, new_n31407_, new_n31400_ );
or   ( new_n31409_, new_n753_, new_n591_ );
or   ( new_n31410_, new_n757_, new_n612_ );
and  ( new_n31411_, new_n31410_, new_n31409_ );
and  ( new_n31412_, new_n31411_, new_n734_ );
and  ( new_n31413_, new_n766_, RI2b1c4342d6c0_69 );
and  ( new_n31414_, new_n751_, RI2b1c4342d648_68 );
or   ( new_n31415_, new_n31414_, new_n31413_ );
and  ( new_n31416_, new_n31415_, new_n762_ );
or   ( new_n31417_, new_n31416_, new_n31412_ );
and  ( new_n31418_, new_n31417_, new_n31408_ );
and  ( new_n31419_, new_n31403_, new_n31399_ );
and  ( new_n31420_, new_n31406_, new_n31390_ );
or   ( new_n31421_, new_n31420_, new_n31419_ );
and  ( new_n31422_, new_n31415_, new_n734_ );
and  ( new_n31423_, new_n31411_, new_n762_ );
or   ( new_n31424_, new_n31423_, new_n31422_ );
and  ( new_n31425_, new_n31424_, new_n31421_ );
or   ( new_n31426_, new_n31425_, new_n31418_ );
or   ( new_n31427_, new_n15396_, new_n428_ );
and  ( new_n31428_, new_n31427_, new_n15406_ );
or   ( new_n31429_, new_n31428_, new_n15397_ );
or   ( new_n31430_, new_n15353_, new_n15344_ );
and  ( new_n31431_, new_n31430_, new_n15335_ );
or   ( new_n31432_, new_n31431_, new_n15354_ );
and  ( new_n31433_, new_n31432_, new_n31429_ );
or   ( new_n31434_, new_n15360_, new_n15357_ );
and  ( new_n31435_, new_n31434_, new_n15366_ );
or   ( new_n31436_, new_n31435_, new_n15361_ );
or   ( new_n31437_, new_n15400_, new_n457_ );
and  ( new_n31438_, new_n31437_, new_n15387_ );
or   ( new_n31439_, new_n31438_, new_n15401_ );
and  ( new_n31440_, new_n31439_, new_n31436_ );
or   ( new_n31441_, new_n31440_, new_n31433_ );
and  ( new_n31442_, new_n31441_, new_n31426_ );
and  ( new_n31443_, new_n31421_, new_n31417_ );
and  ( new_n31444_, new_n31424_, new_n31408_ );
or   ( new_n31445_, new_n31444_, new_n31443_ );
and  ( new_n31446_, new_n31439_, new_n31432_ );
and  ( new_n31447_, new_n31436_, new_n31429_ );
or   ( new_n31448_, new_n31447_, new_n31446_ );
and  ( new_n31449_, new_n31448_, new_n31445_ );
or   ( new_n31450_, new_n31449_, new_n31442_ );
or   ( new_n31451_, new_n15426_, new_n15423_ );
and  ( new_n31452_, new_n31451_, new_n15420_ );
or   ( new_n31453_, new_n31452_, new_n15427_ );
and  ( new_n31454_, new_n31453_, new_n31450_ );
and  ( new_n31455_, new_n31445_, new_n31441_ );
and  ( new_n31456_, new_n31448_, new_n31426_ );
or   ( new_n31457_, new_n31456_, new_n31455_ );
or   ( new_n31458_, new_n15433_, new_n15430_ );
or   ( new_n31459_, new_n15439_, new_n15434_ );
and  ( new_n31460_, new_n31459_, new_n31458_ );
and  ( new_n31461_, new_n31460_, new_n31457_ );
or   ( new_n31462_, new_n31461_, new_n31454_ );
or   ( new_n31463_, new_n15450_, new_n15447_ );
and  ( new_n31464_, new_n31463_, new_n887_ );
or   ( new_n31465_, new_n31464_, new_n15451_ );
or   ( new_n31466_, new_n15371_, new_n15326_ );
and  ( new_n31467_, new_n31466_, new_n15411_ );
or   ( new_n31468_, new_n31467_, new_n15372_ );
and  ( new_n31469_, new_n31468_, new_n31465_ );
or   ( new_n31470_, new_n15457_, new_n15454_ );
or   ( new_n31471_, new_n15458_, new_n721_ );
and  ( new_n31472_, new_n31471_, new_n31470_ );
or   ( new_n31473_, new_n15376_, new_n15373_ );
and  ( new_n31474_, new_n31473_, new_n15418_ );
or   ( new_n31475_, new_n31474_, new_n15377_ );
and  ( new_n31476_, new_n31475_, new_n31472_ );
or   ( new_n31477_, new_n31476_, new_n31469_ );
or   ( new_n31478_, new_n804_, new_n110_ );
or   ( new_n31479_, new_n808_, new_n755_ );
and  ( new_n31480_, new_n31479_, new_n31478_ );
and  ( new_n31481_, new_n31480_, new_n785_ );
and  ( new_n31482_, new_n817_, RI2b1c4342d7b0_71 );
and  ( new_n31483_, new_n802_, RI2b1c4342d738_70 );
or   ( new_n31484_, new_n31483_, new_n31482_ );
and  ( new_n31485_, new_n31484_, new_n813_ );
or   ( new_n31486_, new_n31485_, new_n31481_ );
or   ( new_n31487_, new_n857_, new_n105_ );
or   ( new_n31488_, new_n861_, new_n806_ );
and  ( new_n31489_, new_n31488_, new_n31487_ );
and  ( new_n31490_, new_n31489_, new_n842_ );
and  ( new_n31491_, new_n870_, RI2b1c4342d8a0_73 );
and  ( new_n31492_, new_n855_, RI2b1c4342d828_72 );
or   ( new_n31493_, new_n31492_, new_n31491_ );
and  ( new_n31494_, new_n31493_, new_n866_ );
or   ( new_n31495_, new_n31494_, new_n31490_ );
and  ( new_n31496_, new_n31495_, new_n31486_ );
and  ( new_n31497_, new_n31484_, new_n785_ );
and  ( new_n31498_, new_n31480_, new_n813_ );
or   ( new_n31499_, new_n31498_, new_n31497_ );
and  ( new_n31500_, new_n31493_, new_n842_ );
and  ( new_n31501_, new_n31489_, new_n866_ );
or   ( new_n31502_, new_n31501_, new_n31500_ );
and  ( new_n31503_, new_n31502_, new_n31499_ );
or   ( new_n31504_, new_n31503_, new_n31496_ );
or   ( new_n31505_, new_n841_, new_n859_ );
and  ( new_n31506_, new_n31505_, new_n31504_ );
and  ( new_n31507_, new_n31499_, new_n31495_ );
and  ( new_n31508_, new_n31502_, new_n31486_ );
or   ( new_n31509_, new_n31508_, new_n31507_ );
and  ( new_n31510_, new_n720_, RI2b1c4342d918_74 );
and  ( new_n31511_, new_n31510_, new_n31509_ );
or   ( new_n31512_, new_n31511_, new_n31506_ );
and  ( new_n31513_, new_n31512_, new_n31477_ );
and  ( new_n31514_, new_n31472_, new_n31468_ );
and  ( new_n31515_, new_n31475_, new_n31465_ );
or   ( new_n31516_, new_n31515_, new_n31514_ );
and  ( new_n31517_, new_n31509_, new_n31505_ );
and  ( new_n31518_, new_n31510_, new_n31504_ );
or   ( new_n31519_, new_n31518_, new_n31517_ );
and  ( new_n31520_, new_n31519_, new_n31516_ );
or   ( new_n31521_, new_n31520_, new_n31513_ );
and  ( new_n31522_, new_n31521_, new_n31462_ );
and  ( new_n31523_, new_n31460_, new_n31450_ );
and  ( new_n31524_, new_n31457_, new_n31453_ );
or   ( new_n31525_, new_n31524_, new_n31523_ );
and  ( new_n31526_, new_n31516_, new_n31512_ );
and  ( new_n31527_, new_n31519_, new_n31477_ );
or   ( new_n31528_, new_n31527_, new_n31526_ );
and  ( new_n31529_, new_n31528_, new_n31525_ );
or   ( new_n31530_, new_n31529_, new_n31522_ );
or   ( new_n31531_, new_n15472_, new_n15465_ );
and  ( new_n31532_, new_n31531_, new_n15444_ );
or   ( new_n31533_, new_n31532_, new_n15482_ );
and  ( new_n31534_, new_n31533_, new_n31530_ );
and  ( new_n31535_, new_n31525_, new_n31521_ );
and  ( new_n31536_, new_n31528_, new_n31462_ );
or   ( new_n31537_, new_n31536_, new_n31535_ );
or   ( new_n31538_, new_n15475_, new_n15468_ );
and  ( new_n31539_, new_n31538_, new_n15481_ );
or   ( new_n31540_, new_n31539_, new_n15483_ );
and  ( new_n31541_, new_n31540_, new_n31537_ );
or   ( new_n31542_, new_n31541_, new_n31534_ );
or   ( new_n31543_, new_n15496_, new_n15493_ );
and  ( new_n31544_, new_n31543_, new_n31542_ );
or   ( new_n31545_, new_n31544_, new_n15507_ );
or   ( new_n31546_, new_n31441_, new_n31426_ );
or   ( new_n31547_, new_n31468_, new_n31465_ );
and  ( new_n31548_, new_n31547_, new_n31512_ );
or   ( new_n31549_, new_n31548_, new_n31469_ );
and  ( new_n31550_, new_n31549_, new_n31546_ );
or   ( new_n31551_, new_n31549_, new_n31546_ );
or   ( new_n31552_, new_n610_, new_n526_ );
or   ( new_n31553_, new_n614_, new_n99_ );
and  ( new_n31554_, new_n31553_, new_n31552_ );
and  ( new_n31555_, new_n31554_, new_n590_ );
and  ( new_n31556_, new_n623_, RI2b1c4342d558_66 );
and  ( new_n31557_, new_n608_, RI2b1c4342d4e0_65 );
or   ( new_n31558_, new_n31557_, new_n31556_ );
and  ( new_n31559_, new_n31558_, new_n619_ );
or   ( new_n31560_, new_n31559_, new_n31555_ );
and  ( new_n31561_, new_n31560_, new_n533_ );
and  ( new_n31562_, new_n31558_, new_n590_ );
and  ( new_n31563_, new_n31554_, new_n619_ );
or   ( new_n31564_, new_n31563_, new_n31562_ );
and  ( new_n31565_, new_n31564_, new_n505_ );
or   ( new_n31566_, new_n31565_, new_n31561_ );
or   ( new_n31567_, new_n753_, new_n612_ );
or   ( new_n31568_, new_n757_, new_n112_ );
and  ( new_n31569_, new_n31568_, new_n31567_ );
and  ( new_n31570_, new_n31569_, new_n734_ );
and  ( new_n31571_, new_n766_, RI2b1c4342d648_68 );
and  ( new_n31572_, new_n751_, RI2b1c4342d5d0_67 );
or   ( new_n31573_, new_n31572_, new_n31571_ );
and  ( new_n31574_, new_n31573_, new_n762_ );
or   ( new_n31575_, new_n31574_, new_n31570_ );
and  ( new_n31576_, new_n31575_, new_n31566_ );
and  ( new_n31577_, new_n31560_, new_n505_ );
and  ( new_n31578_, new_n31564_, new_n533_ );
or   ( new_n31579_, new_n31578_, new_n31577_ );
and  ( new_n31580_, new_n31573_, new_n734_ );
and  ( new_n31581_, new_n31569_, new_n762_ );
or   ( new_n31582_, new_n31581_, new_n31580_ );
and  ( new_n31583_, new_n31582_, new_n31579_ );
or   ( new_n31584_, new_n31583_, new_n31576_ );
and  ( new_n31585_, new_n31584_, new_n31446_ );
or   ( new_n31586_, new_n31436_, new_n31429_ );
and  ( new_n31587_, new_n31579_, new_n31575_ );
and  ( new_n31588_, new_n31582_, new_n31566_ );
or   ( new_n31589_, new_n31588_, new_n31587_ );
and  ( new_n31590_, new_n31589_, new_n31586_ );
or   ( new_n31591_, new_n31590_, new_n31585_ );
or   ( new_n31592_, new_n31399_, new_n31390_ );
and  ( new_n31593_, new_n31592_, new_n31417_ );
or   ( new_n31594_, new_n31593_, new_n31400_ );
or   ( new_n31595_, new_n31495_, new_n31486_ );
and  ( new_n31596_, new_n31595_, new_n31505_ );
or   ( new_n31597_, new_n31596_, new_n31496_ );
and  ( new_n31598_, new_n31597_, new_n31594_ );
or   ( new_n31599_, new_n31406_, new_n31403_ );
and  ( new_n31600_, new_n31599_, new_n31424_ );
or   ( new_n31601_, new_n31600_, new_n31407_ );
or   ( new_n31602_, new_n31502_, new_n31499_ );
or   ( new_n31603_, new_n31510_, new_n31503_ );
and  ( new_n31604_, new_n31603_, new_n31602_ );
and  ( new_n31605_, new_n31604_, new_n31601_ );
or   ( new_n31606_, new_n31605_, new_n31598_ );
or   ( new_n31607_, new_n804_, new_n755_ );
or   ( new_n31608_, new_n808_, new_n591_ );
and  ( new_n31609_, new_n31608_, new_n31607_ );
and  ( new_n31610_, new_n31609_, new_n785_ );
and  ( new_n31611_, new_n817_, RI2b1c4342d738_70 );
and  ( new_n31612_, new_n802_, RI2b1c4342d6c0_69 );
or   ( new_n31613_, new_n31612_, new_n31611_ );
and  ( new_n31614_, new_n31613_, new_n813_ );
or   ( new_n31615_, new_n31614_, new_n31610_ );
or   ( new_n31616_, new_n857_, new_n806_ );
or   ( new_n31617_, new_n861_, new_n110_ );
and  ( new_n31618_, new_n31617_, new_n31616_ );
and  ( new_n31619_, new_n31618_, new_n842_ );
and  ( new_n31620_, new_n870_, RI2b1c4342d828_72 );
and  ( new_n31621_, new_n855_, RI2b1c4342d7b0_71 );
or   ( new_n31622_, new_n31621_, new_n31620_ );
and  ( new_n31623_, new_n31622_, new_n866_ );
or   ( new_n31624_, new_n31623_, new_n31619_ );
and  ( new_n31625_, new_n31624_, new_n31615_ );
and  ( new_n31626_, new_n31613_, new_n785_ );
and  ( new_n31627_, new_n31609_, new_n813_ );
or   ( new_n31628_, new_n31627_, new_n31626_ );
and  ( new_n31629_, new_n31622_, new_n842_ );
and  ( new_n31630_, new_n31618_, new_n866_ );
or   ( new_n31631_, new_n31630_, new_n31629_ );
and  ( new_n31632_, new_n31631_, new_n31628_ );
or   ( new_n31633_, new_n31632_, new_n31625_ );
or   ( new_n31634_, new_n841_, new_n105_ );
and  ( new_n31635_, new_n31634_, new_n31633_ );
and  ( new_n31636_, new_n31628_, new_n31624_ );
and  ( new_n31637_, new_n31631_, new_n31615_ );
or   ( new_n31638_, new_n31637_, new_n31636_ );
and  ( new_n31639_, new_n720_, RI2b1c4342d8a0_73 );
and  ( new_n31640_, new_n31639_, new_n31638_ );
or   ( new_n31641_, new_n31640_, new_n31635_ );
and  ( new_n31642_, new_n31641_, new_n31606_ );
and  ( new_n31643_, new_n31601_, new_n31597_ );
and  ( new_n31644_, new_n31604_, new_n31594_ );
or   ( new_n31645_, new_n31644_, new_n31643_ );
and  ( new_n31646_, new_n31638_, new_n31634_ );
and  ( new_n31647_, new_n31639_, new_n31633_ );
or   ( new_n31648_, new_n31647_, new_n31646_ );
and  ( new_n31649_, new_n31648_, new_n31645_ );
or   ( new_n31650_, new_n31649_, new_n31642_ );
and  ( new_n31651_, new_n31650_, new_n31591_ );
and  ( new_n31652_, new_n31586_, new_n31584_ );
and  ( new_n31653_, new_n31589_, new_n31446_ );
or   ( new_n31654_, new_n31653_, new_n31652_ );
and  ( new_n31655_, new_n31645_, new_n31641_ );
and  ( new_n31656_, new_n31648_, new_n31606_ );
or   ( new_n31657_, new_n31656_, new_n31655_ );
and  ( new_n31658_, new_n31657_, new_n31654_ );
or   ( new_n31659_, new_n31658_, new_n31651_ );
and  ( new_n31660_, new_n31659_, new_n31551_ );
or   ( new_n31661_, new_n31660_, new_n31550_ );
or   ( new_n31662_, new_n31584_, new_n31446_ );
and  ( new_n31663_, new_n31662_, new_n31650_ );
or   ( new_n31664_, new_n31663_, new_n31585_ );
and  ( new_n31665_, new_n31664_, new_n31661_ );
or   ( new_n31666_, new_n31589_, new_n31586_ );
and  ( new_n31667_, new_n31666_, new_n31657_ );
or   ( new_n31668_, new_n31667_, new_n31590_ );
or   ( new_n31669_, new_n31475_, new_n31472_ );
and  ( new_n31670_, new_n31669_, new_n31519_ );
or   ( new_n31671_, new_n31670_, new_n31476_ );
and  ( new_n31672_, new_n31671_, new_n31449_ );
or   ( new_n31673_, new_n31671_, new_n31449_ );
and  ( new_n31674_, new_n31654_, new_n31650_ );
and  ( new_n31675_, new_n31657_, new_n31591_ );
or   ( new_n31676_, new_n31675_, new_n31674_ );
and  ( new_n31677_, new_n31676_, new_n31673_ );
or   ( new_n31678_, new_n31677_, new_n31672_ );
and  ( new_n31679_, new_n31678_, new_n31668_ );
or   ( new_n31680_, new_n31679_, new_n31665_ );
or   ( new_n31681_, new_n610_, new_n99_ );
and  ( new_n31682_, new_n31681_, new_n590_ );
and  ( new_n31683_, new_n623_, RI2b1c4342d4e0_65 );
and  ( new_n31684_, new_n31683_, new_n619_ );
or   ( new_n31685_, new_n31684_, new_n31682_ );
or   ( new_n31686_, new_n753_, new_n112_ );
or   ( new_n31687_, new_n757_, new_n526_ );
and  ( new_n31688_, new_n31687_, new_n31686_ );
and  ( new_n31689_, new_n31688_, new_n734_ );
and  ( new_n31690_, new_n766_, RI2b1c4342d5d0_67 );
and  ( new_n31691_, new_n751_, RI2b1c4342d558_66 );
or   ( new_n31692_, new_n31691_, new_n31690_ );
and  ( new_n31693_, new_n31692_, new_n762_ );
or   ( new_n31694_, new_n31693_, new_n31689_ );
and  ( new_n31695_, new_n31694_, new_n31685_ );
and  ( new_n31696_, new_n31683_, new_n590_ );
and  ( new_n31697_, new_n31681_, new_n619_ );
or   ( new_n31698_, new_n31697_, new_n31696_ );
and  ( new_n31699_, new_n31692_, new_n734_ );
and  ( new_n31700_, new_n31688_, new_n762_ );
or   ( new_n31701_, new_n31700_, new_n31699_ );
and  ( new_n31702_, new_n31701_, new_n31698_ );
or   ( new_n31703_, new_n31702_, new_n31695_ );
or   ( new_n31704_, new_n804_, new_n591_ );
or   ( new_n31705_, new_n808_, new_n612_ );
and  ( new_n31706_, new_n31705_, new_n31704_ );
and  ( new_n31707_, new_n31706_, new_n785_ );
and  ( new_n31708_, new_n817_, RI2b1c4342d6c0_69 );
and  ( new_n31709_, new_n802_, RI2b1c4342d648_68 );
or   ( new_n31710_, new_n31709_, new_n31708_ );
and  ( new_n31711_, new_n31710_, new_n813_ );
or   ( new_n31712_, new_n31711_, new_n31707_ );
and  ( new_n31713_, new_n31712_, new_n31703_ );
and  ( new_n31714_, new_n31698_, new_n31694_ );
and  ( new_n31715_, new_n31701_, new_n31685_ );
or   ( new_n31716_, new_n31715_, new_n31714_ );
and  ( new_n31717_, new_n31710_, new_n785_ );
and  ( new_n31718_, new_n31706_, new_n813_ );
or   ( new_n31719_, new_n31718_, new_n31717_ );
and  ( new_n31720_, new_n31719_, new_n31716_ );
or   ( new_n31721_, new_n31720_, new_n31713_ );
or   ( new_n31722_, new_n31597_, new_n31594_ );
and  ( new_n31723_, new_n31722_, new_n31641_ );
or   ( new_n31724_, new_n31723_, new_n31598_ );
and  ( new_n31725_, new_n31724_, new_n31721_ );
and  ( new_n31726_, new_n31716_, new_n31712_ );
and  ( new_n31727_, new_n31719_, new_n31703_ );
or   ( new_n31728_, new_n31727_, new_n31726_ );
or   ( new_n31729_, new_n31604_, new_n31601_ );
or   ( new_n31730_, new_n31648_, new_n31605_ );
and  ( new_n31731_, new_n31730_, new_n31729_ );
and  ( new_n31732_, new_n31731_, new_n31728_ );
or   ( new_n31733_, new_n31732_, new_n31725_ );
or   ( new_n31734_, new_n31624_, new_n31615_ );
and  ( new_n31735_, new_n31734_, new_n31634_ );
or   ( new_n31736_, new_n31735_, new_n31625_ );
or   ( new_n31737_, new_n31560_, new_n533_ );
and  ( new_n31738_, new_n31737_, new_n31575_ );
or   ( new_n31739_, new_n31738_, new_n31561_ );
and  ( new_n31740_, new_n31739_, new_n31736_ );
or   ( new_n31741_, new_n31564_, new_n505_ );
and  ( new_n31742_, new_n31741_, new_n31582_ );
or   ( new_n31743_, new_n31742_, new_n31565_ );
or   ( new_n31744_, new_n31631_, new_n31628_ );
or   ( new_n31745_, new_n31639_, new_n31632_ );
and  ( new_n31746_, new_n31745_, new_n31744_ );
and  ( new_n31747_, new_n31746_, new_n31743_ );
or   ( new_n31748_, new_n31747_, new_n31740_ );
and  ( new_n31749_, new_n870_, RI2b1c4342d7b0_71 );
and  ( new_n31750_, new_n855_, RI2b1c4342d738_70 );
or   ( new_n31751_, new_n31750_, new_n31749_ );
and  ( new_n31752_, new_n31751_, new_n842_ );
or   ( new_n31753_, new_n857_, new_n110_ );
or   ( new_n31754_, new_n861_, new_n755_ );
and  ( new_n31755_, new_n31754_, new_n31753_ );
and  ( new_n31756_, new_n31755_, new_n866_ );
or   ( new_n31757_, new_n31756_, new_n31752_ );
or   ( new_n31758_, new_n841_, new_n806_ );
and  ( new_n31759_, new_n31758_, new_n31757_ );
and  ( new_n31760_, new_n31755_, new_n842_ );
and  ( new_n31761_, new_n31751_, new_n866_ );
or   ( new_n31762_, new_n31761_, new_n31760_ );
and  ( new_n31763_, new_n720_, RI2b1c4342d828_72 );
and  ( new_n31764_, new_n31763_, new_n31762_ );
or   ( new_n31765_, new_n31764_, new_n31759_ );
and  ( new_n31766_, new_n31765_, new_n31748_ );
and  ( new_n31767_, new_n31743_, new_n31736_ );
and  ( new_n31768_, new_n31746_, new_n31739_ );
or   ( new_n31769_, new_n31768_, new_n31767_ );
and  ( new_n31770_, new_n31762_, new_n31758_ );
and  ( new_n31771_, new_n31763_, new_n31757_ );
or   ( new_n31772_, new_n31771_, new_n31770_ );
and  ( new_n31773_, new_n31772_, new_n31769_ );
or   ( new_n31774_, new_n31773_, new_n31766_ );
and  ( new_n31775_, new_n31774_, new_n31733_ );
and  ( new_n31776_, new_n31731_, new_n31721_ );
and  ( new_n31777_, new_n31728_, new_n31724_ );
or   ( new_n31778_, new_n31777_, new_n31776_ );
and  ( new_n31779_, new_n31769_, new_n31765_ );
and  ( new_n31780_, new_n31772_, new_n31748_ );
or   ( new_n31781_, new_n31780_, new_n31779_ );
and  ( new_n31782_, new_n31781_, new_n31778_ );
or   ( new_n31783_, new_n31782_, new_n31775_ );
and  ( new_n31784_, new_n31783_, new_n31680_ );
and  ( new_n31785_, new_n31678_, new_n31664_ );
and  ( new_n31786_, new_n31668_, new_n31661_ );
or   ( new_n31787_, new_n31786_, new_n31785_ );
and  ( new_n31788_, new_n31778_, new_n31774_ );
and  ( new_n31789_, new_n31781_, new_n31733_ );
or   ( new_n31790_, new_n31789_, new_n31788_ );
and  ( new_n31791_, new_n31790_, new_n31787_ );
or   ( new_n31792_, new_n31791_, new_n31784_ );
or   ( new_n31793_, new_n31672_, new_n31550_ );
and  ( new_n31794_, new_n31793_, new_n31659_ );
and  ( new_n31795_, new_n31671_, new_n31546_ );
and  ( new_n31796_, new_n31549_, new_n31449_ );
or   ( new_n31797_, new_n31796_, new_n31795_ );
and  ( new_n31798_, new_n31797_, new_n31676_ );
or   ( new_n31799_, new_n31798_, new_n31794_ );
or   ( new_n31800_, new_n31453_, new_n31450_ );
and  ( new_n31801_, new_n31800_, new_n31521_ );
or   ( new_n31802_, new_n31801_, new_n31454_ );
or   ( new_n31803_, new_n31802_, new_n31799_ );
and  ( new_n31804_, new_n31803_, new_n31792_ );
and  ( new_n31805_, new_n31797_, new_n31659_ );
and  ( new_n31806_, new_n31793_, new_n31676_ );
or   ( new_n31807_, new_n31806_, new_n31805_ );
or   ( new_n31808_, new_n31460_, new_n31457_ );
or   ( new_n31809_, new_n31528_, new_n31461_ );
and  ( new_n31810_, new_n31809_, new_n31808_ );
and  ( new_n31811_, new_n31810_, new_n31807_ );
and  ( new_n31812_, new_n31802_, new_n31799_ );
or   ( new_n31813_, new_n31812_, new_n31811_ );
or   ( new_n31814_, new_n31533_, new_n31530_ );
and  ( new_n31815_, new_n31814_, new_n31813_ );
or   ( new_n31816_, new_n31815_, new_n31804_ );
or   ( new_n31817_, new_n31816_, new_n31545_ );
or   ( new_n31818_, new_n841_, new_n110_ );
or   ( new_n31819_, new_n31352_, new_n31285_ );
and  ( new_n31820_, new_n31819_, new_n31294_ );
and  ( new_n31821_, new_n31284_, new_n590_ );
and  ( new_n31822_, new_n31351_, new_n619_ );
or   ( new_n31823_, new_n31822_, new_n31821_ );
and  ( new_n31824_, new_n31823_, new_n31355_ );
or   ( new_n31825_, new_n31824_, new_n31820_ );
and  ( new_n31826_, new_n31825_, new_n31818_ );
and  ( new_n31827_, new_n720_, RI2b1c4342d7b0_71 );
and  ( new_n31828_, new_n31823_, new_n31294_ );
and  ( new_n31829_, new_n31819_, new_n31355_ );
or   ( new_n31830_, new_n31829_, new_n31828_ );
and  ( new_n31831_, new_n31830_, new_n31827_ );
or   ( new_n31832_, new_n31831_, new_n31826_ );
or   ( new_n31833_, new_n31739_, new_n31736_ );
and  ( new_n31834_, new_n31833_, new_n31765_ );
or   ( new_n31835_, new_n31834_, new_n31740_ );
and  ( new_n31836_, new_n31835_, new_n31832_ );
and  ( new_n31837_, new_n31827_, new_n31825_ );
and  ( new_n31838_, new_n31830_, new_n31818_ );
or   ( new_n31839_, new_n31838_, new_n31837_ );
or   ( new_n31840_, new_n31746_, new_n31743_ );
or   ( new_n31841_, new_n31772_, new_n31747_ );
and  ( new_n31842_, new_n31841_, new_n31840_ );
and  ( new_n31843_, new_n31842_, new_n31839_ );
or   ( new_n31844_, new_n31843_, new_n31836_ );
or   ( new_n31845_, new_n31694_, new_n31685_ );
and  ( new_n31846_, new_n31845_, new_n31712_ );
or   ( new_n31847_, new_n31846_, new_n31695_ );
and  ( new_n31848_, new_n31847_, new_n31770_ );
or   ( new_n31849_, new_n31763_, new_n31757_ );
or   ( new_n31850_, new_n31701_, new_n31698_ );
and  ( new_n31851_, new_n31850_, new_n31719_ );
or   ( new_n31852_, new_n31851_, new_n31702_ );
and  ( new_n31853_, new_n31852_, new_n31849_ );
or   ( new_n31854_, new_n31853_, new_n31848_ );
or   ( new_n31855_, new_n857_, new_n755_ );
or   ( new_n31856_, new_n861_, new_n591_ );
and  ( new_n31857_, new_n31856_, new_n31855_ );
and  ( new_n31858_, new_n31857_, new_n842_ );
and  ( new_n31859_, new_n870_, RI2b1c4342d738_70 );
and  ( new_n31860_, new_n855_, RI2b1c4342d6c0_69 );
or   ( new_n31861_, new_n31860_, new_n31859_ );
and  ( new_n31862_, new_n31861_, new_n866_ );
or   ( new_n31863_, new_n31862_, new_n31858_ );
and  ( new_n31864_, new_n31863_, new_n31854_ );
and  ( new_n31865_, new_n31852_, new_n31770_ );
and  ( new_n31866_, new_n31849_, new_n31847_ );
or   ( new_n31867_, new_n31866_, new_n31865_ );
and  ( new_n31868_, new_n31861_, new_n842_ );
and  ( new_n31869_, new_n31857_, new_n866_ );
or   ( new_n31870_, new_n31869_, new_n31868_ );
and  ( new_n31871_, new_n31870_, new_n31867_ );
or   ( new_n31872_, new_n31871_, new_n31864_ );
and  ( new_n31873_, new_n31872_, new_n31844_ );
and  ( new_n31874_, new_n31842_, new_n31832_ );
and  ( new_n31875_, new_n31839_, new_n31835_ );
or   ( new_n31876_, new_n31875_, new_n31874_ );
and  ( new_n31877_, new_n31867_, new_n31863_ );
and  ( new_n31878_, new_n31870_, new_n31854_ );
or   ( new_n31879_, new_n31878_, new_n31877_ );
and  ( new_n31880_, new_n31879_, new_n31876_ );
or   ( new_n31881_, new_n31880_, new_n31873_ );
or   ( new_n31882_, new_n31724_, new_n31721_ );
and  ( new_n31883_, new_n31882_, new_n31774_ );
or   ( new_n31884_, new_n31883_, new_n31725_ );
and  ( new_n31885_, new_n31884_, new_n31881_ );
and  ( new_n31886_, new_n31876_, new_n31872_ );
and  ( new_n31887_, new_n31879_, new_n31844_ );
or   ( new_n31888_, new_n31887_, new_n31886_ );
or   ( new_n31889_, new_n31731_, new_n31728_ );
or   ( new_n31890_, new_n31781_, new_n31732_ );
and  ( new_n31891_, new_n31890_, new_n31889_ );
and  ( new_n31892_, new_n31891_, new_n31888_ );
or   ( new_n31893_, new_n31892_, new_n31885_ );
or   ( new_n31894_, new_n31664_, new_n31661_ );
and  ( new_n31895_, new_n31894_, new_n31783_ );
or   ( new_n31896_, new_n31895_, new_n31665_ );
and  ( new_n31897_, new_n31896_, new_n31893_ );
or   ( new_n31898_, new_n31825_, new_n31818_ );
or   ( new_n31899_, new_n31847_, new_n31770_ );
and  ( new_n31900_, new_n31899_, new_n31863_ );
or   ( new_n31901_, new_n31900_, new_n31848_ );
and  ( new_n31902_, new_n31901_, new_n31898_ );
or   ( new_n31903_, new_n31852_, new_n31849_ );
and  ( new_n31904_, new_n31903_, new_n31870_ );
or   ( new_n31905_, new_n31904_, new_n31853_ );
and  ( new_n31906_, new_n31905_, new_n31831_ );
or   ( new_n31907_, new_n31906_, new_n31902_ );
or   ( new_n31908_, new_n31359_, new_n31298_ );
and  ( new_n31909_, new_n31908_, new_n31315_ );
and  ( new_n31910_, new_n31358_, new_n31275_ );
and  ( new_n31911_, new_n31297_, new_n31235_ );
or   ( new_n31912_, new_n31911_, new_n31910_ );
and  ( new_n31913_, new_n31912_, new_n31362_ );
or   ( new_n31914_, new_n31913_, new_n31909_ );
and  ( new_n31915_, new_n31914_, new_n31907_ );
and  ( new_n31916_, new_n31905_, new_n31898_ );
and  ( new_n31917_, new_n31901_, new_n31831_ );
or   ( new_n31918_, new_n31917_, new_n31916_ );
and  ( new_n31919_, new_n31912_, new_n31315_ );
and  ( new_n31920_, new_n31908_, new_n31362_ );
or   ( new_n31921_, new_n31920_, new_n31919_ );
and  ( new_n31922_, new_n31921_, new_n31918_ );
or   ( new_n31923_, new_n31922_, new_n31915_ );
or   ( new_n31924_, new_n31835_, new_n31832_ );
and  ( new_n31925_, new_n31924_, new_n31872_ );
or   ( new_n31926_, new_n31925_, new_n31836_ );
and  ( new_n31927_, new_n31926_, new_n31923_ );
and  ( new_n31928_, new_n31918_, new_n31914_ );
and  ( new_n31929_, new_n31921_, new_n31907_ );
or   ( new_n31930_, new_n31929_, new_n31928_ );
or   ( new_n31931_, new_n31842_, new_n31839_ );
or   ( new_n31932_, new_n31879_, new_n31843_ );
and  ( new_n31933_, new_n31932_, new_n31931_ );
and  ( new_n31934_, new_n31933_, new_n31930_ );
or   ( new_n31935_, new_n31934_, new_n31927_ );
or   ( new_n31936_, new_n31884_, new_n31881_ );
and  ( new_n31937_, new_n31936_, new_n31935_ );
or   ( new_n31938_, new_n31937_, new_n31897_ );
or   ( new_n31939_, new_n31366_, new_n31319_ );
and  ( new_n31940_, new_n31939_, new_n31331_ );
and  ( new_n31941_, new_n31365_, new_n31274_ );
and  ( new_n31942_, new_n31348_, new_n31318_ );
or   ( new_n31943_, new_n31942_, new_n31941_ );
and  ( new_n31944_, new_n31943_, new_n31369_ );
or   ( new_n31945_, new_n31944_, new_n31940_ );
or   ( new_n31946_, new_n31901_, new_n31898_ );
and  ( new_n31947_, new_n31946_, new_n31914_ );
or   ( new_n31948_, new_n31947_, new_n31902_ );
and  ( new_n31949_, new_n31948_, new_n31945_ );
and  ( new_n31950_, new_n31943_, new_n31331_ );
and  ( new_n31951_, new_n31939_, new_n31369_ );
or   ( new_n31952_, new_n31951_, new_n31950_ );
or   ( new_n31953_, new_n31905_, new_n31831_ );
or   ( new_n31954_, new_n31921_, new_n31906_ );
and  ( new_n31955_, new_n31954_, new_n31953_ );
and  ( new_n31956_, new_n31955_, new_n31952_ );
or   ( new_n31957_, new_n31956_, new_n31949_ );
or   ( new_n31958_, new_n31926_, new_n31923_ );
and  ( new_n31959_, new_n31958_, new_n31957_ );
or   ( new_n31960_, new_n31376_, new_n31335_ );
and  ( new_n31961_, new_n31960_, new_n31338_ );
and  ( new_n31962_, new_n31372_, new_n31267_ );
and  ( new_n31963_, new_n31375_, new_n31334_ );
or   ( new_n31964_, new_n31963_, new_n31962_ );
and  ( new_n31965_, new_n31964_, new_n31378_ );
or   ( new_n31966_, new_n31965_, new_n31961_ );
or   ( new_n31967_, new_n31948_, new_n31945_ );
and  ( new_n31968_, new_n31967_, new_n31966_ );
or   ( new_n31969_, new_n31968_, new_n31959_ );
or   ( new_n31970_, new_n31969_, new_n31938_ );
or   ( new_n31971_, new_n31970_, new_n31817_ );
or   ( new_n31972_, new_n31971_, new_n4382_ );
or   ( new_n31973_, new_n31972_, new_n31385_ );
or   ( new_n31974_, new_n31971_, new_n4378_ );
or   ( new_n31975_, new_n15321_, new_n15316_ );
or   ( new_n31976_, new_n31975_, new_n31972_ );
or   ( new_n31977_, new_n31814_, new_n31813_ );
or   ( new_n31978_, new_n31803_, new_n31792_ );
and  ( new_n31979_, new_n31978_, new_n31977_ );
or   ( new_n31980_, new_n31979_, new_n31804_ );
or   ( new_n31981_, new_n31543_, new_n31542_ );
and  ( new_n31982_, new_n31981_, new_n15500_ );
or   ( new_n31983_, new_n31982_, new_n31544_ );
or   ( new_n31984_, new_n31983_, new_n31816_ );
and  ( new_n31985_, new_n31984_, new_n31980_ );
or   ( new_n31986_, new_n31985_, new_n31970_ );
or   ( new_n31987_, new_n31958_, new_n31957_ );
or   ( new_n31988_, new_n31967_, new_n31966_ );
and  ( new_n31989_, new_n31988_, new_n31987_ );
or   ( new_n31990_, new_n31989_, new_n31968_ );
or   ( new_n31991_, new_n31896_, new_n31893_ );
or   ( new_n31992_, new_n31936_, new_n31935_ );
and  ( new_n31993_, new_n31992_, new_n31991_ );
or   ( new_n31994_, new_n31993_, new_n31937_ );
or   ( new_n31995_, new_n31994_, new_n31969_ );
and  ( new_n31996_, new_n31995_, new_n31990_ );
and  ( new_n31997_, new_n31996_, new_n31986_ );
and  ( new_n31998_, new_n31997_, new_n31976_ );
and  ( new_n31999_, new_n31998_, new_n31974_ );
and  ( new_n32000_, new_n31999_, new_n31973_ );
and  ( new_n32001_, new_n32000_, new_n31383_ );
and  ( new_n32002_, new_n31341_, new_n31234_ );
and  ( new_n32003_, new_n31381_, new_n31345_ );
or   ( new_n32004_, new_n32003_, new_n32002_ );
and  ( new_n32005_, new_n15994_, new_n15729_ );
or   ( new_n32006_, new_n32005_, new_n15648_ );
and  ( new_n32007_, new_n31540_, new_n31530_ );
and  ( new_n32008_, new_n31537_, new_n31533_ );
or   ( new_n32009_, new_n32008_, new_n32007_ );
or   ( new_n32010_, new_n32009_, new_n15490_ );
and  ( new_n32011_, new_n32010_, new_n15504_ );
and  ( new_n32012_, new_n31787_, new_n31783_ );
and  ( new_n32013_, new_n31790_, new_n31680_ );
or   ( new_n32014_, new_n32013_, new_n32012_ );
or   ( new_n32015_, new_n32014_, new_n31811_ );
and  ( new_n32016_, new_n31810_, new_n31799_ );
and  ( new_n32017_, new_n31807_, new_n31802_ );
or   ( new_n32018_, new_n32017_, new_n32016_ );
or   ( new_n32019_, new_n32018_, new_n31541_ );
and  ( new_n32020_, new_n32019_, new_n32015_ );
and  ( new_n32021_, new_n32020_, new_n32011_ );
and  ( new_n32022_, new_n31891_, new_n31881_ );
and  ( new_n32023_, new_n31888_, new_n31884_ );
or   ( new_n32024_, new_n32023_, new_n32022_ );
or   ( new_n32025_, new_n31678_, new_n31668_ );
and  ( new_n32026_, new_n32025_, new_n31790_ );
or   ( new_n32027_, new_n32026_, new_n31679_ );
or   ( new_n32028_, new_n32027_, new_n32024_ );
and  ( new_n32029_, new_n31933_, new_n31923_ );
and  ( new_n32030_, new_n31930_, new_n31926_ );
or   ( new_n32031_, new_n32030_, new_n32029_ );
or   ( new_n32032_, new_n32031_, new_n31892_ );
and  ( new_n32033_, new_n32032_, new_n32028_ );
and  ( new_n32034_, new_n31955_, new_n31945_ );
and  ( new_n32035_, new_n31952_, new_n31948_ );
or   ( new_n32036_, new_n32035_, new_n32034_ );
or   ( new_n32037_, new_n32036_, new_n31934_ );
and  ( new_n32038_, new_n31964_, new_n31338_ );
and  ( new_n32039_, new_n31960_, new_n31378_ );
or   ( new_n32040_, new_n32039_, new_n32038_ );
or   ( new_n32041_, new_n32040_, new_n31956_ );
and  ( new_n32042_, new_n32041_, new_n32037_ );
and  ( new_n32043_, new_n32042_, new_n32033_ );
and  ( new_n32044_, new_n32043_, new_n32021_ );
and  ( new_n32045_, new_n32044_, new_n15573_ );
and  ( new_n32046_, new_n32045_, new_n32006_ );
and  ( new_n32047_, new_n32044_, new_n15569_ );
and  ( new_n32048_, new_n15994_, new_n15989_ );
and  ( new_n32049_, new_n32048_, new_n32045_ );
and  ( new_n32050_, new_n32014_, new_n31811_ );
and  ( new_n32051_, new_n32018_, new_n31541_ );
and  ( new_n32052_, new_n32051_, new_n32015_ );
or   ( new_n32053_, new_n32052_, new_n32050_ );
and  ( new_n32054_, new_n32009_, new_n15490_ );
and  ( new_n32055_, new_n32010_, new_n15508_ );
or   ( new_n32056_, new_n32055_, new_n32054_ );
and  ( new_n32057_, new_n32056_, new_n32020_ );
or   ( new_n32058_, new_n32057_, new_n32053_ );
and  ( new_n32059_, new_n32058_, new_n32043_ );
and  ( new_n32060_, new_n32040_, new_n31956_ );
and  ( new_n32061_, new_n32036_, new_n31934_ );
and  ( new_n32062_, new_n32061_, new_n32041_ );
or   ( new_n32063_, new_n32062_, new_n32060_ );
and  ( new_n32064_, new_n32031_, new_n31892_ );
and  ( new_n32065_, new_n32027_, new_n32024_ );
and  ( new_n32066_, new_n32065_, new_n32032_ );
or   ( new_n32067_, new_n32066_, new_n32064_ );
and  ( new_n32068_, new_n32067_, new_n32042_ );
or   ( new_n32069_, new_n32068_, new_n32063_ );
or   ( new_n32070_, new_n32069_, new_n32059_ );
or   ( new_n32071_, new_n32070_, new_n32049_ );
or   ( new_n32072_, new_n32071_, new_n32047_ );
or   ( new_n32073_, new_n32072_, new_n32046_ );
and  ( new_n32074_, new_n32073_, new_n32004_ );
or   ( new_n32075_, new_n32074_, new_n32001_ );
and  ( new_n32076_, new_n16102_, RI2b1c4342d5d0_67 );
or   ( new_n32077_, new_n16119_, new_n526_ );
or   ( new_n32078_, new_n16123_, new_n99_ );
and  ( new_n32079_, new_n32078_, new_n32077_ );
or   ( new_n32080_, new_n32079_, new_n16108_ );
and  ( new_n32081_, new_n16132_, RI2b1c4342d558_66 );
and  ( new_n32082_, new_n16114_, RI2b1c4342d4e0_65 );
or   ( new_n32083_, new_n32082_, new_n32081_ );
or   ( new_n32084_, new_n32083_, new_n16128_ );
and  ( new_n32085_, new_n32084_, new_n32080_ );
or   ( new_n32086_, new_n32085_, new_n16151_ );
or   ( new_n32087_, new_n32083_, new_n16108_ );
or   ( new_n32088_, new_n32079_, new_n16128_ );
and  ( new_n32089_, new_n32088_, new_n32087_ );
or   ( new_n32090_, new_n32089_, new_n16170_ );
and  ( new_n32091_, new_n32090_, new_n32086_ );
or   ( new_n32092_, new_n32091_, new_n32076_ );
or   ( new_n32093_, new_n16115_, new_n112_ );
or   ( new_n32094_, new_n32089_, new_n16151_ );
or   ( new_n32095_, new_n32085_, new_n16170_ );
and  ( new_n32096_, new_n32095_, new_n32094_ );
or   ( new_n32097_, new_n32096_, new_n32093_ );
and  ( new_n32098_, new_n32097_, new_n32092_ );
and  ( new_n32099_, new_n16162_, RI2b1c4342d4e0_65 );
or   ( new_n32100_, new_n32099_, new_n16151_ );
or   ( new_n32101_, new_n16174_, new_n99_ );
or   ( new_n32102_, new_n32101_, new_n16170_ );
and  ( new_n32103_, new_n32102_, new_n32100_ );
and  ( new_n32104_, new_n16132_, RI2b1c4342d5d0_67 );
and  ( new_n32105_, new_n16114_, RI2b1c4342d558_66 );
or   ( new_n32106_, new_n32105_, new_n32104_ );
or   ( new_n32107_, new_n32106_, new_n16108_ );
or   ( new_n32108_, new_n16119_, new_n112_ );
or   ( new_n32109_, new_n16123_, new_n526_ );
and  ( new_n32110_, new_n32109_, new_n32108_ );
or   ( new_n32111_, new_n32110_, new_n16128_ );
and  ( new_n32112_, new_n32111_, new_n32107_ );
or   ( new_n32113_, new_n32112_, new_n32103_ );
or   ( new_n32114_, new_n32101_, new_n16151_ );
or   ( new_n32115_, new_n32099_, new_n16170_ );
and  ( new_n32116_, new_n32115_, new_n32114_ );
or   ( new_n32117_, new_n32110_, new_n16108_ );
or   ( new_n32118_, new_n32106_, new_n16128_ );
and  ( new_n32119_, new_n32118_, new_n32117_ );
or   ( new_n32120_, new_n32119_, new_n32116_ );
and  ( new_n32121_, new_n32120_, new_n32113_ );
and  ( new_n32122_, new_n16102_, RI2b1c4342d648_68 );
or   ( new_n32123_, new_n32122_, new_n32121_ );
or   ( new_n32124_, new_n32116_, new_n32112_ );
or   ( new_n32125_, new_n32119_, new_n32103_ );
and  ( new_n32126_, new_n32125_, new_n32124_ );
or   ( new_n32127_, new_n16115_, new_n612_ );
or   ( new_n32128_, new_n32127_, new_n32126_ );
and  ( new_n32129_, new_n32128_, new_n32123_ );
and  ( new_n32130_, new_n16162_, RI2b1c4342d558_66 );
and  ( new_n32131_, new_n16165_, RI2b1c4342d4e0_65 );
or   ( new_n32132_, new_n32131_, new_n32130_ );
or   ( new_n32133_, new_n32132_, new_n16151_ );
or   ( new_n32134_, new_n16174_, new_n526_ );
or   ( new_n32135_, new_n16160_, new_n99_ );
and  ( new_n32136_, new_n32135_, new_n32134_ );
or   ( new_n32137_, new_n32136_, new_n16170_ );
and  ( new_n32138_, new_n32137_, new_n32133_ );
or   ( new_n32139_, new_n32138_, new_n16234_ );
and  ( new_n32140_, new_n16132_, RI2b1c4342d648_68 );
and  ( new_n32141_, new_n16114_, RI2b1c4342d5d0_67 );
or   ( new_n32142_, new_n32141_, new_n32140_ );
or   ( new_n32143_, new_n32142_, new_n16108_ );
or   ( new_n32144_, new_n16119_, new_n612_ );
or   ( new_n32145_, new_n16123_, new_n112_ );
and  ( new_n32146_, new_n32145_, new_n32144_ );
or   ( new_n32147_, new_n32146_, new_n16128_ );
and  ( new_n32148_, new_n32147_, new_n32143_ );
and  ( new_n32149_, new_n32138_, new_n16234_ );
or   ( new_n32150_, new_n32149_, new_n32148_ );
and  ( new_n32151_, new_n32150_, new_n32139_ );
or   ( new_n32152_, new_n32151_, new_n32129_ );
and  ( new_n32153_, new_n32112_, new_n32103_ );
or   ( new_n32154_, new_n32153_, new_n32122_ );
and  ( new_n32155_, new_n32154_, new_n32113_ );
or   ( new_n32156_, new_n32155_, new_n32152_ );
or   ( new_n32157_, new_n32126_, new_n32122_ );
or   ( new_n32158_, new_n32127_, new_n32121_ );
and  ( new_n32159_, new_n32158_, new_n32157_ );
or   ( new_n32160_, new_n32136_, new_n16151_ );
or   ( new_n32161_, new_n32132_, new_n16170_ );
and  ( new_n32162_, new_n32161_, new_n32160_ );
or   ( new_n32163_, new_n32162_, new_n16217_ );
or   ( new_n32164_, new_n32146_, new_n16108_ );
or   ( new_n32165_, new_n32142_, new_n16128_ );
and  ( new_n32166_, new_n32165_, new_n32164_ );
and  ( new_n32167_, new_n32162_, new_n16217_ );
or   ( new_n32168_, new_n32167_, new_n32166_ );
and  ( new_n32169_, new_n32168_, new_n32163_ );
and  ( new_n32170_, new_n32169_, new_n32159_ );
and  ( new_n32171_, new_n32119_, new_n32116_ );
and  ( new_n32172_, new_n32127_, new_n32120_ );
or   ( new_n32173_, new_n32172_, new_n32171_ );
or   ( new_n32174_, new_n32173_, new_n32170_ );
and  ( new_n32175_, new_n32174_, new_n32156_ );
or   ( new_n32176_, new_n32175_, new_n32098_ );
or   ( new_n32177_, new_n32170_, new_n32155_ );
or   ( new_n32178_, new_n32173_, new_n32152_ );
and  ( new_n32179_, new_n32178_, new_n32177_ );
or   ( new_n32180_, new_n32096_, new_n32076_ );
or   ( new_n32181_, new_n32093_, new_n32091_ );
and  ( new_n32182_, new_n32181_, new_n32180_ );
or   ( new_n32183_, new_n32182_, new_n32179_ );
and  ( new_n32184_, new_n32183_, new_n32176_ );
and  ( new_n32185_, new_n16102_, RI2b1c4342d738_70 );
and  ( new_n32186_, new_n16226_, RI2b1c4342d4e0_65 );
or   ( new_n32187_, new_n32186_, new_n16217_ );
or   ( new_n32188_, new_n16238_, new_n99_ );
or   ( new_n32189_, new_n32188_, new_n16234_ );
and  ( new_n32190_, new_n32189_, new_n32187_ );
and  ( new_n32191_, new_n16162_, RI2b1c4342d5d0_67 );
and  ( new_n32192_, new_n16165_, RI2b1c4342d558_66 );
or   ( new_n32193_, new_n32192_, new_n32191_ );
or   ( new_n32194_, new_n32193_, new_n16151_ );
or   ( new_n32195_, new_n16174_, new_n112_ );
or   ( new_n32196_, new_n16160_, new_n526_ );
and  ( new_n32197_, new_n32196_, new_n32195_ );
or   ( new_n32198_, new_n32197_, new_n16170_ );
and  ( new_n32199_, new_n32198_, new_n32194_ );
or   ( new_n32200_, new_n32199_, new_n32190_ );
and  ( new_n32201_, new_n16132_, RI2b1c4342d6c0_69 );
and  ( new_n32202_, new_n16114_, RI2b1c4342d648_68 );
or   ( new_n32203_, new_n32202_, new_n32201_ );
or   ( new_n32204_, new_n32203_, new_n16108_ );
or   ( new_n32205_, new_n16119_, new_n591_ );
or   ( new_n32206_, new_n16123_, new_n612_ );
and  ( new_n32207_, new_n32206_, new_n32205_ );
or   ( new_n32208_, new_n32207_, new_n16128_ );
and  ( new_n32209_, new_n32208_, new_n32204_ );
and  ( new_n32210_, new_n32199_, new_n32190_ );
or   ( new_n32211_, new_n32210_, new_n32209_ );
and  ( new_n32212_, new_n32211_, new_n32200_ );
or   ( new_n32213_, new_n32212_, new_n32185_ );
and  ( new_n32214_, new_n16102_, RI2b1c4342d6c0_69 );
and  ( new_n32215_, new_n32212_, new_n32185_ );
or   ( new_n32216_, new_n32215_, new_n32214_ );
and  ( new_n32217_, new_n32216_, new_n32213_ );
and  ( new_n32218_, new_n32163_, new_n32139_ );
or   ( new_n32219_, new_n32218_, new_n32148_ );
or   ( new_n32220_, new_n32138_, new_n16217_ );
or   ( new_n32221_, new_n32162_, new_n16234_ );
and  ( new_n32222_, new_n32221_, new_n32220_ );
or   ( new_n32223_, new_n32222_, new_n32166_ );
and  ( new_n32224_, new_n32223_, new_n32219_ );
or   ( new_n32225_, new_n16115_, new_n755_ );
and  ( new_n32226_, new_n16226_, RI2b1c4342d558_66 );
and  ( new_n32227_, new_n16229_, RI2b1c4342d4e0_65 );
or   ( new_n32228_, new_n32227_, new_n32226_ );
or   ( new_n32229_, new_n32228_, new_n16217_ );
or   ( new_n32230_, new_n16238_, new_n526_ );
or   ( new_n32231_, new_n16224_, new_n99_ );
and  ( new_n32232_, new_n32231_, new_n32230_ );
or   ( new_n32233_, new_n32232_, new_n16234_ );
and  ( new_n32234_, new_n32233_, new_n32229_ );
or   ( new_n32235_, new_n32234_, new_n16204_ );
and  ( new_n32236_, new_n16162_, RI2b1c4342d648_68 );
and  ( new_n32237_, new_n16165_, RI2b1c4342d5d0_67 );
or   ( new_n32238_, new_n32237_, new_n32236_ );
or   ( new_n32239_, new_n32238_, new_n16151_ );
or   ( new_n32240_, new_n16174_, new_n612_ );
or   ( new_n32241_, new_n16160_, new_n112_ );
and  ( new_n32242_, new_n32241_, new_n32240_ );
or   ( new_n32243_, new_n32242_, new_n16170_ );
and  ( new_n32244_, new_n32243_, new_n32239_ );
and  ( new_n32245_, new_n32234_, new_n16204_ );
or   ( new_n32246_, new_n32245_, new_n32244_ );
and  ( new_n32247_, new_n32246_, new_n32235_ );
or   ( new_n32248_, new_n32247_, new_n32225_ );
or   ( new_n32249_, new_n32188_, new_n16217_ );
or   ( new_n32250_, new_n32186_, new_n16234_ );
and  ( new_n32251_, new_n32250_, new_n32249_ );
or   ( new_n32252_, new_n32197_, new_n16151_ );
or   ( new_n32253_, new_n32193_, new_n16170_ );
and  ( new_n32254_, new_n32253_, new_n32252_ );
or   ( new_n32255_, new_n32254_, new_n32251_ );
and  ( new_n32256_, new_n32255_, new_n32200_ );
or   ( new_n32257_, new_n32256_, new_n32209_ );
or   ( new_n32258_, new_n32251_, new_n32199_ );
or   ( new_n32259_, new_n32254_, new_n32190_ );
and  ( new_n32260_, new_n32259_, new_n32258_ );
or   ( new_n32261_, new_n32207_, new_n16108_ );
or   ( new_n32262_, new_n32203_, new_n16128_ );
and  ( new_n32263_, new_n32262_, new_n32261_ );
or   ( new_n32264_, new_n32263_, new_n32260_ );
and  ( new_n32265_, new_n32264_, new_n32257_ );
and  ( new_n32266_, new_n32247_, new_n32225_ );
or   ( new_n32267_, new_n32266_, new_n32265_ );
and  ( new_n32268_, new_n32267_, new_n32248_ );
or   ( new_n32269_, new_n32268_, new_n32224_ );
and  ( new_n32270_, new_n32254_, new_n32251_ );
or   ( new_n32271_, new_n32270_, new_n32263_ );
and  ( new_n32272_, new_n32271_, new_n32255_ );
or   ( new_n32273_, new_n32272_, new_n32225_ );
and  ( new_n32274_, new_n32273_, new_n32213_ );
or   ( new_n32275_, new_n32274_, new_n32214_ );
or   ( new_n32276_, new_n32272_, new_n32185_ );
or   ( new_n32277_, new_n32225_, new_n32212_ );
and  ( new_n32278_, new_n32277_, new_n32276_ );
or   ( new_n32279_, new_n16115_, new_n591_ );
or   ( new_n32280_, new_n32279_, new_n32278_ );
and  ( new_n32281_, new_n32280_, new_n32275_ );
and  ( new_n32282_, new_n32268_, new_n32224_ );
or   ( new_n32283_, new_n32282_, new_n32281_ );
and  ( new_n32284_, new_n32283_, new_n32269_ );
or   ( new_n32285_, new_n32284_, new_n32217_ );
or   ( new_n32286_, new_n32169_, new_n32129_ );
or   ( new_n32287_, new_n32159_, new_n32151_ );
and  ( new_n32288_, new_n32287_, new_n32286_ );
and  ( new_n32289_, new_n32284_, new_n32217_ );
or   ( new_n32290_, new_n32289_, new_n32288_ );
and  ( new_n32291_, new_n32290_, new_n32285_ );
and  ( new_n32292_, new_n32291_, new_n32184_ );
or   ( new_n32293_, new_n32179_, new_n32098_ );
or   ( new_n32294_, new_n32182_, new_n32175_ );
and  ( new_n32295_, new_n32294_, new_n32293_ );
or   ( new_n32296_, new_n32222_, new_n32148_ );
or   ( new_n32297_, new_n32218_, new_n32166_ );
and  ( new_n32298_, new_n32297_, new_n32296_ );
or   ( new_n32299_, new_n32232_, new_n16217_ );
or   ( new_n32300_, new_n32228_, new_n16234_ );
and  ( new_n32301_, new_n32300_, new_n32299_ );
or   ( new_n32302_, new_n32301_, new_n16186_ );
or   ( new_n32303_, new_n32242_, new_n16151_ );
or   ( new_n32304_, new_n32238_, new_n16170_ );
and  ( new_n32305_, new_n32304_, new_n32303_ );
and  ( new_n32306_, new_n32301_, new_n16186_ );
or   ( new_n32307_, new_n32306_, new_n32305_ );
and  ( new_n32308_, new_n32307_, new_n32302_ );
or   ( new_n32309_, new_n32308_, new_n32185_ );
or   ( new_n32310_, new_n32260_, new_n32209_ );
or   ( new_n32311_, new_n32263_, new_n32256_ );
and  ( new_n32312_, new_n32311_, new_n32310_ );
and  ( new_n32313_, new_n32308_, new_n32185_ );
or   ( new_n32314_, new_n32313_, new_n32312_ );
and  ( new_n32315_, new_n32314_, new_n32309_ );
or   ( new_n32316_, new_n32315_, new_n32298_ );
or   ( new_n32317_, new_n32278_, new_n32214_ );
or   ( new_n32318_, new_n32279_, new_n32274_ );
and  ( new_n32319_, new_n32318_, new_n32317_ );
and  ( new_n32320_, new_n32315_, new_n32298_ );
or   ( new_n32321_, new_n32320_, new_n32319_ );
and  ( new_n32322_, new_n32321_, new_n32316_ );
and  ( new_n32323_, new_n32272_, new_n32225_ );
or   ( new_n32324_, new_n32323_, new_n32279_ );
and  ( new_n32325_, new_n32324_, new_n32273_ );
or   ( new_n32326_, new_n32325_, new_n32322_ );
or   ( new_n32327_, new_n32169_, new_n32159_ );
and  ( new_n32328_, new_n32327_, new_n32152_ );
and  ( new_n32329_, new_n32325_, new_n32322_ );
or   ( new_n32330_, new_n32329_, new_n32328_ );
and  ( new_n32331_, new_n32330_, new_n32326_ );
and  ( new_n32332_, new_n32331_, new_n32295_ );
or   ( new_n32333_, new_n32332_, new_n32292_ );
and  ( new_n32334_, new_n16021_, RI2b1c4342d4e0_65 );
or   ( new_n32335_, new_n32334_, new_n16009_ );
or   ( new_n32336_, new_n16033_, new_n99_ );
or   ( new_n32337_, new_n32336_, new_n16029_ );
and  ( new_n32338_, new_n32337_, new_n32335_ );
and  ( new_n32339_, new_n16196_, RI2b1c4342d5d0_67 );
and  ( new_n32340_, new_n16199_, RI2b1c4342d558_66 );
or   ( new_n32341_, new_n32340_, new_n32339_ );
or   ( new_n32342_, new_n32341_, new_n16186_ );
or   ( new_n32343_, new_n16208_, new_n112_ );
or   ( new_n32344_, new_n16194_, new_n526_ );
and  ( new_n32345_, new_n32344_, new_n32343_ );
or   ( new_n32346_, new_n32345_, new_n16204_ );
and  ( new_n32347_, new_n32346_, new_n32342_ );
or   ( new_n32348_, new_n32347_, new_n32338_ );
or   ( new_n32349_, new_n32336_, new_n16009_ );
or   ( new_n32350_, new_n32334_, new_n16029_ );
and  ( new_n32351_, new_n32350_, new_n32349_ );
or   ( new_n32352_, new_n32345_, new_n16186_ );
or   ( new_n32353_, new_n32341_, new_n16204_ );
and  ( new_n32354_, new_n32353_, new_n32352_ );
or   ( new_n32355_, new_n32354_, new_n32351_ );
and  ( new_n32356_, new_n32355_, new_n32348_ );
and  ( new_n32357_, new_n16226_, RI2b1c4342d6c0_69 );
and  ( new_n32358_, new_n16229_, RI2b1c4342d648_68 );
or   ( new_n32359_, new_n32358_, new_n32357_ );
or   ( new_n32360_, new_n32359_, new_n16217_ );
or   ( new_n32361_, new_n16238_, new_n591_ );
or   ( new_n32362_, new_n16224_, new_n612_ );
and  ( new_n32363_, new_n32362_, new_n32361_ );
or   ( new_n32364_, new_n32363_, new_n16234_ );
and  ( new_n32365_, new_n32364_, new_n32360_ );
or   ( new_n32366_, new_n32365_, new_n32356_ );
or   ( new_n32367_, new_n32351_, new_n32347_ );
or   ( new_n32368_, new_n32354_, new_n32338_ );
and  ( new_n32369_, new_n32368_, new_n32367_ );
or   ( new_n32370_, new_n32363_, new_n16217_ );
or   ( new_n32371_, new_n32359_, new_n16234_ );
and  ( new_n32372_, new_n32371_, new_n32370_ );
or   ( new_n32373_, new_n32372_, new_n32369_ );
and  ( new_n32374_, new_n32373_, new_n32366_ );
and  ( new_n32375_, new_n30471_, new_n16052_ );
or   ( new_n32376_, new_n32375_, new_n30481_ );
and  ( new_n32377_, new_n32376_, new_n30472_ );
and  ( new_n32378_, new_n30514_, new_n30505_ );
or   ( new_n32379_, new_n32378_, new_n30496_ );
and  ( new_n32380_, new_n32379_, new_n30515_ );
or   ( new_n32381_, new_n32380_, new_n32377_ );
and  ( new_n32382_, new_n30521_, new_n30518_ );
or   ( new_n32383_, new_n32382_, new_n30527_ );
and  ( new_n32384_, new_n32383_, new_n30522_ );
and  ( new_n32385_, new_n30475_, new_n16071_ );
or   ( new_n32386_, new_n32385_, new_n30462_ );
and  ( new_n32387_, new_n32386_, new_n30476_ );
or   ( new_n32388_, new_n32387_, new_n32384_ );
and  ( new_n32389_, new_n32388_, new_n32381_ );
and  ( new_n32390_, new_n32389_, new_n32374_ );
and  ( new_n32391_, new_n30578_, new_n30575_ );
or   ( new_n32392_, new_n32391_, new_n17014_ );
and  ( new_n32393_, new_n32392_, new_n30579_ );
and  ( new_n32394_, new_n30532_, new_n30487_ );
or   ( new_n32395_, new_n32394_, new_n30486_ );
and  ( new_n32396_, new_n32395_, new_n30533_ );
or   ( new_n32397_, new_n32396_, new_n32393_ );
and  ( new_n32398_, new_n16162_, RI2b1c4342d7b0_71 );
and  ( new_n32399_, new_n16165_, RI2b1c4342d738_70 );
or   ( new_n32400_, new_n32399_, new_n32398_ );
or   ( new_n32401_, new_n32400_, new_n16151_ );
or   ( new_n32402_, new_n16174_, new_n110_ );
or   ( new_n32403_, new_n16160_, new_n755_ );
and  ( new_n32404_, new_n32403_, new_n32402_ );
or   ( new_n32405_, new_n32404_, new_n16170_ );
and  ( new_n32406_, new_n32405_, new_n32401_ );
and  ( new_n32407_, new_n16132_, RI2b1c4342d8a0_73 );
and  ( new_n32408_, new_n16114_, RI2b1c4342d828_72 );
or   ( new_n32409_, new_n32408_, new_n32407_ );
or   ( new_n32410_, new_n32409_, new_n16108_ );
or   ( new_n32411_, new_n16119_, new_n105_ );
or   ( new_n32412_, new_n16123_, new_n806_ );
and  ( new_n32413_, new_n32412_, new_n32411_ );
or   ( new_n32414_, new_n32413_, new_n16128_ );
and  ( new_n32415_, new_n32414_, new_n32410_ );
or   ( new_n32416_, new_n32415_, new_n32406_ );
or   ( new_n32417_, new_n32404_, new_n16151_ );
or   ( new_n32418_, new_n32400_, new_n16170_ );
and  ( new_n32419_, new_n32418_, new_n32417_ );
or   ( new_n32420_, new_n32413_, new_n16108_ );
or   ( new_n32421_, new_n32409_, new_n16128_ );
and  ( new_n32422_, new_n32421_, new_n32420_ );
or   ( new_n32423_, new_n32422_, new_n32419_ );
and  ( new_n32424_, new_n32423_, new_n32416_ );
and  ( new_n32425_, new_n16102_, RI2b1c4342d918_74 );
or   ( new_n32426_, new_n32425_, new_n32424_ );
or   ( new_n32427_, new_n32419_, new_n32415_ );
or   ( new_n32428_, new_n32422_, new_n32406_ );
and  ( new_n32429_, new_n32428_, new_n32427_ );
or   ( new_n32430_, new_n16115_, new_n859_ );
or   ( new_n32431_, new_n32430_, new_n32429_ );
and  ( new_n32432_, new_n32431_, new_n32426_ );
and  ( new_n32433_, new_n32396_, new_n32393_ );
or   ( new_n32434_, new_n32433_, new_n32432_ );
and  ( new_n32435_, new_n32434_, new_n32397_ );
or   ( new_n32436_, new_n32435_, new_n32390_ );
and  ( new_n32437_, new_n32435_, new_n32390_ );
or   ( new_n32438_, new_n32387_, new_n32380_ );
and  ( new_n32439_, new_n16196_, RI2b1c4342d558_66 );
and  ( new_n32440_, new_n16199_, RI2b1c4342d4e0_65 );
or   ( new_n32441_, new_n32440_, new_n32439_ );
or   ( new_n32442_, new_n32441_, new_n16186_ );
or   ( new_n32443_, new_n16208_, new_n526_ );
or   ( new_n32444_, new_n16194_, new_n99_ );
and  ( new_n32445_, new_n32444_, new_n32443_ );
or   ( new_n32446_, new_n32445_, new_n16204_ );
and  ( new_n32447_, new_n32446_, new_n32442_ );
or   ( new_n32448_, new_n32447_, new_n16029_ );
or   ( new_n32449_, new_n32445_, new_n16186_ );
or   ( new_n32450_, new_n32441_, new_n16204_ );
and  ( new_n32451_, new_n32450_, new_n32449_ );
or   ( new_n32452_, new_n32451_, new_n16009_ );
and  ( new_n32453_, new_n32452_, new_n32448_ );
and  ( new_n32454_, new_n16226_, RI2b1c4342d648_68 );
and  ( new_n32455_, new_n16229_, RI2b1c4342d5d0_67 );
or   ( new_n32456_, new_n32455_, new_n32454_ );
or   ( new_n32457_, new_n32456_, new_n16217_ );
or   ( new_n32458_, new_n16238_, new_n612_ );
or   ( new_n32459_, new_n16224_, new_n112_ );
and  ( new_n32460_, new_n32459_, new_n32458_ );
or   ( new_n32461_, new_n32460_, new_n16234_ );
and  ( new_n32462_, new_n32461_, new_n32457_ );
or   ( new_n32463_, new_n32462_, new_n32453_ );
or   ( new_n32464_, new_n32447_, new_n16009_ );
or   ( new_n32465_, new_n32451_, new_n16029_ );
and  ( new_n32466_, new_n32465_, new_n32464_ );
or   ( new_n32467_, new_n32460_, new_n16217_ );
or   ( new_n32468_, new_n32456_, new_n16234_ );
and  ( new_n32469_, new_n32468_, new_n32467_ );
or   ( new_n32470_, new_n32469_, new_n32466_ );
and  ( new_n32471_, new_n32470_, new_n32463_ );
or   ( new_n32472_, new_n32471_, new_n32438_ );
and  ( new_n32473_, new_n32384_, new_n32377_ );
or   ( new_n32474_, new_n32466_, new_n32462_ );
or   ( new_n32475_, new_n32469_, new_n32453_ );
and  ( new_n32476_, new_n32475_, new_n32474_ );
or   ( new_n32477_, new_n32476_, new_n32473_ );
and  ( new_n32478_, new_n32477_, new_n32472_ );
and  ( new_n32479_, new_n32347_, new_n32338_ );
or   ( new_n32480_, new_n32479_, new_n32365_ );
and  ( new_n32481_, new_n32480_, new_n32348_ );
and  ( new_n32482_, new_n32415_, new_n32406_ );
or   ( new_n32483_, new_n32482_, new_n32425_ );
and  ( new_n32484_, new_n32483_, new_n32416_ );
or   ( new_n32485_, new_n32484_, new_n32481_ );
and  ( new_n32486_, new_n32354_, new_n32351_ );
or   ( new_n32487_, new_n32486_, new_n32372_ );
and  ( new_n32488_, new_n32487_, new_n32355_ );
and  ( new_n32489_, new_n32422_, new_n32419_ );
and  ( new_n32490_, new_n32430_, new_n32423_ );
or   ( new_n32491_, new_n32490_, new_n32489_ );
or   ( new_n32492_, new_n32491_, new_n32488_ );
and  ( new_n32493_, new_n32492_, new_n32485_ );
and  ( new_n32494_, new_n16162_, RI2b1c4342d738_70 );
and  ( new_n32495_, new_n16165_, RI2b1c4342d6c0_69 );
or   ( new_n32496_, new_n32495_, new_n32494_ );
or   ( new_n32497_, new_n32496_, new_n16151_ );
or   ( new_n32498_, new_n16174_, new_n755_ );
or   ( new_n32499_, new_n16160_, new_n591_ );
and  ( new_n32500_, new_n32499_, new_n32498_ );
or   ( new_n32501_, new_n32500_, new_n16170_ );
and  ( new_n32502_, new_n32501_, new_n32497_ );
and  ( new_n32503_, new_n16132_, RI2b1c4342d828_72 );
and  ( new_n32504_, new_n16114_, RI2b1c4342d7b0_71 );
or   ( new_n32505_, new_n32504_, new_n32503_ );
or   ( new_n32506_, new_n32505_, new_n16108_ );
or   ( new_n32507_, new_n16119_, new_n806_ );
or   ( new_n32508_, new_n16123_, new_n110_ );
and  ( new_n32509_, new_n32508_, new_n32507_ );
or   ( new_n32510_, new_n32509_, new_n16128_ );
and  ( new_n32511_, new_n32510_, new_n32506_ );
or   ( new_n32512_, new_n32511_, new_n32502_ );
or   ( new_n32513_, new_n32500_, new_n16151_ );
or   ( new_n32514_, new_n32496_, new_n16170_ );
and  ( new_n32515_, new_n32514_, new_n32513_ );
or   ( new_n32516_, new_n32509_, new_n16108_ );
or   ( new_n32517_, new_n32505_, new_n16128_ );
and  ( new_n32518_, new_n32517_, new_n32516_ );
or   ( new_n32519_, new_n32518_, new_n32515_ );
and  ( new_n32520_, new_n32519_, new_n32512_ );
and  ( new_n32521_, new_n16102_, RI2b1c4342d8a0_73 );
or   ( new_n32522_, new_n32521_, new_n32520_ );
or   ( new_n32523_, new_n32515_, new_n32511_ );
or   ( new_n32524_, new_n32518_, new_n32502_ );
and  ( new_n32525_, new_n32524_, new_n32523_ );
or   ( new_n32526_, new_n16115_, new_n105_ );
or   ( new_n32527_, new_n32526_, new_n32525_ );
and  ( new_n32528_, new_n32527_, new_n32522_ );
or   ( new_n32529_, new_n32528_, new_n32493_ );
or   ( new_n32530_, new_n32488_, new_n32484_ );
or   ( new_n32531_, new_n32491_, new_n32481_ );
and  ( new_n32532_, new_n32531_, new_n32530_ );
or   ( new_n32533_, new_n32525_, new_n32521_ );
or   ( new_n32534_, new_n32526_, new_n32520_ );
and  ( new_n32535_, new_n32534_, new_n32533_ );
or   ( new_n32536_, new_n32535_, new_n32532_ );
and  ( new_n32537_, new_n32536_, new_n32529_ );
or   ( new_n32538_, new_n32537_, new_n32478_ );
or   ( new_n32539_, new_n32473_, new_n32471_ );
or   ( new_n32540_, new_n32476_, new_n32438_ );
and  ( new_n32541_, new_n32540_, new_n32539_ );
or   ( new_n32542_, new_n32532_, new_n32528_ );
or   ( new_n32543_, new_n32535_, new_n32493_ );
and  ( new_n32544_, new_n32543_, new_n32542_ );
or   ( new_n32545_, new_n32544_, new_n32541_ );
and  ( new_n32546_, new_n32545_, new_n32538_ );
or   ( new_n32547_, new_n32546_, new_n32437_ );
and  ( new_n32548_, new_n32547_, new_n32436_ );
and  ( new_n32549_, new_n32471_, new_n32438_ );
or   ( new_n32550_, new_n32549_, new_n32537_ );
and  ( new_n32551_, new_n32550_, new_n32472_ );
or   ( new_n32552_, new_n32551_, new_n32548_ );
and  ( new_n32553_, new_n32476_, new_n32473_ );
or   ( new_n32554_, new_n32553_, new_n32544_ );
and  ( new_n32555_, new_n32554_, new_n32477_ );
or   ( new_n32556_, new_n32369_, new_n32365_ );
or   ( new_n32557_, new_n32372_, new_n32356_ );
and  ( new_n32558_, new_n32557_, new_n32556_ );
or   ( new_n32559_, new_n32384_, new_n32377_ );
and  ( new_n32560_, new_n32559_, new_n32438_ );
or   ( new_n32561_, new_n32560_, new_n32558_ );
and  ( new_n32562_, new_n30585_, new_n30582_ );
and  ( new_n32563_, new_n30586_, new_n16967_ );
or   ( new_n32564_, new_n32563_, new_n32562_ );
and  ( new_n32565_, new_n30537_, new_n30534_ );
or   ( new_n32566_, new_n32565_, new_n30543_ );
and  ( new_n32567_, new_n32566_, new_n30538_ );
or   ( new_n32568_, new_n32567_, new_n32564_ );
or   ( new_n32569_, new_n32429_, new_n32425_ );
or   ( new_n32570_, new_n32430_, new_n32424_ );
and  ( new_n32571_, new_n32570_, new_n32569_ );
and  ( new_n32572_, new_n32567_, new_n32564_ );
or   ( new_n32573_, new_n32572_, new_n32571_ );
and  ( new_n32574_, new_n32573_, new_n32568_ );
or   ( new_n32575_, new_n32574_, new_n32561_ );
and  ( new_n32576_, new_n32574_, new_n32561_ );
or   ( new_n32577_, new_n32541_, new_n32537_ );
or   ( new_n32578_, new_n32544_, new_n32478_ );
and  ( new_n32579_, new_n32578_, new_n32577_ );
or   ( new_n32580_, new_n32579_, new_n32576_ );
and  ( new_n32581_, new_n32580_, new_n32575_ );
or   ( new_n32582_, new_n32581_, new_n32555_ );
and  ( new_n32583_, new_n32582_, new_n32552_ );
and  ( new_n32584_, new_n16196_, RI2b1c4342d4e0_65 );
or   ( new_n32585_, new_n32584_, new_n16186_ );
or   ( new_n32586_, new_n16208_, new_n99_ );
or   ( new_n32587_, new_n32586_, new_n16204_ );
and  ( new_n32588_, new_n32587_, new_n32585_ );
and  ( new_n32589_, new_n16226_, RI2b1c4342d5d0_67 );
and  ( new_n32590_, new_n16229_, RI2b1c4342d558_66 );
or   ( new_n32591_, new_n32590_, new_n32589_ );
or   ( new_n32592_, new_n32591_, new_n16217_ );
or   ( new_n32593_, new_n16238_, new_n112_ );
or   ( new_n32594_, new_n16224_, new_n526_ );
and  ( new_n32595_, new_n32594_, new_n32593_ );
or   ( new_n32596_, new_n32595_, new_n16234_ );
and  ( new_n32597_, new_n32596_, new_n32592_ );
or   ( new_n32598_, new_n32597_, new_n32588_ );
or   ( new_n32599_, new_n32586_, new_n16186_ );
or   ( new_n32600_, new_n32584_, new_n16204_ );
and  ( new_n32601_, new_n32600_, new_n32599_ );
or   ( new_n32602_, new_n32595_, new_n16217_ );
or   ( new_n32603_, new_n32591_, new_n16234_ );
and  ( new_n32604_, new_n32603_, new_n32602_ );
or   ( new_n32605_, new_n32604_, new_n32601_ );
and  ( new_n32606_, new_n32605_, new_n32598_ );
and  ( new_n32607_, new_n16162_, RI2b1c4342d6c0_69 );
and  ( new_n32608_, new_n16165_, RI2b1c4342d648_68 );
or   ( new_n32609_, new_n32608_, new_n32607_ );
or   ( new_n32610_, new_n32609_, new_n16151_ );
or   ( new_n32611_, new_n16174_, new_n591_ );
or   ( new_n32612_, new_n16160_, new_n612_ );
and  ( new_n32613_, new_n32612_, new_n32611_ );
or   ( new_n32614_, new_n32613_, new_n16170_ );
and  ( new_n32615_, new_n32614_, new_n32610_ );
or   ( new_n32616_, new_n32615_, new_n32606_ );
or   ( new_n32617_, new_n32601_, new_n32597_ );
or   ( new_n32618_, new_n32604_, new_n32588_ );
and  ( new_n32619_, new_n32618_, new_n32617_ );
or   ( new_n32620_, new_n32613_, new_n16151_ );
or   ( new_n32621_, new_n32609_, new_n16170_ );
and  ( new_n32622_, new_n32621_, new_n32620_ );
or   ( new_n32623_, new_n32622_, new_n32619_ );
and  ( new_n32624_, new_n32623_, new_n32616_ );
and  ( new_n32625_, new_n32484_, new_n32481_ );
or   ( new_n32626_, new_n32625_, new_n32528_ );
and  ( new_n32627_, new_n32626_, new_n32485_ );
or   ( new_n32628_, new_n32627_, new_n32624_ );
or   ( new_n32629_, new_n32619_, new_n32615_ );
or   ( new_n32630_, new_n32622_, new_n32606_ );
and  ( new_n32631_, new_n32630_, new_n32629_ );
and  ( new_n32632_, new_n32491_, new_n32488_ );
and  ( new_n32633_, new_n32535_, new_n32492_ );
or   ( new_n32634_, new_n32633_, new_n32632_ );
or   ( new_n32635_, new_n32634_, new_n32631_ );
and  ( new_n32636_, new_n32635_, new_n32628_ );
and  ( new_n32637_, new_n32511_, new_n32502_ );
or   ( new_n32638_, new_n32637_, new_n32521_ );
and  ( new_n32639_, new_n32638_, new_n32512_ );
and  ( new_n32640_, new_n32447_, new_n16029_ );
or   ( new_n32641_, new_n32640_, new_n32462_ );
and  ( new_n32642_, new_n32641_, new_n32448_ );
or   ( new_n32643_, new_n32642_, new_n32639_ );
and  ( new_n32644_, new_n32451_, new_n16009_ );
or   ( new_n32645_, new_n32644_, new_n32469_ );
and  ( new_n32646_, new_n32645_, new_n32452_ );
and  ( new_n32647_, new_n32518_, new_n32515_ );
and  ( new_n32648_, new_n32526_, new_n32519_ );
or   ( new_n32649_, new_n32648_, new_n32647_ );
or   ( new_n32650_, new_n32649_, new_n32646_ );
and  ( new_n32651_, new_n32650_, new_n32643_ );
or   ( new_n32652_, new_n16119_, new_n110_ );
or   ( new_n32653_, new_n16123_, new_n755_ );
and  ( new_n32654_, new_n32653_, new_n32652_ );
or   ( new_n32655_, new_n32654_, new_n16108_ );
and  ( new_n32656_, new_n16132_, RI2b1c4342d7b0_71 );
and  ( new_n32657_, new_n16114_, RI2b1c4342d738_70 );
or   ( new_n32658_, new_n32657_, new_n32656_ );
or   ( new_n32659_, new_n32658_, new_n16128_ );
and  ( new_n32660_, new_n32659_, new_n32655_ );
and  ( new_n32661_, new_n16102_, RI2b1c4342d828_72 );
or   ( new_n32662_, new_n32661_, new_n32660_ );
or   ( new_n32663_, new_n32658_, new_n16108_ );
or   ( new_n32664_, new_n32654_, new_n16128_ );
and  ( new_n32665_, new_n32664_, new_n32663_ );
or   ( new_n32666_, new_n16115_, new_n806_ );
or   ( new_n32667_, new_n32666_, new_n32665_ );
and  ( new_n32668_, new_n32667_, new_n32662_ );
or   ( new_n32669_, new_n32668_, new_n32651_ );
or   ( new_n32670_, new_n32646_, new_n32639_ );
or   ( new_n32671_, new_n32649_, new_n32642_ );
and  ( new_n32672_, new_n32671_, new_n32670_ );
or   ( new_n32673_, new_n32665_, new_n32661_ );
or   ( new_n32674_, new_n32666_, new_n32660_ );
and  ( new_n32675_, new_n32674_, new_n32673_ );
or   ( new_n32676_, new_n32675_, new_n32672_ );
and  ( new_n32677_, new_n32676_, new_n32669_ );
or   ( new_n32678_, new_n32677_, new_n32636_ );
or   ( new_n32679_, new_n32634_, new_n32624_ );
or   ( new_n32680_, new_n32631_, new_n32627_ );
and  ( new_n32681_, new_n32680_, new_n32679_ );
or   ( new_n32682_, new_n32672_, new_n32668_ );
or   ( new_n32683_, new_n32675_, new_n32651_ );
and  ( new_n32684_, new_n32683_, new_n32682_ );
or   ( new_n32685_, new_n32684_, new_n32681_ );
and  ( new_n32686_, new_n32685_, new_n32678_ );
or   ( new_n32687_, new_n32686_, new_n32583_ );
or   ( new_n32688_, new_n32581_, new_n32551_ );
or   ( new_n32689_, new_n32555_, new_n32548_ );
and  ( new_n32690_, new_n32689_, new_n32688_ );
or   ( new_n32691_, new_n32681_, new_n32677_ );
or   ( new_n32692_, new_n32684_, new_n32636_ );
and  ( new_n32693_, new_n32692_, new_n32691_ );
or   ( new_n32694_, new_n32693_, new_n32690_ );
and  ( new_n32695_, new_n32694_, new_n32687_ );
and  ( new_n32696_, new_n32575_, new_n32436_ );
or   ( new_n32697_, new_n32696_, new_n32546_ );
or   ( new_n32698_, new_n32574_, new_n32390_ );
or   ( new_n32699_, new_n32561_, new_n32435_ );
and  ( new_n32700_, new_n32699_, new_n32698_ );
or   ( new_n32701_, new_n32700_, new_n32579_ );
and  ( new_n32702_, new_n32701_, new_n32697_ );
or   ( new_n32703_, new_n32389_, new_n32374_ );
and  ( new_n32704_, new_n32703_, new_n32561_ );
and  ( new_n32705_, new_n30554_, new_n30551_ );
or   ( new_n32706_, new_n32705_, new_n30548_ );
and  ( new_n32707_, new_n32706_, new_n30555_ );
or   ( new_n32708_, new_n32707_, new_n32704_ );
and  ( new_n32709_, new_n32568_, new_n32397_ );
or   ( new_n32710_, new_n32709_, new_n32432_ );
or   ( new_n32711_, new_n32564_, new_n32396_ );
or   ( new_n32712_, new_n32567_, new_n32393_ );
and  ( new_n32713_, new_n32712_, new_n32711_ );
or   ( new_n32714_, new_n32713_, new_n32571_ );
and  ( new_n32715_, new_n32714_, new_n32710_ );
and  ( new_n32716_, new_n32707_, new_n32704_ );
or   ( new_n32717_, new_n32716_, new_n32715_ );
and  ( new_n32718_, new_n32717_, new_n32708_ );
and  ( new_n32719_, new_n32718_, new_n32702_ );
or   ( new_n32720_, new_n32719_, new_n32695_ );
or   ( new_n32721_, new_n32700_, new_n32546_ );
or   ( new_n32722_, new_n32696_, new_n32579_ );
and  ( new_n32723_, new_n32722_, new_n32721_ );
or   ( new_n32724_, new_n32558_, new_n32389_ );
or   ( new_n32725_, new_n32560_, new_n32374_ );
and  ( new_n32726_, new_n32725_, new_n32724_ );
and  ( new_n32727_, new_n30561_, new_n30558_ );
and  ( new_n32728_, new_n30567_, new_n30562_ );
or   ( new_n32729_, new_n32728_, new_n32727_ );
and  ( new_n32730_, new_n32729_, new_n32726_ );
or   ( new_n32731_, new_n32729_, new_n32726_ );
or   ( new_n32732_, new_n32713_, new_n32432_ );
or   ( new_n32733_, new_n32709_, new_n32571_ );
and  ( new_n32734_, new_n32733_, new_n32732_ );
and  ( new_n32735_, new_n32734_, new_n32731_ );
or   ( new_n32736_, new_n32735_, new_n32730_ );
or   ( new_n32737_, new_n32736_, new_n32723_ );
or   ( new_n32738_, new_n32718_, new_n32702_ );
and  ( new_n32739_, new_n32738_, new_n32737_ );
and  ( new_n32740_, new_n32731_, new_n32708_ );
or   ( new_n32741_, new_n32740_, new_n32715_ );
or   ( new_n32742_, new_n32729_, new_n32704_ );
or   ( new_n32743_, new_n32726_, new_n32707_ );
and  ( new_n32744_, new_n32743_, new_n32742_ );
or   ( new_n32745_, new_n32744_, new_n32734_ );
and  ( new_n32746_, new_n32745_, new_n32741_ );
and  ( new_n32747_, new_n30600_, new_n30593_ );
or   ( new_n32748_, new_n32747_, new_n30572_ );
and  ( new_n32749_, new_n32748_, new_n30610_ );
and  ( new_n32750_, new_n32749_, new_n32746_ );
or   ( new_n32751_, new_n32750_, new_n32739_ );
and  ( new_n32752_, new_n32751_, new_n32720_ );
or   ( new_n32753_, new_n32749_, new_n32746_ );
or   ( new_n32754_, new_n32744_, new_n32715_ );
or   ( new_n32755_, new_n32740_, new_n32734_ );
and  ( new_n32756_, new_n32755_, new_n32754_ );
and  ( new_n32757_, new_n30603_, new_n30596_ );
or   ( new_n32758_, new_n32757_, new_n30609_ );
and  ( new_n32759_, new_n32758_, new_n30611_ );
or   ( new_n32760_, new_n32759_, new_n32756_ );
and  ( new_n32761_, new_n32760_, new_n32753_ );
and  ( new_n32762_, new_n30624_, new_n30621_ );
or   ( new_n32763_, new_n32762_, new_n32761_ );
and  ( new_n32764_, new_n32763_, new_n30628_ );
and  ( new_n32765_, new_n32764_, new_n32752_ );
and  ( new_n32766_, new_n16102_, RI2b1c4342d7b0_71 );
and  ( new_n32767_, new_n32302_, new_n32235_ );
or   ( new_n32768_, new_n32767_, new_n32244_ );
or   ( new_n32769_, new_n32234_, new_n16186_ );
or   ( new_n32770_, new_n32301_, new_n16204_ );
and  ( new_n32771_, new_n32770_, new_n32769_ );
or   ( new_n32772_, new_n32771_, new_n32305_ );
and  ( new_n32773_, new_n32772_, new_n32768_ );
or   ( new_n32774_, new_n32773_, new_n32766_ );
or   ( new_n32775_, new_n16115_, new_n110_ );
or   ( new_n32776_, new_n32771_, new_n32244_ );
or   ( new_n32777_, new_n32767_, new_n32305_ );
and  ( new_n32778_, new_n32777_, new_n32776_ );
or   ( new_n32779_, new_n32778_, new_n32775_ );
and  ( new_n32780_, new_n32779_, new_n32774_ );
and  ( new_n32781_, new_n32642_, new_n32639_ );
or   ( new_n32782_, new_n32781_, new_n32668_ );
and  ( new_n32783_, new_n32782_, new_n32643_ );
or   ( new_n32784_, new_n32783_, new_n32780_ );
or   ( new_n32785_, new_n32775_, new_n32773_ );
or   ( new_n32786_, new_n32778_, new_n32766_ );
and  ( new_n32787_, new_n32786_, new_n32785_ );
and  ( new_n32788_, new_n32649_, new_n32646_ );
and  ( new_n32789_, new_n32675_, new_n32650_ );
or   ( new_n32790_, new_n32789_, new_n32788_ );
or   ( new_n32791_, new_n32790_, new_n32787_ );
and  ( new_n32792_, new_n32791_, new_n32784_ );
and  ( new_n32793_, new_n32597_, new_n32588_ );
or   ( new_n32794_, new_n32793_, new_n32615_ );
and  ( new_n32795_, new_n32794_, new_n32598_ );
or   ( new_n32796_, new_n32795_, new_n32673_ );
and  ( new_n32797_, new_n32666_, new_n32660_ );
and  ( new_n32798_, new_n32604_, new_n32601_ );
or   ( new_n32799_, new_n32798_, new_n32622_ );
and  ( new_n32800_, new_n32799_, new_n32605_ );
or   ( new_n32801_, new_n32800_, new_n32797_ );
and  ( new_n32802_, new_n32801_, new_n32796_ );
and  ( new_n32803_, new_n16132_, RI2b1c4342d738_70 );
and  ( new_n32804_, new_n16114_, RI2b1c4342d6c0_69 );
or   ( new_n32805_, new_n32804_, new_n32803_ );
or   ( new_n32806_, new_n32805_, new_n16108_ );
or   ( new_n32807_, new_n16119_, new_n755_ );
or   ( new_n32808_, new_n16123_, new_n591_ );
and  ( new_n32809_, new_n32808_, new_n32807_ );
or   ( new_n32810_, new_n32809_, new_n16128_ );
and  ( new_n32811_, new_n32810_, new_n32806_ );
or   ( new_n32812_, new_n32811_, new_n32802_ );
or   ( new_n32813_, new_n32800_, new_n32673_ );
or   ( new_n32814_, new_n32797_, new_n32795_ );
and  ( new_n32815_, new_n32814_, new_n32813_ );
or   ( new_n32816_, new_n32809_, new_n16108_ );
or   ( new_n32817_, new_n32805_, new_n16128_ );
and  ( new_n32818_, new_n32817_, new_n32816_ );
or   ( new_n32819_, new_n32818_, new_n32815_ );
and  ( new_n32820_, new_n32819_, new_n32812_ );
or   ( new_n32821_, new_n32820_, new_n32792_ );
or   ( new_n32822_, new_n32790_, new_n32780_ );
or   ( new_n32823_, new_n32787_, new_n32783_ );
and  ( new_n32824_, new_n32823_, new_n32822_ );
or   ( new_n32825_, new_n32815_, new_n32811_ );
or   ( new_n32826_, new_n32818_, new_n32802_ );
and  ( new_n32827_, new_n32826_, new_n32825_ );
or   ( new_n32828_, new_n32827_, new_n32824_ );
and  ( new_n32829_, new_n32828_, new_n32821_ );
and  ( new_n32830_, new_n32627_, new_n32624_ );
or   ( new_n32831_, new_n32830_, new_n32677_ );
and  ( new_n32832_, new_n32831_, new_n32628_ );
or   ( new_n32833_, new_n32832_, new_n32829_ );
or   ( new_n32834_, new_n32824_, new_n32820_ );
or   ( new_n32835_, new_n32827_, new_n32792_ );
and  ( new_n32836_, new_n32835_, new_n32834_ );
and  ( new_n32837_, new_n32634_, new_n32631_ );
and  ( new_n32838_, new_n32684_, new_n32635_ );
or   ( new_n32839_, new_n32838_, new_n32837_ );
or   ( new_n32840_, new_n32839_, new_n32836_ );
and  ( new_n32841_, new_n32840_, new_n32833_ );
and  ( new_n32842_, new_n32551_, new_n32548_ );
or   ( new_n32843_, new_n32842_, new_n32686_ );
and  ( new_n32844_, new_n32843_, new_n32552_ );
or   ( new_n32845_, new_n32844_, new_n32841_ );
and  ( new_n32846_, new_n32773_, new_n32766_ );
and  ( new_n32847_, new_n32795_, new_n32673_ );
or   ( new_n32848_, new_n32847_, new_n32811_ );
and  ( new_n32849_, new_n32848_, new_n32796_ );
or   ( new_n32850_, new_n32849_, new_n32846_ );
and  ( new_n32851_, new_n32800_, new_n32797_ );
or   ( new_n32852_, new_n32851_, new_n32818_ );
and  ( new_n32853_, new_n32852_, new_n32801_ );
or   ( new_n32854_, new_n32853_, new_n32779_ );
and  ( new_n32855_, new_n32854_, new_n32850_ );
and  ( new_n32856_, new_n32309_, new_n32248_ );
or   ( new_n32857_, new_n32856_, new_n32265_ );
or   ( new_n32858_, new_n32308_, new_n32225_ );
or   ( new_n32859_, new_n32247_, new_n32185_ );
and  ( new_n32860_, new_n32859_, new_n32858_ );
or   ( new_n32861_, new_n32860_, new_n32312_ );
and  ( new_n32862_, new_n32861_, new_n32857_ );
or   ( new_n32863_, new_n32862_, new_n32855_ );
or   ( new_n32864_, new_n32853_, new_n32846_ );
or   ( new_n32865_, new_n32849_, new_n32779_ );
and  ( new_n32866_, new_n32865_, new_n32864_ );
or   ( new_n32867_, new_n32860_, new_n32265_ );
or   ( new_n32868_, new_n32856_, new_n32312_ );
and  ( new_n32869_, new_n32868_, new_n32867_ );
or   ( new_n32870_, new_n32869_, new_n32866_ );
and  ( new_n32871_, new_n32870_, new_n32863_ );
and  ( new_n32872_, new_n32783_, new_n32780_ );
or   ( new_n32873_, new_n32872_, new_n32820_ );
and  ( new_n32874_, new_n32873_, new_n32784_ );
or   ( new_n32875_, new_n32874_, new_n32871_ );
or   ( new_n32876_, new_n32866_, new_n32862_ );
or   ( new_n32877_, new_n32869_, new_n32855_ );
and  ( new_n32878_, new_n32877_, new_n32876_ );
and  ( new_n32879_, new_n32790_, new_n32787_ );
and  ( new_n32880_, new_n32827_, new_n32791_ );
or   ( new_n32881_, new_n32880_, new_n32879_ );
or   ( new_n32882_, new_n32881_, new_n32878_ );
and  ( new_n32883_, new_n32882_, new_n32875_ );
and  ( new_n32884_, new_n32832_, new_n32829_ );
or   ( new_n32885_, new_n32884_, new_n32883_ );
and  ( new_n32886_, new_n32885_, new_n32845_ );
and  ( new_n32887_, new_n32316_, new_n32269_ );
or   ( new_n32888_, new_n32887_, new_n32281_ );
or   ( new_n32889_, new_n32315_, new_n32224_ );
or   ( new_n32890_, new_n32298_, new_n32268_ );
and  ( new_n32891_, new_n32890_, new_n32889_ );
or   ( new_n32892_, new_n32891_, new_n32319_ );
and  ( new_n32893_, new_n32892_, new_n32888_ );
and  ( new_n32894_, new_n32849_, new_n32846_ );
or   ( new_n32895_, new_n32894_, new_n32862_ );
and  ( new_n32896_, new_n32895_, new_n32850_ );
or   ( new_n32897_, new_n32896_, new_n32893_ );
or   ( new_n32898_, new_n32891_, new_n32281_ );
or   ( new_n32899_, new_n32887_, new_n32319_ );
and  ( new_n32900_, new_n32899_, new_n32898_ );
and  ( new_n32901_, new_n32853_, new_n32779_ );
and  ( new_n32902_, new_n32869_, new_n32854_ );
or   ( new_n32903_, new_n32902_, new_n32901_ );
or   ( new_n32904_, new_n32903_, new_n32900_ );
and  ( new_n32905_, new_n32904_, new_n32897_ );
and  ( new_n32906_, new_n32874_, new_n32871_ );
or   ( new_n32907_, new_n32906_, new_n32905_ );
and  ( new_n32908_, new_n32326_, new_n32285_ );
or   ( new_n32909_, new_n32908_, new_n32288_ );
or   ( new_n32910_, new_n32322_, new_n32217_ );
or   ( new_n32911_, new_n32325_, new_n32284_ );
and  ( new_n32912_, new_n32911_, new_n32910_ );
or   ( new_n32913_, new_n32912_, new_n32328_ );
and  ( new_n32914_, new_n32913_, new_n32909_ );
and  ( new_n32915_, new_n32896_, new_n32893_ );
or   ( new_n32916_, new_n32915_, new_n32914_ );
and  ( new_n32917_, new_n32916_, new_n32907_ );
and  ( new_n32918_, new_n32917_, new_n32886_ );
and  ( new_n32919_, new_n32918_, new_n32765_ );
and  ( new_n32920_, new_n32919_, new_n31122_ );
and  ( new_n32921_, new_n32750_, new_n32739_ );
and  ( new_n32922_, new_n32719_, new_n32695_ );
or   ( new_n32923_, new_n32922_, new_n32921_ );
and  ( new_n32924_, new_n32923_, new_n32720_ );
and  ( new_n32925_, new_n32762_, new_n32761_ );
or   ( new_n32926_, new_n32925_, new_n30636_ );
and  ( new_n32927_, new_n32926_, new_n32763_ );
and  ( new_n32928_, new_n32927_, new_n32752_ );
or   ( new_n32929_, new_n32928_, new_n32924_ );
and  ( new_n32930_, new_n32929_, new_n32918_ );
and  ( new_n32931_, new_n32906_, new_n32905_ );
and  ( new_n32932_, new_n32915_, new_n32914_ );
or   ( new_n32933_, new_n32932_, new_n32931_ );
and  ( new_n32934_, new_n32933_, new_n32916_ );
and  ( new_n32935_, new_n32844_, new_n32841_ );
and  ( new_n32936_, new_n32884_, new_n32883_ );
or   ( new_n32937_, new_n32936_, new_n32935_ );
and  ( new_n32938_, new_n32937_, new_n32885_ );
and  ( new_n32939_, new_n32938_, new_n32917_ );
or   ( new_n32940_, new_n32939_, new_n32934_ );
or   ( new_n32941_, new_n32940_, new_n32930_ );
or   ( new_n32942_, new_n32941_, new_n32920_ );
or   ( new_n32943_, new_n32942_, new_n32333_ );
or   ( new_n32944_, new_n32291_, new_n32184_ );
or   ( new_n32945_, new_n32331_, new_n32295_ );
and  ( new_n32946_, new_n32945_, new_n32944_ );
or   ( new_n32947_, new_n32690_, new_n32686_ );
or   ( new_n32948_, new_n32693_, new_n32583_ );
and  ( new_n32949_, new_n32948_, new_n32947_ );
and  ( new_n32950_, new_n32949_, new_n32737_ );
or   ( new_n32951_, new_n32736_, new_n32702_ );
or   ( new_n32952_, new_n32723_, new_n32718_ );
and  ( new_n32953_, new_n32952_, new_n32951_ );
and  ( new_n32954_, new_n32953_, new_n32760_ );
or   ( new_n32955_, new_n32954_, new_n32950_ );
or   ( new_n32956_, new_n32759_, new_n32746_ );
or   ( new_n32957_, new_n32756_, new_n32749_ );
and  ( new_n32958_, new_n32957_, new_n32956_ );
and  ( new_n32959_, new_n32958_, new_n30618_ );
or   ( new_n32960_, new_n32959_, new_n30637_ );
or   ( new_n32961_, new_n32960_, new_n32955_ );
or   ( new_n32962_, new_n32839_, new_n32829_ );
or   ( new_n32963_, new_n32836_, new_n32832_ );
and  ( new_n32964_, new_n32963_, new_n32962_ );
and  ( new_n32965_, new_n32581_, new_n32555_ );
or   ( new_n32966_, new_n32965_, new_n32693_ );
and  ( new_n32967_, new_n32966_, new_n32582_ );
and  ( new_n32968_, new_n32967_, new_n32964_ );
or   ( new_n32969_, new_n32881_, new_n32871_ );
or   ( new_n32970_, new_n32878_, new_n32874_ );
and  ( new_n32971_, new_n32970_, new_n32969_ );
and  ( new_n32972_, new_n32971_, new_n32840_ );
or   ( new_n32973_, new_n32972_, new_n32968_ );
or   ( new_n32974_, new_n32903_, new_n32893_ );
or   ( new_n32975_, new_n32900_, new_n32896_ );
and  ( new_n32976_, new_n32975_, new_n32974_ );
and  ( new_n32977_, new_n32976_, new_n32882_ );
or   ( new_n32978_, new_n32912_, new_n32288_ );
or   ( new_n32979_, new_n32908_, new_n32328_ );
and  ( new_n32980_, new_n32979_, new_n32978_ );
and  ( new_n32981_, new_n32980_, new_n32904_ );
or   ( new_n32982_, new_n32981_, new_n32977_ );
or   ( new_n32983_, new_n32982_, new_n32973_ );
or   ( new_n32984_, new_n32983_, new_n32961_ );
or   ( new_n32985_, new_n32984_, new_n30453_ );
or   ( new_n32986_, new_n32949_, new_n32737_ );
or   ( new_n32987_, new_n32953_, new_n32760_ );
or   ( new_n32988_, new_n32987_, new_n32950_ );
and  ( new_n32989_, new_n32988_, new_n32986_ );
or   ( new_n32990_, new_n32958_, new_n30618_ );
or   ( new_n32991_, new_n32959_, new_n30633_ );
and  ( new_n32992_, new_n32991_, new_n32990_ );
or   ( new_n32993_, new_n32992_, new_n32955_ );
and  ( new_n32994_, new_n32993_, new_n32989_ );
or   ( new_n32995_, new_n32994_, new_n32983_ );
or   ( new_n32996_, new_n32980_, new_n32904_ );
or   ( new_n32997_, new_n32976_, new_n32882_ );
or   ( new_n32998_, new_n32997_, new_n32981_ );
and  ( new_n32999_, new_n32998_, new_n32996_ );
or   ( new_n33000_, new_n32971_, new_n32840_ );
or   ( new_n33001_, new_n32967_, new_n32964_ );
or   ( new_n33002_, new_n33001_, new_n32972_ );
and  ( new_n33003_, new_n33002_, new_n33000_ );
or   ( new_n33004_, new_n33003_, new_n32982_ );
and  ( new_n33005_, new_n33004_, new_n32999_ );
and  ( new_n33006_, new_n33005_, new_n32995_ );
and  ( new_n33007_, new_n33006_, new_n32985_ );
or   ( new_n33008_, new_n33007_, new_n32946_ );
and  ( new_n33009_, new_n33008_, new_n32943_ );
and  ( new_n33010_, new_n33009_, new_n32075_ );
or   ( new_n33011_, new_n33010_, new_n31125_ );
and  ( new_n33012_, new_n32004_, new_n32000_ );
and  ( new_n33013_, new_n32073_, new_n31383_ );
or   ( new_n33014_, new_n33013_, new_n33012_ );
or   ( new_n33015_, new_n32946_, new_n32942_ );
or   ( new_n33016_, new_n33007_, new_n32333_ );
and  ( new_n33017_, new_n33016_, new_n33015_ );
and  ( new_n33018_, new_n33017_, new_n33014_ );
and  ( new_n33019_, new_n6464_, new_n5987_ );
or   ( new_n33020_, new_n33019_, new_n5992_ );
or   ( new_n33021_, new_n6463_, new_n5992_ );
and  ( new_n33022_, new_n7407_, new_n6903_ );
or   ( new_n33023_, new_n33022_, new_n6906_ );
or   ( new_n33024_, new_n33023_, new_n33021_ );
and  ( new_n33025_, new_n33024_, new_n33020_ );
or   ( new_n33026_, new_n7406_, new_n6906_ );
or   ( new_n33027_, new_n33026_, new_n33021_ );
or   ( new_n33028_, new_n15318_, new_n8293_ );
or   ( new_n33029_, new_n9205_, new_n8766_ );
or   ( new_n33030_, new_n33029_, new_n33028_ );
and  ( new_n33031_, new_n9999_, new_n9585_ );
or   ( new_n33032_, new_n33031_, new_n9590_ );
or   ( new_n33033_, new_n9998_, new_n9590_ );
and  ( new_n33034_, new_n10786_, new_n10379_ );
or   ( new_n33035_, new_n33034_, new_n10382_ );
or   ( new_n33036_, new_n33035_, new_n33033_ );
and  ( new_n33037_, new_n33036_, new_n33032_ );
or   ( new_n33038_, new_n10785_, new_n10382_ );
or   ( new_n33039_, new_n33038_, new_n33033_ );
and  ( new_n33040_, new_n11530_, new_n11166_ );
or   ( new_n33041_, new_n33040_, new_n11173_ );
or   ( new_n33042_, new_n11529_, new_n11173_ );
and  ( new_n33043_, new_n11858_, new_n11660_ );
or   ( new_n33044_, new_n33043_, new_n11663_ );
or   ( new_n33045_, new_n33044_, new_n33042_ );
and  ( new_n33046_, new_n33045_, new_n33041_ );
or   ( new_n33047_, new_n11857_, new_n11663_ );
or   ( new_n33048_, new_n33047_, new_n33042_ );
or   ( new_n33049_, new_n12466_, new_n12180_ );
or   ( new_n33050_, new_n12985_, new_n12732_ );
or   ( new_n33051_, new_n33050_, new_n33049_ );
or   ( new_n33052_, new_n13509_, new_n13259_ );
or   ( new_n33053_, new_n13959_, new_n13740_ );
or   ( new_n33054_, new_n33053_, new_n33052_ );
or   ( new_n33055_, new_n14119_, new_n13948_ );
or   ( new_n33056_, new_n14605_, new_n14309_ );
or   ( new_n33057_, new_n14744_, new_n14587_ );
or   ( new_n33058_, new_n14979_, new_n14810_ );
or   ( new_n33059_, new_n15026_, new_n14966_ );
or   ( new_n33060_, new_n15254_, new_n15207_ );
and  ( new_n33061_, new_n15208_, new_n15174_ );
or   ( new_n33062_, new_n33061_, new_n15177_ );
and  ( new_n33063_, new_n33062_, new_n33060_ );
or   ( new_n33064_, new_n33063_, new_n15143_ );
or   ( new_n33065_, new_n33064_, new_n15084_ );
or   ( new_n33066_, new_n33065_, new_n33059_ );
and  ( new_n33067_, new_n15268_, new_n15027_ );
or   ( new_n33068_, new_n33067_, new_n14966_ );
and  ( new_n33069_, new_n15144_, new_n15081_ );
or   ( new_n33070_, new_n33069_, new_n15084_ );
or   ( new_n33071_, new_n33070_, new_n33059_ );
and  ( new_n33072_, new_n33071_, new_n33068_ );
and  ( new_n33073_, new_n33072_, new_n33066_ );
or   ( new_n33074_, new_n33073_, new_n33058_ );
or   ( new_n33075_, new_n33074_, new_n33057_ );
and  ( new_n33076_, new_n15281_, new_n15263_ );
or   ( new_n33077_, new_n33076_, new_n14587_ );
and  ( new_n33078_, new_n15267_, new_n15264_ );
or   ( new_n33079_, new_n33078_, new_n14810_ );
or   ( new_n33080_, new_n33079_, new_n33057_ );
and  ( new_n33081_, new_n33080_, new_n33077_ );
and  ( new_n33082_, new_n33081_, new_n33075_ );
or   ( new_n33083_, new_n33082_, new_n33056_ );
or   ( new_n33084_, new_n33083_, new_n33055_ );
and  ( new_n33085_, new_n15294_, new_n15276_ );
or   ( new_n33086_, new_n33085_, new_n13948_ );
and  ( new_n33087_, new_n15280_, new_n15277_ );
or   ( new_n33088_, new_n33087_, new_n14309_ );
or   ( new_n33089_, new_n33088_, new_n33055_ );
and  ( new_n33090_, new_n33089_, new_n33086_ );
and  ( new_n33091_, new_n33090_, new_n33084_ );
or   ( new_n33092_, new_n33091_, new_n33054_ );
or   ( new_n33093_, new_n33092_, new_n33051_ );
and  ( new_n33094_, new_n15302_, new_n12175_ );
or   ( new_n33095_, new_n33094_, new_n12180_ );
and  ( new_n33096_, new_n15306_, new_n15303_ );
or   ( new_n33097_, new_n33096_, new_n12732_ );
or   ( new_n33098_, new_n33097_, new_n33049_ );
and  ( new_n33099_, new_n33098_, new_n33095_ );
and  ( new_n33100_, new_n15307_, new_n15289_ );
or   ( new_n33101_, new_n33100_, new_n13259_ );
and  ( new_n33102_, new_n15293_, new_n15290_ );
or   ( new_n33103_, new_n33102_, new_n13740_ );
or   ( new_n33104_, new_n33103_, new_n33052_ );
and  ( new_n33105_, new_n33104_, new_n33101_ );
or   ( new_n33106_, new_n33105_, new_n33051_ );
and  ( new_n33107_, new_n33106_, new_n33099_ );
and  ( new_n33108_, new_n33107_, new_n33093_ );
or   ( new_n33109_, new_n33108_, new_n33048_ );
and  ( new_n33110_, new_n33109_, new_n33046_ );
or   ( new_n33111_, new_n33110_, new_n33039_ );
and  ( new_n33112_, new_n33111_, new_n33037_ );
or   ( new_n33113_, new_n33112_, new_n33030_ );
or   ( new_n33114_, new_n33113_, new_n33027_ );
and  ( new_n33115_, new_n8294_, new_n7854_ );
or   ( new_n33116_, new_n33115_, new_n15318_ );
and  ( new_n33117_, new_n9206_, new_n8763_ );
or   ( new_n33118_, new_n33117_, new_n8766_ );
or   ( new_n33119_, new_n33118_, new_n33028_ );
and  ( new_n33120_, new_n33119_, new_n33116_ );
or   ( new_n33121_, new_n33120_, new_n33027_ );
and  ( new_n33122_, new_n33121_, new_n33114_ );
and  ( new_n33123_, new_n33122_, new_n33025_ );
or   ( new_n33124_, new_n4374_, new_n3316_ );
or   ( new_n33125_, new_n4370_, new_n4014_ );
or   ( new_n33126_, new_n33125_, new_n33124_ );
or   ( new_n33127_, new_n4762_, new_n4379_ );
or   ( new_n33128_, new_n5576_, new_n5151_ );
or   ( new_n33129_, new_n33128_, new_n33127_ );
or   ( new_n33130_, new_n33129_, new_n33126_ );
or   ( new_n33131_, new_n33130_, new_n33123_ );
or   ( new_n33132_, new_n31815_, new_n31544_ );
or   ( new_n33133_, new_n31897_, new_n31804_ );
or   ( new_n33134_, new_n33133_, new_n33132_ );
or   ( new_n33135_, new_n2635_, new_n2309_ );
or   ( new_n33136_, new_n15507_, new_n1798_ );
or   ( new_n33137_, new_n33136_, new_n33135_ );
or   ( new_n33138_, new_n33137_, new_n33134_ );
or   ( new_n33139_, new_n33138_, new_n33131_ );
and  ( new_n33140_, new_n3317_, new_n2968_ );
or   ( new_n33141_, new_n33140_, new_n4374_ );
and  ( new_n33142_, new_n4015_, new_n3658_ );
or   ( new_n33143_, new_n33142_, new_n4370_ );
or   ( new_n33144_, new_n33143_, new_n33124_ );
and  ( new_n33145_, new_n33144_, new_n33141_ );
and  ( new_n33146_, new_n4763_, new_n4367_ );
or   ( new_n33147_, new_n33146_, new_n4379_ );
and  ( new_n33148_, new_n5577_, new_n5148_ );
or   ( new_n33149_, new_n33148_, new_n5151_ );
or   ( new_n33150_, new_n33149_, new_n33127_ );
and  ( new_n33151_, new_n33150_, new_n33147_ );
or   ( new_n33152_, new_n33151_, new_n33126_ );
and  ( new_n33153_, new_n33152_, new_n33145_ );
or   ( new_n33154_, new_n33153_, new_n33138_ );
and  ( new_n33155_, new_n31991_, new_n31978_ );
or   ( new_n33156_, new_n33155_, new_n31897_ );
and  ( new_n33157_, new_n31981_, new_n31977_ );
or   ( new_n33158_, new_n33157_, new_n31815_ );
or   ( new_n33159_, new_n33158_, new_n33133_ );
and  ( new_n33160_, new_n33159_, new_n33156_ );
and  ( new_n33161_, new_n15500_, new_n2306_ );
or   ( new_n33162_, new_n33161_, new_n15507_ );
and  ( new_n33163_, new_n2636_, new_n2305_ );
or   ( new_n33164_, new_n33163_, new_n2309_ );
or   ( new_n33165_, new_n33164_, new_n33136_ );
and  ( new_n33166_, new_n33165_, new_n33162_ );
or   ( new_n33167_, new_n33166_, new_n33134_ );
and  ( new_n33168_, new_n33167_, new_n33160_ );
and  ( new_n33169_, new_n33168_, new_n33154_ );
and  ( new_n33170_, new_n33169_, new_n33139_ );
or   ( new_n33171_, new_n32064_, new_n31937_ );
and  ( new_n33172_, new_n33171_, new_n33170_ );
and  ( new_n33173_, new_n32032_, new_n31992_ );
and  ( new_n33174_, new_n15615_, new_n15606_ );
and  ( new_n33175_, new_n15635_, new_n15626_ );
or   ( new_n33176_, new_n33175_, new_n15623_ );
and  ( new_n33177_, new_n33176_, new_n33174_ );
and  ( new_n33178_, new_n15616_, new_n15606_ );
or   ( new_n33179_, new_n33178_, new_n15601_ );
or   ( new_n33180_, new_n33179_, new_n33177_ );
and  ( new_n33181_, new_n15634_, new_n15626_ );
and  ( new_n33182_, new_n33181_, new_n33174_ );
and  ( new_n33183_, new_n15991_, new_n15655_ );
and  ( new_n33184_, new_n15674_, new_n15666_ );
and  ( new_n33185_, new_n33184_, new_n33183_ );
and  ( new_n33186_, new_n15696_, new_n15687_ );
and  ( new_n33187_, new_n15716_, new_n15707_ );
or   ( new_n33188_, new_n33187_, new_n15704_ );
and  ( new_n33189_, new_n33188_, new_n33186_ );
and  ( new_n33190_, new_n15697_, new_n15687_ );
or   ( new_n33191_, new_n33190_, new_n15682_ );
or   ( new_n33192_, new_n33191_, new_n33189_ );
and  ( new_n33193_, new_n15715_, new_n15707_ );
and  ( new_n33194_, new_n33193_, new_n33186_ );
and  ( new_n33195_, new_n15737_, new_n15730_ );
and  ( new_n33196_, new_n15752_, new_n15744_ );
or   ( new_n33197_, new_n33196_, new_n15741_ );
and  ( new_n33198_, new_n33197_, new_n33195_ );
and  ( new_n33199_, new_n15736_, new_n15730_ );
or   ( new_n33200_, new_n33199_, new_n15723_ );
or   ( new_n33201_, new_n33200_, new_n33198_ );
and  ( new_n33202_, new_n15753_, new_n15744_ );
and  ( new_n33203_, new_n33202_, new_n33195_ );
and  ( new_n33204_, new_n15774_, new_n15765_ );
and  ( new_n33205_, new_n15789_, new_n15781_ );
and  ( new_n33206_, new_n33205_, new_n33204_ );
and  ( new_n33207_, new_n15804_, new_n15796_ );
and  ( new_n33208_, new_n15820_, new_n15808_ );
and  ( new_n33209_, new_n33208_, new_n33207_ );
and  ( new_n33210_, new_n15828_, new_n15816_ );
and  ( new_n33211_, new_n15847_, new_n15835_ );
and  ( new_n33212_, new_n15852_, new_n15840_ );
and  ( new_n33213_, new_n15868_, new_n15856_ );
and  ( new_n33214_, new_n15874_, new_n15861_ );
and  ( new_n33215_, new_n15897_, new_n15893_ );
or   ( new_n33216_, new_n33215_, new_n15928_ );
and  ( new_n33217_, new_n15898_, new_n15893_ );
and  ( new_n33218_, new_n33217_, new_n15922_ );
or   ( new_n33219_, new_n33218_, new_n33216_ );
and  ( new_n33220_, new_n15889_, new_n15884_ );
and  ( new_n33221_, new_n33220_, new_n33219_ );
and  ( new_n33222_, new_n33221_, new_n33214_ );
and  ( new_n33223_, new_n15927_, new_n15884_ );
or   ( new_n33224_, new_n33223_, new_n15881_ );
and  ( new_n33225_, new_n33224_, new_n33214_ );
and  ( new_n33226_, new_n15873_, new_n15861_ );
or   ( new_n33227_, new_n33226_, new_n15941_ );
or   ( new_n33228_, new_n33227_, new_n33225_ );
or   ( new_n33229_, new_n33228_, new_n33222_ );
and  ( new_n33230_, new_n33229_, new_n33213_ );
and  ( new_n33231_, new_n33230_, new_n33212_ );
and  ( new_n33232_, new_n15940_, new_n15856_ );
or   ( new_n33233_, new_n33232_, new_n15937_ );
and  ( new_n33234_, new_n33233_, new_n33212_ );
and  ( new_n33235_, new_n15936_, new_n15840_ );
or   ( new_n33236_, new_n33235_, new_n15954_ );
or   ( new_n33237_, new_n33236_, new_n33234_ );
or   ( new_n33238_, new_n33237_, new_n33231_ );
and  ( new_n33239_, new_n33238_, new_n33211_ );
and  ( new_n33240_, new_n33239_, new_n33210_ );
and  ( new_n33241_, new_n15953_, new_n15835_ );
or   ( new_n33242_, new_n33241_, new_n15950_ );
and  ( new_n33243_, new_n33242_, new_n33210_ );
and  ( new_n33244_, new_n15949_, new_n15816_ );
or   ( new_n33245_, new_n33244_, new_n15967_ );
or   ( new_n33246_, new_n33245_, new_n33243_ );
or   ( new_n33247_, new_n33246_, new_n33240_ );
and  ( new_n33248_, new_n33247_, new_n33209_ );
and  ( new_n33249_, new_n33248_, new_n33206_ );
or   ( new_n33250_, new_n15975_, new_n15760_ );
and  ( new_n33251_, new_n33250_, new_n15765_ );
or   ( new_n33252_, new_n15979_, new_n15976_ );
and  ( new_n33253_, new_n33252_, new_n15781_ );
and  ( new_n33254_, new_n33253_, new_n33204_ );
or   ( new_n33255_, new_n33254_, new_n33251_ );
or   ( new_n33256_, new_n15980_, new_n15962_ );
and  ( new_n33257_, new_n33256_, new_n15796_ );
and  ( new_n33258_, new_n15966_, new_n15808_ );
or   ( new_n33259_, new_n33258_, new_n15963_ );
and  ( new_n33260_, new_n33259_, new_n33207_ );
or   ( new_n33261_, new_n33260_, new_n33257_ );
and  ( new_n33262_, new_n33261_, new_n33206_ );
or   ( new_n33263_, new_n33262_, new_n33255_ );
or   ( new_n33264_, new_n33263_, new_n33249_ );
and  ( new_n33265_, new_n33264_, new_n33203_ );
or   ( new_n33266_, new_n33265_, new_n33201_ );
and  ( new_n33267_, new_n33266_, new_n33194_ );
or   ( new_n33268_, new_n33267_, new_n33192_ );
and  ( new_n33269_, new_n33268_, new_n33185_ );
and  ( new_n33270_, new_n33269_, new_n33182_ );
and  ( new_n33271_, new_n15675_, new_n15666_ );
or   ( new_n33272_, new_n33271_, new_n15663_ );
and  ( new_n33273_, new_n33272_, new_n33183_ );
and  ( new_n33274_, new_n15991_, new_n15656_ );
or   ( new_n33275_, new_n33274_, new_n15642_ );
or   ( new_n33276_, new_n33275_, new_n33273_ );
and  ( new_n33277_, new_n33276_, new_n33182_ );
or   ( new_n33278_, new_n33277_, new_n33270_ );
or   ( new_n33279_, new_n33278_, new_n33180_ );
and  ( new_n33280_, new_n15565_, new_n15543_ );
and  ( new_n33281_, new_n15561_, new_n15554_ );
and  ( new_n33282_, new_n33281_, new_n33280_ );
and  ( new_n33283_, new_n15578_, new_n15570_ );
and  ( new_n33284_, new_n15594_, new_n15588_ );
and  ( new_n33285_, new_n33284_, new_n33283_ );
and  ( new_n33286_, new_n33285_, new_n33282_ );
and  ( new_n33287_, new_n33286_, new_n33279_ );
and  ( new_n33288_, new_n15530_, new_n15524_ );
and  ( new_n33289_, new_n15514_, new_n15504_ );
and  ( new_n33290_, new_n33289_, new_n33288_ );
and  ( new_n33291_, new_n32019_, new_n32010_ );
and  ( new_n33292_, new_n32028_, new_n32015_ );
and  ( new_n33293_, new_n33292_, new_n33291_ );
and  ( new_n33294_, new_n33293_, new_n33290_ );
and  ( new_n33295_, new_n33294_, new_n33287_ );
and  ( new_n33296_, new_n15561_, new_n15553_ );
or   ( new_n33297_, new_n33296_, new_n15547_ );
and  ( new_n33298_, new_n33297_, new_n33280_ );
and  ( new_n33299_, new_n15565_, new_n15542_ );
or   ( new_n33300_, new_n33299_, new_n15534_ );
or   ( new_n33301_, new_n33300_, new_n33298_ );
or   ( new_n33302_, new_n15593_, new_n15585_ );
and  ( new_n33303_, new_n33302_, new_n15588_ );
and  ( new_n33304_, new_n33303_, new_n33283_ );
and  ( new_n33305_, new_n15577_, new_n15570_ );
or   ( new_n33306_, new_n33305_, new_n15558_ );
or   ( new_n33307_, new_n33306_, new_n33304_ );
and  ( new_n33308_, new_n33307_, new_n33282_ );
or   ( new_n33309_, new_n33308_, new_n33301_ );
and  ( new_n33310_, new_n33309_, new_n33294_ );
and  ( new_n33311_, new_n32054_, new_n32019_ );
or   ( new_n33312_, new_n33311_, new_n32051_ );
and  ( new_n33313_, new_n33312_, new_n33292_ );
and  ( new_n33314_, new_n32050_, new_n32028_ );
or   ( new_n33315_, new_n33314_, new_n32065_ );
or   ( new_n33316_, new_n33315_, new_n33313_ );
and  ( new_n33317_, new_n15529_, new_n15524_ );
or   ( new_n33318_, new_n33317_, new_n15521_ );
and  ( new_n33319_, new_n33318_, new_n33289_ );
and  ( new_n33320_, new_n15513_, new_n15504_ );
or   ( new_n33321_, new_n33320_, new_n15508_ );
or   ( new_n33322_, new_n33321_, new_n33319_ );
and  ( new_n33323_, new_n33322_, new_n33293_ );
or   ( new_n33324_, new_n33323_, new_n33316_ );
or   ( new_n33325_, new_n33324_, new_n33310_ );
or   ( new_n33326_, new_n33325_, new_n33295_ );
and  ( new_n33327_, new_n33326_, new_n33173_ );
or   ( new_n33328_, new_n33327_, new_n33172_ );
or   ( new_n33329_, new_n32972_, new_n32936_ );
or   ( new_n33330_, new_n21656_, new_n21194_ );
or   ( new_n33331_, new_n22564_, new_n22101_ );
and  ( new_n33332_, new_n33331_, new_n22098_ );
or   ( new_n33333_, new_n33332_, new_n33330_ );
or   ( new_n33334_, new_n21657_, new_n21194_ );
and  ( new_n33335_, new_n33334_, new_n21189_ );
and  ( new_n33336_, new_n33335_, new_n33333_ );
or   ( new_n33337_, new_n22563_, new_n22101_ );
or   ( new_n33338_, new_n33337_, new_n33330_ );
or   ( new_n33339_, new_n23451_, new_n23017_ );
or   ( new_n33340_, new_n24360_, new_n23923_ );
or   ( new_n33341_, new_n33340_, new_n33339_ );
or   ( new_n33342_, new_n25151_, new_n24745_ );
or   ( new_n33343_, new_n25937_, new_n25536_ );
and  ( new_n33344_, new_n33343_, new_n25533_ );
or   ( new_n33345_, new_n33344_, new_n33342_ );
or   ( new_n33346_, new_n25152_, new_n24745_ );
and  ( new_n33347_, new_n33346_, new_n24740_ );
and  ( new_n33348_, new_n33347_, new_n33345_ );
or   ( new_n33349_, new_n25936_, new_n25536_ );
or   ( new_n33350_, new_n33349_, new_n33342_ );
or   ( new_n33351_, new_n26678_, new_n26324_ );
or   ( new_n33352_, new_n27006_, new_n26811_ );
and  ( new_n33353_, new_n33352_, new_n26808_ );
or   ( new_n33354_, new_n33353_, new_n33351_ );
or   ( new_n33355_, new_n26677_, new_n26324_ );
and  ( new_n33356_, new_n33355_, new_n26318_ );
and  ( new_n33357_, new_n33356_, new_n33354_ );
or   ( new_n33358_, new_n27007_, new_n26811_ );
or   ( new_n33359_, new_n33358_, new_n33351_ );
or   ( new_n33360_, new_n27611_, new_n27327_ );
or   ( new_n33361_, new_n28130_, new_n27876_ );
or   ( new_n33362_, new_n33361_, new_n33360_ );
or   ( new_n33363_, new_n28651_, new_n28401_ );
or   ( new_n33364_, new_n29099_, new_n28881_ );
or   ( new_n33365_, new_n33364_, new_n33363_ );
or   ( new_n33366_, new_n29258_, new_n29088_ );
or   ( new_n33367_, new_n29740_, new_n29446_ );
or   ( new_n33368_, new_n29878_, new_n29721_ );
or   ( new_n33369_, new_n30111_, new_n29944_ );
or   ( new_n33370_, new_n30159_, new_n30098_ );
or   ( new_n33371_, new_n30378_, new_n30327_ );
or   ( new_n33372_, new_n33371_, new_n30316_ );
or   ( new_n33373_, new_n33371_, new_n30325_ );
or   ( new_n33374_, new_n30378_, new_n30282_ );
and  ( new_n33375_, new_n33374_, new_n30382_ );
and  ( new_n33376_, new_n33375_, new_n33373_ );
and  ( new_n33377_, new_n33376_, new_n33372_ );
or   ( new_n33378_, new_n30367_, new_n30216_ );
or   ( new_n33379_, new_n33378_, new_n33377_ );
or   ( new_n33380_, new_n33379_, new_n33370_ );
or   ( new_n33381_, new_n30381_, new_n30216_ );
and  ( new_n33382_, new_n33381_, new_n30213_ );
or   ( new_n33383_, new_n33382_, new_n33370_ );
or   ( new_n33384_, new_n30158_, new_n30098_ );
and  ( new_n33385_, new_n33384_, new_n30395_ );
and  ( new_n33386_, new_n33385_, new_n33383_ );
and  ( new_n33387_, new_n33386_, new_n33380_ );
or   ( new_n33388_, new_n33387_, new_n33369_ );
or   ( new_n33389_, new_n33388_, new_n33368_ );
or   ( new_n33390_, new_n30394_, new_n29944_ );
and  ( new_n33391_, new_n33390_, new_n30391_ );
or   ( new_n33392_, new_n33391_, new_n33368_ );
or   ( new_n33393_, new_n30390_, new_n29721_ );
and  ( new_n33394_, new_n33393_, new_n30408_ );
and  ( new_n33395_, new_n33394_, new_n33392_ );
and  ( new_n33396_, new_n33395_, new_n33389_ );
or   ( new_n33397_, new_n33396_, new_n33367_ );
or   ( new_n33398_, new_n33397_, new_n33366_ );
or   ( new_n33399_, new_n30407_, new_n29446_ );
and  ( new_n33400_, new_n33399_, new_n30404_ );
or   ( new_n33401_, new_n33400_, new_n33366_ );
or   ( new_n33402_, new_n30403_, new_n29088_ );
and  ( new_n33403_, new_n33402_, new_n30421_ );
and  ( new_n33404_, new_n33403_, new_n33401_ );
and  ( new_n33405_, new_n33404_, new_n33398_ );
or   ( new_n33406_, new_n33405_, new_n33365_ );
or   ( new_n33407_, new_n33406_, new_n33362_ );
and  ( new_n33408_, new_n30429_, new_n27322_ );
or   ( new_n33409_, new_n33408_, new_n27327_ );
and  ( new_n33410_, new_n30433_, new_n30430_ );
or   ( new_n33411_, new_n33410_, new_n27876_ );
or   ( new_n33412_, new_n33411_, new_n33360_ );
and  ( new_n33413_, new_n33412_, new_n33409_ );
and  ( new_n33414_, new_n30434_, new_n30416_ );
or   ( new_n33415_, new_n33414_, new_n28401_ );
or   ( new_n33416_, new_n30420_, new_n28881_ );
and  ( new_n33417_, new_n33416_, new_n30417_ );
or   ( new_n33418_, new_n33417_, new_n33363_ );
and  ( new_n33419_, new_n33418_, new_n33415_ );
or   ( new_n33420_, new_n33419_, new_n33362_ );
and  ( new_n33421_, new_n33420_, new_n33413_ );
and  ( new_n33422_, new_n33421_, new_n33407_ );
or   ( new_n33423_, new_n33422_, new_n33359_ );
and  ( new_n33424_, new_n33423_, new_n33357_ );
or   ( new_n33425_, new_n33424_, new_n33350_ );
and  ( new_n33426_, new_n33425_, new_n33348_ );
or   ( new_n33427_, new_n33426_, new_n33341_ );
or   ( new_n33428_, new_n33427_, new_n33338_ );
or   ( new_n33429_, new_n24361_, new_n23923_ );
and  ( new_n33430_, new_n33429_, new_n23920_ );
or   ( new_n33431_, new_n33430_, new_n33339_ );
or   ( new_n33432_, new_n23452_, new_n23017_ );
and  ( new_n33433_, new_n33432_, new_n23012_ );
and  ( new_n33434_, new_n33433_, new_n33431_ );
or   ( new_n33435_, new_n33434_, new_n33338_ );
and  ( new_n33436_, new_n33435_, new_n33428_ );
and  ( new_n33437_, new_n33436_, new_n33336_ );
or   ( new_n33438_, new_n18589_, new_n18247_ );
or   ( new_n33439_, new_n19614_, new_n19268_ );
or   ( new_n33440_, new_n33439_, new_n33438_ );
or   ( new_n33441_, new_n19995_, new_n19618_ );
or   ( new_n33442_, new_n20793_, new_n20373_ );
or   ( new_n33443_, new_n33442_, new_n33441_ );
or   ( new_n33444_, new_n33443_, new_n33440_ );
or   ( new_n33445_, new_n33444_, new_n33437_ );
or   ( new_n33446_, new_n32959_, new_n32954_ );
or   ( new_n33447_, new_n32968_, new_n32950_ );
or   ( new_n33448_, new_n33447_, new_n33446_ );
or   ( new_n33449_, new_n30637_, new_n17109_ );
or   ( new_n33450_, new_n17923_, new_n17601_ );
or   ( new_n33451_, new_n33450_, new_n33449_ );
or   ( new_n33452_, new_n33451_, new_n33448_ );
or   ( new_n33453_, new_n33452_, new_n33445_ );
or   ( new_n33454_, new_n19614_, new_n19267_ );
and  ( new_n33455_, new_n33454_, new_n18920_ );
or   ( new_n33456_, new_n33455_, new_n33438_ );
or   ( new_n33457_, new_n18588_, new_n18247_ );
and  ( new_n33458_, new_n33457_, new_n18242_ );
and  ( new_n33459_, new_n33458_, new_n33456_ );
and  ( new_n33460_, new_n20792_, new_n20370_ );
or   ( new_n33461_, new_n33460_, new_n20373_ );
or   ( new_n33462_, new_n33461_, new_n33441_ );
or   ( new_n33463_, new_n19994_, new_n19618_ );
and  ( new_n33464_, new_n33463_, new_n19611_ );
and  ( new_n33465_, new_n33464_, new_n33462_ );
or   ( new_n33466_, new_n33465_, new_n33440_ );
and  ( new_n33467_, new_n33466_, new_n33459_ );
or   ( new_n33468_, new_n33467_, new_n33452_ );
or   ( new_n33469_, new_n32986_, new_n32968_ );
and  ( new_n33470_, new_n33469_, new_n33001_ );
or   ( new_n33471_, new_n32990_, new_n32954_ );
and  ( new_n33472_, new_n33471_, new_n32987_ );
or   ( new_n33473_, new_n33472_, new_n33447_ );
and  ( new_n33474_, new_n33473_, new_n33470_ );
or   ( new_n33475_, new_n30637_, new_n17108_ );
and  ( new_n33476_, new_n33475_, new_n30633_ );
or   ( new_n33477_, new_n17922_, new_n17601_ );
and  ( new_n33478_, new_n33477_, new_n17598_ );
or   ( new_n33479_, new_n33478_, new_n33449_ );
and  ( new_n33480_, new_n33479_, new_n33476_ );
or   ( new_n33481_, new_n33480_, new_n33448_ );
and  ( new_n33482_, new_n33481_, new_n33474_ );
and  ( new_n33483_, new_n33482_, new_n33468_ );
and  ( new_n33484_, new_n33483_, new_n33453_ );
or   ( new_n33485_, new_n33484_, new_n33329_ );
and  ( new_n33486_, new_n30822_, new_n30813_ );
and  ( new_n33487_, new_n30841_, new_n30833_ );
and  ( new_n33488_, new_n33487_, new_n33486_ );
and  ( new_n33489_, new_n30899_, new_n30890_ );
and  ( new_n33490_, new_n30914_, new_n30906_ );
and  ( new_n33491_, new_n33490_, new_n33489_ );
and  ( new_n33492_, new_n30929_, new_n30921_ );
and  ( new_n33493_, new_n30945_, new_n30934_ );
and  ( new_n33494_, new_n33493_, new_n33492_ );
and  ( new_n33495_, new_n30953_, new_n30941_ );
and  ( new_n33496_, new_n30973_, new_n30960_ );
and  ( new_n33497_, new_n30978_, new_n30966_ );
and  ( new_n33498_, new_n30994_, new_n30982_ );
and  ( new_n33499_, new_n30999_, new_n30988_ );
and  ( new_n33500_, new_n31051_, new_n31047_ );
or   ( new_n33501_, new_n31026_, new_n31020_ );
and  ( new_n33502_, new_n33501_, new_n31049_ );
or   ( new_n33503_, new_n33502_, new_n33500_ );
and  ( new_n33504_, new_n31015_, new_n31009_ );
and  ( new_n33505_, new_n33504_, new_n33503_ );
and  ( new_n33506_, new_n33505_, new_n33499_ );
or   ( new_n33507_, new_n31064_, new_n31000_ );
and  ( new_n33508_, new_n33507_, new_n30988_ );
or   ( new_n33509_, new_n31016_, new_n31006_ );
and  ( new_n33510_, new_n33509_, new_n31009_ );
and  ( new_n33511_, new_n33510_, new_n33499_ );
or   ( new_n33512_, new_n33511_, new_n33508_ );
or   ( new_n33513_, new_n33512_, new_n33506_ );
and  ( new_n33514_, new_n33513_, new_n33498_ );
and  ( new_n33515_, new_n33514_, new_n33497_ );
or   ( new_n33516_, new_n31077_, new_n31059_ );
and  ( new_n33517_, new_n33516_, new_n30966_ );
or   ( new_n33518_, new_n31063_, new_n31060_ );
and  ( new_n33519_, new_n33518_, new_n30982_ );
and  ( new_n33520_, new_n33519_, new_n33497_ );
or   ( new_n33521_, new_n33520_, new_n33517_ );
or   ( new_n33522_, new_n33521_, new_n33515_ );
and  ( new_n33523_, new_n33522_, new_n33496_ );
and  ( new_n33524_, new_n33523_, new_n33495_ );
or   ( new_n33525_, new_n31090_, new_n31072_ );
and  ( new_n33526_, new_n33525_, new_n30941_ );
or   ( new_n33527_, new_n31076_, new_n31073_ );
and  ( new_n33528_, new_n33527_, new_n30960_ );
and  ( new_n33529_, new_n33528_, new_n33495_ );
or   ( new_n33530_, new_n33529_, new_n33526_ );
or   ( new_n33531_, new_n33530_, new_n33524_ );
and  ( new_n33532_, new_n33531_, new_n33494_ );
and  ( new_n33533_, new_n33532_, new_n33491_ );
or   ( new_n33534_, new_n31098_, new_n30885_ );
and  ( new_n33535_, new_n33534_, new_n30890_ );
or   ( new_n33536_, new_n31102_, new_n31099_ );
and  ( new_n33537_, new_n33536_, new_n30906_ );
and  ( new_n33538_, new_n33537_, new_n33489_ );
or   ( new_n33539_, new_n33538_, new_n33535_ );
or   ( new_n33540_, new_n31103_, new_n31085_ );
and  ( new_n33541_, new_n33540_, new_n30921_ );
or   ( new_n33542_, new_n31089_, new_n31086_ );
and  ( new_n33543_, new_n33542_, new_n30934_ );
and  ( new_n33544_, new_n33543_, new_n33492_ );
or   ( new_n33545_, new_n33544_, new_n33541_ );
and  ( new_n33546_, new_n33545_, new_n33491_ );
or   ( new_n33547_, new_n33546_, new_n33539_ );
or   ( new_n33548_, new_n33547_, new_n33533_ );
and  ( new_n33549_, new_n30862_, new_n30855_ );
and  ( new_n33550_, new_n30877_, new_n30870_ );
and  ( new_n33551_, new_n33550_, new_n33549_ );
and  ( new_n33552_, new_n33551_, new_n33548_ );
and  ( new_n33553_, new_n33552_, new_n33488_ );
or   ( new_n33554_, new_n30823_, new_n30808_ );
and  ( new_n33555_, new_n33554_, new_n30813_ );
or   ( new_n33556_, new_n30842_, new_n30830_ );
and  ( new_n33557_, new_n33556_, new_n30833_ );
and  ( new_n33558_, new_n33557_, new_n33486_ );
or   ( new_n33559_, new_n33558_, new_n33555_ );
or   ( new_n33560_, new_n30863_, new_n30849_ );
and  ( new_n33561_, new_n33560_, new_n30855_ );
or   ( new_n33562_, new_n30878_, new_n30867_ );
and  ( new_n33563_, new_n33562_, new_n30870_ );
and  ( new_n33564_, new_n33563_, new_n33549_ );
or   ( new_n33565_, new_n33564_, new_n33561_ );
and  ( new_n33566_, new_n33565_, new_n33488_ );
or   ( new_n33567_, new_n33566_, new_n33559_ );
or   ( new_n33568_, new_n33567_, new_n33553_ );
and  ( new_n33569_, new_n30740_, new_n30731_ );
and  ( new_n33570_, new_n30759_, new_n30751_ );
and  ( new_n33571_, new_n33570_, new_n33569_ );
and  ( new_n33572_, new_n30781_, new_n30772_ );
and  ( new_n33573_, new_n30800_, new_n30792_ );
and  ( new_n33574_, new_n33573_, new_n33572_ );
and  ( new_n33575_, new_n33574_, new_n33571_ );
and  ( new_n33576_, new_n33575_, new_n33568_ );
or   ( new_n33577_, new_n30741_, new_n30726_ );
and  ( new_n33578_, new_n33577_, new_n30731_ );
or   ( new_n33579_, new_n30760_, new_n30748_ );
and  ( new_n33580_, new_n33579_, new_n30751_ );
and  ( new_n33581_, new_n33580_, new_n33569_ );
or   ( new_n33582_, new_n33581_, new_n33578_ );
or   ( new_n33583_, new_n30782_, new_n30767_ );
and  ( new_n33584_, new_n33583_, new_n30772_ );
or   ( new_n33585_, new_n30801_, new_n30789_ );
and  ( new_n33586_, new_n33585_, new_n30792_ );
and  ( new_n33587_, new_n33586_, new_n33572_ );
or   ( new_n33588_, new_n33587_, new_n33584_ );
and  ( new_n33589_, new_n33588_, new_n33571_ );
or   ( new_n33590_, new_n33589_, new_n33582_ );
or   ( new_n33591_, new_n33590_, new_n33576_ );
and  ( new_n33592_, new_n30674_, new_n30668_ );
and  ( new_n33593_, new_n30693_, new_n30685_ );
and  ( new_n33594_, new_n33593_, new_n33592_ );
and  ( new_n33595_, new_n30703_, new_n30697_ );
and  ( new_n33596_, new_n30719_, new_n30713_ );
and  ( new_n33597_, new_n33596_, new_n33595_ );
and  ( new_n33598_, new_n33597_, new_n33594_ );
and  ( new_n33599_, new_n33598_, new_n33591_ );
or   ( new_n33600_, new_n30675_, new_n30663_ );
and  ( new_n33601_, new_n33600_, new_n30668_ );
or   ( new_n33602_, new_n30686_, new_n30679_ );
and  ( new_n33603_, new_n33602_, new_n30693_ );
and  ( new_n33604_, new_n33603_, new_n33592_ );
or   ( new_n33605_, new_n33604_, new_n33601_ );
or   ( new_n33606_, new_n30704_, new_n30690_ );
and  ( new_n33607_, new_n33606_, new_n30697_ );
or   ( new_n33608_, new_n30720_, new_n30710_ );
and  ( new_n33609_, new_n33608_, new_n30713_ );
and  ( new_n33610_, new_n33609_, new_n33595_ );
or   ( new_n33611_, new_n33610_, new_n33607_ );
and  ( new_n33612_, new_n33611_, new_n33594_ );
or   ( new_n33613_, new_n33612_, new_n33605_ );
or   ( new_n33614_, new_n33613_, new_n33599_ );
and  ( new_n33615_, new_n32763_, new_n32751_ );
and  ( new_n33616_, new_n32845_, new_n32720_ );
and  ( new_n33617_, new_n33616_, new_n33615_ );
and  ( new_n33618_, new_n30642_, new_n30628_ );
and  ( new_n33619_, new_n30658_, new_n30652_ );
and  ( new_n33620_, new_n33619_, new_n33618_ );
and  ( new_n33621_, new_n33620_, new_n33617_ );
and  ( new_n33622_, new_n33621_, new_n33614_ );
or   ( new_n33623_, new_n32935_, new_n32922_ );
and  ( new_n33624_, new_n33623_, new_n32845_ );
or   ( new_n33625_, new_n32925_, new_n32921_ );
and  ( new_n33626_, new_n33625_, new_n32751_ );
and  ( new_n33627_, new_n33626_, new_n33616_ );
or   ( new_n33628_, new_n33627_, new_n33624_ );
or   ( new_n33629_, new_n30649_, new_n30636_ );
and  ( new_n33630_, new_n33629_, new_n30628_ );
or   ( new_n33631_, new_n30659_, new_n30648_ );
and  ( new_n33632_, new_n33631_, new_n30652_ );
and  ( new_n33633_, new_n33632_, new_n33618_ );
or   ( new_n33634_, new_n33633_, new_n33630_ );
and  ( new_n33635_, new_n33634_, new_n33617_ );
or   ( new_n33636_, new_n33635_, new_n33628_ );
or   ( new_n33637_, new_n33636_, new_n33622_ );
and  ( new_n33638_, new_n33000_, new_n32885_ );
or   ( new_n33639_, new_n33638_, new_n33637_ );
and  ( new_n33640_, new_n33639_, new_n33485_ );
and  ( new_n33641_, new_n33640_, new_n33328_ );
or   ( new_n33642_, new_n33641_, new_n33018_ );
or   ( new_n33643_, new_n33642_, new_n33011_ );
or   ( new_n33644_, new_n5150_, new_n4380_ );
and  ( new_n33645_, new_n33644_, new_n4369_ );
or   ( new_n33646_, new_n5152_, new_n4380_ );
or   ( new_n33647_, new_n6905_, new_n5993_ );
and  ( new_n33648_, new_n33647_, new_n5989_ );
or   ( new_n33649_, new_n6907_, new_n5993_ );
or   ( new_n33650_, new_n15319_, new_n8767_ );
or   ( new_n33651_, new_n10383_, new_n9591_ );
or   ( new_n33652_, new_n11662_, new_n11174_ );
and  ( new_n33653_, new_n33652_, new_n11168_ );
or   ( new_n33654_, new_n15259_, new_n14980_ );
or   ( new_n33655_, new_n15083_, new_n14980_ );
and  ( new_n33656_, new_n33655_, new_n15270_ );
and  ( new_n33657_, new_n33656_, new_n33654_ );
or   ( new_n33658_, new_n33657_, new_n14811_ );
or   ( new_n33659_, new_n33658_, new_n14606_ );
or   ( new_n33660_, new_n15266_, new_n14606_ );
and  ( new_n33661_, new_n33660_, new_n15283_ );
and  ( new_n33662_, new_n33661_, new_n33659_ );
or   ( new_n33663_, new_n33662_, new_n14310_ );
or   ( new_n33664_, new_n33663_, new_n13960_ );
or   ( new_n33665_, new_n15279_, new_n13960_ );
and  ( new_n33666_, new_n33665_, new_n15296_ );
and  ( new_n33667_, new_n33666_, new_n33664_ );
or   ( new_n33668_, new_n33667_, new_n13741_ );
or   ( new_n33669_, new_n33668_, new_n13260_ );
or   ( new_n33670_, new_n15292_, new_n13260_ );
and  ( new_n33671_, new_n33670_, new_n15309_ );
and  ( new_n33672_, new_n33671_, new_n33669_ );
or   ( new_n33673_, new_n33672_, new_n12733_ );
or   ( new_n33674_, new_n33673_, new_n12181_ );
or   ( new_n33675_, new_n15305_, new_n12181_ );
and  ( new_n33676_, new_n33675_, new_n12177_ );
and  ( new_n33677_, new_n33676_, new_n33674_ );
or   ( new_n33678_, new_n33677_, new_n11664_ );
or   ( new_n33679_, new_n33678_, new_n11174_ );
and  ( new_n33680_, new_n33679_, new_n33653_ );
or   ( new_n33681_, new_n33680_, new_n33651_ );
or   ( new_n33682_, new_n33681_, new_n33650_ );
or   ( new_n33683_, new_n15319_, new_n8765_ );
and  ( new_n33684_, new_n33683_, new_n7856_ );
or   ( new_n33685_, new_n10381_, new_n9591_ );
and  ( new_n33686_, new_n33685_, new_n9587_ );
or   ( new_n33687_, new_n33686_, new_n33650_ );
and  ( new_n33688_, new_n33687_, new_n33684_ );
and  ( new_n33689_, new_n33688_, new_n33682_ );
or   ( new_n33690_, new_n33689_, new_n33649_ );
and  ( new_n33691_, new_n33690_, new_n33648_ );
or   ( new_n33692_, new_n33691_, new_n33646_ );
and  ( new_n33693_, new_n33692_, new_n33645_ );
and  ( new_n33694_, new_n15561_, new_n3658_ );
and  ( new_n33695_, new_n33694_, new_n33693_ );
and  ( new_n33696_, new_n15587_, new_n15571_ );
or   ( new_n33697_, new_n33696_, new_n15560_ );
and  ( new_n33698_, new_n15589_, new_n15571_ );
and  ( new_n33699_, new_n15625_, new_n15607_ );
or   ( new_n33700_, new_n33699_, new_n15603_ );
and  ( new_n33701_, new_n15627_, new_n15607_ );
and  ( new_n33702_, new_n15992_, new_n15667_ );
and  ( new_n33703_, new_n15708_, new_n15688_ );
and  ( new_n33704_, new_n15743_, new_n15731_ );
or   ( new_n33705_, new_n33704_, new_n15725_ );
and  ( new_n33706_, new_n15932_, new_n15869_ );
and  ( new_n33707_, new_n15883_, new_n15869_ );
or   ( new_n33708_, new_n33707_, new_n15943_ );
or   ( new_n33709_, new_n33708_, new_n33706_ );
and  ( new_n33710_, new_n33709_, new_n15857_ );
and  ( new_n33711_, new_n33710_, new_n15848_ );
and  ( new_n33712_, new_n15939_, new_n15848_ );
or   ( new_n33713_, new_n33712_, new_n15956_ );
or   ( new_n33714_, new_n33713_, new_n33711_ );
and  ( new_n33715_, new_n33714_, new_n15836_ );
and  ( new_n33716_, new_n33715_, new_n15821_ );
and  ( new_n33717_, new_n15952_, new_n15821_ );
or   ( new_n33718_, new_n33717_, new_n15969_ );
or   ( new_n33719_, new_n33718_, new_n33716_ );
and  ( new_n33720_, new_n33719_, new_n15809_ );
and  ( new_n33721_, new_n33720_, new_n15797_ );
and  ( new_n33722_, new_n15965_, new_n15797_ );
or   ( new_n33723_, new_n33722_, new_n15982_ );
or   ( new_n33724_, new_n33723_, new_n33721_ );
and  ( new_n33725_, new_n33724_, new_n15782_ );
and  ( new_n33726_, new_n33725_, new_n15766_ );
and  ( new_n33727_, new_n15978_, new_n15766_ );
or   ( new_n33728_, new_n33727_, new_n15762_ );
or   ( new_n33729_, new_n33728_, new_n33726_ );
and  ( new_n33730_, new_n33729_, new_n15745_ );
and  ( new_n33731_, new_n33730_, new_n15731_ );
or   ( new_n33732_, new_n33731_, new_n33705_ );
and  ( new_n33733_, new_n33732_, new_n33703_ );
and  ( new_n33734_, new_n33733_, new_n33702_ );
and  ( new_n33735_, new_n15992_, new_n15665_ );
or   ( new_n33736_, new_n33735_, new_n15644_ );
and  ( new_n33737_, new_n15706_, new_n15688_ );
or   ( new_n33738_, new_n33737_, new_n15684_ );
and  ( new_n33739_, new_n33738_, new_n33702_ );
or   ( new_n33740_, new_n33739_, new_n33736_ );
or   ( new_n33741_, new_n33740_, new_n33734_ );
and  ( new_n33742_, new_n33741_, new_n33701_ );
or   ( new_n33743_, new_n33742_, new_n33700_ );
and  ( new_n33744_, new_n33743_, new_n33698_ );
or   ( new_n33745_, new_n33744_, new_n33697_ );
or   ( new_n33746_, new_n15547_, new_n4370_ );
and  ( new_n33747_, new_n33746_, new_n33745_ );
or   ( new_n33748_, new_n33747_, new_n33695_ );
or   ( new_n33749_, new_n20372_, new_n19619_ );
and  ( new_n33750_, new_n33749_, new_n19613_ );
or   ( new_n33751_, new_n20374_, new_n19619_ );
or   ( new_n33752_, new_n22100_, new_n21195_ );
and  ( new_n33753_, new_n33752_, new_n21191_ );
or   ( new_n33754_, new_n22102_, new_n21195_ );
or   ( new_n33755_, new_n23924_, new_n23018_ );
or   ( new_n33756_, new_n25537_, new_n24746_ );
or   ( new_n33757_, new_n30386_, new_n30112_ );
or   ( new_n33758_, new_n30215_, new_n30112_ );
and  ( new_n33759_, new_n33758_, new_n30397_ );
and  ( new_n33760_, new_n33759_, new_n33757_ );
or   ( new_n33761_, new_n33760_, new_n29945_ );
or   ( new_n33762_, new_n33761_, new_n29741_ );
or   ( new_n33763_, new_n30393_, new_n29741_ );
and  ( new_n33764_, new_n33763_, new_n30410_ );
and  ( new_n33765_, new_n33764_, new_n33762_ );
or   ( new_n33766_, new_n33765_, new_n29447_ );
or   ( new_n33767_, new_n33766_, new_n29100_ );
or   ( new_n33768_, new_n30406_, new_n29100_ );
and  ( new_n33769_, new_n33768_, new_n30423_ );
and  ( new_n33770_, new_n33769_, new_n33767_ );
or   ( new_n33771_, new_n33770_, new_n28882_ );
or   ( new_n33772_, new_n33771_, new_n28402_ );
or   ( new_n33773_, new_n30419_, new_n28402_ );
and  ( new_n33774_, new_n33773_, new_n30436_ );
and  ( new_n33775_, new_n33774_, new_n33772_ );
or   ( new_n33776_, new_n33775_, new_n27877_ );
or   ( new_n33777_, new_n33776_, new_n27328_ );
or   ( new_n33778_, new_n30432_, new_n27328_ );
and  ( new_n33779_, new_n33778_, new_n27324_ );
and  ( new_n33780_, new_n33779_, new_n33777_ );
or   ( new_n33781_, new_n33780_, new_n26812_ );
or   ( new_n33782_, new_n33781_, new_n26325_ );
or   ( new_n33783_, new_n26810_, new_n26325_ );
and  ( new_n33784_, new_n33783_, new_n26320_ );
and  ( new_n33785_, new_n33784_, new_n33782_ );
or   ( new_n33786_, new_n33785_, new_n33756_ );
or   ( new_n33787_, new_n33786_, new_n33755_ );
or   ( new_n33788_, new_n23922_, new_n23018_ );
and  ( new_n33789_, new_n33788_, new_n23014_ );
or   ( new_n33790_, new_n25535_, new_n24746_ );
and  ( new_n33791_, new_n33790_, new_n24742_ );
or   ( new_n33792_, new_n33791_, new_n33755_ );
and  ( new_n33793_, new_n33792_, new_n33789_ );
and  ( new_n33794_, new_n33793_, new_n33787_ );
or   ( new_n33795_, new_n33794_, new_n33754_ );
and  ( new_n33796_, new_n33795_, new_n33753_ );
or   ( new_n33797_, new_n33796_, new_n33751_ );
and  ( new_n33798_, new_n33797_, new_n33750_ );
and  ( new_n33799_, new_n30693_, new_n18920_ );
or   ( new_n33800_, new_n33799_, new_n33798_ );
and  ( new_n33801_, new_n30712_, new_n30698_ );
or   ( new_n33802_, new_n33801_, new_n30692_ );
and  ( new_n33803_, new_n30714_, new_n30698_ );
and  ( new_n33804_, new_n30750_, new_n30732_ );
or   ( new_n33805_, new_n33804_, new_n30728_ );
and  ( new_n33806_, new_n30752_, new_n30732_ );
and  ( new_n33807_, new_n30793_, new_n30773_ );
and  ( new_n33808_, new_n30834_, new_n30814_ );
and  ( new_n33809_, new_n31055_, new_n30995_ );
and  ( new_n33810_, new_n31008_, new_n30995_ );
or   ( new_n33811_, new_n33810_, new_n31066_ );
or   ( new_n33812_, new_n33811_, new_n33809_ );
and  ( new_n33813_, new_n33812_, new_n30983_ );
and  ( new_n33814_, new_n33813_, new_n30974_ );
and  ( new_n33815_, new_n31062_, new_n30974_ );
or   ( new_n33816_, new_n33815_, new_n31079_ );
or   ( new_n33817_, new_n33816_, new_n33814_ );
and  ( new_n33818_, new_n33817_, new_n30961_ );
and  ( new_n33819_, new_n33818_, new_n30946_ );
and  ( new_n33820_, new_n31075_, new_n30946_ );
or   ( new_n33821_, new_n33820_, new_n31092_ );
or   ( new_n33822_, new_n33821_, new_n33819_ );
and  ( new_n33823_, new_n33822_, new_n30935_ );
and  ( new_n33824_, new_n33823_, new_n30922_ );
and  ( new_n33825_, new_n31088_, new_n30922_ );
or   ( new_n33826_, new_n33825_, new_n31105_ );
or   ( new_n33827_, new_n33826_, new_n33824_ );
and  ( new_n33828_, new_n33827_, new_n30907_ );
and  ( new_n33829_, new_n33828_, new_n30891_ );
and  ( new_n33830_, new_n31101_, new_n30891_ );
or   ( new_n33831_, new_n33830_, new_n30887_ );
or   ( new_n33832_, new_n33831_, new_n33829_ );
and  ( new_n33833_, new_n33832_, new_n30871_ );
and  ( new_n33834_, new_n33833_, new_n30856_ );
and  ( new_n33835_, new_n30869_, new_n30856_ );
or   ( new_n33836_, new_n33835_, new_n30851_ );
or   ( new_n33837_, new_n33836_, new_n33834_ );
and  ( new_n33838_, new_n33837_, new_n33808_ );
and  ( new_n33839_, new_n33838_, new_n33807_ );
and  ( new_n33840_, new_n30791_, new_n30773_ );
or   ( new_n33841_, new_n33840_, new_n30769_ );
and  ( new_n33842_, new_n30832_, new_n30814_ );
or   ( new_n33843_, new_n33842_, new_n30810_ );
and  ( new_n33844_, new_n33843_, new_n33807_ );
or   ( new_n33845_, new_n33844_, new_n33841_ );
or   ( new_n33846_, new_n33845_, new_n33839_ );
and  ( new_n33847_, new_n33846_, new_n33806_ );
or   ( new_n33848_, new_n33847_, new_n33805_ );
and  ( new_n33849_, new_n33848_, new_n33803_ );
or   ( new_n33850_, new_n33849_, new_n33802_ );
or   ( new_n33851_, new_n30679_, new_n19614_ );
or   ( new_n33852_, new_n33851_, new_n33850_ );
and  ( new_n33853_, new_n33852_, new_n33800_ );
and  ( new_n33854_, new_n33853_, new_n33748_ );
and  ( new_n33855_, new_n33746_, new_n33693_ );
and  ( new_n33856_, new_n33745_, new_n33694_ );
or   ( new_n33857_, new_n33856_, new_n33855_ );
or   ( new_n33858_, new_n33851_, new_n33798_ );
or   ( new_n33859_, new_n33850_, new_n33799_ );
and  ( new_n33860_, new_n33859_, new_n33858_ );
and  ( new_n33861_, new_n33860_, new_n33857_ );
or   ( new_n33862_, new_n33861_, new_n33854_ );
and  ( new_n33863_, new_n33173_, new_n33170_ );
and  ( new_n33864_, new_n33326_, new_n33171_ );
or   ( new_n33865_, new_n33864_, new_n33863_ );
or   ( new_n33866_, new_n33637_, new_n33329_ );
or   ( new_n33867_, new_n33638_, new_n33484_ );
and  ( new_n33868_, new_n33867_, new_n33866_ );
and  ( new_n33869_, new_n33868_, new_n33865_ );
and  ( new_n33870_, new_n15509_, new_n15325_ );
and  ( new_n33871_, new_n15998_, new_n15505_ );
or   ( new_n33872_, new_n33871_, new_n33870_ );
or   ( new_n33873_, new_n30638_, new_n30453_ );
or   ( new_n33874_, new_n31122_, new_n30634_ );
and  ( new_n33875_, new_n33874_, new_n33873_ );
and  ( new_n33876_, new_n33875_, new_n33872_ );
or   ( new_n33877_, new_n33876_, new_n33869_ );
or   ( new_n33878_, new_n33877_, new_n33862_ );
or   ( new_n33879_, new_n33878_, new_n33643_ );
or   ( new_n33880_, new_n4375_, new_n4371_ );
or   ( new_n33881_, new_n31545_, new_n2310_ );
or   ( new_n33882_, new_n33881_, new_n33880_ );
or   ( new_n33883_, new_n33882_, new_n33693_ );
or   ( new_n33884_, new_n4375_, new_n3660_ );
and  ( new_n33885_, new_n33884_, new_n2970_ );
or   ( new_n33886_, new_n33885_, new_n33881_ );
or   ( new_n33887_, new_n31545_, new_n2308_ );
and  ( new_n33888_, new_n33887_, new_n31983_ );
and  ( new_n33889_, new_n33888_, new_n33886_ );
and  ( new_n33890_, new_n33889_, new_n33883_ );
or   ( new_n33891_, new_n32051_, new_n31815_ );
and  ( new_n33892_, new_n33891_, new_n33890_ );
and  ( new_n33893_, new_n32019_, new_n31977_ );
and  ( new_n33894_, new_n15566_, new_n15562_ );
and  ( new_n33895_, new_n32011_, new_n15525_ );
and  ( new_n33896_, new_n33895_, new_n33894_ );
and  ( new_n33897_, new_n33896_, new_n33745_ );
and  ( new_n33898_, new_n15566_, new_n15549_ );
or   ( new_n33899_, new_n33898_, new_n15536_ );
and  ( new_n33900_, new_n33899_, new_n33895_ );
and  ( new_n33901_, new_n32011_, new_n15523_ );
or   ( new_n33902_, new_n33901_, new_n32056_ );
or   ( new_n33903_, new_n33902_, new_n33900_ );
or   ( new_n33904_, new_n33903_, new_n33897_ );
and  ( new_n33905_, new_n33904_, new_n33893_ );
or   ( new_n33906_, new_n33905_, new_n33892_ );
or   ( new_n33907_, new_n32954_, new_n32921_ );
or   ( new_n33908_, new_n32960_, new_n17602_ );
or   ( new_n33909_, new_n19615_, new_n18248_ );
or   ( new_n33910_, new_n33909_, new_n33908_ );
or   ( new_n33911_, new_n33910_, new_n33798_ );
or   ( new_n33912_, new_n18922_, new_n18248_ );
and  ( new_n33913_, new_n33912_, new_n18244_ );
or   ( new_n33914_, new_n33913_, new_n33908_ );
or   ( new_n33915_, new_n32960_, new_n17600_ );
and  ( new_n33916_, new_n33915_, new_n32992_ );
and  ( new_n33917_, new_n33916_, new_n33914_ );
and  ( new_n33918_, new_n33917_, new_n33911_ );
or   ( new_n33919_, new_n33918_, new_n33907_ );
and  ( new_n33920_, new_n32764_, new_n30653_ );
and  ( new_n33921_, new_n30694_, new_n30669_ );
and  ( new_n33922_, new_n33921_, new_n33920_ );
and  ( new_n33923_, new_n33922_, new_n33850_ );
and  ( new_n33924_, new_n30681_, new_n30669_ );
or   ( new_n33925_, new_n33924_, new_n30665_ );
and  ( new_n33926_, new_n33925_, new_n33920_ );
and  ( new_n33927_, new_n32764_, new_n30651_ );
or   ( new_n33928_, new_n33927_, new_n32927_ );
or   ( new_n33929_, new_n33928_, new_n33926_ );
or   ( new_n33930_, new_n33929_, new_n33923_ );
and  ( new_n33931_, new_n32987_, new_n32751_ );
or   ( new_n33932_, new_n33931_, new_n33930_ );
and  ( new_n33933_, new_n33932_, new_n33919_ );
and  ( new_n33934_, new_n33933_, new_n33906_ );
and  ( new_n33935_, new_n33893_, new_n33890_ );
and  ( new_n33936_, new_n33904_, new_n33891_ );
or   ( new_n33937_, new_n33936_, new_n33935_ );
or   ( new_n33938_, new_n33930_, new_n33907_ );
or   ( new_n33939_, new_n33931_, new_n33918_ );
and  ( new_n33940_, new_n33939_, new_n33938_ );
and  ( new_n33941_, new_n33940_, new_n33937_ );
or   ( new_n33942_, new_n33941_, new_n33934_ );
or   ( new_n33943_, new_n33942_, new_n33879_ );
and  ( new_n33944_, new_n33105_, new_n33092_ );
or   ( new_n33945_, new_n33944_, new_n33051_ );
or   ( new_n33946_, new_n33945_, new_n33048_ );
or   ( new_n33947_, new_n33099_, new_n33048_ );
and  ( new_n33948_, new_n33947_, new_n33046_ );
and  ( new_n33949_, new_n33948_, new_n33946_ );
or   ( new_n33950_, new_n33949_, new_n33039_ );
and  ( new_n33951_, new_n33950_, new_n33037_ );
or   ( new_n33952_, new_n33951_, new_n33030_ );
and  ( new_n33953_, new_n33952_, new_n33120_ );
or   ( new_n33954_, new_n33953_, new_n33027_ );
and  ( new_n33955_, new_n33954_, new_n33025_ );
or   ( new_n33956_, new_n33955_, new_n33129_ );
and  ( new_n33957_, new_n33956_, new_n33151_ );
or   ( new_n33958_, new_n33137_, new_n33126_ );
or   ( new_n33959_, new_n33958_, new_n33957_ );
or   ( new_n33960_, new_n33145_, new_n33137_ );
and  ( new_n33961_, new_n33960_, new_n33166_ );
and  ( new_n33962_, new_n33961_, new_n33959_ );
and  ( new_n33963_, new_n32010_, new_n31981_ );
and  ( new_n33964_, new_n33963_, new_n33962_ );
or   ( new_n33965_, new_n32054_, new_n31544_ );
or   ( new_n33966_, new_n33261_, new_n33248_ );
and  ( new_n33967_, new_n33966_, new_n33206_ );
and  ( new_n33968_, new_n33967_, new_n33203_ );
and  ( new_n33969_, new_n33255_, new_n33203_ );
or   ( new_n33970_, new_n33969_, new_n33201_ );
or   ( new_n33971_, new_n33970_, new_n33968_ );
and  ( new_n33972_, new_n33971_, new_n33194_ );
or   ( new_n33973_, new_n33972_, new_n33192_ );
and  ( new_n33974_, new_n33973_, new_n33185_ );
or   ( new_n33975_, new_n33974_, new_n33276_ );
and  ( new_n33976_, new_n33975_, new_n33182_ );
or   ( new_n33977_, new_n33976_, new_n33180_ );
and  ( new_n33978_, new_n33977_, new_n33285_ );
or   ( new_n33979_, new_n33978_, new_n33307_ );
and  ( new_n33980_, new_n33290_, new_n33282_ );
and  ( new_n33981_, new_n33980_, new_n33979_ );
and  ( new_n33982_, new_n33301_, new_n33290_ );
or   ( new_n33983_, new_n33982_, new_n33322_ );
or   ( new_n33984_, new_n33983_, new_n33981_ );
and  ( new_n33985_, new_n33984_, new_n33965_ );
or   ( new_n33986_, new_n33985_, new_n33964_ );
and  ( new_n33987_, new_n32990_, new_n32763_ );
and  ( new_n33988_, new_n33419_, new_n33406_ );
or   ( new_n33989_, new_n33988_, new_n33362_ );
or   ( new_n33990_, new_n33989_, new_n33359_ );
or   ( new_n33991_, new_n33413_, new_n33359_ );
and  ( new_n33992_, new_n33991_, new_n33357_ );
and  ( new_n33993_, new_n33992_, new_n33990_ );
or   ( new_n33994_, new_n33993_, new_n33350_ );
and  ( new_n33995_, new_n33994_, new_n33348_ );
or   ( new_n33996_, new_n33995_, new_n33341_ );
and  ( new_n33997_, new_n33996_, new_n33434_ );
or   ( new_n33998_, new_n33997_, new_n33338_ );
and  ( new_n33999_, new_n33998_, new_n33336_ );
or   ( new_n34000_, new_n33999_, new_n33443_ );
and  ( new_n34001_, new_n34000_, new_n33465_ );
or   ( new_n34002_, new_n33451_, new_n33440_ );
or   ( new_n34003_, new_n34002_, new_n34001_ );
or   ( new_n34004_, new_n33459_, new_n33451_ );
and  ( new_n34005_, new_n34004_, new_n33480_ );
and  ( new_n34006_, new_n34005_, new_n34003_ );
or   ( new_n34007_, new_n34006_, new_n33987_ );
or   ( new_n34008_, new_n33545_, new_n33532_ );
and  ( new_n34009_, new_n34008_, new_n33491_ );
and  ( new_n34010_, new_n34009_, new_n33551_ );
and  ( new_n34011_, new_n33551_, new_n33539_ );
or   ( new_n34012_, new_n34011_, new_n33565_ );
or   ( new_n34013_, new_n34012_, new_n34010_ );
and  ( new_n34014_, new_n34013_, new_n33488_ );
or   ( new_n34015_, new_n34014_, new_n33559_ );
and  ( new_n34016_, new_n34015_, new_n33574_ );
or   ( new_n34017_, new_n34016_, new_n33588_ );
and  ( new_n34018_, new_n34017_, new_n33571_ );
or   ( new_n34019_, new_n34018_, new_n33582_ );
and  ( new_n34020_, new_n34019_, new_n33597_ );
or   ( new_n34021_, new_n34020_, new_n33611_ );
and  ( new_n34022_, new_n33620_, new_n33594_ );
and  ( new_n34023_, new_n34022_, new_n34021_ );
and  ( new_n34024_, new_n33620_, new_n33605_ );
or   ( new_n34025_, new_n34024_, new_n33634_ );
or   ( new_n34026_, new_n34025_, new_n34023_ );
or   ( new_n34027_, new_n32959_, new_n32925_ );
or   ( new_n34028_, new_n34027_, new_n34026_ );
and  ( new_n34029_, new_n34028_, new_n34007_ );
and  ( new_n34030_, new_n34029_, new_n33986_ );
and  ( new_n34031_, new_n33965_, new_n33962_ );
and  ( new_n34032_, new_n33984_, new_n33963_ );
or   ( new_n34033_, new_n34032_, new_n34031_ );
or   ( new_n34034_, new_n34026_, new_n33987_ );
or   ( new_n34035_, new_n34027_, new_n34006_ );
and  ( new_n34036_, new_n34035_, new_n34034_ );
and  ( new_n34037_, new_n34036_, new_n34033_ );
or   ( new_n34038_, new_n33135_, new_n33124_ );
or   ( new_n34039_, new_n33147_, new_n33125_ );
and  ( new_n34040_, new_n34039_, new_n33143_ );
or   ( new_n34041_, new_n34040_, new_n34038_ );
or   ( new_n34042_, new_n33141_, new_n33135_ );
and  ( new_n34043_, new_n34042_, new_n33164_ );
and  ( new_n34044_, new_n34043_, new_n34041_ );
or   ( new_n34045_, new_n33127_, new_n33125_ );
or   ( new_n34046_, new_n34045_, new_n34038_ );
or   ( new_n34047_, new_n33128_, new_n33021_ );
or   ( new_n34048_, new_n33116_, new_n33026_ );
and  ( new_n34049_, new_n34048_, new_n33023_ );
or   ( new_n34050_, new_n34049_, new_n34047_ );
or   ( new_n34051_, new_n33128_, new_n33020_ );
and  ( new_n34052_, new_n34051_, new_n33149_ );
and  ( new_n34053_, new_n34052_, new_n34050_ );
or   ( new_n34054_, new_n33028_, new_n33026_ );
or   ( new_n34055_, new_n34054_, new_n34047_ );
or   ( new_n34056_, new_n33033_, new_n33029_ );
or   ( new_n34057_, new_n33041_, new_n33038_ );
and  ( new_n34058_, new_n34057_, new_n33035_ );
or   ( new_n34059_, new_n34058_, new_n34056_ );
or   ( new_n34060_, new_n33032_, new_n33029_ );
and  ( new_n34061_, new_n34060_, new_n33118_ );
and  ( new_n34062_, new_n34061_, new_n34059_ );
and  ( new_n34063_, new_n33070_, new_n33065_ );
or   ( new_n34064_, new_n34063_, new_n33059_ );
or   ( new_n34065_, new_n34064_, new_n33058_ );
or   ( new_n34066_, new_n33068_, new_n33058_ );
and  ( new_n34067_, new_n34066_, new_n33079_ );
and  ( new_n34068_, new_n34067_, new_n34065_ );
or   ( new_n34069_, new_n34068_, new_n33057_ );
or   ( new_n34070_, new_n34069_, new_n33056_ );
or   ( new_n34071_, new_n33077_, new_n33056_ );
and  ( new_n34072_, new_n34071_, new_n33088_ );
and  ( new_n34073_, new_n34072_, new_n34070_ );
or   ( new_n34074_, new_n34073_, new_n33055_ );
or   ( new_n34075_, new_n34074_, new_n33053_ );
or   ( new_n34076_, new_n33086_, new_n33053_ );
and  ( new_n34077_, new_n34076_, new_n33103_ );
and  ( new_n34078_, new_n34077_, new_n34075_ );
or   ( new_n34079_, new_n34078_, new_n33052_ );
or   ( new_n34080_, new_n34079_, new_n33050_ );
or   ( new_n34081_, new_n33101_, new_n33050_ );
and  ( new_n34082_, new_n34081_, new_n33097_ );
and  ( new_n34083_, new_n34082_, new_n34080_ );
or   ( new_n34084_, new_n34083_, new_n33049_ );
and  ( new_n34085_, new_n34084_, new_n33095_ );
or   ( new_n34086_, new_n34085_, new_n33047_ );
and  ( new_n34087_, new_n34086_, new_n33044_ );
or   ( new_n34088_, new_n34087_, new_n33042_ );
or   ( new_n34089_, new_n34088_, new_n33038_ );
or   ( new_n34090_, new_n34089_, new_n34056_ );
and  ( new_n34091_, new_n34090_, new_n34062_ );
or   ( new_n34092_, new_n34091_, new_n34055_ );
and  ( new_n34093_, new_n34092_, new_n34053_ );
or   ( new_n34094_, new_n34093_, new_n34046_ );
and  ( new_n34095_, new_n34094_, new_n34044_ );
or   ( new_n34096_, new_n15513_, new_n1798_ );
and  ( new_n34097_, new_n34096_, new_n34095_ );
and  ( new_n34098_, new_n15514_, new_n2306_ );
and  ( new_n34099_, new_n33288_, new_n33280_ );
and  ( new_n34100_, new_n33306_, new_n33281_ );
or   ( new_n34101_, new_n34100_, new_n33297_ );
and  ( new_n34102_, new_n34101_, new_n34099_ );
and  ( new_n34103_, new_n33300_, new_n33288_ );
or   ( new_n34104_, new_n34103_, new_n33318_ );
or   ( new_n34105_, new_n34104_, new_n34102_ );
and  ( new_n34106_, new_n33283_, new_n33281_ );
and  ( new_n34107_, new_n34106_, new_n34099_ );
and  ( new_n34108_, new_n33284_, new_n33174_ );
and  ( new_n34109_, new_n33275_, new_n33181_ );
or   ( new_n34110_, new_n34109_, new_n33176_ );
and  ( new_n34111_, new_n34110_, new_n34108_ );
and  ( new_n34112_, new_n33284_, new_n33179_ );
or   ( new_n34113_, new_n34112_, new_n33303_ );
or   ( new_n34114_, new_n34113_, new_n34111_ );
and  ( new_n34115_, new_n33183_, new_n33181_ );
and  ( new_n34116_, new_n34115_, new_n34108_ );
and  ( new_n34117_, new_n33200_, new_n33193_ );
or   ( new_n34118_, new_n34117_, new_n33188_ );
and  ( new_n34119_, new_n33186_, new_n33184_ );
and  ( new_n34120_, new_n34119_, new_n34118_ );
and  ( new_n34121_, new_n33191_, new_n33184_ );
or   ( new_n34122_, new_n34121_, new_n33272_ );
or   ( new_n34123_, new_n34122_, new_n34120_ );
or   ( new_n34124_, new_n33224_, new_n33221_ );
and  ( new_n34125_, new_n34124_, new_n33214_ );
and  ( new_n34126_, new_n34125_, new_n33213_ );
and  ( new_n34127_, new_n33227_, new_n33213_ );
or   ( new_n34128_, new_n34127_, new_n33233_ );
or   ( new_n34129_, new_n34128_, new_n34126_ );
and  ( new_n34130_, new_n34129_, new_n33212_ );
and  ( new_n34131_, new_n34130_, new_n33211_ );
and  ( new_n34132_, new_n33236_, new_n33211_ );
or   ( new_n34133_, new_n34132_, new_n33242_ );
or   ( new_n34134_, new_n34133_, new_n34131_ );
and  ( new_n34135_, new_n34134_, new_n33210_ );
and  ( new_n34136_, new_n34135_, new_n33208_ );
and  ( new_n34137_, new_n33245_, new_n33208_ );
or   ( new_n34138_, new_n34137_, new_n33259_ );
or   ( new_n34139_, new_n34138_, new_n34136_ );
and  ( new_n34140_, new_n34139_, new_n33207_ );
and  ( new_n34141_, new_n34140_, new_n33205_ );
and  ( new_n34142_, new_n33257_, new_n33205_ );
or   ( new_n34143_, new_n34142_, new_n33253_ );
or   ( new_n34144_, new_n34143_, new_n34141_ );
and  ( new_n34145_, new_n34144_, new_n33204_ );
and  ( new_n34146_, new_n34145_, new_n33202_ );
and  ( new_n34147_, new_n33251_, new_n33202_ );
or   ( new_n34148_, new_n34147_, new_n33197_ );
or   ( new_n34149_, new_n34148_, new_n34146_ );
and  ( new_n34150_, new_n34149_, new_n33195_ );
and  ( new_n34151_, new_n34150_, new_n33193_ );
and  ( new_n34152_, new_n34151_, new_n34119_ );
or   ( new_n34153_, new_n34152_, new_n34123_ );
and  ( new_n34154_, new_n34153_, new_n34116_ );
or   ( new_n34155_, new_n34154_, new_n34114_ );
and  ( new_n34156_, new_n34155_, new_n34107_ );
or   ( new_n34157_, new_n34156_, new_n34105_ );
and  ( new_n34158_, new_n34157_, new_n34098_ );
or   ( new_n34159_, new_n34158_, new_n34097_ );
or   ( new_n34160_, new_n33442_, new_n33330_ );
and  ( new_n34161_, new_n30382_, new_n30329_ );
or   ( new_n34162_, new_n34161_, new_n30378_ );
or   ( new_n34163_, new_n34162_, new_n33378_ );
and  ( new_n34164_, new_n34163_, new_n33382_ );
or   ( new_n34165_, new_n34164_, new_n33370_ );
or   ( new_n34166_, new_n34165_, new_n33369_ );
or   ( new_n34167_, new_n33385_, new_n33369_ );
and  ( new_n34168_, new_n34167_, new_n33391_ );
and  ( new_n34169_, new_n34168_, new_n34166_ );
or   ( new_n34170_, new_n34169_, new_n33368_ );
or   ( new_n34171_, new_n34170_, new_n33367_ );
or   ( new_n34172_, new_n33394_, new_n33367_ );
and  ( new_n34173_, new_n34172_, new_n33400_ );
and  ( new_n34174_, new_n34173_, new_n34171_ );
or   ( new_n34175_, new_n34174_, new_n33366_ );
or   ( new_n34176_, new_n34175_, new_n33364_ );
or   ( new_n34177_, new_n33403_, new_n33364_ );
and  ( new_n34178_, new_n34177_, new_n33417_ );
and  ( new_n34179_, new_n34178_, new_n34176_ );
or   ( new_n34180_, new_n34179_, new_n33363_ );
or   ( new_n34181_, new_n34180_, new_n33361_ );
or   ( new_n34182_, new_n33415_, new_n33361_ );
and  ( new_n34183_, new_n34182_, new_n33411_ );
and  ( new_n34184_, new_n34183_, new_n34181_ );
or   ( new_n34185_, new_n34184_, new_n33360_ );
and  ( new_n34186_, new_n34185_, new_n33409_ );
or   ( new_n34187_, new_n34186_, new_n33358_ );
and  ( new_n34188_, new_n34187_, new_n33353_ );
or   ( new_n34189_, new_n34188_, new_n33351_ );
or   ( new_n34190_, new_n34189_, new_n33349_ );
or   ( new_n34191_, new_n33356_, new_n33349_ );
and  ( new_n34192_, new_n34191_, new_n33344_ );
and  ( new_n34193_, new_n34192_, new_n34190_ );
or   ( new_n34194_, new_n34193_, new_n33342_ );
or   ( new_n34195_, new_n34194_, new_n33340_ );
or   ( new_n34196_, new_n33347_, new_n33340_ );
and  ( new_n34197_, new_n34196_, new_n33430_ );
and  ( new_n34198_, new_n34197_, new_n34195_ );
or   ( new_n34199_, new_n33339_, new_n33337_ );
or   ( new_n34200_, new_n34199_, new_n34198_ );
or   ( new_n34201_, new_n34200_, new_n34160_ );
or   ( new_n34202_, new_n33433_, new_n33337_ );
and  ( new_n34203_, new_n34202_, new_n33332_ );
or   ( new_n34204_, new_n34203_, new_n34160_ );
or   ( new_n34205_, new_n33442_, new_n33335_ );
and  ( new_n34206_, new_n34205_, new_n33461_ );
and  ( new_n34207_, new_n34206_, new_n34204_ );
and  ( new_n34208_, new_n34207_, new_n34201_ );
or   ( new_n34209_, new_n33450_, new_n33438_ );
or   ( new_n34210_, new_n33441_, new_n33439_ );
or   ( new_n34211_, new_n34210_, new_n34209_ );
or   ( new_n34212_, new_n34211_, new_n34208_ );
or   ( new_n34213_, new_n33464_, new_n33439_ );
and  ( new_n34214_, new_n34213_, new_n33455_ );
or   ( new_n34215_, new_n34214_, new_n34209_ );
or   ( new_n34216_, new_n33458_, new_n33450_ );
and  ( new_n34217_, new_n34216_, new_n33478_ );
and  ( new_n34218_, new_n34217_, new_n34215_ );
and  ( new_n34219_, new_n34218_, new_n34212_ );
or   ( new_n34220_, new_n30649_, new_n17109_ );
or   ( new_n34221_, new_n34220_, new_n34219_ );
and  ( new_n34222_, new_n33596_, new_n33569_ );
or   ( new_n34223_, new_n33510_, new_n33505_ );
and  ( new_n34224_, new_n34223_, new_n33499_ );
and  ( new_n34225_, new_n34224_, new_n33498_ );
and  ( new_n34226_, new_n33508_, new_n33498_ );
or   ( new_n34227_, new_n34226_, new_n33519_ );
or   ( new_n34228_, new_n34227_, new_n34225_ );
and  ( new_n34229_, new_n34228_, new_n33497_ );
and  ( new_n34230_, new_n34229_, new_n33496_ );
and  ( new_n34231_, new_n33517_, new_n33496_ );
or   ( new_n34232_, new_n34231_, new_n33528_ );
or   ( new_n34233_, new_n34232_, new_n34230_ );
and  ( new_n34234_, new_n34233_, new_n33495_ );
and  ( new_n34235_, new_n34234_, new_n33493_ );
and  ( new_n34236_, new_n33526_, new_n33493_ );
or   ( new_n34237_, new_n34236_, new_n33543_ );
or   ( new_n34238_, new_n34237_, new_n34235_ );
and  ( new_n34239_, new_n34238_, new_n33492_ );
and  ( new_n34240_, new_n34239_, new_n33490_ );
and  ( new_n34241_, new_n33541_, new_n33490_ );
or   ( new_n34242_, new_n34241_, new_n33537_ );
or   ( new_n34243_, new_n34242_, new_n34240_ );
and  ( new_n34244_, new_n34243_, new_n33489_ );
or   ( new_n34245_, new_n34244_, new_n33535_ );
and  ( new_n34246_, new_n34245_, new_n33550_ );
or   ( new_n34247_, new_n34246_, new_n33563_ );
and  ( new_n34248_, new_n34247_, new_n33549_ );
and  ( new_n34249_, new_n34248_, new_n33487_ );
and  ( new_n34250_, new_n33561_, new_n33487_ );
or   ( new_n34251_, new_n34250_, new_n33557_ );
or   ( new_n34252_, new_n34251_, new_n34249_ );
and  ( new_n34253_, new_n34252_, new_n33486_ );
and  ( new_n34254_, new_n34253_, new_n33573_ );
and  ( new_n34255_, new_n33573_, new_n33555_ );
or   ( new_n34256_, new_n34255_, new_n33586_ );
or   ( new_n34257_, new_n34256_, new_n34254_ );
and  ( new_n34258_, new_n33572_, new_n33570_ );
and  ( new_n34259_, new_n34258_, new_n34257_ );
and  ( new_n34260_, new_n34259_, new_n34222_ );
and  ( new_n34261_, new_n33584_, new_n33570_ );
or   ( new_n34262_, new_n34261_, new_n33580_ );
and  ( new_n34263_, new_n34262_, new_n34222_ );
and  ( new_n34264_, new_n33596_, new_n33578_ );
or   ( new_n34265_, new_n34264_, new_n33609_ );
or   ( new_n34266_, new_n34265_, new_n34263_ );
or   ( new_n34267_, new_n34266_, new_n34260_ );
and  ( new_n34268_, new_n33619_, new_n33592_ );
and  ( new_n34269_, new_n33595_, new_n33593_ );
and  ( new_n34270_, new_n34269_, new_n34268_ );
and  ( new_n34271_, new_n34270_, new_n34267_ );
and  ( new_n34272_, new_n33607_, new_n33593_ );
or   ( new_n34273_, new_n34272_, new_n33603_ );
and  ( new_n34274_, new_n34273_, new_n34268_ );
and  ( new_n34275_, new_n33619_, new_n33601_ );
or   ( new_n34276_, new_n34275_, new_n33632_ );
or   ( new_n34277_, new_n34276_, new_n34274_ );
or   ( new_n34278_, new_n34277_, new_n34271_ );
and  ( new_n34279_, new_n30642_, new_n17108_ );
or   ( new_n34280_, new_n34279_, new_n34278_ );
and  ( new_n34281_, new_n34280_, new_n34221_ );
and  ( new_n34282_, new_n34281_, new_n34159_ );
or   ( new_n34283_, new_n15553_, new_n4014_ );
and  ( new_n34284_, new_n34283_, new_n33957_ );
and  ( new_n34285_, new_n15554_, new_n4015_ );
and  ( new_n34286_, new_n34285_, new_n33979_ );
or   ( new_n34287_, new_n34286_, new_n34284_ );
or   ( new_n34288_, new_n30686_, new_n19268_ );
or   ( new_n34289_, new_n34288_, new_n34001_ );
and  ( new_n34290_, new_n30685_, new_n19267_ );
or   ( new_n34291_, new_n34290_, new_n34021_ );
and  ( new_n34292_, new_n34291_, new_n34289_ );
and  ( new_n34293_, new_n34292_, new_n34287_ );
or   ( new_n34294_, new_n33880_, new_n33645_ );
and  ( new_n34295_, new_n34294_, new_n33885_ );
or   ( new_n34296_, new_n33880_, new_n33646_ );
or   ( new_n34297_, new_n33684_, new_n33649_ );
and  ( new_n34298_, new_n34297_, new_n33648_ );
or   ( new_n34299_, new_n33650_, new_n33649_ );
or   ( new_n34300_, new_n33679_, new_n33651_ );
or   ( new_n34301_, new_n33653_, new_n33651_ );
and  ( new_n34302_, new_n34301_, new_n33686_ );
and  ( new_n34303_, new_n34302_, new_n34300_ );
or   ( new_n34304_, new_n34303_, new_n34299_ );
and  ( new_n34305_, new_n34304_, new_n34298_ );
or   ( new_n34306_, new_n34305_, new_n34296_ );
and  ( new_n34307_, new_n34306_, new_n34295_ );
and  ( new_n34308_, new_n15524_, new_n2305_ );
and  ( new_n34309_, new_n34308_, new_n34307_ );
or   ( new_n34310_, new_n15521_, new_n2309_ );
and  ( new_n34311_, new_n33894_, new_n33697_ );
or   ( new_n34312_, new_n34311_, new_n33899_ );
and  ( new_n34313_, new_n33894_, new_n33698_ );
and  ( new_n34314_, new_n33736_, new_n33701_ );
or   ( new_n34315_, new_n34314_, new_n33700_ );
and  ( new_n34316_, new_n33702_, new_n33701_ );
and  ( new_n34317_, new_n33705_, new_n33703_ );
or   ( new_n34318_, new_n34317_, new_n33738_ );
and  ( new_n34319_, new_n33731_, new_n33703_ );
or   ( new_n34320_, new_n34319_, new_n34318_ );
and  ( new_n34321_, new_n34320_, new_n34316_ );
or   ( new_n34322_, new_n34321_, new_n34315_ );
and  ( new_n34323_, new_n34322_, new_n34313_ );
or   ( new_n34324_, new_n34323_, new_n34312_ );
and  ( new_n34325_, new_n34324_, new_n34310_ );
or   ( new_n34326_, new_n34325_, new_n34309_ );
or   ( new_n34327_, new_n33843_, new_n33838_ );
and  ( new_n34328_, new_n33807_, new_n33806_ );
and  ( new_n34329_, new_n34328_, new_n34327_ );
and  ( new_n34330_, new_n33841_, new_n33806_ );
or   ( new_n34331_, new_n34330_, new_n33805_ );
or   ( new_n34332_, new_n34331_, new_n34329_ );
and  ( new_n34333_, new_n34332_, new_n33803_ );
or   ( new_n34334_, new_n34333_, new_n33802_ );
and  ( new_n34335_, new_n34334_, new_n33921_ );
or   ( new_n34336_, new_n34335_, new_n33925_ );
or   ( new_n34337_, new_n30648_, new_n17601_ );
or   ( new_n34338_, new_n34337_, new_n34336_ );
and  ( new_n34339_, new_n33791_, new_n33786_ );
or   ( new_n34340_, new_n33755_, new_n33754_ );
or   ( new_n34341_, new_n34340_, new_n34339_ );
or   ( new_n34342_, new_n33789_, new_n33754_ );
and  ( new_n34343_, new_n34342_, new_n33753_ );
and  ( new_n34344_, new_n34343_, new_n34341_ );
or   ( new_n34345_, new_n34344_, new_n33751_ );
and  ( new_n34346_, new_n34345_, new_n33750_ );
or   ( new_n34347_, new_n34346_, new_n33909_ );
and  ( new_n34348_, new_n34347_, new_n33913_ );
and  ( new_n34349_, new_n30652_, new_n17598_ );
or   ( new_n34350_, new_n34349_, new_n34348_ );
and  ( new_n34351_, new_n34350_, new_n34338_ );
and  ( new_n34352_, new_n34351_, new_n34326_ );
or   ( new_n34353_, new_n34352_, new_n34293_ );
or   ( new_n34354_, new_n34353_, new_n34282_ );
or   ( new_n34355_, new_n34354_, new_n34037_ );
or   ( new_n34356_, new_n34355_, new_n34030_ );
and  ( new_n34357_, new_n34089_, new_n34058_ );
or   ( new_n34358_, new_n34357_, new_n34056_ );
or   ( new_n34359_, new_n34358_, new_n34054_ );
or   ( new_n34360_, new_n34061_, new_n34054_ );
and  ( new_n34361_, new_n34360_, new_n34049_ );
and  ( new_n34362_, new_n34361_, new_n34359_ );
or   ( new_n34363_, new_n15616_, new_n6463_ );
and  ( new_n34364_, new_n34363_, new_n34362_ );
or   ( new_n34365_, new_n34151_, new_n34118_ );
and  ( new_n34366_, new_n34365_, new_n34119_ );
and  ( new_n34367_, new_n34366_, new_n34115_ );
and  ( new_n34368_, new_n34122_, new_n34115_ );
or   ( new_n34369_, new_n34368_, new_n34110_ );
or   ( new_n34370_, new_n34369_, new_n34367_ );
and  ( new_n34371_, new_n15615_, new_n6464_ );
and  ( new_n34372_, new_n34371_, new_n34370_ );
or   ( new_n34373_, new_n34372_, new_n34364_ );
and  ( new_n34374_, new_n34203_, new_n34200_ );
or   ( new_n34375_, new_n30741_, new_n21656_ );
or   ( new_n34376_, new_n34375_, new_n34374_ );
or   ( new_n34377_, new_n34262_, new_n34259_ );
and  ( new_n34378_, new_n30740_, new_n21657_ );
or   ( new_n34379_, new_n34378_, new_n34377_ );
and  ( new_n34380_, new_n34379_, new_n34376_ );
and  ( new_n34381_, new_n34380_, new_n34373_ );
and  ( new_n34382_, new_n15626_, new_n6903_ );
and  ( new_n34383_, new_n34382_, new_n33689_ );
or   ( new_n34384_, new_n15623_, new_n6906_ );
and  ( new_n34385_, new_n34384_, new_n33741_ );
or   ( new_n34386_, new_n34385_, new_n34383_ );
and  ( new_n34387_, new_n30751_, new_n22098_ );
or   ( new_n34388_, new_n34387_, new_n33794_ );
or   ( new_n34389_, new_n30748_, new_n22101_ );
or   ( new_n34390_, new_n34389_, new_n33846_ );
and  ( new_n34391_, new_n34390_, new_n34388_ );
and  ( new_n34392_, new_n34391_, new_n34386_ );
or   ( new_n34393_, new_n34392_, new_n34381_ );
and  ( new_n34394_, new_n15991_, new_n7854_ );
and  ( new_n34395_, new_n34394_, new_n15317_ );
or   ( new_n34396_, new_n15642_, new_n15318_ );
and  ( new_n34397_, new_n34396_, new_n15990_ );
or   ( new_n34398_, new_n34397_, new_n34395_ );
and  ( new_n34399_, new_n30772_, new_n23012_ );
or   ( new_n34400_, new_n34399_, new_n30445_ );
or   ( new_n34401_, new_n30767_, new_n23017_ );
or   ( new_n34402_, new_n34401_, new_n31114_ );
and  ( new_n34403_, new_n34402_, new_n34400_ );
and  ( new_n34404_, new_n34403_, new_n34398_ );
and  ( new_n34405_, new_n34384_, new_n33689_ );
and  ( new_n34406_, new_n34382_, new_n33741_ );
or   ( new_n34407_, new_n34406_, new_n34405_ );
or   ( new_n34408_, new_n34389_, new_n33794_ );
or   ( new_n34409_, new_n34387_, new_n33846_ );
and  ( new_n34410_, new_n34409_, new_n34408_ );
and  ( new_n34411_, new_n34410_, new_n34407_ );
or   ( new_n34412_, new_n34411_, new_n34404_ );
or   ( new_n34413_, new_n34412_, new_n34393_ );
or   ( new_n34414_, new_n15313_, new_n11175_ );
or   ( new_n34415_, new_n12179_, new_n11175_ );
and  ( new_n34416_, new_n34415_, new_n11170_ );
and  ( new_n34417_, new_n34416_, new_n34414_ );
or   ( new_n34418_, new_n34417_, new_n9592_ );
or   ( new_n34419_, new_n34418_, new_n15320_ );
or   ( new_n34420_, new_n15320_, new_n9589_ );
and  ( new_n34421_, new_n34420_, new_n34419_ );
and  ( new_n34422_, new_n34421_, new_n7858_ );
or   ( new_n34423_, new_n5994_, new_n4381_ );
or   ( new_n34424_, new_n34423_, new_n34422_ );
or   ( new_n34425_, new_n5991_, new_n4381_ );
and  ( new_n34426_, new_n34425_, new_n4373_ );
or   ( new_n34427_, new_n15534_, new_n4374_ );
and  ( new_n34428_, new_n30730_, new_n30699_ );
or   ( new_n34429_, new_n34428_, new_n30696_ );
and  ( new_n34430_, new_n31109_, new_n30857_ );
and  ( new_n34431_, new_n30889_, new_n30857_ );
or   ( new_n34432_, new_n34431_, new_n30853_ );
or   ( new_n34433_, new_n34432_, new_n34430_ );
and  ( new_n34434_, new_n34433_, new_n30815_ );
and  ( new_n34435_, new_n34434_, new_n30774_ );
and  ( new_n34436_, new_n30812_, new_n30774_ );
or   ( new_n34437_, new_n34436_, new_n34435_ );
or   ( new_n34438_, new_n34437_, new_n30771_ );
and  ( new_n34439_, new_n30733_, new_n30699_ );
and  ( new_n34440_, new_n34439_, new_n34438_ );
or   ( new_n34441_, new_n34440_, new_n34429_ );
and  ( new_n34442_, new_n30668_, new_n18242_ );
or   ( new_n34443_, new_n34442_, new_n34441_ );
or   ( new_n34444_, new_n30663_, new_n18247_ );
or   ( new_n34445_, new_n21193_, new_n19620_ );
and  ( new_n34446_, new_n34445_, new_n19617_ );
or   ( new_n34447_, new_n30440_, new_n26326_ );
or   ( new_n34448_, new_n27326_, new_n26326_ );
and  ( new_n34449_, new_n34448_, new_n26322_ );
and  ( new_n34450_, new_n34449_, new_n34447_ );
or   ( new_n34451_, new_n34450_, new_n24747_ );
or   ( new_n34452_, new_n34451_, new_n23019_ );
or   ( new_n34453_, new_n24744_, new_n23019_ );
and  ( new_n34454_, new_n34453_, new_n34452_ );
and  ( new_n34455_, new_n34454_, new_n23016_ );
or   ( new_n34456_, new_n21196_, new_n19620_ );
or   ( new_n34457_, new_n34456_, new_n34455_ );
and  ( new_n34458_, new_n34457_, new_n34446_ );
or   ( new_n34459_, new_n34458_, new_n34444_ );
and  ( new_n34460_, new_n34459_, new_n34443_ );
and  ( new_n34461_, new_n34460_, new_n34427_ );
or   ( new_n34462_, new_n34444_, new_n34441_ );
or   ( new_n34463_, new_n34458_, new_n34442_ );
and  ( new_n34464_, new_n34463_, new_n34462_ );
and  ( new_n34465_, new_n15565_, new_n2968_ );
and  ( new_n34466_, new_n34465_, new_n34464_ );
or   ( new_n34467_, new_n34466_, new_n34461_ );
and  ( new_n34468_, new_n34467_, new_n34426_ );
and  ( new_n34469_, new_n34468_, new_n34424_ );
and  ( new_n34470_, new_n34396_, new_n15317_ );
and  ( new_n34471_, new_n34394_, new_n15990_ );
or   ( new_n34472_, new_n34471_, new_n34470_ );
or   ( new_n34473_, new_n34401_, new_n30445_ );
or   ( new_n34474_, new_n34399_, new_n31114_ );
and  ( new_n34475_, new_n34474_, new_n34473_ );
and  ( new_n34476_, new_n34475_, new_n34472_ );
or   ( new_n34477_, new_n34476_, new_n34469_ );
and  ( new_n34478_, new_n34371_, new_n34362_ );
and  ( new_n34479_, new_n34370_, new_n34363_ );
or   ( new_n34480_, new_n34479_, new_n34478_ );
or   ( new_n34481_, new_n34378_, new_n34374_ );
or   ( new_n34482_, new_n34377_, new_n34375_ );
and  ( new_n34483_, new_n34482_, new_n34481_ );
and  ( new_n34484_, new_n34483_, new_n34480_ );
or   ( new_n34485_, new_n34047_, new_n34045_ );
or   ( new_n34486_, new_n34485_, new_n34362_ );
or   ( new_n34487_, new_n33136_, new_n33132_ );
or   ( new_n34488_, new_n34487_, new_n34038_ );
or   ( new_n34489_, new_n34488_, new_n34486_ );
or   ( new_n34490_, new_n34052_, new_n34045_ );
and  ( new_n34491_, new_n34490_, new_n34040_ );
or   ( new_n34492_, new_n34491_, new_n34488_ );
or   ( new_n34493_, new_n34487_, new_n34043_ );
or   ( new_n34494_, new_n33162_, new_n33132_ );
and  ( new_n34495_, new_n34494_, new_n33158_ );
and  ( new_n34496_, new_n32015_, new_n31978_ );
and  ( new_n34497_, new_n34269_, new_n34222_ );
and  ( new_n34498_, new_n34497_, new_n34377_ );
and  ( new_n34499_, new_n33618_, new_n33615_ );
and  ( new_n34500_, new_n34499_, new_n34268_ );
and  ( new_n34501_, new_n34500_, new_n34498_ );
and  ( new_n34502_, new_n34269_, new_n34265_ );
or   ( new_n34503_, new_n34502_, new_n34273_ );
and  ( new_n34504_, new_n34503_, new_n34500_ );
and  ( new_n34505_, new_n33630_, new_n33615_ );
or   ( new_n34506_, new_n34505_, new_n33626_ );
and  ( new_n34507_, new_n34499_, new_n34276_ );
or   ( new_n34508_, new_n34507_, new_n34506_ );
or   ( new_n34509_, new_n34508_, new_n34504_ );
or   ( new_n34510_, new_n34509_, new_n34501_ );
or   ( new_n34511_, new_n32950_, new_n32922_ );
or   ( new_n34512_, new_n34511_, new_n34510_ );
and  ( new_n34513_, new_n32986_, new_n32720_ );
or   ( new_n34514_, new_n34210_, new_n34160_ );
or   ( new_n34515_, new_n34514_, new_n34374_ );
or   ( new_n34516_, new_n33449_, new_n33446_ );
or   ( new_n34517_, new_n34516_, new_n34209_ );
or   ( new_n34518_, new_n34517_, new_n34515_ );
or   ( new_n34519_, new_n34210_, new_n34206_ );
and  ( new_n34520_, new_n34519_, new_n34214_ );
or   ( new_n34521_, new_n34520_, new_n34517_ );
or   ( new_n34522_, new_n33476_, new_n33446_ );
and  ( new_n34523_, new_n34522_, new_n33472_ );
or   ( new_n34524_, new_n34516_, new_n34217_ );
and  ( new_n34525_, new_n34524_, new_n34523_ );
and  ( new_n34526_, new_n34525_, new_n34521_ );
and  ( new_n34527_, new_n34526_, new_n34518_ );
or   ( new_n34528_, new_n34527_, new_n34513_ );
and  ( new_n34529_, new_n34528_, new_n34512_ );
and  ( new_n34530_, new_n34529_, new_n34496_ );
or   ( new_n34531_, new_n34513_, new_n34510_ );
or   ( new_n34532_, new_n34527_, new_n34511_ );
and  ( new_n34533_, new_n34532_, new_n34531_ );
or   ( new_n34534_, new_n32050_, new_n31804_ );
and  ( new_n34535_, new_n34534_, new_n34533_ );
or   ( new_n34536_, new_n34535_, new_n34530_ );
and  ( new_n34537_, new_n34536_, new_n34495_ );
and  ( new_n34538_, new_n34537_, new_n34493_ );
and  ( new_n34539_, new_n34538_, new_n34492_ );
and  ( new_n34540_, new_n34539_, new_n34489_ );
or   ( new_n34541_, new_n34540_, new_n34484_ );
or   ( new_n34542_, new_n34541_, new_n34477_ );
or   ( new_n34543_, new_n34542_, new_n34413_ );
and  ( new_n34544_, new_n34491_, new_n34486_ );
and  ( new_n34545_, new_n15543_, new_n3317_ );
and  ( new_n34546_, new_n34545_, new_n34544_ );
or   ( new_n34547_, new_n15542_, new_n3316_ );
and  ( new_n34548_, new_n34113_, new_n34106_ );
or   ( new_n34549_, new_n34548_, new_n34101_ );
and  ( new_n34550_, new_n34108_, new_n34106_ );
and  ( new_n34551_, new_n34550_, new_n34370_ );
or   ( new_n34552_, new_n34551_, new_n34549_ );
and  ( new_n34553_, new_n34552_, new_n34547_ );
or   ( new_n34554_, new_n34553_, new_n34546_ );
or   ( new_n34555_, new_n34503_, new_n34498_ );
or   ( new_n34556_, new_n30675_, new_n18589_ );
or   ( new_n34557_, new_n34556_, new_n34555_ );
and  ( new_n34558_, new_n30674_, new_n18588_ );
and  ( new_n34559_, new_n34520_, new_n34515_ );
or   ( new_n34560_, new_n34559_, new_n34558_ );
and  ( new_n34561_, new_n34560_, new_n34557_ );
and  ( new_n34562_, new_n34561_, new_n34554_ );
or   ( new_n34563_, new_n32065_, new_n31897_ );
or   ( new_n34564_, new_n32968_, new_n32935_ );
and  ( new_n34565_, new_n32765_, new_n30670_ );
and  ( new_n34566_, new_n34565_, new_n34440_ );
and  ( new_n34567_, new_n34565_, new_n34429_ );
and  ( new_n34568_, new_n32765_, new_n30667_ );
or   ( new_n34569_, new_n34568_, new_n32929_ );
or   ( new_n34570_, new_n34569_, new_n34567_ );
or   ( new_n34571_, new_n34570_, new_n34566_ );
or   ( new_n34572_, new_n34571_, new_n34564_ );
and  ( new_n34573_, new_n33001_, new_n32845_ );
or   ( new_n34574_, new_n32961_, new_n18249_ );
or   ( new_n34575_, new_n34574_, new_n34457_ );
or   ( new_n34576_, new_n34574_, new_n34446_ );
or   ( new_n34577_, new_n32961_, new_n18246_ );
and  ( new_n34578_, new_n34577_, new_n32994_ );
and  ( new_n34579_, new_n34578_, new_n34576_ );
and  ( new_n34580_, new_n34579_, new_n34575_ );
or   ( new_n34581_, new_n34580_, new_n34573_ );
and  ( new_n34582_, new_n34581_, new_n34572_ );
and  ( new_n34583_, new_n34582_, new_n34563_ );
and  ( new_n34584_, new_n32028_, new_n31991_ );
or   ( new_n34585_, new_n34573_, new_n34571_ );
or   ( new_n34586_, new_n34580_, new_n34564_ );
and  ( new_n34587_, new_n34586_, new_n34585_ );
and  ( new_n34588_, new_n34587_, new_n34584_ );
or   ( new_n34589_, new_n34588_, new_n34583_ );
and  ( new_n34590_, new_n15986_, new_n15732_ );
and  ( new_n34591_, new_n15764_, new_n15732_ );
or   ( new_n34592_, new_n34591_, new_n15727_ );
or   ( new_n34593_, new_n34592_, new_n34590_ );
and  ( new_n34594_, new_n34593_, new_n15689_ );
and  ( new_n34595_, new_n34594_, new_n15993_ );
and  ( new_n34596_, new_n15993_, new_n15686_ );
or   ( new_n34597_, new_n34596_, new_n34595_ );
or   ( new_n34598_, new_n34597_, new_n15646_ );
and  ( new_n34599_, new_n15608_, new_n15572_ );
and  ( new_n34600_, new_n34599_, new_n34598_ );
and  ( new_n34601_, new_n32021_, new_n15567_ );
and  ( new_n34602_, new_n34601_, new_n34600_ );
and  ( new_n34603_, new_n15605_, new_n15572_ );
or   ( new_n34604_, new_n34603_, new_n15564_ );
and  ( new_n34605_, new_n34604_, new_n34601_ );
and  ( new_n34606_, new_n32021_, new_n15538_ );
or   ( new_n34607_, new_n34606_, new_n32058_ );
or   ( new_n34608_, new_n34607_, new_n34605_ );
or   ( new_n34609_, new_n34608_, new_n34602_ );
and  ( new_n34610_, new_n34609_, new_n34589_ );
or   ( new_n34611_, new_n34610_, new_n34562_ );
or   ( new_n34612_, new_n34611_, new_n34543_ );
or   ( new_n34613_, new_n32060_, new_n31968_ );
and  ( new_n34614_, new_n32907_, new_n32885_ );
and  ( new_n34615_, new_n34614_, new_n33616_ );
and  ( new_n34616_, new_n34615_, new_n34499_ );
and  ( new_n34617_, new_n34616_, new_n34278_ );
and  ( new_n34618_, new_n34615_, new_n34506_ );
and  ( new_n34619_, new_n34614_, new_n33624_ );
or   ( new_n34620_, new_n32936_, new_n32931_ );
and  ( new_n34621_, new_n34620_, new_n32907_ );
or   ( new_n34622_, new_n34621_, new_n34619_ );
or   ( new_n34623_, new_n34622_, new_n34618_ );
or   ( new_n34624_, new_n34623_, new_n34617_ );
or   ( new_n34625_, new_n32981_, new_n32932_ );
or   ( new_n34626_, new_n34625_, new_n34624_ );
and  ( new_n34627_, new_n32996_, new_n32916_ );
or   ( new_n34628_, new_n32977_, new_n32972_ );
or   ( new_n34629_, new_n34628_, new_n33447_ );
or   ( new_n34630_, new_n34629_, new_n34516_ );
or   ( new_n34631_, new_n34630_, new_n34219_ );
or   ( new_n34632_, new_n34629_, new_n34523_ );
or   ( new_n34633_, new_n34628_, new_n33470_ );
or   ( new_n34634_, new_n33000_, new_n32977_ );
and  ( new_n34635_, new_n34634_, new_n32997_ );
and  ( new_n34636_, new_n34635_, new_n34633_ );
and  ( new_n34637_, new_n34636_, new_n34632_ );
and  ( new_n34638_, new_n34637_, new_n34631_ );
or   ( new_n34639_, new_n34638_, new_n34627_ );
and  ( new_n34640_, new_n34639_, new_n34626_ );
and  ( new_n34641_, new_n34640_, new_n34613_ );
or   ( new_n34642_, new_n34627_, new_n34624_ );
or   ( new_n34643_, new_n34638_, new_n34625_ );
and  ( new_n34644_, new_n34643_, new_n34642_ );
and  ( new_n34645_, new_n32041_, new_n31988_ );
and  ( new_n34646_, new_n34645_, new_n34644_ );
or   ( new_n34647_, new_n34646_, new_n34641_ );
and  ( new_n34648_, new_n34123_, new_n34116_ );
or   ( new_n34649_, new_n34648_, new_n34114_ );
and  ( new_n34650_, new_n33291_, new_n33289_ );
and  ( new_n34651_, new_n32037_, new_n32032_ );
and  ( new_n34652_, new_n34651_, new_n33292_ );
and  ( new_n34653_, new_n34652_, new_n34650_ );
and  ( new_n34654_, new_n34653_, new_n34107_ );
and  ( new_n34655_, new_n34654_, new_n34649_ );
and  ( new_n34656_, new_n34653_, new_n34105_ );
and  ( new_n34657_, new_n34152_, new_n34116_ );
and  ( new_n34658_, new_n34657_, new_n34654_ );
and  ( new_n34659_, new_n33321_, new_n33291_ );
or   ( new_n34660_, new_n34659_, new_n33312_ );
and  ( new_n34661_, new_n34660_, new_n34652_ );
and  ( new_n34662_, new_n32064_, new_n32037_ );
or   ( new_n34663_, new_n34662_, new_n32061_ );
and  ( new_n34664_, new_n34651_, new_n33315_ );
or   ( new_n34665_, new_n34664_, new_n34663_ );
or   ( new_n34666_, new_n34665_, new_n34661_ );
or   ( new_n34667_, new_n34666_, new_n34658_ );
or   ( new_n34668_, new_n34667_, new_n34656_ );
or   ( new_n34669_, new_n34668_, new_n34655_ );
and  ( new_n34670_, new_n34669_, new_n34647_ );
or   ( new_n34671_, new_n34604_, new_n34600_ );
and  ( new_n34672_, new_n34464_, new_n34427_ );
and  ( new_n34673_, new_n34465_, new_n34460_ );
or   ( new_n34674_, new_n34673_, new_n34672_ );
and  ( new_n34675_, new_n34674_, new_n34671_ );
or   ( new_n34676_, new_n34675_, new_n34670_ );
or   ( new_n34677_, new_n15585_, new_n5151_ );
and  ( new_n34678_, new_n34677_, new_n34305_ );
and  ( new_n34679_, new_n15588_, new_n5148_ );
and  ( new_n34680_, new_n34679_, new_n34322_ );
or   ( new_n34681_, new_n34680_, new_n34678_ );
or   ( new_n34682_, new_n30710_, new_n20373_ );
or   ( new_n34683_, new_n34682_, new_n34344_ );
and  ( new_n34684_, new_n30713_, new_n20370_ );
or   ( new_n34685_, new_n34684_, new_n34332_ );
and  ( new_n34686_, new_n34685_, new_n34683_ );
and  ( new_n34687_, new_n34686_, new_n34681_ );
and  ( new_n34688_, new_n15578_, new_n4763_ );
and  ( new_n34689_, new_n34688_, new_n34093_ );
or   ( new_n34690_, new_n15577_, new_n4762_ );
and  ( new_n34691_, new_n34690_, new_n34155_ );
or   ( new_n34692_, new_n34691_, new_n34689_ );
and  ( new_n34693_, new_n30703_, new_n19994_ );
or   ( new_n34694_, new_n34693_, new_n34208_ );
or   ( new_n34695_, new_n30704_, new_n19995_ );
or   ( new_n34696_, new_n34695_, new_n34267_ );
and  ( new_n34697_, new_n34696_, new_n34694_ );
and  ( new_n34698_, new_n34697_, new_n34692_ );
or   ( new_n34699_, new_n34698_, new_n34687_ );
or   ( new_n34700_, new_n34699_, new_n34676_ );
or   ( new_n34701_, new_n15663_, new_n8766_ );
and  ( new_n34702_, new_n34701_, new_n34303_ );
and  ( new_n34703_, new_n15666_, new_n8763_ );
and  ( new_n34704_, new_n34703_, new_n34320_ );
or   ( new_n34705_, new_n34704_, new_n34702_ );
or   ( new_n34706_, new_n30789_, new_n23923_ );
or   ( new_n34707_, new_n34706_, new_n34339_ );
and  ( new_n34708_, new_n30792_, new_n23920_ );
or   ( new_n34709_, new_n34708_, new_n34327_ );
and  ( new_n34710_, new_n34709_, new_n34707_ );
and  ( new_n34711_, new_n34710_, new_n34705_ );
or   ( new_n34712_, new_n15682_, new_n9590_ );
and  ( new_n34713_, new_n34712_, new_n34417_ );
and  ( new_n34714_, new_n15687_, new_n9585_ );
and  ( new_n34715_, new_n34714_, new_n34593_ );
or   ( new_n34716_, new_n34715_, new_n34713_ );
or   ( new_n34717_, new_n30808_, new_n24745_ );
or   ( new_n34718_, new_n34717_, new_n34450_ );
and  ( new_n34719_, new_n30813_, new_n24740_ );
or   ( new_n34720_, new_n34719_, new_n34433_ );
and  ( new_n34721_, new_n34720_, new_n34718_ );
and  ( new_n34722_, new_n34721_, new_n34716_ );
and  ( new_n34723_, new_n34714_, new_n34417_ );
and  ( new_n34724_, new_n34712_, new_n34593_ );
or   ( new_n34725_, new_n34724_, new_n34723_ );
or   ( new_n34726_, new_n34719_, new_n34450_ );
or   ( new_n34727_, new_n34717_, new_n34433_ );
and  ( new_n34728_, new_n34727_, new_n34726_ );
and  ( new_n34729_, new_n34728_, new_n34725_ );
and  ( new_n34730_, new_n15715_, new_n10786_ );
and  ( new_n34731_, new_n34730_, new_n33949_ );
or   ( new_n34732_, new_n15716_, new_n10785_ );
and  ( new_n34733_, new_n34732_, new_n33971_ );
or   ( new_n34734_, new_n34733_, new_n34731_ );
and  ( new_n34735_, new_n30841_, new_n25937_ );
or   ( new_n34736_, new_n34735_, new_n33993_ );
or   ( new_n34737_, new_n30842_, new_n25936_ );
or   ( new_n34738_, new_n34737_, new_n34013_ );
and  ( new_n34739_, new_n34738_, new_n34736_ );
and  ( new_n34740_, new_n34739_, new_n34734_ );
and  ( new_n34741_, new_n34732_, new_n33949_ );
and  ( new_n34742_, new_n34730_, new_n33971_ );
or   ( new_n34743_, new_n34742_, new_n34741_ );
or   ( new_n34744_, new_n34737_, new_n33993_ );
or   ( new_n34745_, new_n34735_, new_n34013_ );
and  ( new_n34746_, new_n34745_, new_n34744_ );
and  ( new_n34747_, new_n34746_, new_n34743_ );
and  ( new_n34748_, new_n15737_, new_n11530_ );
and  ( new_n34749_, new_n34748_, new_n34087_ );
or   ( new_n34750_, new_n15736_, new_n11529_ );
and  ( new_n34751_, new_n34750_, new_n34149_ );
or   ( new_n34752_, new_n34751_, new_n34749_ );
and  ( new_n34753_, new_n30862_, new_n26677_ );
or   ( new_n34754_, new_n34753_, new_n34188_ );
or   ( new_n34755_, new_n30863_, new_n26678_ );
or   ( new_n34756_, new_n34755_, new_n34247_ );
and  ( new_n34757_, new_n34756_, new_n34754_ );
and  ( new_n34758_, new_n34757_, new_n34752_ );
and  ( new_n34759_, new_n34750_, new_n34087_ );
and  ( new_n34760_, new_n34748_, new_n34149_ );
or   ( new_n34761_, new_n34760_, new_n34759_ );
or   ( new_n34762_, new_n34755_, new_n34188_ );
or   ( new_n34763_, new_n34753_, new_n34247_ );
and  ( new_n34764_, new_n34763_, new_n34762_ );
and  ( new_n34765_, new_n34764_, new_n34761_ );
and  ( new_n34766_, new_n15744_, new_n11660_ );
and  ( new_n34767_, new_n34766_, new_n33677_ );
or   ( new_n34768_, new_n15741_, new_n11663_ );
and  ( new_n34769_, new_n34768_, new_n33729_ );
or   ( new_n34770_, new_n34769_, new_n34767_ );
and  ( new_n34771_, new_n30870_, new_n26808_ );
or   ( new_n34772_, new_n34771_, new_n33780_ );
or   ( new_n34773_, new_n30867_, new_n26811_ );
or   ( new_n34774_, new_n34773_, new_n33832_ );
and  ( new_n34775_, new_n34774_, new_n34772_ );
and  ( new_n34776_, new_n34775_, new_n34770_ );
and  ( new_n34777_, new_n34768_, new_n33677_ );
and  ( new_n34778_, new_n34766_, new_n33729_ );
or   ( new_n34779_, new_n34778_, new_n34777_ );
or   ( new_n34780_, new_n34773_, new_n33780_ );
or   ( new_n34781_, new_n34771_, new_n33832_ );
and  ( new_n34782_, new_n34781_, new_n34780_ );
and  ( new_n34783_, new_n34782_, new_n34779_ );
or   ( new_n34784_, new_n15760_, new_n12180_ );
and  ( new_n34785_, new_n34784_, new_n15312_ );
and  ( new_n34786_, new_n15765_, new_n12175_ );
and  ( new_n34787_, new_n34786_, new_n15985_ );
or   ( new_n34788_, new_n34787_, new_n34785_ );
or   ( new_n34789_, new_n30885_, new_n27327_ );
or   ( new_n34790_, new_n34789_, new_n30439_ );
and  ( new_n34791_, new_n30890_, new_n27322_ );
or   ( new_n34792_, new_n34791_, new_n31108_ );
and  ( new_n34793_, new_n34792_, new_n34790_ );
and  ( new_n34794_, new_n34793_, new_n34788_ );
and  ( new_n34795_, new_n34786_, new_n15312_ );
and  ( new_n34796_, new_n34784_, new_n15985_ );
or   ( new_n34797_, new_n34796_, new_n34795_ );
or   ( new_n34798_, new_n34791_, new_n30439_ );
or   ( new_n34799_, new_n34789_, new_n31108_ );
and  ( new_n34800_, new_n34799_, new_n34798_ );
and  ( new_n34801_, new_n34800_, new_n34797_ );
and  ( new_n34802_, new_n15774_, new_n15302_ );
and  ( new_n34803_, new_n34802_, new_n34083_ );
or   ( new_n34804_, new_n15975_, new_n12466_ );
and  ( new_n34805_, new_n34804_, new_n34144_ );
or   ( new_n34806_, new_n34805_, new_n34803_ );
and  ( new_n34807_, new_n30899_, new_n30429_ );
or   ( new_n34808_, new_n34807_, new_n34184_ );
or   ( new_n34809_, new_n31098_, new_n27611_ );
or   ( new_n34810_, new_n34809_, new_n34243_ );
and  ( new_n34811_, new_n34810_, new_n34808_ );
and  ( new_n34812_, new_n34811_, new_n34806_ );
and  ( new_n34813_, new_n34804_, new_n34083_ );
and  ( new_n34814_, new_n34802_, new_n34144_ );
or   ( new_n34815_, new_n34814_, new_n34813_ );
or   ( new_n34816_, new_n34809_, new_n34184_ );
or   ( new_n34817_, new_n34807_, new_n34243_ );
and  ( new_n34818_, new_n34817_, new_n34816_ );
and  ( new_n34819_, new_n34818_, new_n34815_ );
or   ( new_n34820_, new_n15976_, new_n12732_ );
and  ( new_n34821_, new_n34820_, new_n33672_ );
and  ( new_n34822_, new_n15781_, new_n15303_ );
and  ( new_n34823_, new_n34822_, new_n33724_ );
or   ( new_n34824_, new_n34823_, new_n34821_ );
or   ( new_n34825_, new_n31099_, new_n27876_ );
or   ( new_n34826_, new_n34825_, new_n33775_ );
and  ( new_n34827_, new_n30906_, new_n30430_ );
or   ( new_n34828_, new_n34827_, new_n33827_ );
and  ( new_n34829_, new_n34828_, new_n34826_ );
and  ( new_n34830_, new_n34829_, new_n34824_ );
and  ( new_n34831_, new_n34822_, new_n33672_ );
and  ( new_n34832_, new_n34820_, new_n33724_ );
or   ( new_n34833_, new_n34832_, new_n34831_ );
or   ( new_n34834_, new_n34827_, new_n33775_ );
or   ( new_n34835_, new_n34825_, new_n33827_ );
and  ( new_n34836_, new_n34835_, new_n34834_ );
and  ( new_n34837_, new_n34836_, new_n34833_ );
or   ( new_n34838_, new_n15980_, new_n13259_ );
and  ( new_n34839_, new_n34838_, new_n15299_ );
and  ( new_n34840_, new_n15796_, new_n15307_ );
and  ( new_n34841_, new_n34840_, new_n15972_ );
or   ( new_n34842_, new_n34841_, new_n34839_ );
or   ( new_n34843_, new_n31103_, new_n28401_ );
or   ( new_n34844_, new_n34843_, new_n30426_ );
and  ( new_n34845_, new_n30921_, new_n30434_ );
or   ( new_n34846_, new_n34845_, new_n31095_ );
and  ( new_n34847_, new_n34846_, new_n34844_ );
and  ( new_n34848_, new_n34847_, new_n34842_ );
and  ( new_n34849_, new_n34840_, new_n15299_ );
and  ( new_n34850_, new_n34838_, new_n15972_ );
or   ( new_n34851_, new_n34850_, new_n34849_ );
or   ( new_n34852_, new_n34845_, new_n30426_ );
or   ( new_n34853_, new_n34843_, new_n31095_ );
and  ( new_n34854_, new_n34853_, new_n34852_ );
and  ( new_n34855_, new_n34854_, new_n34851_ );
and  ( new_n34856_, new_n15804_, new_n15289_ );
and  ( new_n34857_, new_n34856_, new_n34078_ );
or   ( new_n34858_, new_n15962_, new_n13509_ );
and  ( new_n34859_, new_n34858_, new_n34139_ );
or   ( new_n34860_, new_n34859_, new_n34857_ );
and  ( new_n34861_, new_n30929_, new_n30416_ );
or   ( new_n34862_, new_n34861_, new_n34179_ );
or   ( new_n34863_, new_n31085_, new_n28651_ );
or   ( new_n34864_, new_n34863_, new_n34238_ );
and  ( new_n34865_, new_n34864_, new_n34862_ );
and  ( new_n34866_, new_n34865_, new_n34860_ );
and  ( new_n34867_, new_n34858_, new_n34078_ );
and  ( new_n34868_, new_n34856_, new_n34139_ );
or   ( new_n34869_, new_n34868_, new_n34867_ );
or   ( new_n34870_, new_n34863_, new_n34179_ );
or   ( new_n34871_, new_n34861_, new_n34238_ );
and  ( new_n34872_, new_n34871_, new_n34870_ );
and  ( new_n34873_, new_n34872_, new_n34869_ );
or   ( new_n34874_, new_n15963_, new_n13740_ );
and  ( new_n34875_, new_n34874_, new_n33667_ );
and  ( new_n34876_, new_n15808_, new_n15290_ );
and  ( new_n34877_, new_n34876_, new_n33719_ );
or   ( new_n34878_, new_n34877_, new_n34875_ );
or   ( new_n34879_, new_n31086_, new_n28881_ );
or   ( new_n34880_, new_n34879_, new_n33770_ );
and  ( new_n34881_, new_n30934_, new_n30417_ );
or   ( new_n34882_, new_n34881_, new_n33822_ );
and  ( new_n34883_, new_n34882_, new_n34880_ );
and  ( new_n34884_, new_n34883_, new_n34878_ );
and  ( new_n34885_, new_n34876_, new_n33667_ );
and  ( new_n34886_, new_n34874_, new_n33719_ );
or   ( new_n34887_, new_n34886_, new_n34885_ );
or   ( new_n34888_, new_n34881_, new_n33770_ );
or   ( new_n34889_, new_n34879_, new_n33822_ );
and  ( new_n34890_, new_n34889_, new_n34888_ );
and  ( new_n34891_, new_n34890_, new_n34887_ );
or   ( new_n34892_, new_n15966_, new_n13959_ );
and  ( new_n34893_, new_n34892_, new_n33091_ );
and  ( new_n34894_, new_n15820_, new_n15293_ );
and  ( new_n34895_, new_n34894_, new_n33247_ );
or   ( new_n34896_, new_n34895_, new_n34893_ );
or   ( new_n34897_, new_n31089_, new_n29099_ );
or   ( new_n34898_, new_n34897_, new_n33405_ );
and  ( new_n34899_, new_n30945_, new_n30420_ );
or   ( new_n34900_, new_n34899_, new_n33531_ );
and  ( new_n34901_, new_n34900_, new_n34898_ );
and  ( new_n34902_, new_n34901_, new_n34896_ );
and  ( new_n34903_, new_n34894_, new_n33091_ );
and  ( new_n34904_, new_n34892_, new_n33247_ );
or   ( new_n34905_, new_n34904_, new_n34903_ );
or   ( new_n34906_, new_n34899_, new_n33405_ );
or   ( new_n34907_, new_n34897_, new_n33531_ );
and  ( new_n34908_, new_n34907_, new_n34906_ );
and  ( new_n34909_, new_n34908_, new_n34905_ );
or   ( new_n34910_, new_n15967_, new_n13948_ );
and  ( new_n34911_, new_n34910_, new_n15286_ );
and  ( new_n34912_, new_n15816_, new_n15294_ );
and  ( new_n34913_, new_n34912_, new_n15959_ );
or   ( new_n34914_, new_n34913_, new_n34911_ );
or   ( new_n34915_, new_n31090_, new_n29088_ );
or   ( new_n34916_, new_n34915_, new_n30413_ );
and  ( new_n34917_, new_n30941_, new_n30421_ );
or   ( new_n34918_, new_n34917_, new_n31082_ );
and  ( new_n34919_, new_n34918_, new_n34916_ );
and  ( new_n34920_, new_n34919_, new_n34914_ );
and  ( new_n34921_, new_n34912_, new_n15286_ );
and  ( new_n34922_, new_n34910_, new_n15959_ );
or   ( new_n34923_, new_n34922_, new_n34921_ );
or   ( new_n34924_, new_n34917_, new_n30413_ );
or   ( new_n34925_, new_n34915_, new_n31082_ );
and  ( new_n34926_, new_n34925_, new_n34924_ );
and  ( new_n34927_, new_n34926_, new_n34923_ );
and  ( new_n34928_, new_n15828_, new_n15276_ );
and  ( new_n34929_, new_n34928_, new_n34073_ );
or   ( new_n34930_, new_n15949_, new_n14119_ );
and  ( new_n34931_, new_n34930_, new_n34134_ );
or   ( new_n34932_, new_n34931_, new_n34929_ );
and  ( new_n34933_, new_n30953_, new_n30403_ );
or   ( new_n34934_, new_n34933_, new_n34174_ );
or   ( new_n34935_, new_n31072_, new_n29258_ );
or   ( new_n34936_, new_n34935_, new_n34233_ );
and  ( new_n34937_, new_n34936_, new_n34934_ );
and  ( new_n34938_, new_n34937_, new_n34932_ );
and  ( new_n34939_, new_n34930_, new_n34073_ );
and  ( new_n34940_, new_n34928_, new_n34134_ );
or   ( new_n34941_, new_n34940_, new_n34939_ );
or   ( new_n34942_, new_n34935_, new_n34174_ );
or   ( new_n34943_, new_n34933_, new_n34233_ );
and  ( new_n34944_, new_n34943_, new_n34942_ );
and  ( new_n34945_, new_n34944_, new_n34941_ );
and  ( new_n34946_, new_n15835_, new_n15277_ );
and  ( new_n34947_, new_n34946_, new_n33662_ );
or   ( new_n34948_, new_n15950_, new_n14309_ );
and  ( new_n34949_, new_n34948_, new_n33714_ );
or   ( new_n34950_, new_n34949_, new_n34947_ );
and  ( new_n34951_, new_n30960_, new_n30404_ );
or   ( new_n34952_, new_n34951_, new_n33765_ );
or   ( new_n34953_, new_n31073_, new_n29446_ );
or   ( new_n34954_, new_n34953_, new_n33817_ );
and  ( new_n34955_, new_n34954_, new_n34952_ );
and  ( new_n34956_, new_n34955_, new_n34950_ );
and  ( new_n34957_, new_n34948_, new_n33662_ );
and  ( new_n34958_, new_n34946_, new_n33714_ );
or   ( new_n34959_, new_n34958_, new_n34957_ );
or   ( new_n34960_, new_n34953_, new_n33765_ );
or   ( new_n34961_, new_n34951_, new_n33817_ );
and  ( new_n34962_, new_n34961_, new_n34960_ );
and  ( new_n34963_, new_n34962_, new_n34959_ );
or   ( new_n34964_, new_n15953_, new_n14605_ );
and  ( new_n34965_, new_n34964_, new_n33082_ );
and  ( new_n34966_, new_n15847_, new_n15280_ );
and  ( new_n34967_, new_n34966_, new_n33238_ );
or   ( new_n34968_, new_n34967_, new_n34965_ );
or   ( new_n34969_, new_n31076_, new_n29740_ );
or   ( new_n34970_, new_n34969_, new_n33396_ );
and  ( new_n34971_, new_n30973_, new_n30407_ );
or   ( new_n34972_, new_n34971_, new_n33522_ );
and  ( new_n34973_, new_n34972_, new_n34970_ );
and  ( new_n34974_, new_n34973_, new_n34968_ );
and  ( new_n34975_, new_n34966_, new_n33082_ );
and  ( new_n34976_, new_n34964_, new_n33238_ );
or   ( new_n34977_, new_n34976_, new_n34975_ );
or   ( new_n34978_, new_n34971_, new_n33396_ );
or   ( new_n34979_, new_n34969_, new_n33522_ );
and  ( new_n34980_, new_n34979_, new_n34978_ );
and  ( new_n34981_, new_n34980_, new_n34977_ );
or   ( new_n34982_, new_n15954_, new_n14587_ );
and  ( new_n34983_, new_n34982_, new_n15273_ );
and  ( new_n34984_, new_n15840_, new_n15281_ );
and  ( new_n34985_, new_n34984_, new_n15946_ );
or   ( new_n34986_, new_n34985_, new_n34983_ );
or   ( new_n34987_, new_n31077_, new_n29721_ );
or   ( new_n34988_, new_n34987_, new_n30400_ );
and  ( new_n34989_, new_n30966_, new_n30408_ );
or   ( new_n34990_, new_n34989_, new_n31069_ );
and  ( new_n34991_, new_n34990_, new_n34988_ );
and  ( new_n34992_, new_n34991_, new_n34986_ );
and  ( new_n34993_, new_n34984_, new_n15273_ );
and  ( new_n34994_, new_n34982_, new_n15946_ );
or   ( new_n34995_, new_n34994_, new_n34993_ );
or   ( new_n34996_, new_n34989_, new_n30400_ );
or   ( new_n34997_, new_n34987_, new_n31069_ );
and  ( new_n34998_, new_n34997_, new_n34996_ );
and  ( new_n34999_, new_n34998_, new_n34995_ );
and  ( new_n35000_, new_n15852_, new_n15263_ );
and  ( new_n35001_, new_n35000_, new_n34068_ );
or   ( new_n35002_, new_n15936_, new_n14744_ );
and  ( new_n35003_, new_n35002_, new_n34129_ );
or   ( new_n35004_, new_n35003_, new_n35001_ );
or   ( new_n35005_, new_n31059_, new_n29878_ );
or   ( new_n35006_, new_n35005_, new_n34228_ );
and  ( new_n35007_, new_n30978_, new_n30390_ );
or   ( new_n35008_, new_n35007_, new_n34169_ );
and  ( new_n35009_, new_n35008_, new_n35006_ );
and  ( new_n35010_, new_n35009_, new_n35004_ );
and  ( new_n35011_, new_n35002_, new_n34068_ );
and  ( new_n35012_, new_n35000_, new_n34129_ );
or   ( new_n35013_, new_n35012_, new_n35011_ );
or   ( new_n35014_, new_n35007_, new_n34228_ );
or   ( new_n35015_, new_n35005_, new_n34169_ );
and  ( new_n35016_, new_n35015_, new_n35014_ );
and  ( new_n35017_, new_n35016_, new_n35013_ );
and  ( new_n35018_, new_n15856_, new_n15264_ );
and  ( new_n35019_, new_n35018_, new_n33657_ );
or   ( new_n35020_, new_n15937_, new_n14810_ );
and  ( new_n35021_, new_n35020_, new_n33709_ );
or   ( new_n35022_, new_n35021_, new_n35019_ );
or   ( new_n35023_, new_n31060_, new_n29944_ );
or   ( new_n35024_, new_n35023_, new_n33812_ );
and  ( new_n35025_, new_n30982_, new_n30391_ );
or   ( new_n35026_, new_n35025_, new_n33760_ );
and  ( new_n35027_, new_n35026_, new_n35024_ );
and  ( new_n35028_, new_n35027_, new_n35022_ );
and  ( new_n35029_, new_n35020_, new_n33657_ );
and  ( new_n35030_, new_n35018_, new_n33709_ );
or   ( new_n35031_, new_n35030_, new_n35029_ );
or   ( new_n35032_, new_n35025_, new_n33812_ );
or   ( new_n35033_, new_n35023_, new_n33760_ );
and  ( new_n35034_, new_n35033_, new_n35032_ );
and  ( new_n35035_, new_n35034_, new_n35031_ );
and  ( new_n35036_, new_n15868_, new_n15267_ );
and  ( new_n35037_, new_n35036_, new_n33073_ );
or   ( new_n35038_, new_n15940_, new_n14979_ );
and  ( new_n35039_, new_n35038_, new_n33229_ );
or   ( new_n35040_, new_n35039_, new_n35037_ );
or   ( new_n35041_, new_n31063_, new_n30111_ );
or   ( new_n35042_, new_n35041_, new_n33513_ );
and  ( new_n35043_, new_n30994_, new_n30394_ );
or   ( new_n35044_, new_n35043_, new_n33387_ );
and  ( new_n35045_, new_n35044_, new_n35042_ );
and  ( new_n35046_, new_n35045_, new_n35040_ );
and  ( new_n35047_, new_n35038_, new_n33073_ );
and  ( new_n35048_, new_n35036_, new_n33229_ );
or   ( new_n35049_, new_n35048_, new_n35047_ );
or   ( new_n35050_, new_n35043_, new_n33513_ );
or   ( new_n35051_, new_n35041_, new_n33387_ );
and  ( new_n35052_, new_n35051_, new_n35050_ );
and  ( new_n35053_, new_n35052_, new_n35049_ );
and  ( new_n35054_, new_n15861_, new_n15268_ );
and  ( new_n35055_, new_n35054_, new_n15260_ );
or   ( new_n35056_, new_n15941_, new_n14966_ );
and  ( new_n35057_, new_n35056_, new_n15933_ );
or   ( new_n35058_, new_n35057_, new_n35055_ );
or   ( new_n35059_, new_n31064_, new_n30098_ );
or   ( new_n35060_, new_n35059_, new_n31056_ );
and  ( new_n35061_, new_n30988_, new_n30395_ );
or   ( new_n35062_, new_n35061_, new_n30387_ );
and  ( new_n35063_, new_n35062_, new_n35060_ );
and  ( new_n35064_, new_n35063_, new_n35058_ );
and  ( new_n35065_, new_n35056_, new_n15260_ );
and  ( new_n35066_, new_n35054_, new_n15933_ );
or   ( new_n35067_, new_n35066_, new_n35065_ );
or   ( new_n35068_, new_n35061_, new_n31056_ );
or   ( new_n35069_, new_n35059_, new_n30387_ );
and  ( new_n35070_, new_n35069_, new_n35068_ );
and  ( new_n35071_, new_n35070_, new_n35067_ );
or   ( new_n35072_, new_n31000_, new_n30159_ );
or   ( new_n35073_, new_n35072_, new_n34164_ );
and  ( new_n35074_, new_n30999_, new_n30158_ );
or   ( new_n35075_, new_n35074_, new_n34223_ );
and  ( new_n35076_, new_n35075_, new_n35073_ );
and  ( new_n35077_, new_n35076_, new_n34124_ );
or   ( new_n35078_, new_n35074_, new_n34164_ );
or   ( new_n35079_, new_n35072_, new_n34223_ );
and  ( new_n35080_, new_n35079_, new_n35078_ );
and  ( new_n35081_, new_n35080_, new_n34063_ );
or   ( new_n35082_, new_n35081_, new_n35077_ );
and  ( new_n35083_, new_n35082_, new_n15027_ );
and  ( new_n35084_, new_n35083_, new_n15874_ );
or   ( new_n35085_, new_n15873_, new_n15026_ );
and  ( new_n35086_, new_n35080_, new_n34124_ );
and  ( new_n35087_, new_n35076_, new_n34063_ );
or   ( new_n35088_, new_n35087_, new_n35086_ );
and  ( new_n35089_, new_n35088_, new_n35085_ );
or   ( new_n35090_, new_n15881_, new_n15084_ );
and  ( new_n35091_, new_n35090_, new_n15258_ );
and  ( new_n35092_, new_n15884_, new_n15081_ );
and  ( new_n35093_, new_n35092_, new_n15931_ );
or   ( new_n35094_, new_n35093_, new_n35091_ );
and  ( new_n35095_, new_n31009_, new_n30213_ );
or   ( new_n35096_, new_n35095_, new_n31054_ );
or   ( new_n35097_, new_n31006_, new_n30216_ );
or   ( new_n35098_, new_n35097_, new_n30385_ );
and  ( new_n35099_, new_n35098_, new_n35096_ );
and  ( new_n35100_, new_n35099_, new_n35094_ );
and  ( new_n35101_, new_n35092_, new_n15258_ );
and  ( new_n35102_, new_n35090_, new_n15931_ );
or   ( new_n35103_, new_n35102_, new_n35101_ );
or   ( new_n35104_, new_n35097_, new_n31054_ );
or   ( new_n35105_, new_n35095_, new_n30385_ );
and  ( new_n35106_, new_n35105_, new_n35104_ );
and  ( new_n35107_, new_n35106_, new_n35103_ );
and  ( new_n35108_, new_n15889_, new_n15144_ );
and  ( new_n35109_, new_n35108_, new_n33063_ );
or   ( new_n35110_, new_n15927_, new_n15143_ );
and  ( new_n35111_, new_n35110_, new_n33219_ );
or   ( new_n35112_, new_n35111_, new_n35109_ );
or   ( new_n35113_, new_n31016_, new_n30367_ );
or   ( new_n35114_, new_n35113_, new_n33503_ );
and  ( new_n35115_, new_n31015_, new_n30381_ );
or   ( new_n35116_, new_n35115_, new_n33377_ );
and  ( new_n35117_, new_n35116_, new_n35114_ );
and  ( new_n35118_, new_n35117_, new_n35112_ );
and  ( new_n35119_, new_n35110_, new_n33063_ );
and  ( new_n35120_, new_n35108_, new_n33219_ );
or   ( new_n35121_, new_n35120_, new_n35119_ );
or   ( new_n35122_, new_n35115_, new_n33503_ );
or   ( new_n35123_, new_n35113_, new_n33377_ );
and  ( new_n35124_, new_n35123_, new_n35122_ );
and  ( new_n35125_, new_n35124_, new_n35121_ );
and  ( new_n35126_, new_n15893_, new_n15174_ );
or   ( new_n35127_, new_n15255_, new_n15206_ );
and  ( new_n35128_, new_n35127_, new_n35126_ );
or   ( new_n35129_, new_n15928_, new_n15177_ );
and  ( new_n35130_, new_n35129_, new_n15924_ );
or   ( new_n35131_, new_n35130_, new_n35128_ );
or   ( new_n35132_, new_n31020_, new_n30378_ );
and  ( new_n35133_, new_n31050_, new_n31048_ );
or   ( new_n35134_, new_n35133_, new_n35132_ );
and  ( new_n35135_, new_n31049_, new_n30382_ );
or   ( new_n35136_, new_n35135_, new_n30329_ );
and  ( new_n35137_, new_n35136_, new_n35134_ );
and  ( new_n35138_, new_n35137_, new_n35131_ );
and  ( new_n35139_, new_n35129_, new_n35127_ );
and  ( new_n35140_, new_n35126_, new_n15924_ );
or   ( new_n35141_, new_n35140_, new_n35139_ );
or   ( new_n35142_, new_n35135_, new_n35133_ );
or   ( new_n35143_, new_n35132_, new_n30329_ );
and  ( new_n35144_, new_n35143_, new_n35142_ );
and  ( new_n35145_, new_n35144_, new_n35141_ );
or   ( new_n35146_, new_n35145_, new_n35138_ );
or   ( new_n35147_, new_n35146_, new_n35125_ );
or   ( new_n35148_, new_n35147_, new_n35118_ );
or   ( new_n35149_, new_n35148_, new_n35107_ );
or   ( new_n35150_, new_n35149_, new_n35100_ );
or   ( new_n35151_, new_n35150_, new_n35089_ );
or   ( new_n35152_, new_n35151_, new_n35084_ );
or   ( new_n35153_, new_n35152_, new_n35071_ );
or   ( new_n35154_, new_n35153_, new_n35064_ );
or   ( new_n35155_, new_n35154_, new_n35053_ );
or   ( new_n35156_, new_n35155_, new_n35046_ );
or   ( new_n35157_, new_n35156_, new_n35035_ );
or   ( new_n35158_, new_n35157_, new_n35028_ );
or   ( new_n35159_, new_n35158_, new_n35017_ );
or   ( new_n35160_, new_n35159_, new_n35010_ );
or   ( new_n35161_, new_n35160_, new_n34999_ );
or   ( new_n35162_, new_n35161_, new_n34992_ );
or   ( new_n35163_, new_n35162_, new_n34981_ );
or   ( new_n35164_, new_n35163_, new_n34974_ );
or   ( new_n35165_, new_n35164_, new_n34963_ );
or   ( new_n35166_, new_n35165_, new_n34956_ );
or   ( new_n35167_, new_n35166_, new_n34945_ );
or   ( new_n35168_, new_n35167_, new_n34938_ );
or   ( new_n35169_, new_n35168_, new_n34927_ );
or   ( new_n35170_, new_n35169_, new_n34920_ );
or   ( new_n35171_, new_n35170_, new_n34909_ );
or   ( new_n35172_, new_n35171_, new_n34902_ );
or   ( new_n35173_, new_n35172_, new_n34891_ );
or   ( new_n35174_, new_n35173_, new_n34884_ );
or   ( new_n35175_, new_n35174_, new_n34873_ );
or   ( new_n35176_, new_n35175_, new_n34866_ );
or   ( new_n35177_, new_n35176_, new_n34855_ );
or   ( new_n35178_, new_n35177_, new_n34848_ );
or   ( new_n35179_, new_n15979_, new_n12985_ );
and  ( new_n35180_, new_n35179_, new_n33944_ );
and  ( new_n35181_, new_n15789_, new_n15306_ );
and  ( new_n35182_, new_n35181_, new_n33966_ );
or   ( new_n35183_, new_n35182_, new_n35180_ );
or   ( new_n35184_, new_n31102_, new_n28130_ );
or   ( new_n35185_, new_n35184_, new_n33988_ );
and  ( new_n35186_, new_n30914_, new_n30433_ );
or   ( new_n35187_, new_n35186_, new_n34008_ );
and  ( new_n35188_, new_n35187_, new_n35185_ );
and  ( new_n35189_, new_n35188_, new_n35183_ );
and  ( new_n35190_, new_n35181_, new_n33944_ );
and  ( new_n35191_, new_n35179_, new_n33966_ );
or   ( new_n35192_, new_n35191_, new_n35190_ );
or   ( new_n35193_, new_n35186_, new_n33988_ );
or   ( new_n35194_, new_n35184_, new_n34008_ );
and  ( new_n35195_, new_n35194_, new_n35193_ );
and  ( new_n35196_, new_n35195_, new_n35192_ );
or   ( new_n35197_, new_n35196_, new_n35189_ );
or   ( new_n35198_, new_n35197_, new_n35178_ );
or   ( new_n35199_, new_n35198_, new_n34837_ );
or   ( new_n35200_, new_n35199_, new_n34830_ );
or   ( new_n35201_, new_n35200_, new_n34819_ );
or   ( new_n35202_, new_n35201_, new_n34812_ );
or   ( new_n35203_, new_n35202_, new_n34801_ );
or   ( new_n35204_, new_n35203_, new_n34794_ );
or   ( new_n35205_, new_n15752_, new_n11857_ );
and  ( new_n35206_, new_n35205_, new_n33108_ );
and  ( new_n35207_, new_n15753_, new_n11858_ );
and  ( new_n35208_, new_n35207_, new_n33264_ );
or   ( new_n35209_, new_n35208_, new_n35206_ );
or   ( new_n35210_, new_n30878_, new_n27007_ );
or   ( new_n35211_, new_n35210_, new_n33422_ );
and  ( new_n35212_, new_n30877_, new_n27006_ );
or   ( new_n35213_, new_n35212_, new_n33548_ );
and  ( new_n35214_, new_n35213_, new_n35211_ );
and  ( new_n35215_, new_n35214_, new_n35209_ );
and  ( new_n35216_, new_n35207_, new_n33108_ );
and  ( new_n35217_, new_n35205_, new_n33264_ );
or   ( new_n35218_, new_n35217_, new_n35216_ );
or   ( new_n35219_, new_n35212_, new_n33422_ );
or   ( new_n35220_, new_n35210_, new_n33548_ );
and  ( new_n35221_, new_n35220_, new_n35219_ );
and  ( new_n35222_, new_n35221_, new_n35218_ );
or   ( new_n35223_, new_n35222_, new_n35215_ );
or   ( new_n35224_, new_n35223_, new_n35204_ );
or   ( new_n35225_, new_n35224_, new_n34783_ );
or   ( new_n35226_, new_n35225_, new_n34776_ );
or   ( new_n35227_, new_n35226_, new_n34765_ );
or   ( new_n35228_, new_n35227_, new_n34758_ );
and  ( new_n35229_, new_n15730_, new_n11166_ );
and  ( new_n35230_, new_n35229_, new_n15314_ );
or   ( new_n35231_, new_n15723_, new_n11173_ );
and  ( new_n35232_, new_n35231_, new_n15987_ );
or   ( new_n35233_, new_n35232_, new_n35230_ );
and  ( new_n35234_, new_n30855_, new_n26318_ );
or   ( new_n35235_, new_n35234_, new_n30441_ );
or   ( new_n35236_, new_n30849_, new_n26324_ );
or   ( new_n35237_, new_n35236_, new_n31110_ );
and  ( new_n35238_, new_n35237_, new_n35235_ );
and  ( new_n35239_, new_n35238_, new_n35233_ );
and  ( new_n35240_, new_n35231_, new_n15314_ );
and  ( new_n35241_, new_n35229_, new_n15987_ );
or   ( new_n35242_, new_n35241_, new_n35240_ );
or   ( new_n35243_, new_n35236_, new_n30441_ );
or   ( new_n35244_, new_n35234_, new_n31110_ );
and  ( new_n35245_, new_n35244_, new_n35243_ );
and  ( new_n35246_, new_n35245_, new_n35242_ );
or   ( new_n35247_, new_n35246_, new_n35239_ );
or   ( new_n35248_, new_n35247_, new_n35228_ );
or   ( new_n35249_, new_n35248_, new_n34747_ );
or   ( new_n35250_, new_n35249_, new_n34740_ );
or   ( new_n35251_, new_n15704_, new_n10382_ );
and  ( new_n35252_, new_n35251_, new_n33680_ );
and  ( new_n35253_, new_n15707_, new_n10379_ );
and  ( new_n35254_, new_n35253_, new_n33732_ );
or   ( new_n35255_, new_n35254_, new_n35252_ );
or   ( new_n35256_, new_n30830_, new_n25536_ );
or   ( new_n35257_, new_n35256_, new_n33785_ );
and  ( new_n35258_, new_n30833_, new_n25533_ );
or   ( new_n35259_, new_n35258_, new_n33837_ );
and  ( new_n35260_, new_n35259_, new_n35257_ );
and  ( new_n35261_, new_n35260_, new_n35255_ );
and  ( new_n35262_, new_n35253_, new_n33680_ );
and  ( new_n35263_, new_n35251_, new_n33732_ );
or   ( new_n35264_, new_n35263_, new_n35262_ );
or   ( new_n35265_, new_n35258_, new_n33785_ );
or   ( new_n35266_, new_n35256_, new_n33837_ );
and  ( new_n35267_, new_n35266_, new_n35265_ );
and  ( new_n35268_, new_n35267_, new_n35264_ );
or   ( new_n35269_, new_n35268_, new_n35261_ );
or   ( new_n35270_, new_n35269_, new_n35250_ );
or   ( new_n35271_, new_n15697_, new_n9998_ );
and  ( new_n35272_, new_n35271_, new_n34357_ );
and  ( new_n35273_, new_n15696_, new_n9999_ );
and  ( new_n35274_, new_n35273_, new_n34365_ );
or   ( new_n35275_, new_n35274_, new_n35272_ );
or   ( new_n35276_, new_n30823_, new_n25151_ );
or   ( new_n35277_, new_n35276_, new_n34193_ );
and  ( new_n35278_, new_n30822_, new_n25152_ );
or   ( new_n35279_, new_n35278_, new_n34252_ );
and  ( new_n35280_, new_n35279_, new_n35277_ );
and  ( new_n35281_, new_n35280_, new_n35275_ );
and  ( new_n35282_, new_n35273_, new_n34357_ );
and  ( new_n35283_, new_n35271_, new_n34365_ );
or   ( new_n35284_, new_n35283_, new_n35282_ );
or   ( new_n35285_, new_n35278_, new_n34193_ );
or   ( new_n35286_, new_n35276_, new_n34252_ );
and  ( new_n35287_, new_n35286_, new_n35285_ );
and  ( new_n35288_, new_n35287_, new_n35284_ );
or   ( new_n35289_, new_n35288_, new_n35281_ );
or   ( new_n35290_, new_n35289_, new_n35270_ );
or   ( new_n35291_, new_n35290_, new_n34729_ );
or   ( new_n35292_, new_n35291_, new_n34722_ );
or   ( new_n35293_, new_n15675_, new_n9205_ );
and  ( new_n35294_, new_n35293_, new_n33112_ );
and  ( new_n35295_, new_n15674_, new_n9206_ );
and  ( new_n35296_, new_n35295_, new_n33268_ );
or   ( new_n35297_, new_n35296_, new_n35294_ );
or   ( new_n35298_, new_n30801_, new_n24360_ );
or   ( new_n35299_, new_n35298_, new_n33426_ );
and  ( new_n35300_, new_n30800_, new_n24361_ );
or   ( new_n35301_, new_n35300_, new_n33568_ );
and  ( new_n35302_, new_n35301_, new_n35299_ );
and  ( new_n35303_, new_n35302_, new_n35297_ );
and  ( new_n35304_, new_n35295_, new_n33112_ );
and  ( new_n35305_, new_n35293_, new_n33268_ );
or   ( new_n35306_, new_n35305_, new_n35304_ );
or   ( new_n35307_, new_n35300_, new_n33426_ );
or   ( new_n35308_, new_n35298_, new_n33568_ );
and  ( new_n35309_, new_n35308_, new_n35307_ );
and  ( new_n35310_, new_n35309_, new_n35306_ );
or   ( new_n35311_, new_n35310_, new_n35303_ );
or   ( new_n35312_, new_n35311_, new_n35292_ );
or   ( new_n35313_, new_n35312_, new_n34711_ );
and  ( new_n35314_, new_n15655_, new_n8294_ );
and  ( new_n35315_, new_n35314_, new_n34091_ );
or   ( new_n35316_, new_n15656_, new_n8293_ );
and  ( new_n35317_, new_n35316_, new_n34153_ );
or   ( new_n35318_, new_n35317_, new_n35315_ );
and  ( new_n35319_, new_n30781_, new_n23452_ );
or   ( new_n35320_, new_n35319_, new_n34198_ );
or   ( new_n35321_, new_n30782_, new_n23451_ );
or   ( new_n35322_, new_n35321_, new_n34257_ );
and  ( new_n35323_, new_n35322_, new_n35320_ );
and  ( new_n35324_, new_n35323_, new_n35318_ );
and  ( new_n35325_, new_n15634_, new_n7407_ );
and  ( new_n35326_, new_n35325_, new_n33953_ );
or   ( new_n35327_, new_n15635_, new_n7406_ );
and  ( new_n35328_, new_n35327_, new_n33975_ );
or   ( new_n35329_, new_n35328_, new_n35326_ );
and  ( new_n35330_, new_n30759_, new_n22564_ );
or   ( new_n35331_, new_n35330_, new_n33997_ );
or   ( new_n35332_, new_n30760_, new_n22563_ );
or   ( new_n35333_, new_n35332_, new_n34017_ );
and  ( new_n35334_, new_n35333_, new_n35331_ );
and  ( new_n35335_, new_n35334_, new_n35329_ );
or   ( new_n35336_, new_n35335_, new_n35324_ );
or   ( new_n35337_, new_n35336_, new_n35313_ );
or   ( new_n35338_, new_n31938_, new_n31816_ );
or   ( new_n35339_, new_n35338_, new_n33881_ );
or   ( new_n35340_, new_n35339_, new_n34296_ );
or   ( new_n35341_, new_n34302_, new_n34299_ );
and  ( new_n35342_, new_n35341_, new_n34298_ );
or   ( new_n35343_, new_n35342_, new_n35340_ );
or   ( new_n35344_, new_n35339_, new_n34295_ );
or   ( new_n35345_, new_n34300_, new_n34299_ );
or   ( new_n35346_, new_n35345_, new_n35340_ );
or   ( new_n35347_, new_n32061_, new_n31959_ );
and  ( new_n35348_, new_n32997_, new_n32907_ );
and  ( new_n35349_, new_n32924_, new_n32886_ );
or   ( new_n35350_, new_n35349_, new_n32938_ );
and  ( new_n35351_, new_n32886_, new_n32752_ );
and  ( new_n35352_, new_n34336_, new_n33920_ );
or   ( new_n35353_, new_n35352_, new_n33928_ );
and  ( new_n35354_, new_n35353_, new_n35351_ );
or   ( new_n35355_, new_n35354_, new_n35350_ );
or   ( new_n35356_, new_n35355_, new_n35348_ );
or   ( new_n35357_, new_n32977_, new_n32931_ );
or   ( new_n35358_, new_n32989_, new_n32973_ );
and  ( new_n35359_, new_n35358_, new_n33003_ );
or   ( new_n35360_, new_n32973_, new_n32955_ );
or   ( new_n35361_, new_n34348_, new_n33908_ );
and  ( new_n35362_, new_n35361_, new_n33916_ );
or   ( new_n35363_, new_n35362_, new_n35360_ );
and  ( new_n35364_, new_n35363_, new_n35359_ );
or   ( new_n35365_, new_n35364_, new_n35357_ );
and  ( new_n35366_, new_n35365_, new_n35356_ );
and  ( new_n35367_, new_n35366_, new_n35347_ );
and  ( new_n35368_, new_n32037_, new_n31987_ );
or   ( new_n35369_, new_n35357_, new_n35355_ );
or   ( new_n35370_, new_n35364_, new_n35348_ );
and  ( new_n35371_, new_n35370_, new_n35369_ );
and  ( new_n35372_, new_n35371_, new_n35368_ );
or   ( new_n35373_, new_n35372_, new_n35367_ );
or   ( new_n35374_, new_n31980_, new_n31938_ );
and  ( new_n35375_, new_n35374_, new_n31994_ );
or   ( new_n35376_, new_n35338_, new_n33888_ );
and  ( new_n35377_, new_n35376_, new_n35375_ );
and  ( new_n35378_, new_n35377_, new_n35373_ );
and  ( new_n35379_, new_n35378_, new_n35346_ );
and  ( new_n35380_, new_n35379_, new_n35344_ );
and  ( new_n35381_, new_n35380_, new_n35343_ );
or   ( new_n35382_, new_n31959_, new_n31937_ );
or   ( new_n35383_, new_n35382_, new_n33133_ );
or   ( new_n35384_, new_n35383_, new_n34487_ );
or   ( new_n35385_, new_n35384_, new_n34046_ );
or   ( new_n35386_, new_n34062_, new_n34055_ );
and  ( new_n35387_, new_n35386_, new_n34053_ );
or   ( new_n35388_, new_n35387_, new_n35385_ );
or   ( new_n35389_, new_n35384_, new_n34044_ );
or   ( new_n35390_, new_n35385_, new_n34090_ );
or   ( new_n35391_, new_n35390_, new_n34055_ );
or   ( new_n35392_, new_n35383_, new_n34495_ );
and  ( new_n35393_, new_n34644_, new_n34613_ );
and  ( new_n35394_, new_n34645_, new_n34640_ );
or   ( new_n35395_, new_n35394_, new_n35393_ );
or   ( new_n35396_, new_n35382_, new_n33156_ );
and  ( new_n35397_, new_n31992_, new_n31987_ );
or   ( new_n35398_, new_n35397_, new_n31959_ );
and  ( new_n35399_, new_n35398_, new_n35396_ );
and  ( new_n35400_, new_n35399_, new_n35395_ );
and  ( new_n35401_, new_n35400_, new_n35392_ );
and  ( new_n35402_, new_n35401_, new_n35391_ );
and  ( new_n35403_, new_n35402_, new_n35389_ );
and  ( new_n35404_, new_n35403_, new_n35388_ );
or   ( new_n35405_, new_n35404_, new_n35381_ );
or   ( new_n35406_, new_n35405_, new_n35337_ );
and  ( new_n35407_, new_n34318_, new_n34316_ );
or   ( new_n35408_, new_n35407_, new_n34315_ );
and  ( new_n35409_, new_n32033_, new_n32020_ );
and  ( new_n35410_, new_n35409_, new_n33895_ );
and  ( new_n35411_, new_n35410_, new_n34313_ );
and  ( new_n35412_, new_n35411_, new_n35408_ );
and  ( new_n35413_, new_n35410_, new_n34312_ );
and  ( new_n35414_, new_n34319_, new_n34316_ );
and  ( new_n35415_, new_n35414_, new_n35411_ );
and  ( new_n35416_, new_n32053_, new_n32033_ );
or   ( new_n35417_, new_n35416_, new_n32067_ );
and  ( new_n35418_, new_n35409_, new_n33902_ );
or   ( new_n35419_, new_n35418_, new_n35417_ );
or   ( new_n35420_, new_n35419_, new_n35415_ );
or   ( new_n35421_, new_n35420_, new_n35413_ );
or   ( new_n35422_, new_n35421_, new_n35412_ );
and  ( new_n35423_, new_n35371_, new_n35347_ );
and  ( new_n35424_, new_n35368_, new_n35366_ );
or   ( new_n35425_, new_n35424_, new_n35423_ );
and  ( new_n35426_, new_n35425_, new_n35422_ );
and  ( new_n35427_, new_n35327_, new_n33953_ );
and  ( new_n35428_, new_n35325_, new_n33975_ );
or   ( new_n35429_, new_n35428_, new_n35427_ );
or   ( new_n35430_, new_n35332_, new_n33997_ );
or   ( new_n35431_, new_n35330_, new_n34017_ );
and  ( new_n35432_, new_n35431_, new_n35430_ );
and  ( new_n35433_, new_n35432_, new_n35429_ );
and  ( new_n35434_, new_n34703_, new_n34303_ );
and  ( new_n35435_, new_n34701_, new_n34320_ );
or   ( new_n35436_, new_n35435_, new_n35434_ );
or   ( new_n35437_, new_n34708_, new_n34339_ );
or   ( new_n35438_, new_n34706_, new_n34327_ );
and  ( new_n35439_, new_n35438_, new_n35437_ );
and  ( new_n35440_, new_n35439_, new_n35436_ );
and  ( new_n35441_, new_n35316_, new_n34091_ );
and  ( new_n35442_, new_n35314_, new_n34153_ );
or   ( new_n35443_, new_n35442_, new_n35441_ );
or   ( new_n35444_, new_n35321_, new_n34198_ );
or   ( new_n35445_, new_n35319_, new_n34257_ );
and  ( new_n35446_, new_n35445_, new_n35444_ );
and  ( new_n35447_, new_n35446_, new_n35443_ );
or   ( new_n35448_, new_n35447_, new_n35440_ );
or   ( new_n35449_, new_n35448_, new_n35433_ );
or   ( new_n35450_, new_n35449_, new_n35426_ );
or   ( new_n35451_, new_n35450_, new_n35406_ );
or   ( new_n35452_, new_n35451_, new_n34700_ );
or   ( new_n35453_, new_n35452_, new_n34612_ );
or   ( new_n35454_, new_n857_, new_n99_ );
and  ( new_n35455_, new_n35454_, new_n842_ );
and  ( new_n35456_, new_n870_, RI2b1c4342d4e0_65 );
and  ( new_n35457_, new_n35456_, new_n866_ );
or   ( new_n35458_, new_n35457_, new_n35455_ );
or   ( new_n35459_, new_n841_, new_n526_ );
and  ( new_n35460_, new_n35459_, new_n35458_ );
and  ( new_n35461_, new_n35456_, new_n842_ );
and  ( new_n35462_, new_n35454_, new_n866_ );
or   ( new_n35463_, new_n35462_, new_n35461_ );
and  ( new_n35464_, new_n720_, RI2b1c4342d558_66 );
and  ( new_n35465_, new_n35464_, new_n35463_ );
or   ( new_n35466_, new_n35465_, new_n35460_ );
or   ( new_n35467_, new_n31135_, new_n785_ );
or   ( new_n35468_, new_n31143_, new_n31136_ );
and  ( new_n35469_, new_n35468_, new_n35467_ );
and  ( new_n35470_, new_n35469_, new_n35466_ );
and  ( new_n35471_, new_n35463_, new_n35459_ );
and  ( new_n35472_, new_n35464_, new_n35458_ );
or   ( new_n35473_, new_n35472_, new_n35471_ );
or   ( new_n35474_, new_n31139_, new_n813_ );
and  ( new_n35475_, new_n35474_, new_n31126_ );
or   ( new_n35476_, new_n35475_, new_n31140_ );
and  ( new_n35477_, new_n35476_, new_n35473_ );
or   ( new_n35478_, new_n35477_, new_n35470_ );
or   ( new_n35479_, new_n31205_, new_n31202_ );
and  ( new_n35480_, new_n35479_, new_n31148_ );
or   ( new_n35481_, new_n35480_, new_n31206_ );
or   ( new_n35482_, new_n35481_, new_n35478_ );
and  ( new_n35483_, new_n35473_, new_n35469_ );
and  ( new_n35484_, new_n35476_, new_n35466_ );
or   ( new_n35485_, new_n35484_, new_n35483_ );
or   ( new_n35486_, new_n31223_, new_n31220_ );
or   ( new_n35487_, new_n31229_, new_n31224_ );
and  ( new_n35488_, new_n35487_, new_n35486_ );
or   ( new_n35489_, new_n35488_, new_n35485_ );
and  ( new_n35490_, new_n35489_, new_n35482_ );
and  ( new_n35491_, new_n16132_, RI2b1c4342d4e0_65 );
or   ( new_n35492_, new_n35491_, new_n16108_ );
or   ( new_n35493_, new_n16119_, new_n99_ );
or   ( new_n35494_, new_n35493_, new_n16128_ );
and  ( new_n35495_, new_n35494_, new_n35492_ );
and  ( new_n35496_, new_n16102_, RI2b1c4342d558_66 );
or   ( new_n35497_, new_n35496_, new_n35495_ );
or   ( new_n35498_, new_n35493_, new_n16108_ );
or   ( new_n35499_, new_n35491_, new_n16128_ );
and  ( new_n35500_, new_n35499_, new_n35498_ );
or   ( new_n35501_, new_n16115_, new_n526_ );
or   ( new_n35502_, new_n35501_, new_n35500_ );
and  ( new_n35503_, new_n35502_, new_n35497_ );
and  ( new_n35504_, new_n32085_, new_n16151_ );
and  ( new_n35505_, new_n32093_, new_n32086_ );
or   ( new_n35506_, new_n35505_, new_n35504_ );
or   ( new_n35507_, new_n35506_, new_n35503_ );
or   ( new_n35508_, new_n35500_, new_n35496_ );
or   ( new_n35509_, new_n35501_, new_n35495_ );
and  ( new_n35510_, new_n35509_, new_n35508_ );
and  ( new_n35511_, new_n32089_, new_n16170_ );
or   ( new_n35512_, new_n35511_, new_n32076_ );
and  ( new_n35513_, new_n35512_, new_n32090_ );
or   ( new_n35514_, new_n35513_, new_n35510_ );
and  ( new_n35515_, new_n35514_, new_n35507_ );
and  ( new_n35516_, new_n32155_, new_n32152_ );
or   ( new_n35517_, new_n35516_, new_n32098_ );
and  ( new_n35518_, new_n35517_, new_n32156_ );
or   ( new_n35519_, new_n35518_, new_n35515_ );
or   ( new_n35520_, new_n35510_, new_n35506_ );
or   ( new_n35521_, new_n35513_, new_n35503_ );
and  ( new_n35522_, new_n35521_, new_n35520_ );
and  ( new_n35523_, new_n32173_, new_n32170_ );
and  ( new_n35524_, new_n32182_, new_n32174_ );
or   ( new_n35525_, new_n35524_, new_n35523_ );
or   ( new_n35526_, new_n35525_, new_n35522_ );
and  ( new_n35527_, new_n35526_, new_n35519_ );
and  ( new_n35528_, new_n32944_, new_n32916_ );
and  ( new_n35529_, new_n35528_, new_n34614_ );
and  ( new_n35530_, new_n35529_, new_n33617_ );
and  ( new_n35531_, new_n35530_, new_n34023_ );
and  ( new_n35532_, new_n35530_, new_n34025_ );
and  ( new_n35533_, new_n35529_, new_n33628_ );
and  ( new_n35534_, new_n35528_, new_n34621_ );
and  ( new_n35535_, new_n32944_, new_n32932_ );
or   ( new_n35536_, new_n35535_, new_n32292_ );
or   ( new_n35537_, new_n35536_, new_n35534_ );
or   ( new_n35538_, new_n35537_, new_n35533_ );
or   ( new_n35539_, new_n35538_, new_n35532_ );
or   ( new_n35540_, new_n35539_, new_n35531_ );
or   ( new_n35541_, new_n35540_, new_n35527_ );
and  ( new_n35542_, new_n35518_, new_n35515_ );
and  ( new_n35543_, new_n35525_, new_n35522_ );
or   ( new_n35544_, new_n35543_, new_n35542_ );
or   ( new_n35545_, new_n32981_, new_n32332_ );
or   ( new_n35546_, new_n35545_, new_n34628_ );
or   ( new_n35547_, new_n35546_, new_n33448_ );
or   ( new_n35548_, new_n35547_, new_n34003_ );
or   ( new_n35549_, new_n35547_, new_n34005_ );
or   ( new_n35550_, new_n35546_, new_n33474_ );
or   ( new_n35551_, new_n35545_, new_n34635_ );
or   ( new_n35552_, new_n32996_, new_n32332_ );
and  ( new_n35553_, new_n35552_, new_n32945_ );
and  ( new_n35554_, new_n35553_, new_n35551_ );
and  ( new_n35555_, new_n35554_, new_n35550_ );
and  ( new_n35556_, new_n35555_, new_n35549_ );
and  ( new_n35557_, new_n35556_, new_n35548_ );
or   ( new_n35558_, new_n35557_, new_n35544_ );
and  ( new_n35559_, new_n35558_, new_n35541_ );
and  ( new_n35560_, new_n35559_, new_n35490_ );
and  ( new_n35561_, new_n35481_, new_n35478_ );
and  ( new_n35562_, new_n35488_, new_n35485_ );
or   ( new_n35563_, new_n35562_, new_n35561_ );
or   ( new_n35564_, new_n35544_, new_n35540_ );
or   ( new_n35565_, new_n35557_, new_n35527_ );
and  ( new_n35566_, new_n35565_, new_n35564_ );
and  ( new_n35567_, new_n35566_, new_n35563_ );
or   ( new_n35568_, new_n35567_, new_n35560_ );
and  ( new_n35569_, new_n32041_, new_n31382_ );
and  ( new_n35570_, new_n35569_, new_n34651_ );
and  ( new_n35571_, new_n35570_, new_n33293_ );
and  ( new_n35572_, new_n35571_, new_n33981_ );
and  ( new_n35573_, new_n35571_, new_n33983_ );
and  ( new_n35574_, new_n35570_, new_n33316_ );
and  ( new_n35575_, new_n35569_, new_n34663_ );
and  ( new_n35576_, new_n32060_, new_n31382_ );
or   ( new_n35577_, new_n35576_, new_n32003_ );
or   ( new_n35578_, new_n35577_, new_n35575_ );
or   ( new_n35579_, new_n35578_, new_n35574_ );
or   ( new_n35580_, new_n35579_, new_n35573_ );
or   ( new_n35581_, new_n35580_, new_n35572_ );
and  ( new_n35582_, new_n35581_, new_n35568_ );
and  ( new_n35583_, new_n15570_, new_n4367_ );
and  ( new_n35584_, new_n35583_, new_n15323_ );
or   ( new_n35585_, new_n15558_, new_n4379_ );
and  ( new_n35586_, new_n35585_, new_n15996_ );
or   ( new_n35587_, new_n35586_, new_n35584_ );
and  ( new_n35588_, new_n30697_, new_n19611_ );
or   ( new_n35589_, new_n35588_, new_n30449_ );
or   ( new_n35590_, new_n30690_, new_n19618_ );
or   ( new_n35591_, new_n35590_, new_n31118_ );
and  ( new_n35592_, new_n35591_, new_n35589_ );
and  ( new_n35593_, new_n35592_, new_n35587_ );
and  ( new_n35594_, new_n34547_, new_n34544_ );
and  ( new_n35595_, new_n34552_, new_n34545_ );
or   ( new_n35596_, new_n35595_, new_n35594_ );
or   ( new_n35597_, new_n34558_, new_n34555_ );
or   ( new_n35598_, new_n34559_, new_n34556_ );
and  ( new_n35599_, new_n35598_, new_n35597_ );
and  ( new_n35600_, new_n35599_, new_n35596_ );
and  ( new_n35601_, new_n35585_, new_n15323_ );
and  ( new_n35602_, new_n35583_, new_n15996_ );
or   ( new_n35603_, new_n35602_, new_n35601_ );
or   ( new_n35604_, new_n35590_, new_n30449_ );
or   ( new_n35605_, new_n35588_, new_n31118_ );
and  ( new_n35606_, new_n35605_, new_n35604_ );
and  ( new_n35607_, new_n35606_, new_n35603_ );
or   ( new_n35608_, new_n35607_, new_n35600_ );
or   ( new_n35609_, new_n35608_, new_n35593_ );
or   ( new_n35610_, new_n35609_, new_n35582_ );
or   ( new_n35611_, new_n35610_, new_n35453_ );
and  ( new_n35612_, new_n34285_, new_n33957_ );
and  ( new_n35613_, new_n34283_, new_n33979_ );
or   ( new_n35614_, new_n35613_, new_n35612_ );
or   ( new_n35615_, new_n34288_, new_n34021_ );
or   ( new_n35616_, new_n34290_, new_n34001_ );
and  ( new_n35617_, new_n35616_, new_n35615_ );
and  ( new_n35618_, new_n35617_, new_n35614_ );
and  ( new_n35619_, new_n34310_, new_n34307_ );
and  ( new_n35620_, new_n34324_, new_n34308_ );
or   ( new_n35621_, new_n35620_, new_n35619_ );
or   ( new_n35622_, new_n34348_, new_n34337_ );
or   ( new_n35623_, new_n34349_, new_n34336_ );
and  ( new_n35624_, new_n35623_, new_n35622_ );
and  ( new_n35625_, new_n35624_, new_n35621_ );
or   ( new_n35626_, new_n35625_, new_n35618_ );
and  ( new_n35627_, new_n33153_, new_n33131_ );
or   ( new_n35628_, new_n15529_, new_n2635_ );
and  ( new_n35629_, new_n35628_, new_n35627_ );
and  ( new_n35630_, new_n15530_, new_n2636_ );
or   ( new_n35631_, new_n33309_, new_n33287_ );
and  ( new_n35632_, new_n35631_, new_n35630_ );
or   ( new_n35633_, new_n35632_, new_n35629_ );
and  ( new_n35634_, new_n30658_, new_n17922_ );
or   ( new_n35635_, new_n35634_, new_n33614_ );
and  ( new_n35636_, new_n33467_, new_n33445_ );
or   ( new_n35637_, new_n30659_, new_n17923_ );
or   ( new_n35638_, new_n35637_, new_n35636_ );
and  ( new_n35639_, new_n35638_, new_n35635_ );
and  ( new_n35640_, new_n35639_, new_n35633_ );
and  ( new_n35641_, new_n34098_, new_n34095_ );
and  ( new_n35642_, new_n34157_, new_n34096_ );
or   ( new_n35643_, new_n35642_, new_n35641_ );
or   ( new_n35644_, new_n34279_, new_n34219_ );
or   ( new_n35645_, new_n34278_, new_n34220_ );
and  ( new_n35646_, new_n35645_, new_n35644_ );
and  ( new_n35647_, new_n35646_, new_n35643_ );
or   ( new_n35648_, new_n35647_, new_n35640_ );
or   ( new_n35649_, new_n35648_, new_n35626_ );
and  ( new_n35650_, new_n34690_, new_n34093_ );
and  ( new_n35651_, new_n34688_, new_n34155_ );
or   ( new_n35652_, new_n35651_, new_n35650_ );
or   ( new_n35653_, new_n34695_, new_n34208_ );
or   ( new_n35654_, new_n34693_, new_n34267_ );
and  ( new_n35655_, new_n35654_, new_n35653_ );
and  ( new_n35656_, new_n35655_, new_n35652_ );
or   ( new_n35657_, new_n15593_, new_n5576_ );
and  ( new_n35658_, new_n35657_, new_n33123_ );
and  ( new_n35659_, new_n15594_, new_n5577_ );
and  ( new_n35660_, new_n35659_, new_n33279_ );
or   ( new_n35661_, new_n35660_, new_n35658_ );
or   ( new_n35662_, new_n30720_, new_n20793_ );
or   ( new_n35663_, new_n35662_, new_n33437_ );
and  ( new_n35664_, new_n30719_, new_n20792_ );
or   ( new_n35665_, new_n35664_, new_n33591_ );
and  ( new_n35666_, new_n35665_, new_n35663_ );
and  ( new_n35667_, new_n35666_, new_n35661_ );
or   ( new_n35668_, new_n35667_, new_n35656_ );
and  ( new_n35669_, new_n34679_, new_n34305_ );
and  ( new_n35670_, new_n34677_, new_n34322_ );
or   ( new_n35671_, new_n35670_, new_n35669_ );
or   ( new_n35672_, new_n34684_, new_n34344_ );
or   ( new_n35673_, new_n34682_, new_n34332_ );
and  ( new_n35674_, new_n35673_, new_n35672_ );
and  ( new_n35675_, new_n35674_, new_n35671_ );
and  ( new_n35676_, new_n35659_, new_n33123_ );
and  ( new_n35677_, new_n35657_, new_n33279_ );
or   ( new_n35678_, new_n35677_, new_n35676_ );
or   ( new_n35679_, new_n35664_, new_n33437_ );
or   ( new_n35680_, new_n35662_, new_n33591_ );
and  ( new_n35681_, new_n35680_, new_n35679_ );
and  ( new_n35682_, new_n35681_, new_n35678_ );
or   ( new_n35683_, new_n35682_, new_n35675_ );
or   ( new_n35684_, new_n35683_, new_n35668_ );
and  ( new_n35685_, new_n34533_, new_n34496_ );
and  ( new_n35686_, new_n34534_, new_n34529_ );
or   ( new_n35687_, new_n35686_, new_n35685_ );
and  ( new_n35688_, new_n34650_, new_n34099_ );
and  ( new_n35689_, new_n35688_, new_n34551_ );
and  ( new_n35690_, new_n35688_, new_n34549_ );
and  ( new_n35691_, new_n34650_, new_n34104_ );
or   ( new_n35692_, new_n35691_, new_n34660_ );
or   ( new_n35693_, new_n35692_, new_n35690_ );
or   ( new_n35694_, new_n35693_, new_n35689_ );
and  ( new_n35695_, new_n35694_, new_n35687_ );
or   ( new_n35696_, new_n31817_, new_n4376_ );
or   ( new_n35697_, new_n35696_, new_n34424_ );
or   ( new_n35698_, new_n35696_, new_n34426_ );
or   ( new_n35699_, new_n31817_, new_n2972_ );
and  ( new_n35700_, new_n34587_, new_n34563_ );
and  ( new_n35701_, new_n34584_, new_n34582_ );
or   ( new_n35702_, new_n35701_, new_n35700_ );
and  ( new_n35703_, new_n35702_, new_n31985_ );
and  ( new_n35704_, new_n35703_, new_n35699_ );
and  ( new_n35705_, new_n35704_, new_n35698_ );
and  ( new_n35706_, new_n35705_, new_n35697_ );
or   ( new_n35707_, new_n35706_, new_n35695_ );
and  ( new_n35708_, new_n15606_, new_n5987_ );
and  ( new_n35709_, new_n35708_, new_n34422_ );
or   ( new_n35710_, new_n15601_, new_n5992_ );
and  ( new_n35711_, new_n35710_, new_n34598_ );
or   ( new_n35712_, new_n35711_, new_n35709_ );
and  ( new_n35713_, new_n30731_, new_n21189_ );
or   ( new_n35714_, new_n35713_, new_n34455_ );
or   ( new_n35715_, new_n30726_, new_n21194_ );
or   ( new_n35716_, new_n35715_, new_n34438_ );
and  ( new_n35717_, new_n35716_, new_n35714_ );
and  ( new_n35718_, new_n35717_, new_n35712_ );
and  ( new_n35719_, new_n35710_, new_n34422_ );
and  ( new_n35720_, new_n35708_, new_n34598_ );
or   ( new_n35721_, new_n35720_, new_n35719_ );
or   ( new_n35722_, new_n35715_, new_n34455_ );
or   ( new_n35723_, new_n35713_, new_n34438_ );
and  ( new_n35724_, new_n35723_, new_n35722_ );
and  ( new_n35725_, new_n35724_, new_n35721_ );
or   ( new_n35726_, new_n35725_, new_n35718_ );
or   ( new_n35727_, new_n35726_, new_n35707_ );
or   ( new_n35728_, new_n35727_, new_n35684_ );
and  ( new_n35729_, new_n35630_, new_n35627_ );
and  ( new_n35730_, new_n35631_, new_n35628_ );
or   ( new_n35731_, new_n35730_, new_n35729_ );
or   ( new_n35732_, new_n35636_, new_n35634_ );
or   ( new_n35733_, new_n35637_, new_n33614_ );
and  ( new_n35734_, new_n35733_, new_n35732_ );
and  ( new_n35735_, new_n35734_, new_n35731_ );
or   ( new_n35736_, new_n32002_, new_n31968_ );
or   ( new_n35737_, new_n35736_, new_n35382_ );
or   ( new_n35738_, new_n35737_, new_n33134_ );
or   ( new_n35739_, new_n35738_, new_n33959_ );
or   ( new_n35740_, new_n35738_, new_n33961_ );
and  ( new_n35741_, new_n35566_, new_n35490_ );
and  ( new_n35742_, new_n35563_, new_n35559_ );
or   ( new_n35743_, new_n35742_, new_n35741_ );
or   ( new_n35744_, new_n35737_, new_n33160_ );
or   ( new_n35745_, new_n35736_, new_n35398_ );
or   ( new_n35746_, new_n32002_, new_n31988_ );
and  ( new_n35747_, new_n35746_, new_n31342_ );
and  ( new_n35748_, new_n35747_, new_n35745_ );
and  ( new_n35749_, new_n35748_, new_n35744_ );
and  ( new_n35750_, new_n35749_, new_n35743_ );
and  ( new_n35751_, new_n35750_, new_n35740_ );
and  ( new_n35752_, new_n35751_, new_n35739_ );
or   ( new_n35753_, new_n35752_, new_n35735_ );
or   ( new_n35754_, new_n35753_, new_n35728_ );
or   ( new_n35755_, new_n35754_, new_n35649_ );
or   ( new_n35756_, new_n35755_, new_n35611_ );
or   ( new_n35757_, new_n35756_, new_n34356_ );
or   ( new_n35758_, new_n841_, new_n99_ );
or   ( new_n35759_, new_n35464_, new_n35463_ );
and  ( new_n35760_, new_n35759_, new_n866_ );
and  ( new_n35761_, new_n35460_, new_n842_ );
or   ( new_n35762_, new_n35761_, new_n35760_ );
and  ( new_n35763_, new_n35762_, new_n35758_ );
and  ( new_n35764_, new_n35460_, new_n866_ );
and  ( new_n35765_, new_n35759_, new_n842_ );
or   ( new_n35766_, new_n35765_, new_n35764_ );
and  ( new_n35767_, new_n720_, RI2b1c4342d4e0_65 );
and  ( new_n35768_, new_n35767_, new_n35766_ );
or   ( new_n35769_, new_n35768_, new_n35763_ );
and  ( new_n35770_, new_n35769_, new_n35470_ );
and  ( new_n35771_, new_n35766_, new_n35758_ );
and  ( new_n35772_, new_n35767_, new_n35762_ );
or   ( new_n35773_, new_n35772_, new_n35771_ );
or   ( new_n35774_, new_n35476_, new_n35473_ );
and  ( new_n35775_, new_n35774_, new_n35773_ );
or   ( new_n35776_, new_n35775_, new_n35770_ );
or   ( new_n35777_, new_n35561_, new_n32002_ );
or   ( new_n35778_, new_n35777_, new_n31969_ );
or   ( new_n35779_, new_n35778_, new_n35338_ );
or   ( new_n35780_, new_n35779_, new_n33883_ );
or   ( new_n35781_, new_n35779_, new_n33889_ );
or   ( new_n35782_, new_n35778_, new_n35375_ );
or   ( new_n35783_, new_n35777_, new_n31990_ );
or   ( new_n35784_, new_n35561_, new_n31342_ );
and  ( new_n35785_, new_n35784_, new_n35482_ );
and  ( new_n35786_, new_n35785_, new_n35783_ );
and  ( new_n35787_, new_n35786_, new_n35782_ );
and  ( new_n35788_, new_n35787_, new_n35781_ );
and  ( new_n35789_, new_n35788_, new_n35780_ );
and  ( new_n35790_, new_n35789_, new_n35776_ );
or   ( new_n35791_, new_n35774_, new_n35773_ );
or   ( new_n35792_, new_n35769_, new_n35470_ );
and  ( new_n35793_, new_n35792_, new_n35791_ );
and  ( new_n35794_, new_n35489_, new_n31382_ );
and  ( new_n35795_, new_n35794_, new_n32042_ );
and  ( new_n35796_, new_n35795_, new_n35409_ );
and  ( new_n35797_, new_n35796_, new_n33897_ );
and  ( new_n35798_, new_n35796_, new_n33903_ );
and  ( new_n35799_, new_n35795_, new_n35417_ );
and  ( new_n35800_, new_n35794_, new_n32063_ );
and  ( new_n35801_, new_n35489_, new_n32003_ );
or   ( new_n35802_, new_n35801_, new_n35562_ );
or   ( new_n35803_, new_n35802_, new_n35800_ );
or   ( new_n35804_, new_n35803_, new_n35799_ );
or   ( new_n35805_, new_n35804_, new_n35798_ );
or   ( new_n35806_, new_n35805_, new_n35797_ );
and  ( new_n35807_, new_n35806_, new_n35793_ );
or   ( new_n35808_, new_n35807_, new_n35790_ );
and  ( new_n35809_, new_n16102_, RI2b1c4342d4e0_65 );
and  ( new_n35810_, new_n35501_, new_n35500_ );
or   ( new_n35811_, new_n35810_, new_n16128_ );
or   ( new_n35812_, new_n35497_, new_n16108_ );
and  ( new_n35813_, new_n35812_, new_n35811_ );
or   ( new_n35814_, new_n35813_, new_n35809_ );
or   ( new_n35815_, new_n35497_, new_n16128_ );
or   ( new_n35816_, new_n35810_, new_n16108_ );
and  ( new_n35817_, new_n35816_, new_n35815_ );
or   ( new_n35818_, new_n16115_, new_n99_ );
or   ( new_n35819_, new_n35818_, new_n35817_ );
and  ( new_n35820_, new_n35819_, new_n35814_ );
or   ( new_n35821_, new_n35820_, new_n35507_ );
or   ( new_n35822_, new_n35817_, new_n35809_ );
or   ( new_n35823_, new_n35818_, new_n35813_ );
and  ( new_n35824_, new_n35823_, new_n35822_ );
and  ( new_n35825_, new_n35513_, new_n35510_ );
or   ( new_n35826_, new_n35825_, new_n35824_ );
and  ( new_n35827_, new_n35826_, new_n35821_ );
and  ( new_n35828_, new_n35519_, new_n32944_ );
and  ( new_n35829_, new_n35828_, new_n32917_ );
and  ( new_n35830_, new_n35829_, new_n35351_ );
and  ( new_n35831_, new_n35830_, new_n33923_ );
and  ( new_n35832_, new_n35830_, new_n33929_ );
and  ( new_n35833_, new_n35829_, new_n35350_ );
and  ( new_n35834_, new_n35828_, new_n32934_ );
and  ( new_n35835_, new_n35519_, new_n32292_ );
or   ( new_n35836_, new_n35835_, new_n35542_ );
or   ( new_n35837_, new_n35836_, new_n35834_ );
or   ( new_n35838_, new_n35837_, new_n35833_ );
or   ( new_n35839_, new_n35838_, new_n35832_ );
or   ( new_n35840_, new_n35839_, new_n35831_ );
or   ( new_n35841_, new_n35840_, new_n35827_ );
and  ( new_n35842_, new_n35825_, new_n35824_ );
and  ( new_n35843_, new_n35820_, new_n35507_ );
or   ( new_n35844_, new_n35843_, new_n35842_ );
or   ( new_n35845_, new_n35543_, new_n32332_ );
or   ( new_n35846_, new_n35845_, new_n32982_ );
or   ( new_n35847_, new_n35846_, new_n35360_ );
or   ( new_n35848_, new_n35847_, new_n33911_ );
or   ( new_n35849_, new_n35847_, new_n33917_ );
or   ( new_n35850_, new_n35846_, new_n35359_ );
or   ( new_n35851_, new_n35845_, new_n32999_ );
or   ( new_n35852_, new_n35543_, new_n32945_ );
and  ( new_n35853_, new_n35852_, new_n35526_ );
and  ( new_n35854_, new_n35853_, new_n35851_ );
and  ( new_n35855_, new_n35854_, new_n35850_ );
and  ( new_n35856_, new_n35855_, new_n35849_ );
and  ( new_n35857_, new_n35856_, new_n35848_ );
or   ( new_n35858_, new_n35857_, new_n35844_ );
and  ( new_n35859_, new_n35858_, new_n35841_ );
and  ( new_n35860_, new_n35859_, new_n35808_ );
and  ( new_n35861_, new_n35793_, new_n35789_ );
and  ( new_n35862_, new_n35806_, new_n35776_ );
or   ( new_n35863_, new_n35862_, new_n35861_ );
or   ( new_n35864_, new_n35857_, new_n35827_ );
or   ( new_n35865_, new_n35844_, new_n35840_ );
and  ( new_n35866_, new_n35865_, new_n35864_ );
and  ( new_n35867_, new_n35866_, new_n35863_ );
or   ( new_n35868_, new_n35867_, new_n35860_ );
or   ( new_n35869_, new_n35868_, new_n35757_ );
or   ( eq, new_n35869_, new_n33943_ );
endmodule


