module miter ( 
    RIbb2f070_13, RIbb2eff8_14, RIbb2ef80_15, RIbb2d798_66, RIbb2f160_11,
    RIbb2f0e8_12, RIbb2d810_65, RIbb2d6a8_68, RIbb2f250_9, RIbb2f1d8_10,
    RIbb2d720_67, RIbb2d5b8_70, RIbb2f340_7, RIbb2f2c8_8, RIbb2d630_69,
    RIbb2d4c8_72, RIbb2f430_5, RIbb2f3b8_6, RIbb2d540_71, RIbb2d3d8_74,
    RIbb2f520_3, RIbb2f4a8_4, RIbb2d450_73, RIbb2d2e8_76, RIbb2f610_1,
    RIbb2f598_2, RIbb2d360_75, RIbb2d270_77, RIbb2d1f8_78, RIbb2ef08_16,
    RIbb2ee90_17, RIbb2d180_79, RIbb2d108_80, RIbb2ee18_18, RIbb2eda0_19,
    RIbb2d090_81, RIbb2ed28_20, RIbb2ecb0_21, RIbb2d018_82, RIbb2cfa0_83,
    RIbb2cf28_84, RIbb2ec38_22, RIbb2ebc0_23, RIbb2ceb0_85, RIbb2ce38_86,
    RIbb2eb48_24, RIbb2ead0_25, RIbb2cdc0_87, RIbb2cd48_88, RIbb2ea58_26,
    RIbb2e9e0_27, RIbb2ccd0_89, RIbb2cc58_90, RIbb2e968_28, RIbb2e8f0_29,
    RIbb2cbe0_91, RIbb2cb68_92, RIbb2e878_30, RIbb2e800_31, RIbb2caf0_93,
    RIbb2ca78_94, RIbb2e788_32, RIbb2e710_33, RIbb2ca00_95, RIbb2c988_96,
    RIbb2e698_34, RIbb2e620_35, RIbb2c910_97, RIbb2c898_98, RIbb2e5a8_36,
    RIbb2e530_37, RIbb2c820_99, RIbb2e4b8_38, RIbb2e440_39, RIbb2c7a8_100,
    RIbb2c730_101, RIbb2c6b8_102, RIbb2e3c8_40, RIbb2e350_41,
    RIbb2c640_103, RIbb2c5c8_104, RIbb2e2d8_42, RIbb2e260_43,
    RIbb2c550_105, RIbb2c4d8_106, RIbb2e1e8_44, RIbb2e170_45,
    RIbb2c460_107, RIbb2c3e8_108, RIbb2e0f8_46, RIbb2e080_47,
    RIbb2c370_109, RIbb2c2f8_110, RIbb2e008_48, RIbb2df90_49,
    RIbb2c280_111, RIbb2c208_112, RIbb2df18_50, RIbb2dea0_51,
    RIbb2c190_113, RIbb2c118_114, RIbb2de28_52, RIbb2ddb0_53,
    RIbb2c0a0_115, RIbb2c028_116, RIbb2dd38_54, RIbb2dcc0_55,
    RIbb2bfb0_117, RIbb2dc48_56, RIbb2dbd0_57, RIbb2bf38_118,
    RIbb2bec0_119, RIbb2be48_120, RIbb2db58_58, RIbb2dae0_59,
    RIbb2bdd0_121, RIbb2bd58_122, RIbb2da68_60, RIbb2d9f0_61,
    RIbb2bce0_123, RIbb2bc68_124, RIbb2d978_62, RIbb2d900_63,
    RIbb2bbf0_125, RIbb2bb78_126, RIbb31500_127, RIbb2d888_64,
    RIbb31578_128, RIbb31668_130, RIbb315f0_129, RIbb31758_132,
    RIbb316e0_131, RIbb31848_134, RIbb317d0_133, RIbb31938_136,
    RIbb318c0_135, RIbb31a28_138, RIbb319b0_137, RIbb31b18_140,
    RIbb31aa0_139, RIbb31b90_141, RIbb31c08_142, RIbb31c80_143,
    RIbb31cf8_144, RIbb31d70_145, RIbb31de8_146, RIbb31e60_147,
    RIbb31ed8_148, RIbb31f50_149, RIbb31fc8_150, RIbb32040_151,
    RIbb320b8_152, RIbb32130_153, RIbb321a8_154, RIbb32220_155,
    RIbb32298_156, RIbb32310_157, RIbb32388_158, RIbb32400_159,
    RIbb32478_160, RIbb324f0_161, RIbb32568_162, RIbb325e0_163,
    RIbb32658_164, RIbb326d0_165, RIbb32748_166, RIbb327c0_167,
    RIbb32838_168, RIbb328b0_169, RIbb32928_170, RIbb329a0_171,
    RIbb32a18_172, RIbb32a90_173, RIbb32b08_174, RIbb32b80_175,
    RIbb32bf8_176, RIbb32c70_177, RIbb32ce8_178, RIbb32d60_179,
    RIbb32dd8_180, RIbb32e50_181, RIbb32ec8_182, RIbb32f40_183,
    RIbb32fb8_184, RIbb33030_185, RIbb330a8_186, RIbb33120_187,
    RIbb33198_188, RIbb33210_189, RIbb33288_190, RIbb33300_191,
    RIbb33378_192, RIbb333f0_193, RIbb33468_194, RIbb334e0_195,
    RIbb33558_196, RIbb335d0_197, RIbb33648_198, RIbb336c0_199,
    RIbb33738_200, RIbb337b0_201, RIbb33828_202, RIbb338a0_203,
    RIbb33918_204, RIbb33990_205, RIbb33a08_206, RIbb33a80_207,
    RIbb33af8_208, RIbb33b70_209, RIbb33be8_210, RIbb33c60_211,
    RIbb33cd8_212, RIbb33d50_213, RIbb33dc8_214, RIbb33e40_215,
    RIbb33eb8_216, RIbb33f30_217, RIbb33fa8_218, RIbb34020_219,
    RIbb34098_220, RIbb34110_221, RIbb34188_222, RIbb34200_223,
    RIbb34278_224, RIbb342f0_225, RIbb34368_226, RIbb343e0_227,
    RIbb34458_228, RIbb344d0_229, RIbb34548_230, RIbb345c0_231,
    RIbb34638_232, RIbb346b0_233, RIbb34728_234, RIbb347a0_235,
    RIbb34818_236, RIbb34890_237, RIbb34908_238, RIbb34980_239,
    RIbb349f8_240, RIbb34a70_241, RIbb34ae8_242, RIbb34b60_243,
    RIbb34bd8_244, RIbb34c50_245, RIbb34cc8_246, RIbb34d40_247,
    RIbb34db8_248, RIbb34e30_249, RIbb34ea8_250, RIbb34f20_251,
    RIbb34f98_252, RIbb35010_253, RIbb35088_254, RIbb35100_255,
    RIbb35178_256,
    eq  );
  input  RIbb2f070_13, RIbb2eff8_14, RIbb2ef80_15, RIbb2d798_66,
    RIbb2f160_11, RIbb2f0e8_12, RIbb2d810_65, RIbb2d6a8_68, RIbb2f250_9,
    RIbb2f1d8_10, RIbb2d720_67, RIbb2d5b8_70, RIbb2f340_7, RIbb2f2c8_8,
    RIbb2d630_69, RIbb2d4c8_72, RIbb2f430_5, RIbb2f3b8_6, RIbb2d540_71,
    RIbb2d3d8_74, RIbb2f520_3, RIbb2f4a8_4, RIbb2d450_73, RIbb2d2e8_76,
    RIbb2f610_1, RIbb2f598_2, RIbb2d360_75, RIbb2d270_77, RIbb2d1f8_78,
    RIbb2ef08_16, RIbb2ee90_17, RIbb2d180_79, RIbb2d108_80, RIbb2ee18_18,
    RIbb2eda0_19, RIbb2d090_81, RIbb2ed28_20, RIbb2ecb0_21, RIbb2d018_82,
    RIbb2cfa0_83, RIbb2cf28_84, RIbb2ec38_22, RIbb2ebc0_23, RIbb2ceb0_85,
    RIbb2ce38_86, RIbb2eb48_24, RIbb2ead0_25, RIbb2cdc0_87, RIbb2cd48_88,
    RIbb2ea58_26, RIbb2e9e0_27, RIbb2ccd0_89, RIbb2cc58_90, RIbb2e968_28,
    RIbb2e8f0_29, RIbb2cbe0_91, RIbb2cb68_92, RIbb2e878_30, RIbb2e800_31,
    RIbb2caf0_93, RIbb2ca78_94, RIbb2e788_32, RIbb2e710_33, RIbb2ca00_95,
    RIbb2c988_96, RIbb2e698_34, RIbb2e620_35, RIbb2c910_97, RIbb2c898_98,
    RIbb2e5a8_36, RIbb2e530_37, RIbb2c820_99, RIbb2e4b8_38, RIbb2e440_39,
    RIbb2c7a8_100, RIbb2c730_101, RIbb2c6b8_102, RIbb2e3c8_40,
    RIbb2e350_41, RIbb2c640_103, RIbb2c5c8_104, RIbb2e2d8_42, RIbb2e260_43,
    RIbb2c550_105, RIbb2c4d8_106, RIbb2e1e8_44, RIbb2e170_45,
    RIbb2c460_107, RIbb2c3e8_108, RIbb2e0f8_46, RIbb2e080_47,
    RIbb2c370_109, RIbb2c2f8_110, RIbb2e008_48, RIbb2df90_49,
    RIbb2c280_111, RIbb2c208_112, RIbb2df18_50, RIbb2dea0_51,
    RIbb2c190_113, RIbb2c118_114, RIbb2de28_52, RIbb2ddb0_53,
    RIbb2c0a0_115, RIbb2c028_116, RIbb2dd38_54, RIbb2dcc0_55,
    RIbb2bfb0_117, RIbb2dc48_56, RIbb2dbd0_57, RIbb2bf38_118,
    RIbb2bec0_119, RIbb2be48_120, RIbb2db58_58, RIbb2dae0_59,
    RIbb2bdd0_121, RIbb2bd58_122, RIbb2da68_60, RIbb2d9f0_61,
    RIbb2bce0_123, RIbb2bc68_124, RIbb2d978_62, RIbb2d900_63,
    RIbb2bbf0_125, RIbb2bb78_126, RIbb31500_127, RIbb2d888_64,
    RIbb31578_128, RIbb31668_130, RIbb315f0_129, RIbb31758_132,
    RIbb316e0_131, RIbb31848_134, RIbb317d0_133, RIbb31938_136,
    RIbb318c0_135, RIbb31a28_138, RIbb319b0_137, RIbb31b18_140,
    RIbb31aa0_139, RIbb31b90_141, RIbb31c08_142, RIbb31c80_143,
    RIbb31cf8_144, RIbb31d70_145, RIbb31de8_146, RIbb31e60_147,
    RIbb31ed8_148, RIbb31f50_149, RIbb31fc8_150, RIbb32040_151,
    RIbb320b8_152, RIbb32130_153, RIbb321a8_154, RIbb32220_155,
    RIbb32298_156, RIbb32310_157, RIbb32388_158, RIbb32400_159,
    RIbb32478_160, RIbb324f0_161, RIbb32568_162, RIbb325e0_163,
    RIbb32658_164, RIbb326d0_165, RIbb32748_166, RIbb327c0_167,
    RIbb32838_168, RIbb328b0_169, RIbb32928_170, RIbb329a0_171,
    RIbb32a18_172, RIbb32a90_173, RIbb32b08_174, RIbb32b80_175,
    RIbb32bf8_176, RIbb32c70_177, RIbb32ce8_178, RIbb32d60_179,
    RIbb32dd8_180, RIbb32e50_181, RIbb32ec8_182, RIbb32f40_183,
    RIbb32fb8_184, RIbb33030_185, RIbb330a8_186, RIbb33120_187,
    RIbb33198_188, RIbb33210_189, RIbb33288_190, RIbb33300_191,
    RIbb33378_192, RIbb333f0_193, RIbb33468_194, RIbb334e0_195,
    RIbb33558_196, RIbb335d0_197, RIbb33648_198, RIbb336c0_199,
    RIbb33738_200, RIbb337b0_201, RIbb33828_202, RIbb338a0_203,
    RIbb33918_204, RIbb33990_205, RIbb33a08_206, RIbb33a80_207,
    RIbb33af8_208, RIbb33b70_209, RIbb33be8_210, RIbb33c60_211,
    RIbb33cd8_212, RIbb33d50_213, RIbb33dc8_214, RIbb33e40_215,
    RIbb33eb8_216, RIbb33f30_217, RIbb33fa8_218, RIbb34020_219,
    RIbb34098_220, RIbb34110_221, RIbb34188_222, RIbb34200_223,
    RIbb34278_224, RIbb342f0_225, RIbb34368_226, RIbb343e0_227,
    RIbb34458_228, RIbb344d0_229, RIbb34548_230, RIbb345c0_231,
    RIbb34638_232, RIbb346b0_233, RIbb34728_234, RIbb347a0_235,
    RIbb34818_236, RIbb34890_237, RIbb34908_238, RIbb34980_239,
    RIbb349f8_240, RIbb34a70_241, RIbb34ae8_242, RIbb34b60_243,
    RIbb34bd8_244, RIbb34c50_245, RIbb34cc8_246, RIbb34d40_247,
    RIbb34db8_248, RIbb34e30_249, RIbb34ea8_250, RIbb34f20_251,
    RIbb34f98_252, RIbb35010_253, RIbb35088_254, RIbb35100_255,
    RIbb35178_256;
  output eq;
  wire new_n258_, new_n259_, new_n260_, new_n261_, new_n262_, new_n263_,
    new_n264_, new_n265_, new_n266_, new_n267_, new_n268_, new_n269_,
    new_n270_, new_n271_, new_n272_, new_n273_, new_n274_, new_n275_,
    new_n276_, new_n277_, new_n278_, new_n279_, new_n280_, new_n281_,
    new_n282_, new_n283_, new_n284_, new_n285_, new_n286_, new_n287_,
    new_n288_, new_n289_, new_n290_, new_n291_, new_n292_, new_n293_,
    new_n294_, new_n295_, new_n296_, new_n297_, new_n298_, new_n299_,
    new_n300_, new_n301_, new_n302_, new_n303_, new_n304_, new_n305_,
    new_n306_, new_n307_, new_n308_, new_n309_, new_n310_, new_n311_,
    new_n312_, new_n313_, new_n314_, new_n315_, new_n316_, new_n317_,
    new_n318_, new_n319_, new_n320_, new_n321_, new_n322_, new_n323_,
    new_n324_, new_n325_, new_n326_, new_n327_, new_n328_, new_n329_,
    new_n330_, new_n331_, new_n332_, new_n333_, new_n334_, new_n335_,
    new_n336_, new_n337_, new_n338_, new_n339_, new_n340_, new_n341_,
    new_n342_, new_n343_, new_n344_, new_n345_, new_n346_, new_n347_,
    new_n348_, new_n349_, new_n350_, new_n351_, new_n352_, new_n353_,
    new_n354_, new_n355_, new_n356_, new_n357_, new_n358_, new_n359_,
    new_n360_, new_n361_, new_n362_, new_n363_, new_n364_, new_n365_,
    new_n366_, new_n367_, new_n368_, new_n369_, new_n370_, new_n371_,
    new_n372_, new_n373_, new_n374_, new_n375_, new_n376_, new_n377_,
    new_n378_, new_n379_, new_n380_, new_n381_, new_n382_, new_n383_,
    new_n384_, new_n385_, new_n386_, new_n387_, new_n388_, new_n389_,
    new_n390_, new_n391_, new_n392_, new_n393_, new_n394_, new_n395_,
    new_n396_, new_n397_, new_n398_, new_n399_, new_n400_, new_n401_,
    new_n402_, new_n403_, new_n404_, new_n405_, new_n406_, new_n407_,
    new_n408_, new_n409_, new_n410_, new_n411_, new_n412_, new_n413_,
    new_n414_, new_n415_, new_n416_, new_n417_, new_n418_, new_n419_,
    new_n420_, new_n421_, new_n422_, new_n423_, new_n424_, new_n425_,
    new_n426_, new_n427_, new_n428_, new_n429_, new_n430_, new_n431_,
    new_n432_, new_n433_, new_n434_, new_n435_, new_n436_, new_n437_,
    new_n438_, new_n439_, new_n440_, new_n441_, new_n442_, new_n443_,
    new_n444_, new_n445_, new_n446_, new_n447_, new_n448_, new_n449_,
    new_n450_, new_n451_, new_n452_, new_n453_, new_n454_, new_n455_,
    new_n456_, new_n457_, new_n458_, new_n459_, new_n460_, new_n461_,
    new_n462_, new_n463_, new_n464_, new_n465_, new_n466_, new_n467_,
    new_n468_, new_n469_, new_n470_, new_n471_, new_n472_, new_n473_,
    new_n474_, new_n475_, new_n476_, new_n477_, new_n478_, new_n479_,
    new_n480_, new_n481_, new_n482_, new_n483_, new_n484_, new_n485_,
    new_n486_, new_n487_, new_n488_, new_n489_, new_n490_, new_n491_,
    new_n492_, new_n493_, new_n494_, new_n495_, new_n496_, new_n497_,
    new_n498_, new_n499_, new_n500_, new_n501_, new_n502_, new_n503_,
    new_n504_, new_n505_, new_n506_, new_n507_, new_n508_, new_n509_,
    new_n510_, new_n511_, new_n512_, new_n513_, new_n514_, new_n515_,
    new_n516_, new_n517_, new_n518_, new_n519_, new_n520_, new_n521_,
    new_n522_, new_n523_, new_n524_, new_n525_, new_n526_, new_n527_,
    new_n528_, new_n529_, new_n530_, new_n531_, new_n532_, new_n533_,
    new_n534_, new_n535_, new_n536_, new_n537_, new_n538_, new_n539_,
    new_n540_, new_n541_, new_n542_, new_n543_, new_n544_, new_n545_,
    new_n546_, new_n547_, new_n548_, new_n549_, new_n550_, new_n551_,
    new_n552_, new_n553_, new_n554_, new_n555_, new_n556_, new_n557_,
    new_n558_, new_n559_, new_n560_, new_n561_, new_n562_, new_n563_,
    new_n564_, new_n565_, new_n566_, new_n567_, new_n568_, new_n569_,
    new_n570_, new_n571_, new_n572_, new_n573_, new_n574_, new_n575_,
    new_n576_, new_n577_, new_n578_, new_n579_, new_n580_, new_n581_,
    new_n582_, new_n583_, new_n584_, new_n585_, new_n586_, new_n587_,
    new_n588_, new_n589_, new_n590_, new_n591_, new_n592_, new_n593_,
    new_n594_, new_n595_, new_n596_, new_n597_, new_n598_, new_n599_,
    new_n600_, new_n601_, new_n602_, new_n603_, new_n604_, new_n605_,
    new_n606_, new_n607_, new_n608_, new_n609_, new_n610_, new_n611_,
    new_n612_, new_n613_, new_n614_, new_n615_, new_n616_, new_n617_,
    new_n618_, new_n619_, new_n620_, new_n621_, new_n622_, new_n623_,
    new_n624_, new_n625_, new_n626_, new_n627_, new_n628_, new_n629_,
    new_n630_, new_n631_, new_n632_, new_n633_, new_n634_, new_n635_,
    new_n636_, new_n637_, new_n638_, new_n639_, new_n640_, new_n641_,
    new_n642_, new_n643_, new_n644_, new_n645_, new_n646_, new_n647_,
    new_n648_, new_n649_, new_n650_, new_n651_, new_n652_, new_n653_,
    new_n654_, new_n655_, new_n656_, new_n657_, new_n658_, new_n659_,
    new_n660_, new_n661_, new_n662_, new_n663_, new_n664_, new_n665_,
    new_n666_, new_n667_, new_n668_, new_n669_, new_n670_, new_n671_,
    new_n672_, new_n673_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n680_, new_n681_, new_n682_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n771_, new_n772_, new_n773_,
    new_n774_, new_n775_, new_n776_, new_n777_, new_n778_, new_n779_,
    new_n780_, new_n781_, new_n782_, new_n783_, new_n784_, new_n785_,
    new_n786_, new_n787_, new_n788_, new_n789_, new_n790_, new_n791_,
    new_n792_, new_n793_, new_n794_, new_n795_, new_n796_, new_n797_,
    new_n798_, new_n799_, new_n800_, new_n801_, new_n802_, new_n803_,
    new_n804_, new_n805_, new_n806_, new_n807_, new_n808_, new_n809_,
    new_n810_, new_n811_, new_n812_, new_n813_, new_n814_, new_n815_,
    new_n816_, new_n817_, new_n818_, new_n819_, new_n820_, new_n821_,
    new_n822_, new_n823_, new_n824_, new_n825_, new_n826_, new_n827_,
    new_n828_, new_n829_, new_n830_, new_n831_, new_n832_, new_n833_,
    new_n834_, new_n835_, new_n836_, new_n837_, new_n838_, new_n839_,
    new_n840_, new_n841_, new_n842_, new_n843_, new_n844_, new_n845_,
    new_n846_, new_n847_, new_n848_, new_n849_, new_n850_, new_n851_,
    new_n852_, new_n853_, new_n854_, new_n855_, new_n856_, new_n857_,
    new_n858_, new_n859_, new_n860_, new_n861_, new_n862_, new_n863_,
    new_n864_, new_n865_, new_n866_, new_n867_, new_n868_, new_n869_,
    new_n870_, new_n871_, new_n872_, new_n873_, new_n874_, new_n875_,
    new_n876_, new_n877_, new_n878_, new_n879_, new_n880_, new_n881_,
    new_n882_, new_n883_, new_n884_, new_n885_, new_n886_, new_n887_,
    new_n888_, new_n889_, new_n890_, new_n891_, new_n892_, new_n893_,
    new_n894_, new_n895_, new_n896_, new_n897_, new_n898_, new_n899_,
    new_n900_, new_n901_, new_n902_, new_n903_, new_n904_, new_n905_,
    new_n906_, new_n907_, new_n908_, new_n909_, new_n910_, new_n911_,
    new_n912_, new_n913_, new_n914_, new_n915_, new_n916_, new_n917_,
    new_n918_, new_n919_, new_n920_, new_n921_, new_n922_, new_n923_,
    new_n924_, new_n925_, new_n926_, new_n927_, new_n928_, new_n929_,
    new_n930_, new_n931_, new_n932_, new_n933_, new_n934_, new_n935_,
    new_n936_, new_n937_, new_n938_, new_n939_, new_n940_, new_n941_,
    new_n942_, new_n943_, new_n944_, new_n945_, new_n946_, new_n947_,
    new_n948_, new_n949_, new_n950_, new_n951_, new_n952_, new_n953_,
    new_n954_, new_n955_, new_n956_, new_n957_, new_n958_, new_n959_,
    new_n960_, new_n961_, new_n962_, new_n963_, new_n964_, new_n965_,
    new_n966_, new_n967_, new_n968_, new_n969_, new_n970_, new_n971_,
    new_n972_, new_n973_, new_n974_, new_n975_, new_n976_, new_n977_,
    new_n978_, new_n979_, new_n980_, new_n981_, new_n982_, new_n983_,
    new_n984_, new_n985_, new_n986_, new_n987_, new_n988_, new_n989_,
    new_n990_, new_n991_, new_n992_, new_n993_, new_n994_, new_n995_,
    new_n996_, new_n997_, new_n998_, new_n999_, new_n1000_, new_n1001_,
    new_n1002_, new_n1003_, new_n1004_, new_n1005_, new_n1006_, new_n1007_,
    new_n1008_, new_n1009_, new_n1010_, new_n1011_, new_n1012_, new_n1013_,
    new_n1014_, new_n1015_, new_n1016_, new_n1017_, new_n1018_, new_n1019_,
    new_n1020_, new_n1021_, new_n1022_, new_n1023_, new_n1024_, new_n1025_,
    new_n1026_, new_n1027_, new_n1028_, new_n1029_, new_n1030_, new_n1031_,
    new_n1032_, new_n1033_, new_n1034_, new_n1035_, new_n1036_, new_n1037_,
    new_n1038_, new_n1039_, new_n1040_, new_n1041_, new_n1042_, new_n1043_,
    new_n1044_, new_n1045_, new_n1046_, new_n1047_, new_n1048_, new_n1049_,
    new_n1050_, new_n1051_, new_n1052_, new_n1053_, new_n1054_, new_n1055_,
    new_n1056_, new_n1057_, new_n1058_, new_n1059_, new_n1060_, new_n1061_,
    new_n1062_, new_n1063_, new_n1064_, new_n1065_, new_n1066_, new_n1067_,
    new_n1068_, new_n1069_, new_n1070_, new_n1071_, new_n1072_, new_n1073_,
    new_n1074_, new_n1075_, new_n1076_, new_n1077_, new_n1078_, new_n1079_,
    new_n1080_, new_n1081_, new_n1082_, new_n1083_, new_n1084_, new_n1085_,
    new_n1086_, new_n1087_, new_n1088_, new_n1089_, new_n1090_, new_n1091_,
    new_n1092_, new_n1093_, new_n1094_, new_n1095_, new_n1096_, new_n1097_,
    new_n1098_, new_n1099_, new_n1100_, new_n1101_, new_n1102_, new_n1103_,
    new_n1104_, new_n1105_, new_n1106_, new_n1107_, new_n1108_, new_n1109_,
    new_n1110_, new_n1111_, new_n1112_, new_n1113_, new_n1114_, new_n1115_,
    new_n1116_, new_n1117_, new_n1118_, new_n1119_, new_n1120_, new_n1121_,
    new_n1122_, new_n1123_, new_n1124_, new_n1125_, new_n1126_, new_n1127_,
    new_n1128_, new_n1129_, new_n1130_, new_n1131_, new_n1132_, new_n1133_,
    new_n1134_, new_n1135_, new_n1136_, new_n1137_, new_n1138_, new_n1139_,
    new_n1140_, new_n1141_, new_n1142_, new_n1143_, new_n1144_, new_n1145_,
    new_n1146_, new_n1147_, new_n1148_, new_n1149_, new_n1150_, new_n1151_,
    new_n1152_, new_n1153_, new_n1154_, new_n1155_, new_n1156_, new_n1157_,
    new_n1158_, new_n1159_, new_n1160_, new_n1161_, new_n1162_, new_n1163_,
    new_n1164_, new_n1165_, new_n1166_, new_n1167_, new_n1168_, new_n1169_,
    new_n1170_, new_n1171_, new_n1172_, new_n1173_, new_n1174_, new_n1175_,
    new_n1176_, new_n1177_, new_n1178_, new_n1179_, new_n1180_, new_n1181_,
    new_n1182_, new_n1183_, new_n1184_, new_n1185_, new_n1186_, new_n1187_,
    new_n1188_, new_n1189_, new_n1190_, new_n1191_, new_n1192_, new_n1193_,
    new_n1194_, new_n1195_, new_n1196_, new_n1197_, new_n1198_, new_n1199_,
    new_n1200_, new_n1201_, new_n1202_, new_n1203_, new_n1204_, new_n1205_,
    new_n1206_, new_n1207_, new_n1208_, new_n1209_, new_n1210_, new_n1211_,
    new_n1212_, new_n1213_, new_n1214_, new_n1215_, new_n1216_, new_n1217_,
    new_n1218_, new_n1219_, new_n1220_, new_n1221_, new_n1222_, new_n1223_,
    new_n1224_, new_n1225_, new_n1226_, new_n1227_, new_n1228_, new_n1229_,
    new_n1230_, new_n1231_, new_n1232_, new_n1233_, new_n1234_, new_n1235_,
    new_n1236_, new_n1237_, new_n1238_, new_n1239_, new_n1240_, new_n1241_,
    new_n1242_, new_n1243_, new_n1244_, new_n1245_, new_n1246_, new_n1247_,
    new_n1248_, new_n1249_, new_n1250_, new_n1251_, new_n1252_, new_n1253_,
    new_n1254_, new_n1255_, new_n1256_, new_n1257_, new_n1258_, new_n1259_,
    new_n1260_, new_n1261_, new_n1262_, new_n1263_, new_n1264_, new_n1265_,
    new_n1266_, new_n1267_, new_n1268_, new_n1269_, new_n1270_, new_n1271_,
    new_n1272_, new_n1273_, new_n1274_, new_n1275_, new_n1276_, new_n1277_,
    new_n1278_, new_n1279_, new_n1280_, new_n1281_, new_n1282_, new_n1283_,
    new_n1284_, new_n1285_, new_n1286_, new_n1287_, new_n1288_, new_n1289_,
    new_n1290_, new_n1291_, new_n1292_, new_n1293_, new_n1294_, new_n1295_,
    new_n1296_, new_n1297_, new_n1298_, new_n1299_, new_n1300_, new_n1301_,
    new_n1302_, new_n1303_, new_n1304_, new_n1305_, new_n1306_, new_n1307_,
    new_n1308_, new_n1309_, new_n1310_, new_n1311_, new_n1312_, new_n1313_,
    new_n1314_, new_n1315_, new_n1316_, new_n1317_, new_n1318_, new_n1319_,
    new_n1320_, new_n1321_, new_n1322_, new_n1323_, new_n1324_, new_n1325_,
    new_n1326_, new_n1327_, new_n1328_, new_n1329_, new_n1330_, new_n1331_,
    new_n1332_, new_n1333_, new_n1334_, new_n1335_, new_n1336_, new_n1337_,
    new_n1338_, new_n1339_, new_n1340_, new_n1341_, new_n1342_, new_n1343_,
    new_n1344_, new_n1345_, new_n1346_, new_n1347_, new_n1348_, new_n1349_,
    new_n1350_, new_n1351_, new_n1352_, new_n1353_, new_n1354_, new_n1355_,
    new_n1356_, new_n1357_, new_n1358_, new_n1359_, new_n1360_, new_n1361_,
    new_n1362_, new_n1363_, new_n1364_, new_n1365_, new_n1366_, new_n1367_,
    new_n1368_, new_n1369_, new_n1370_, new_n1371_, new_n1372_, new_n1373_,
    new_n1374_, new_n1375_, new_n1376_, new_n1377_, new_n1378_, new_n1379_,
    new_n1380_, new_n1381_, new_n1382_, new_n1383_, new_n1384_, new_n1385_,
    new_n1386_, new_n1387_, new_n1388_, new_n1389_, new_n1390_, new_n1391_,
    new_n1392_, new_n1393_, new_n1394_, new_n1395_, new_n1396_, new_n1397_,
    new_n1398_, new_n1399_, new_n1400_, new_n1401_, new_n1402_, new_n1403_,
    new_n1404_, new_n1405_, new_n1406_, new_n1407_, new_n1408_, new_n1409_,
    new_n1410_, new_n1411_, new_n1412_, new_n1413_, new_n1414_, new_n1415_,
    new_n1416_, new_n1417_, new_n1418_, new_n1419_, new_n1420_, new_n1421_,
    new_n1422_, new_n1423_, new_n1424_, new_n1425_, new_n1426_, new_n1427_,
    new_n1428_, new_n1429_, new_n1430_, new_n1431_, new_n1432_, new_n1433_,
    new_n1434_, new_n1435_, new_n1436_, new_n1437_, new_n1438_, new_n1439_,
    new_n1440_, new_n1441_, new_n1442_, new_n1443_, new_n1444_, new_n1445_,
    new_n1446_, new_n1447_, new_n1448_, new_n1449_, new_n1450_, new_n1451_,
    new_n1452_, new_n1453_, new_n1454_, new_n1455_, new_n1456_, new_n1457_,
    new_n1458_, new_n1459_, new_n1460_, new_n1461_, new_n1462_, new_n1463_,
    new_n1464_, new_n1465_, new_n1466_, new_n1467_, new_n1468_, new_n1469_,
    new_n1470_, new_n1471_, new_n1472_, new_n1473_, new_n1474_, new_n1475_,
    new_n1476_, new_n1477_, new_n1478_, new_n1479_, new_n1480_, new_n1481_,
    new_n1482_, new_n1483_, new_n1484_, new_n1485_, new_n1486_, new_n1487_,
    new_n1488_, new_n1489_, new_n1490_, new_n1491_, new_n1492_, new_n1493_,
    new_n1494_, new_n1495_, new_n1496_, new_n1497_, new_n1498_, new_n1499_,
    new_n1500_, new_n1501_, new_n1502_, new_n1503_, new_n1504_, new_n1505_,
    new_n1506_, new_n1507_, new_n1508_, new_n1509_, new_n1510_, new_n1511_,
    new_n1512_, new_n1513_, new_n1514_, new_n1515_, new_n1516_, new_n1517_,
    new_n1518_, new_n1519_, new_n1520_, new_n1521_, new_n1522_, new_n1523_,
    new_n1524_, new_n1525_, new_n1526_, new_n1527_, new_n1528_, new_n1529_,
    new_n1530_, new_n1531_, new_n1532_, new_n1533_, new_n1534_, new_n1535_,
    new_n1536_, new_n1537_, new_n1538_, new_n1539_, new_n1540_, new_n1541_,
    new_n1542_, new_n1543_, new_n1544_, new_n1545_, new_n1546_, new_n1547_,
    new_n1548_, new_n1549_, new_n1550_, new_n1551_, new_n1552_, new_n1553_,
    new_n1554_, new_n1555_, new_n1556_, new_n1557_, new_n1558_, new_n1559_,
    new_n1560_, new_n1561_, new_n1562_, new_n1563_, new_n1564_, new_n1565_,
    new_n1566_, new_n1567_, new_n1568_, new_n1569_, new_n1570_, new_n1571_,
    new_n1572_, new_n1573_, new_n1574_, new_n1575_, new_n1576_, new_n1577_,
    new_n1578_, new_n1579_, new_n1580_, new_n1581_, new_n1582_, new_n1583_,
    new_n1584_, new_n1585_, new_n1586_, new_n1587_, new_n1588_, new_n1589_,
    new_n1590_, new_n1591_, new_n1592_, new_n1593_, new_n1594_, new_n1595_,
    new_n1596_, new_n1597_, new_n1598_, new_n1599_, new_n1600_, new_n1601_,
    new_n1602_, new_n1603_, new_n1604_, new_n1605_, new_n1606_, new_n1607_,
    new_n1608_, new_n1609_, new_n1610_, new_n1611_, new_n1612_, new_n1613_,
    new_n1614_, new_n1615_, new_n1616_, new_n1617_, new_n1618_, new_n1619_,
    new_n1620_, new_n1621_, new_n1622_, new_n1623_, new_n1624_, new_n1625_,
    new_n1626_, new_n1627_, new_n1628_, new_n1629_, new_n1630_, new_n1631_,
    new_n1632_, new_n1633_, new_n1634_, new_n1635_, new_n1636_, new_n1637_,
    new_n1638_, new_n1639_, new_n1640_, new_n1641_, new_n1642_, new_n1643_,
    new_n1644_, new_n1645_, new_n1646_, new_n1647_, new_n1648_, new_n1649_,
    new_n1650_, new_n1651_, new_n1652_, new_n1653_, new_n1654_, new_n1655_,
    new_n1656_, new_n1657_, new_n1658_, new_n1659_, new_n1660_, new_n1661_,
    new_n1662_, new_n1663_, new_n1664_, new_n1665_, new_n1666_, new_n1667_,
    new_n1668_, new_n1669_, new_n1670_, new_n1671_, new_n1672_, new_n1673_,
    new_n1674_, new_n1675_, new_n1676_, new_n1677_, new_n1678_, new_n1679_,
    new_n1680_, new_n1681_, new_n1682_, new_n1683_, new_n1684_, new_n1685_,
    new_n1686_, new_n1687_, new_n1688_, new_n1689_, new_n1690_, new_n1691_,
    new_n1692_, new_n1693_, new_n1694_, new_n1695_, new_n1696_, new_n1697_,
    new_n1698_, new_n1699_, new_n1700_, new_n1701_, new_n1702_, new_n1703_,
    new_n1704_, new_n1705_, new_n1706_, new_n1707_, new_n1708_, new_n1709_,
    new_n1710_, new_n1711_, new_n1712_, new_n1713_, new_n1714_, new_n1715_,
    new_n1716_, new_n1717_, new_n1718_, new_n1719_, new_n1720_, new_n1721_,
    new_n1722_, new_n1723_, new_n1724_, new_n1725_, new_n1726_, new_n1727_,
    new_n1728_, new_n1729_, new_n1730_, new_n1731_, new_n1732_, new_n1733_,
    new_n1734_, new_n1735_, new_n1736_, new_n1737_, new_n1738_, new_n1739_,
    new_n1740_, new_n1741_, new_n1742_, new_n1743_, new_n1744_, new_n1745_,
    new_n1746_, new_n1747_, new_n1748_, new_n1749_, new_n1750_, new_n1751_,
    new_n1752_, new_n1753_, new_n1754_, new_n1755_, new_n1756_, new_n1757_,
    new_n1758_, new_n1759_, new_n1760_, new_n1761_, new_n1762_, new_n1763_,
    new_n1764_, new_n1765_, new_n1766_, new_n1767_, new_n1768_, new_n1769_,
    new_n1770_, new_n1771_, new_n1772_, new_n1773_, new_n1774_, new_n1775_,
    new_n1776_, new_n1777_, new_n1778_, new_n1779_, new_n1780_, new_n1781_,
    new_n1782_, new_n1783_, new_n1784_, new_n1785_, new_n1786_, new_n1787_,
    new_n1788_, new_n1789_, new_n1790_, new_n1791_, new_n1792_, new_n1793_,
    new_n1794_, new_n1795_, new_n1796_, new_n1797_, new_n1798_, new_n1799_,
    new_n1800_, new_n1801_, new_n1802_, new_n1803_, new_n1804_, new_n1805_,
    new_n1806_, new_n1807_, new_n1808_, new_n1809_, new_n1810_, new_n1811_,
    new_n1812_, new_n1813_, new_n1814_, new_n1815_, new_n1816_, new_n1817_,
    new_n1818_, new_n1819_, new_n1820_, new_n1821_, new_n1822_, new_n1823_,
    new_n1824_, new_n1825_, new_n1826_, new_n1827_, new_n1828_, new_n1829_,
    new_n1830_, new_n1831_, new_n1832_, new_n1833_, new_n1834_, new_n1835_,
    new_n1836_, new_n1837_, new_n1838_, new_n1839_, new_n1840_, new_n1841_,
    new_n1842_, new_n1843_, new_n1844_, new_n1845_, new_n1846_, new_n1847_,
    new_n1848_, new_n1849_, new_n1850_, new_n1851_, new_n1852_, new_n1853_,
    new_n1854_, new_n1855_, new_n1856_, new_n1857_, new_n1858_, new_n1859_,
    new_n1860_, new_n1861_, new_n1862_, new_n1863_, new_n1864_, new_n1865_,
    new_n1866_, new_n1867_, new_n1868_, new_n1869_, new_n1870_, new_n1871_,
    new_n1872_, new_n1873_, new_n1874_, new_n1875_, new_n1876_, new_n1877_,
    new_n1878_, new_n1879_, new_n1880_, new_n1881_, new_n1882_, new_n1883_,
    new_n1884_, new_n1885_, new_n1886_, new_n1887_, new_n1888_, new_n1889_,
    new_n1890_, new_n1891_, new_n1892_, new_n1893_, new_n1894_, new_n1895_,
    new_n1896_, new_n1897_, new_n1898_, new_n1899_, new_n1900_, new_n1901_,
    new_n1902_, new_n1903_, new_n1904_, new_n1905_, new_n1906_, new_n1907_,
    new_n1908_, new_n1909_, new_n1910_, new_n1911_, new_n1912_, new_n1913_,
    new_n1914_, new_n1915_, new_n1916_, new_n1917_, new_n1918_, new_n1919_,
    new_n1920_, new_n1921_, new_n1922_, new_n1923_, new_n1924_, new_n1925_,
    new_n1926_, new_n1927_, new_n1928_, new_n1929_, new_n1930_, new_n1931_,
    new_n1932_, new_n1933_, new_n1934_, new_n1935_, new_n1936_, new_n1937_,
    new_n1938_, new_n1939_, new_n1940_, new_n1941_, new_n1942_, new_n1943_,
    new_n1944_, new_n1945_, new_n1946_, new_n1947_, new_n1948_, new_n1949_,
    new_n1950_, new_n1951_, new_n1952_, new_n1953_, new_n1954_, new_n1955_,
    new_n1956_, new_n1957_, new_n1958_, new_n1959_, new_n1960_, new_n1961_,
    new_n1962_, new_n1963_, new_n1964_, new_n1965_, new_n1966_, new_n1967_,
    new_n1968_, new_n1969_, new_n1970_, new_n1971_, new_n1972_, new_n1973_,
    new_n1974_, new_n1975_, new_n1976_, new_n1977_, new_n1978_, new_n1979_,
    new_n1980_, new_n1981_, new_n1982_, new_n1983_, new_n1984_, new_n1985_,
    new_n1986_, new_n1987_, new_n1988_, new_n1989_, new_n1990_, new_n1991_,
    new_n1992_, new_n1993_, new_n1994_, new_n1995_, new_n1996_, new_n1997_,
    new_n1998_, new_n1999_, new_n2000_, new_n2001_, new_n2002_, new_n2003_,
    new_n2004_, new_n2005_, new_n2006_, new_n2007_, new_n2008_, new_n2009_,
    new_n2010_, new_n2011_, new_n2012_, new_n2013_, new_n2014_, new_n2015_,
    new_n2016_, new_n2017_, new_n2018_, new_n2019_, new_n2020_, new_n2021_,
    new_n2022_, new_n2023_, new_n2024_, new_n2025_, new_n2026_, new_n2027_,
    new_n2028_, new_n2029_, new_n2030_, new_n2031_, new_n2032_, new_n2033_,
    new_n2034_, new_n2035_, new_n2036_, new_n2037_, new_n2038_, new_n2039_,
    new_n2040_, new_n2041_, new_n2042_, new_n2043_, new_n2044_, new_n2045_,
    new_n2046_, new_n2047_, new_n2048_, new_n2049_, new_n2050_, new_n2051_,
    new_n2052_, new_n2053_, new_n2054_, new_n2055_, new_n2056_, new_n2057_,
    new_n2058_, new_n2059_, new_n2060_, new_n2061_, new_n2062_, new_n2063_,
    new_n2064_, new_n2065_, new_n2066_, new_n2067_, new_n2068_, new_n2069_,
    new_n2070_, new_n2071_, new_n2072_, new_n2073_, new_n2074_, new_n2075_,
    new_n2076_, new_n2077_, new_n2078_, new_n2079_, new_n2080_, new_n2081_,
    new_n2082_, new_n2083_, new_n2084_, new_n2085_, new_n2086_, new_n2087_,
    new_n2088_, new_n2089_, new_n2090_, new_n2091_, new_n2092_, new_n2093_,
    new_n2094_, new_n2095_, new_n2096_, new_n2097_, new_n2098_, new_n2099_,
    new_n2100_, new_n2101_, new_n2102_, new_n2103_, new_n2104_, new_n2105_,
    new_n2106_, new_n2107_, new_n2108_, new_n2109_, new_n2110_, new_n2111_,
    new_n2112_, new_n2113_, new_n2114_, new_n2115_, new_n2116_, new_n2117_,
    new_n2118_, new_n2119_, new_n2120_, new_n2121_, new_n2122_, new_n2123_,
    new_n2124_, new_n2125_, new_n2126_, new_n2127_, new_n2128_, new_n2129_,
    new_n2130_, new_n2131_, new_n2132_, new_n2133_, new_n2134_, new_n2135_,
    new_n2136_, new_n2137_, new_n2138_, new_n2139_, new_n2140_, new_n2141_,
    new_n2142_, new_n2143_, new_n2144_, new_n2145_, new_n2146_, new_n2147_,
    new_n2148_, new_n2149_, new_n2150_, new_n2151_, new_n2152_, new_n2153_,
    new_n2154_, new_n2155_, new_n2156_, new_n2157_, new_n2158_, new_n2159_,
    new_n2160_, new_n2161_, new_n2162_, new_n2163_, new_n2164_, new_n2165_,
    new_n2166_, new_n2167_, new_n2168_, new_n2169_, new_n2170_, new_n2171_,
    new_n2172_, new_n2173_, new_n2174_, new_n2175_, new_n2176_, new_n2177_,
    new_n2178_, new_n2179_, new_n2180_, new_n2181_, new_n2182_, new_n2183_,
    new_n2184_, new_n2185_, new_n2186_, new_n2187_, new_n2188_, new_n2189_,
    new_n2190_, new_n2191_, new_n2192_, new_n2193_, new_n2194_, new_n2195_,
    new_n2196_, new_n2197_, new_n2198_, new_n2199_, new_n2200_, new_n2201_,
    new_n2202_, new_n2203_, new_n2204_, new_n2205_, new_n2206_, new_n2207_,
    new_n2208_, new_n2209_, new_n2210_, new_n2211_, new_n2212_, new_n2213_,
    new_n2214_, new_n2215_, new_n2216_, new_n2217_, new_n2218_, new_n2219_,
    new_n2220_, new_n2221_, new_n2222_, new_n2223_, new_n2224_, new_n2225_,
    new_n2226_, new_n2227_, new_n2228_, new_n2229_, new_n2230_, new_n2231_,
    new_n2232_, new_n2233_, new_n2234_, new_n2235_, new_n2236_, new_n2237_,
    new_n2238_, new_n2239_, new_n2240_, new_n2241_, new_n2242_, new_n2243_,
    new_n2244_, new_n2245_, new_n2246_, new_n2247_, new_n2248_, new_n2249_,
    new_n2250_, new_n2251_, new_n2252_, new_n2253_, new_n2254_, new_n2255_,
    new_n2256_, new_n2257_, new_n2258_, new_n2259_, new_n2260_, new_n2261_,
    new_n2262_, new_n2263_, new_n2264_, new_n2265_, new_n2266_, new_n2267_,
    new_n2268_, new_n2269_, new_n2270_, new_n2271_, new_n2272_, new_n2273_,
    new_n2274_, new_n2275_, new_n2276_, new_n2277_, new_n2278_, new_n2279_,
    new_n2280_, new_n2281_, new_n2282_, new_n2283_, new_n2284_, new_n2285_,
    new_n2286_, new_n2287_, new_n2288_, new_n2289_, new_n2290_, new_n2291_,
    new_n2292_, new_n2293_, new_n2294_, new_n2295_, new_n2296_, new_n2297_,
    new_n2298_, new_n2299_, new_n2300_, new_n2301_, new_n2302_, new_n2303_,
    new_n2304_, new_n2305_, new_n2306_, new_n2307_, new_n2308_, new_n2309_,
    new_n2310_, new_n2311_, new_n2312_, new_n2313_, new_n2314_, new_n2315_,
    new_n2316_, new_n2317_, new_n2318_, new_n2319_, new_n2320_, new_n2321_,
    new_n2322_, new_n2323_, new_n2324_, new_n2325_, new_n2326_, new_n2327_,
    new_n2328_, new_n2329_, new_n2330_, new_n2331_, new_n2332_, new_n2333_,
    new_n2334_, new_n2335_, new_n2336_, new_n2337_, new_n2338_, new_n2339_,
    new_n2340_, new_n2341_, new_n2342_, new_n2343_, new_n2344_, new_n2345_,
    new_n2346_, new_n2347_, new_n2348_, new_n2349_, new_n2350_, new_n2351_,
    new_n2352_, new_n2353_, new_n2354_, new_n2355_, new_n2356_, new_n2357_,
    new_n2358_, new_n2359_, new_n2360_, new_n2361_, new_n2362_, new_n2363_,
    new_n2364_, new_n2365_, new_n2366_, new_n2367_, new_n2368_, new_n2369_,
    new_n2370_, new_n2371_, new_n2372_, new_n2373_, new_n2374_, new_n2375_,
    new_n2376_, new_n2377_, new_n2378_, new_n2379_, new_n2380_, new_n2381_,
    new_n2382_, new_n2383_, new_n2384_, new_n2385_, new_n2386_, new_n2387_,
    new_n2388_, new_n2389_, new_n2390_, new_n2391_, new_n2392_, new_n2393_,
    new_n2394_, new_n2395_, new_n2396_, new_n2397_, new_n2398_, new_n2399_,
    new_n2400_, new_n2401_, new_n2402_, new_n2403_, new_n2404_, new_n2405_,
    new_n2406_, new_n2407_, new_n2408_, new_n2409_, new_n2410_, new_n2411_,
    new_n2412_, new_n2413_, new_n2414_, new_n2415_, new_n2416_, new_n2417_,
    new_n2418_, new_n2419_, new_n2420_, new_n2421_, new_n2422_, new_n2423_,
    new_n2424_, new_n2425_, new_n2426_, new_n2427_, new_n2428_, new_n2429_,
    new_n2430_, new_n2431_, new_n2432_, new_n2433_, new_n2434_, new_n2435_,
    new_n2436_, new_n2437_, new_n2438_, new_n2439_, new_n2440_, new_n2441_,
    new_n2442_, new_n2443_, new_n2444_, new_n2445_, new_n2446_, new_n2447_,
    new_n2448_, new_n2449_, new_n2450_, new_n2451_, new_n2452_, new_n2453_,
    new_n2454_, new_n2455_, new_n2456_, new_n2457_, new_n2458_, new_n2459_,
    new_n2460_, new_n2461_, new_n2462_, new_n2463_, new_n2464_, new_n2465_,
    new_n2466_, new_n2467_, new_n2468_, new_n2469_, new_n2470_, new_n2471_,
    new_n2472_, new_n2473_, new_n2474_, new_n2475_, new_n2476_, new_n2477_,
    new_n2478_, new_n2479_, new_n2480_, new_n2481_, new_n2482_, new_n2483_,
    new_n2484_, new_n2485_, new_n2486_, new_n2487_, new_n2488_, new_n2489_,
    new_n2490_, new_n2491_, new_n2492_, new_n2493_, new_n2494_, new_n2495_,
    new_n2496_, new_n2497_, new_n2498_, new_n2499_, new_n2500_, new_n2501_,
    new_n2502_, new_n2503_, new_n2504_, new_n2505_, new_n2506_, new_n2507_,
    new_n2508_, new_n2509_, new_n2510_, new_n2511_, new_n2512_, new_n2513_,
    new_n2514_, new_n2515_, new_n2516_, new_n2517_, new_n2518_, new_n2519_,
    new_n2520_, new_n2521_, new_n2522_, new_n2523_, new_n2524_, new_n2525_,
    new_n2526_, new_n2527_, new_n2528_, new_n2529_, new_n2530_, new_n2531_,
    new_n2532_, new_n2533_, new_n2534_, new_n2535_, new_n2536_, new_n2537_,
    new_n2538_, new_n2539_, new_n2540_, new_n2541_, new_n2542_, new_n2543_,
    new_n2544_, new_n2545_, new_n2546_, new_n2547_, new_n2548_, new_n2549_,
    new_n2550_, new_n2551_, new_n2552_, new_n2553_, new_n2554_, new_n2555_,
    new_n2556_, new_n2557_, new_n2558_, new_n2559_, new_n2560_, new_n2561_,
    new_n2562_, new_n2563_, new_n2564_, new_n2565_, new_n2566_, new_n2567_,
    new_n2568_, new_n2569_, new_n2570_, new_n2571_, new_n2572_, new_n2573_,
    new_n2574_, new_n2575_, new_n2576_, new_n2577_, new_n2578_, new_n2579_,
    new_n2580_, new_n2581_, new_n2582_, new_n2583_, new_n2584_, new_n2585_,
    new_n2586_, new_n2587_, new_n2588_, new_n2589_, new_n2590_, new_n2591_,
    new_n2592_, new_n2593_, new_n2594_, new_n2595_, new_n2596_, new_n2597_,
    new_n2598_, new_n2599_, new_n2600_, new_n2601_, new_n2602_, new_n2603_,
    new_n2604_, new_n2605_, new_n2606_, new_n2607_, new_n2608_, new_n2609_,
    new_n2610_, new_n2611_, new_n2612_, new_n2613_, new_n2614_, new_n2615_,
    new_n2616_, new_n2617_, new_n2618_, new_n2619_, new_n2620_, new_n2621_,
    new_n2622_, new_n2623_, new_n2624_, new_n2625_, new_n2626_, new_n2627_,
    new_n2628_, new_n2629_, new_n2630_, new_n2631_, new_n2632_, new_n2633_,
    new_n2634_, new_n2635_, new_n2636_, new_n2637_, new_n2638_, new_n2639_,
    new_n2640_, new_n2641_, new_n2642_, new_n2643_, new_n2644_, new_n2645_,
    new_n2646_, new_n2647_, new_n2648_, new_n2649_, new_n2650_, new_n2651_,
    new_n2652_, new_n2653_, new_n2654_, new_n2655_, new_n2656_, new_n2657_,
    new_n2658_, new_n2659_, new_n2660_, new_n2661_, new_n2662_, new_n2663_,
    new_n2664_, new_n2665_, new_n2666_, new_n2667_, new_n2668_, new_n2669_,
    new_n2670_, new_n2671_, new_n2672_, new_n2673_, new_n2674_, new_n2675_,
    new_n2676_, new_n2677_, new_n2678_, new_n2679_, new_n2680_, new_n2681_,
    new_n2682_, new_n2683_, new_n2684_, new_n2685_, new_n2686_, new_n2687_,
    new_n2688_, new_n2689_, new_n2690_, new_n2691_, new_n2692_, new_n2693_,
    new_n2694_, new_n2695_, new_n2696_, new_n2697_, new_n2698_, new_n2699_,
    new_n2700_, new_n2701_, new_n2702_, new_n2703_, new_n2704_, new_n2705_,
    new_n2706_, new_n2707_, new_n2708_, new_n2709_, new_n2710_, new_n2711_,
    new_n2712_, new_n2713_, new_n2714_, new_n2715_, new_n2716_, new_n2717_,
    new_n2718_, new_n2719_, new_n2720_, new_n2721_, new_n2722_, new_n2723_,
    new_n2724_, new_n2725_, new_n2726_, new_n2727_, new_n2728_, new_n2729_,
    new_n2730_, new_n2731_, new_n2732_, new_n2733_, new_n2734_, new_n2735_,
    new_n2736_, new_n2737_, new_n2738_, new_n2739_, new_n2740_, new_n2741_,
    new_n2742_, new_n2743_, new_n2744_, new_n2745_, new_n2746_, new_n2747_,
    new_n2748_, new_n2749_, new_n2750_, new_n2751_, new_n2752_, new_n2753_,
    new_n2754_, new_n2755_, new_n2756_, new_n2757_, new_n2758_, new_n2759_,
    new_n2760_, new_n2761_, new_n2762_, new_n2763_, new_n2764_, new_n2765_,
    new_n2766_, new_n2767_, new_n2768_, new_n2769_, new_n2770_, new_n2771_,
    new_n2772_, new_n2773_, new_n2774_, new_n2775_, new_n2776_, new_n2777_,
    new_n2778_, new_n2779_, new_n2780_, new_n2781_, new_n2782_, new_n2783_,
    new_n2784_, new_n2785_, new_n2786_, new_n2787_, new_n2788_, new_n2789_,
    new_n2790_, new_n2791_, new_n2792_, new_n2793_, new_n2794_, new_n2795_,
    new_n2796_, new_n2797_, new_n2798_, new_n2799_, new_n2800_, new_n2801_,
    new_n2802_, new_n2803_, new_n2804_, new_n2805_, new_n2806_, new_n2807_,
    new_n2808_, new_n2809_, new_n2810_, new_n2811_, new_n2812_, new_n2813_,
    new_n2814_, new_n2815_, new_n2816_, new_n2817_, new_n2818_, new_n2819_,
    new_n2820_, new_n2821_, new_n2822_, new_n2823_, new_n2824_, new_n2825_,
    new_n2826_, new_n2827_, new_n2828_, new_n2829_, new_n2830_, new_n2831_,
    new_n2832_, new_n2833_, new_n2834_, new_n2835_, new_n2836_, new_n2837_,
    new_n2838_, new_n2839_, new_n2840_, new_n2841_, new_n2842_, new_n2843_,
    new_n2844_, new_n2845_, new_n2846_, new_n2847_, new_n2848_, new_n2849_,
    new_n2850_, new_n2851_, new_n2852_, new_n2853_, new_n2854_, new_n2855_,
    new_n2856_, new_n2857_, new_n2858_, new_n2859_, new_n2860_, new_n2861_,
    new_n2862_, new_n2863_, new_n2864_, new_n2865_, new_n2866_, new_n2867_,
    new_n2868_, new_n2869_, new_n2870_, new_n2871_, new_n2872_, new_n2873_,
    new_n2874_, new_n2875_, new_n2876_, new_n2877_, new_n2878_, new_n2879_,
    new_n2880_, new_n2881_, new_n2882_, new_n2883_, new_n2884_, new_n2885_,
    new_n2886_, new_n2887_, new_n2888_, new_n2889_, new_n2890_, new_n2891_,
    new_n2892_, new_n2893_, new_n2894_, new_n2895_, new_n2896_, new_n2897_,
    new_n2898_, new_n2899_, new_n2900_, new_n2901_, new_n2902_, new_n2903_,
    new_n2904_, new_n2905_, new_n2906_, new_n2907_, new_n2908_, new_n2909_,
    new_n2910_, new_n2911_, new_n2912_, new_n2913_, new_n2914_, new_n2915_,
    new_n2916_, new_n2917_, new_n2918_, new_n2919_, new_n2920_, new_n2921_,
    new_n2922_, new_n2923_, new_n2924_, new_n2925_, new_n2926_, new_n2927_,
    new_n2928_, new_n2929_, new_n2930_, new_n2931_, new_n2932_, new_n2933_,
    new_n2934_, new_n2935_, new_n2936_, new_n2937_, new_n2938_, new_n2939_,
    new_n2940_, new_n2941_, new_n2942_, new_n2943_, new_n2944_, new_n2945_,
    new_n2946_, new_n2947_, new_n2948_, new_n2949_, new_n2950_, new_n2951_,
    new_n2952_, new_n2953_, new_n2954_, new_n2955_, new_n2956_, new_n2957_,
    new_n2958_, new_n2959_, new_n2960_, new_n2961_, new_n2962_, new_n2963_,
    new_n2964_, new_n2965_, new_n2966_, new_n2967_, new_n2968_, new_n2969_,
    new_n2970_, new_n2971_, new_n2972_, new_n2973_, new_n2974_, new_n2975_,
    new_n2976_, new_n2977_, new_n2978_, new_n2979_, new_n2980_, new_n2981_,
    new_n2982_, new_n2983_, new_n2984_, new_n2985_, new_n2986_, new_n2987_,
    new_n2988_, new_n2989_, new_n2990_, new_n2991_, new_n2992_, new_n2993_,
    new_n2994_, new_n2995_, new_n2996_, new_n2997_, new_n2998_, new_n2999_,
    new_n3000_, new_n3001_, new_n3002_, new_n3003_, new_n3004_, new_n3005_,
    new_n3006_, new_n3007_, new_n3008_, new_n3009_, new_n3010_, new_n3011_,
    new_n3012_, new_n3013_, new_n3014_, new_n3015_, new_n3016_, new_n3017_,
    new_n3018_, new_n3019_, new_n3020_, new_n3021_, new_n3022_, new_n3023_,
    new_n3024_, new_n3025_, new_n3026_, new_n3027_, new_n3028_, new_n3029_,
    new_n3030_, new_n3031_, new_n3032_, new_n3033_, new_n3034_, new_n3035_,
    new_n3036_, new_n3037_, new_n3038_, new_n3039_, new_n3040_, new_n3041_,
    new_n3042_, new_n3043_, new_n3044_, new_n3045_, new_n3046_, new_n3047_,
    new_n3048_, new_n3049_, new_n3050_, new_n3051_, new_n3052_, new_n3053_,
    new_n3054_, new_n3055_, new_n3056_, new_n3057_, new_n3058_, new_n3059_,
    new_n3060_, new_n3061_, new_n3062_, new_n3063_, new_n3064_, new_n3065_,
    new_n3066_, new_n3067_, new_n3068_, new_n3069_, new_n3070_, new_n3071_,
    new_n3072_, new_n3073_, new_n3074_, new_n3075_, new_n3076_, new_n3077_,
    new_n3078_, new_n3079_, new_n3080_, new_n3081_, new_n3082_, new_n3083_,
    new_n3084_, new_n3085_, new_n3086_, new_n3087_, new_n3088_, new_n3089_,
    new_n3090_, new_n3091_, new_n3092_, new_n3093_, new_n3094_, new_n3095_,
    new_n3096_, new_n3097_, new_n3098_, new_n3099_, new_n3100_, new_n3101_,
    new_n3102_, new_n3103_, new_n3104_, new_n3105_, new_n3106_, new_n3107_,
    new_n3108_, new_n3109_, new_n3110_, new_n3111_, new_n3112_, new_n3113_,
    new_n3114_, new_n3115_, new_n3116_, new_n3117_, new_n3118_, new_n3119_,
    new_n3120_, new_n3121_, new_n3122_, new_n3123_, new_n3124_, new_n3125_,
    new_n3126_, new_n3127_, new_n3128_, new_n3129_, new_n3130_, new_n3131_,
    new_n3132_, new_n3133_, new_n3134_, new_n3135_, new_n3136_, new_n3137_,
    new_n3138_, new_n3139_, new_n3140_, new_n3141_, new_n3142_, new_n3143_,
    new_n3144_, new_n3145_, new_n3146_, new_n3147_, new_n3148_, new_n3149_,
    new_n3150_, new_n3151_, new_n3152_, new_n3153_, new_n3154_, new_n3155_,
    new_n3156_, new_n3157_, new_n3158_, new_n3159_, new_n3160_, new_n3161_,
    new_n3162_, new_n3163_, new_n3164_, new_n3165_, new_n3166_, new_n3167_,
    new_n3168_, new_n3169_, new_n3170_, new_n3171_, new_n3172_, new_n3173_,
    new_n3174_, new_n3175_, new_n3176_, new_n3177_, new_n3178_, new_n3179_,
    new_n3180_, new_n3181_, new_n3182_, new_n3183_, new_n3184_, new_n3185_,
    new_n3186_, new_n3187_, new_n3188_, new_n3189_, new_n3190_, new_n3191_,
    new_n3192_, new_n3193_, new_n3194_, new_n3195_, new_n3196_, new_n3197_,
    new_n3198_, new_n3199_, new_n3200_, new_n3201_, new_n3202_, new_n3203_,
    new_n3204_, new_n3205_, new_n3206_, new_n3207_, new_n3208_, new_n3209_,
    new_n3210_, new_n3211_, new_n3212_, new_n3213_, new_n3214_, new_n3215_,
    new_n3216_, new_n3217_, new_n3218_, new_n3219_, new_n3220_, new_n3221_,
    new_n3222_, new_n3223_, new_n3224_, new_n3225_, new_n3226_, new_n3227_,
    new_n3228_, new_n3229_, new_n3230_, new_n3231_, new_n3232_, new_n3233_,
    new_n3234_, new_n3235_, new_n3236_, new_n3237_, new_n3238_, new_n3239_,
    new_n3240_, new_n3241_, new_n3242_, new_n3243_, new_n3244_, new_n3245_,
    new_n3246_, new_n3247_, new_n3248_, new_n3249_, new_n3250_, new_n3251_,
    new_n3252_, new_n3253_, new_n3254_, new_n3255_, new_n3256_, new_n3257_,
    new_n3258_, new_n3259_, new_n3260_, new_n3261_, new_n3262_, new_n3263_,
    new_n3264_, new_n3265_, new_n3266_, new_n3267_, new_n3268_, new_n3269_,
    new_n3270_, new_n3271_, new_n3272_, new_n3273_, new_n3274_, new_n3275_,
    new_n3276_, new_n3277_, new_n3278_, new_n3279_, new_n3280_, new_n3281_,
    new_n3282_, new_n3283_, new_n3284_, new_n3285_, new_n3286_, new_n3287_,
    new_n3288_, new_n3289_, new_n3290_, new_n3291_, new_n3292_, new_n3293_,
    new_n3294_, new_n3295_, new_n3296_, new_n3297_, new_n3298_, new_n3299_,
    new_n3300_, new_n3301_, new_n3302_, new_n3303_, new_n3304_, new_n3305_,
    new_n3306_, new_n3307_, new_n3308_, new_n3309_, new_n3310_, new_n3311_,
    new_n3312_, new_n3313_, new_n3314_, new_n3315_, new_n3316_, new_n3317_,
    new_n3318_, new_n3319_, new_n3320_, new_n3321_, new_n3322_, new_n3323_,
    new_n3324_, new_n3325_, new_n3326_, new_n3327_, new_n3328_, new_n3329_,
    new_n3330_, new_n3331_, new_n3332_, new_n3333_, new_n3334_, new_n3335_,
    new_n3336_, new_n3337_, new_n3338_, new_n3339_, new_n3340_, new_n3341_,
    new_n3342_, new_n3343_, new_n3344_, new_n3345_, new_n3346_, new_n3347_,
    new_n3348_, new_n3349_, new_n3350_, new_n3351_, new_n3352_, new_n3353_,
    new_n3354_, new_n3355_, new_n3356_, new_n3357_, new_n3358_, new_n3359_,
    new_n3360_, new_n3361_, new_n3362_, new_n3363_, new_n3364_, new_n3365_,
    new_n3366_, new_n3367_, new_n3368_, new_n3369_, new_n3370_, new_n3371_,
    new_n3372_, new_n3373_, new_n3374_, new_n3375_, new_n3376_, new_n3377_,
    new_n3378_, new_n3379_, new_n3380_, new_n3381_, new_n3382_, new_n3383_,
    new_n3384_, new_n3385_, new_n3386_, new_n3387_, new_n3388_, new_n3389_,
    new_n3390_, new_n3391_, new_n3392_, new_n3393_, new_n3394_, new_n3395_,
    new_n3396_, new_n3397_, new_n3398_, new_n3399_, new_n3400_, new_n3401_,
    new_n3402_, new_n3403_, new_n3404_, new_n3405_, new_n3406_, new_n3407_,
    new_n3408_, new_n3409_, new_n3410_, new_n3411_, new_n3412_, new_n3413_,
    new_n3414_, new_n3415_, new_n3416_, new_n3417_, new_n3418_, new_n3419_,
    new_n3420_, new_n3421_, new_n3422_, new_n3423_, new_n3424_, new_n3425_,
    new_n3426_, new_n3427_, new_n3428_, new_n3429_, new_n3430_, new_n3431_,
    new_n3432_, new_n3433_, new_n3434_, new_n3435_, new_n3436_, new_n3437_,
    new_n3438_, new_n3439_, new_n3440_, new_n3441_, new_n3442_, new_n3443_,
    new_n3444_, new_n3445_, new_n3446_, new_n3447_, new_n3448_, new_n3449_,
    new_n3450_, new_n3451_, new_n3452_, new_n3453_, new_n3454_, new_n3455_,
    new_n3456_, new_n3457_, new_n3458_, new_n3459_, new_n3460_, new_n3461_,
    new_n3462_, new_n3463_, new_n3464_, new_n3465_, new_n3466_, new_n3467_,
    new_n3468_, new_n3469_, new_n3470_, new_n3471_, new_n3472_, new_n3473_,
    new_n3474_, new_n3475_, new_n3476_, new_n3477_, new_n3478_, new_n3479_,
    new_n3480_, new_n3481_, new_n3482_, new_n3483_, new_n3484_, new_n3485_,
    new_n3486_, new_n3487_, new_n3488_, new_n3489_, new_n3490_, new_n3491_,
    new_n3492_, new_n3493_, new_n3494_, new_n3495_, new_n3496_, new_n3497_,
    new_n3498_, new_n3499_, new_n3500_, new_n3501_, new_n3502_, new_n3503_,
    new_n3504_, new_n3505_, new_n3506_, new_n3507_, new_n3508_, new_n3509_,
    new_n3510_, new_n3511_, new_n3512_, new_n3513_, new_n3514_, new_n3515_,
    new_n3516_, new_n3517_, new_n3518_, new_n3519_, new_n3520_, new_n3521_,
    new_n3522_, new_n3523_, new_n3524_, new_n3525_, new_n3526_, new_n3527_,
    new_n3528_, new_n3529_, new_n3530_, new_n3531_, new_n3532_, new_n3533_,
    new_n3534_, new_n3535_, new_n3536_, new_n3537_, new_n3538_, new_n3539_,
    new_n3540_, new_n3541_, new_n3542_, new_n3543_, new_n3544_, new_n3545_,
    new_n3546_, new_n3547_, new_n3548_, new_n3549_, new_n3550_, new_n3551_,
    new_n3552_, new_n3553_, new_n3554_, new_n3555_, new_n3556_, new_n3557_,
    new_n3558_, new_n3559_, new_n3560_, new_n3561_, new_n3562_, new_n3563_,
    new_n3564_, new_n3565_, new_n3566_, new_n3567_, new_n3568_, new_n3569_,
    new_n3570_, new_n3571_, new_n3572_, new_n3573_, new_n3574_, new_n3575_,
    new_n3576_, new_n3577_, new_n3578_, new_n3579_, new_n3580_, new_n3581_,
    new_n3582_, new_n3583_, new_n3584_, new_n3585_, new_n3586_, new_n3587_,
    new_n3588_, new_n3589_, new_n3590_, new_n3591_, new_n3592_, new_n3593_,
    new_n3594_, new_n3595_, new_n3596_, new_n3597_, new_n3598_, new_n3599_,
    new_n3600_, new_n3601_, new_n3602_, new_n3603_, new_n3604_, new_n3605_,
    new_n3606_, new_n3607_, new_n3608_, new_n3609_, new_n3610_, new_n3611_,
    new_n3612_, new_n3613_, new_n3614_, new_n3615_, new_n3616_, new_n3617_,
    new_n3618_, new_n3619_, new_n3620_, new_n3621_, new_n3622_, new_n3623_,
    new_n3624_, new_n3625_, new_n3626_, new_n3627_, new_n3628_, new_n3629_,
    new_n3630_, new_n3631_, new_n3632_, new_n3633_, new_n3634_, new_n3635_,
    new_n3636_, new_n3637_, new_n3638_, new_n3639_, new_n3640_, new_n3641_,
    new_n3642_, new_n3643_, new_n3644_, new_n3645_, new_n3646_, new_n3647_,
    new_n3648_, new_n3649_, new_n3650_, new_n3651_, new_n3652_, new_n3653_,
    new_n3654_, new_n3655_, new_n3656_, new_n3657_, new_n3658_, new_n3659_,
    new_n3660_, new_n3661_, new_n3662_, new_n3663_, new_n3664_, new_n3665_,
    new_n3666_, new_n3667_, new_n3668_, new_n3669_, new_n3670_, new_n3671_,
    new_n3672_, new_n3673_, new_n3674_, new_n3675_, new_n3676_, new_n3677_,
    new_n3678_, new_n3679_, new_n3680_, new_n3681_, new_n3682_, new_n3683_,
    new_n3684_, new_n3685_, new_n3686_, new_n3687_, new_n3688_, new_n3689_,
    new_n3690_, new_n3691_, new_n3692_, new_n3693_, new_n3694_, new_n3695_,
    new_n3696_, new_n3697_, new_n3698_, new_n3699_, new_n3700_, new_n3701_,
    new_n3702_, new_n3703_, new_n3704_, new_n3705_, new_n3706_, new_n3707_,
    new_n3708_, new_n3709_, new_n3710_, new_n3711_, new_n3712_, new_n3713_,
    new_n3714_, new_n3715_, new_n3716_, new_n3717_, new_n3718_, new_n3719_,
    new_n3720_, new_n3721_, new_n3722_, new_n3723_, new_n3724_, new_n3725_,
    new_n3726_, new_n3727_, new_n3728_, new_n3729_, new_n3730_, new_n3731_,
    new_n3732_, new_n3733_, new_n3734_, new_n3735_, new_n3736_, new_n3737_,
    new_n3738_, new_n3739_, new_n3740_, new_n3741_, new_n3742_, new_n3743_,
    new_n3744_, new_n3745_, new_n3746_, new_n3747_, new_n3748_, new_n3749_,
    new_n3750_, new_n3751_, new_n3752_, new_n3753_, new_n3754_, new_n3755_,
    new_n3756_, new_n3757_, new_n3758_, new_n3759_, new_n3760_, new_n3761_,
    new_n3762_, new_n3763_, new_n3764_, new_n3765_, new_n3766_, new_n3767_,
    new_n3768_, new_n3769_, new_n3770_, new_n3771_, new_n3772_, new_n3773_,
    new_n3774_, new_n3775_, new_n3776_, new_n3777_, new_n3778_, new_n3779_,
    new_n3780_, new_n3781_, new_n3782_, new_n3783_, new_n3784_, new_n3785_,
    new_n3786_, new_n3787_, new_n3788_, new_n3789_, new_n3790_, new_n3791_,
    new_n3792_, new_n3793_, new_n3794_, new_n3795_, new_n3796_, new_n3797_,
    new_n3798_, new_n3799_, new_n3800_, new_n3801_, new_n3802_, new_n3803_,
    new_n3804_, new_n3805_, new_n3806_, new_n3807_, new_n3808_, new_n3809_,
    new_n3810_, new_n3811_, new_n3812_, new_n3813_, new_n3814_, new_n3815_,
    new_n3816_, new_n3817_, new_n3818_, new_n3819_, new_n3820_, new_n3821_,
    new_n3822_, new_n3823_, new_n3824_, new_n3825_, new_n3826_, new_n3827_,
    new_n3828_, new_n3829_, new_n3830_, new_n3831_, new_n3832_, new_n3833_,
    new_n3834_, new_n3835_, new_n3836_, new_n3837_, new_n3838_, new_n3839_,
    new_n3840_, new_n3841_, new_n3842_, new_n3843_, new_n3844_, new_n3845_,
    new_n3846_, new_n3847_, new_n3848_, new_n3849_, new_n3850_, new_n3851_,
    new_n3852_, new_n3853_, new_n3854_, new_n3855_, new_n3856_, new_n3857_,
    new_n3858_, new_n3859_, new_n3860_, new_n3861_, new_n3862_, new_n3863_,
    new_n3864_, new_n3865_, new_n3866_, new_n3867_, new_n3868_, new_n3869_,
    new_n3870_, new_n3871_, new_n3872_, new_n3873_, new_n3874_, new_n3875_,
    new_n3876_, new_n3877_, new_n3878_, new_n3879_, new_n3880_, new_n3881_,
    new_n3882_, new_n3883_, new_n3884_, new_n3885_, new_n3886_, new_n3887_,
    new_n3888_, new_n3889_, new_n3890_, new_n3891_, new_n3892_, new_n3893_,
    new_n3894_, new_n3895_, new_n3896_, new_n3897_, new_n3898_, new_n3899_,
    new_n3900_, new_n3901_, new_n3902_, new_n3903_, new_n3904_, new_n3905_,
    new_n3906_, new_n3907_, new_n3908_, new_n3909_, new_n3910_, new_n3911_,
    new_n3912_, new_n3913_, new_n3914_, new_n3915_, new_n3916_, new_n3917_,
    new_n3918_, new_n3919_, new_n3920_, new_n3921_, new_n3922_, new_n3923_,
    new_n3924_, new_n3925_, new_n3926_, new_n3927_, new_n3928_, new_n3929_,
    new_n3930_, new_n3931_, new_n3932_, new_n3933_, new_n3934_, new_n3935_,
    new_n3936_, new_n3937_, new_n3938_, new_n3939_, new_n3940_, new_n3941_,
    new_n3942_, new_n3943_, new_n3944_, new_n3945_, new_n3946_, new_n3947_,
    new_n3948_, new_n3949_, new_n3950_, new_n3951_, new_n3952_, new_n3953_,
    new_n3954_, new_n3955_, new_n3956_, new_n3957_, new_n3958_, new_n3959_,
    new_n3960_, new_n3961_, new_n3962_, new_n3963_, new_n3964_, new_n3965_,
    new_n3966_, new_n3967_, new_n3968_, new_n3969_, new_n3970_, new_n3971_,
    new_n3972_, new_n3973_, new_n3974_, new_n3975_, new_n3976_, new_n3977_,
    new_n3978_, new_n3979_, new_n3980_, new_n3981_, new_n3982_, new_n3983_,
    new_n3984_, new_n3985_, new_n3986_, new_n3987_, new_n3988_, new_n3989_,
    new_n3990_, new_n3991_, new_n3992_, new_n3993_, new_n3994_, new_n3995_,
    new_n3996_, new_n3997_, new_n3998_, new_n3999_, new_n4000_, new_n4001_,
    new_n4002_, new_n4003_, new_n4004_, new_n4005_, new_n4006_, new_n4007_,
    new_n4008_, new_n4009_, new_n4010_, new_n4011_, new_n4012_, new_n4013_,
    new_n4014_, new_n4015_, new_n4016_, new_n4017_, new_n4018_, new_n4019_,
    new_n4020_, new_n4021_, new_n4022_, new_n4023_, new_n4024_, new_n4025_,
    new_n4026_, new_n4027_, new_n4028_, new_n4029_, new_n4030_, new_n4031_,
    new_n4032_, new_n4033_, new_n4034_, new_n4035_, new_n4036_, new_n4037_,
    new_n4038_, new_n4039_, new_n4040_, new_n4041_, new_n4042_, new_n4043_,
    new_n4044_, new_n4045_, new_n4046_, new_n4047_, new_n4048_, new_n4049_,
    new_n4050_, new_n4051_, new_n4052_, new_n4053_, new_n4054_, new_n4055_,
    new_n4056_, new_n4057_, new_n4058_, new_n4059_, new_n4060_, new_n4061_,
    new_n4062_, new_n4063_, new_n4064_, new_n4065_, new_n4066_, new_n4067_,
    new_n4068_, new_n4069_, new_n4070_, new_n4071_, new_n4072_, new_n4073_,
    new_n4074_, new_n4075_, new_n4076_, new_n4077_, new_n4078_, new_n4079_,
    new_n4080_, new_n4081_, new_n4082_, new_n4083_, new_n4084_, new_n4085_,
    new_n4086_, new_n4087_, new_n4088_, new_n4089_, new_n4090_, new_n4091_,
    new_n4092_, new_n4093_, new_n4094_, new_n4095_, new_n4096_, new_n4097_,
    new_n4098_, new_n4099_, new_n4100_, new_n4101_, new_n4102_, new_n4103_,
    new_n4104_, new_n4105_, new_n4106_, new_n4107_, new_n4108_, new_n4109_,
    new_n4110_, new_n4111_, new_n4112_, new_n4113_, new_n4114_, new_n4115_,
    new_n4116_, new_n4117_, new_n4118_, new_n4119_, new_n4120_, new_n4121_,
    new_n4122_, new_n4123_, new_n4124_, new_n4125_, new_n4126_, new_n4127_,
    new_n4128_, new_n4129_, new_n4130_, new_n4131_, new_n4132_, new_n4133_,
    new_n4134_, new_n4135_, new_n4136_, new_n4137_, new_n4138_, new_n4139_,
    new_n4140_, new_n4141_, new_n4142_, new_n4143_, new_n4144_, new_n4145_,
    new_n4146_, new_n4147_, new_n4148_, new_n4149_, new_n4150_, new_n4151_,
    new_n4152_, new_n4153_, new_n4154_, new_n4155_, new_n4156_, new_n4157_,
    new_n4158_, new_n4159_, new_n4160_, new_n4161_, new_n4162_, new_n4163_,
    new_n4164_, new_n4165_, new_n4166_, new_n4167_, new_n4168_, new_n4169_,
    new_n4170_, new_n4171_, new_n4172_, new_n4173_, new_n4174_, new_n4175_,
    new_n4176_, new_n4177_, new_n4178_, new_n4179_, new_n4180_, new_n4181_,
    new_n4182_, new_n4183_, new_n4184_, new_n4185_, new_n4186_, new_n4187_,
    new_n4188_, new_n4189_, new_n4190_, new_n4191_, new_n4192_, new_n4193_,
    new_n4194_, new_n4195_, new_n4196_, new_n4197_, new_n4198_, new_n4199_,
    new_n4200_, new_n4201_, new_n4202_, new_n4203_, new_n4204_, new_n4205_,
    new_n4206_, new_n4207_, new_n4208_, new_n4209_, new_n4210_, new_n4211_,
    new_n4212_, new_n4213_, new_n4214_, new_n4215_, new_n4216_, new_n4217_,
    new_n4218_, new_n4219_, new_n4220_, new_n4221_, new_n4222_, new_n4223_,
    new_n4224_, new_n4225_, new_n4226_, new_n4227_, new_n4228_, new_n4229_,
    new_n4230_, new_n4231_, new_n4232_, new_n4233_, new_n4234_, new_n4235_,
    new_n4236_, new_n4237_, new_n4238_, new_n4239_, new_n4240_, new_n4241_,
    new_n4242_, new_n4243_, new_n4244_, new_n4245_, new_n4246_, new_n4247_,
    new_n4248_, new_n4249_, new_n4250_, new_n4251_, new_n4252_, new_n4253_,
    new_n4254_, new_n4255_, new_n4256_, new_n4257_, new_n4258_, new_n4259_,
    new_n4260_, new_n4261_, new_n4262_, new_n4263_, new_n4264_, new_n4265_,
    new_n4266_, new_n4267_, new_n4268_, new_n4269_, new_n4270_, new_n4271_,
    new_n4272_, new_n4273_, new_n4274_, new_n4275_, new_n4276_, new_n4277_,
    new_n4278_, new_n4279_, new_n4280_, new_n4281_, new_n4282_, new_n4283_,
    new_n4284_, new_n4285_, new_n4286_, new_n4287_, new_n4288_, new_n4289_,
    new_n4290_, new_n4291_, new_n4292_, new_n4293_, new_n4294_, new_n4295_,
    new_n4296_, new_n4297_, new_n4298_, new_n4299_, new_n4300_, new_n4301_,
    new_n4302_, new_n4303_, new_n4304_, new_n4305_, new_n4306_, new_n4307_,
    new_n4308_, new_n4309_, new_n4310_, new_n4311_, new_n4312_, new_n4313_,
    new_n4314_, new_n4315_, new_n4316_, new_n4317_, new_n4318_, new_n4319_,
    new_n4320_, new_n4321_, new_n4322_, new_n4323_, new_n4324_, new_n4325_,
    new_n4326_, new_n4327_, new_n4328_, new_n4329_, new_n4330_, new_n4331_,
    new_n4332_, new_n4333_, new_n4334_, new_n4335_, new_n4336_, new_n4337_,
    new_n4338_, new_n4339_, new_n4340_, new_n4341_, new_n4342_, new_n4343_,
    new_n4344_, new_n4345_, new_n4346_, new_n4347_, new_n4348_, new_n4349_,
    new_n4350_, new_n4351_, new_n4352_, new_n4353_, new_n4354_, new_n4355_,
    new_n4356_, new_n4357_, new_n4358_, new_n4359_, new_n4360_, new_n4361_,
    new_n4362_, new_n4363_, new_n4364_, new_n4365_, new_n4366_, new_n4367_,
    new_n4368_, new_n4369_, new_n4370_, new_n4371_, new_n4372_, new_n4373_,
    new_n4374_, new_n4375_, new_n4376_, new_n4377_, new_n4378_, new_n4379_,
    new_n4380_, new_n4381_, new_n4382_, new_n4383_, new_n4384_, new_n4385_,
    new_n4386_, new_n4387_, new_n4388_, new_n4389_, new_n4390_, new_n4391_,
    new_n4392_, new_n4393_, new_n4394_, new_n4395_, new_n4396_, new_n4397_,
    new_n4398_, new_n4399_, new_n4400_, new_n4401_, new_n4402_, new_n4403_,
    new_n4404_, new_n4405_, new_n4406_, new_n4407_, new_n4408_, new_n4409_,
    new_n4410_, new_n4411_, new_n4412_, new_n4413_, new_n4414_, new_n4415_,
    new_n4416_, new_n4417_, new_n4418_, new_n4419_, new_n4420_, new_n4421_,
    new_n4422_, new_n4423_, new_n4424_, new_n4425_, new_n4426_, new_n4427_,
    new_n4428_, new_n4429_, new_n4430_, new_n4431_, new_n4432_, new_n4433_,
    new_n4434_, new_n4435_, new_n4436_, new_n4437_, new_n4438_, new_n4439_,
    new_n4440_, new_n4441_, new_n4442_, new_n4443_, new_n4444_, new_n4445_,
    new_n4446_, new_n4447_, new_n4448_, new_n4449_, new_n4450_, new_n4451_,
    new_n4452_, new_n4453_, new_n4454_, new_n4455_, new_n4456_, new_n4457_,
    new_n4458_, new_n4459_, new_n4460_, new_n4461_, new_n4462_, new_n4463_,
    new_n4464_, new_n4465_, new_n4466_, new_n4467_, new_n4468_, new_n4469_,
    new_n4470_, new_n4471_, new_n4472_, new_n4473_, new_n4474_, new_n4475_,
    new_n4476_, new_n4477_, new_n4478_, new_n4479_, new_n4480_, new_n4481_,
    new_n4482_, new_n4483_, new_n4484_, new_n4485_, new_n4486_, new_n4487_,
    new_n4488_, new_n4489_, new_n4490_, new_n4491_, new_n4492_, new_n4493_,
    new_n4494_, new_n4495_, new_n4496_, new_n4497_, new_n4498_, new_n4499_,
    new_n4500_, new_n4501_, new_n4502_, new_n4503_, new_n4504_, new_n4505_,
    new_n4506_, new_n4507_, new_n4508_, new_n4509_, new_n4510_, new_n4511_,
    new_n4512_, new_n4513_, new_n4514_, new_n4515_, new_n4516_, new_n4517_,
    new_n4518_, new_n4519_, new_n4520_, new_n4521_, new_n4522_, new_n4523_,
    new_n4524_, new_n4525_, new_n4526_, new_n4527_, new_n4528_, new_n4529_,
    new_n4530_, new_n4531_, new_n4532_, new_n4533_, new_n4534_, new_n4535_,
    new_n4536_, new_n4537_, new_n4538_, new_n4539_, new_n4540_, new_n4541_,
    new_n4542_, new_n4543_, new_n4544_, new_n4545_, new_n4546_, new_n4547_,
    new_n4548_, new_n4549_, new_n4550_, new_n4551_, new_n4552_, new_n4553_,
    new_n4554_, new_n4555_, new_n4556_, new_n4557_, new_n4558_, new_n4559_,
    new_n4560_, new_n4561_, new_n4562_, new_n4563_, new_n4564_, new_n4565_,
    new_n4566_, new_n4567_, new_n4568_, new_n4569_, new_n4570_, new_n4571_,
    new_n4572_, new_n4573_, new_n4574_, new_n4575_, new_n4576_, new_n4577_,
    new_n4578_, new_n4579_, new_n4580_, new_n4581_, new_n4582_, new_n4583_,
    new_n4584_, new_n4585_, new_n4586_, new_n4587_, new_n4588_, new_n4589_,
    new_n4590_, new_n4591_, new_n4592_, new_n4593_, new_n4594_, new_n4595_,
    new_n4596_, new_n4597_, new_n4598_, new_n4599_, new_n4600_, new_n4601_,
    new_n4602_, new_n4603_, new_n4604_, new_n4605_, new_n4606_, new_n4607_,
    new_n4608_, new_n4609_, new_n4610_, new_n4611_, new_n4612_, new_n4613_,
    new_n4614_, new_n4615_, new_n4616_, new_n4617_, new_n4618_, new_n4619_,
    new_n4620_, new_n4621_, new_n4622_, new_n4623_, new_n4624_, new_n4625_,
    new_n4626_, new_n4627_, new_n4628_, new_n4629_, new_n4630_, new_n4631_,
    new_n4632_, new_n4633_, new_n4634_, new_n4635_, new_n4636_, new_n4637_,
    new_n4638_, new_n4639_, new_n4640_, new_n4641_, new_n4642_, new_n4643_,
    new_n4644_, new_n4645_, new_n4646_, new_n4647_, new_n4648_, new_n4649_,
    new_n4650_, new_n4651_, new_n4652_, new_n4653_, new_n4654_, new_n4655_,
    new_n4656_, new_n4657_, new_n4658_, new_n4659_, new_n4660_, new_n4661_,
    new_n4662_, new_n4663_, new_n4664_, new_n4665_, new_n4666_, new_n4667_,
    new_n4668_, new_n4669_, new_n4670_, new_n4671_, new_n4672_, new_n4673_,
    new_n4674_, new_n4675_, new_n4676_, new_n4677_, new_n4678_, new_n4679_,
    new_n4680_, new_n4681_, new_n4682_, new_n4683_, new_n4684_, new_n4685_,
    new_n4686_, new_n4687_, new_n4688_, new_n4689_, new_n4690_, new_n4691_,
    new_n4692_, new_n4693_, new_n4694_, new_n4695_, new_n4696_, new_n4697_,
    new_n4698_, new_n4699_, new_n4700_, new_n4701_, new_n4702_, new_n4703_,
    new_n4704_, new_n4705_, new_n4706_, new_n4707_, new_n4708_, new_n4709_,
    new_n4710_, new_n4711_, new_n4712_, new_n4713_, new_n4714_, new_n4715_,
    new_n4716_, new_n4717_, new_n4718_, new_n4719_, new_n4720_, new_n4721_,
    new_n4722_, new_n4723_, new_n4724_, new_n4725_, new_n4726_, new_n4727_,
    new_n4728_, new_n4729_, new_n4730_, new_n4731_, new_n4732_, new_n4733_,
    new_n4734_, new_n4735_, new_n4736_, new_n4737_, new_n4738_, new_n4739_,
    new_n4740_, new_n4741_, new_n4742_, new_n4743_, new_n4744_, new_n4745_,
    new_n4746_, new_n4747_, new_n4748_, new_n4749_, new_n4750_, new_n4751_,
    new_n4752_, new_n4753_, new_n4754_, new_n4755_, new_n4756_, new_n4757_,
    new_n4758_, new_n4759_, new_n4760_, new_n4761_, new_n4762_, new_n4763_,
    new_n4764_, new_n4765_, new_n4766_, new_n4767_, new_n4768_, new_n4769_,
    new_n4770_, new_n4771_, new_n4772_, new_n4773_, new_n4774_, new_n4775_,
    new_n4776_, new_n4777_, new_n4778_, new_n4779_, new_n4780_, new_n4781_,
    new_n4782_, new_n4783_, new_n4784_, new_n4785_, new_n4786_, new_n4787_,
    new_n4788_, new_n4789_, new_n4790_, new_n4791_, new_n4792_, new_n4793_,
    new_n4794_, new_n4795_, new_n4796_, new_n4797_, new_n4798_, new_n4799_,
    new_n4800_, new_n4801_, new_n4802_, new_n4803_, new_n4804_, new_n4805_,
    new_n4806_, new_n4807_, new_n4808_, new_n4809_, new_n4810_, new_n4811_,
    new_n4812_, new_n4813_, new_n4814_, new_n4815_, new_n4816_, new_n4817_,
    new_n4818_, new_n4819_, new_n4820_, new_n4821_, new_n4822_, new_n4823_,
    new_n4824_, new_n4825_, new_n4826_, new_n4827_, new_n4828_, new_n4829_,
    new_n4830_, new_n4831_, new_n4832_, new_n4833_, new_n4834_, new_n4835_,
    new_n4836_, new_n4837_, new_n4838_, new_n4839_, new_n4840_, new_n4841_,
    new_n4842_, new_n4843_, new_n4844_, new_n4845_, new_n4846_, new_n4847_,
    new_n4848_, new_n4849_, new_n4850_, new_n4851_, new_n4852_, new_n4853_,
    new_n4854_, new_n4855_, new_n4856_, new_n4857_, new_n4858_, new_n4859_,
    new_n4860_, new_n4861_, new_n4862_, new_n4863_, new_n4864_, new_n4865_,
    new_n4866_, new_n4867_, new_n4868_, new_n4869_, new_n4870_, new_n4871_,
    new_n4872_, new_n4873_, new_n4874_, new_n4875_, new_n4876_, new_n4877_,
    new_n4878_, new_n4879_, new_n4880_, new_n4881_, new_n4882_, new_n4883_,
    new_n4884_, new_n4885_, new_n4886_, new_n4887_, new_n4888_, new_n4889_,
    new_n4890_, new_n4891_, new_n4892_, new_n4893_, new_n4894_, new_n4895_,
    new_n4896_, new_n4897_, new_n4898_, new_n4899_, new_n4900_, new_n4901_,
    new_n4902_, new_n4903_, new_n4904_, new_n4905_, new_n4906_, new_n4907_,
    new_n4908_, new_n4909_, new_n4910_, new_n4911_, new_n4912_, new_n4913_,
    new_n4914_, new_n4915_, new_n4916_, new_n4917_, new_n4918_, new_n4919_,
    new_n4920_, new_n4921_, new_n4922_, new_n4923_, new_n4924_, new_n4925_,
    new_n4926_, new_n4927_, new_n4928_, new_n4929_, new_n4930_, new_n4931_,
    new_n4932_, new_n4933_, new_n4934_, new_n4935_, new_n4936_, new_n4937_,
    new_n4938_, new_n4939_, new_n4940_, new_n4941_, new_n4942_, new_n4943_,
    new_n4944_, new_n4945_, new_n4946_, new_n4947_, new_n4948_, new_n4949_,
    new_n4950_, new_n4951_, new_n4952_, new_n4953_, new_n4954_, new_n4955_,
    new_n4956_, new_n4957_, new_n4958_, new_n4959_, new_n4960_, new_n4961_,
    new_n4962_, new_n4963_, new_n4964_, new_n4965_, new_n4966_, new_n4967_,
    new_n4968_, new_n4969_, new_n4970_, new_n4971_, new_n4972_, new_n4973_,
    new_n4974_, new_n4975_, new_n4976_, new_n4977_, new_n4978_, new_n4979_,
    new_n4980_, new_n4981_, new_n4982_, new_n4983_, new_n4984_, new_n4985_,
    new_n4986_, new_n4987_, new_n4988_, new_n4989_, new_n4990_, new_n4991_,
    new_n4992_, new_n4993_, new_n4994_, new_n4995_, new_n4996_, new_n4997_,
    new_n4998_, new_n4999_, new_n5000_, new_n5001_, new_n5002_, new_n5003_,
    new_n5004_, new_n5005_, new_n5006_, new_n5007_, new_n5008_, new_n5009_,
    new_n5010_, new_n5011_, new_n5012_, new_n5013_, new_n5014_, new_n5015_,
    new_n5016_, new_n5017_, new_n5018_, new_n5019_, new_n5020_, new_n5021_,
    new_n5022_, new_n5023_, new_n5024_, new_n5025_, new_n5026_, new_n5027_,
    new_n5028_, new_n5029_, new_n5030_, new_n5031_, new_n5032_, new_n5033_,
    new_n5034_, new_n5035_, new_n5036_, new_n5037_, new_n5038_, new_n5039_,
    new_n5040_, new_n5041_, new_n5042_, new_n5043_, new_n5044_, new_n5045_,
    new_n5046_, new_n5047_, new_n5048_, new_n5049_, new_n5050_, new_n5051_,
    new_n5052_, new_n5053_, new_n5054_, new_n5055_, new_n5056_, new_n5057_,
    new_n5058_, new_n5059_, new_n5060_, new_n5061_, new_n5062_, new_n5063_,
    new_n5064_, new_n5065_, new_n5066_, new_n5067_, new_n5068_, new_n5069_,
    new_n5070_, new_n5071_, new_n5072_, new_n5073_, new_n5074_, new_n5075_,
    new_n5076_, new_n5077_, new_n5078_, new_n5079_, new_n5080_, new_n5081_,
    new_n5082_, new_n5083_, new_n5084_, new_n5085_, new_n5086_, new_n5087_,
    new_n5088_, new_n5089_, new_n5090_, new_n5091_, new_n5092_, new_n5093_,
    new_n5094_, new_n5095_, new_n5096_, new_n5097_, new_n5098_, new_n5099_,
    new_n5100_, new_n5101_, new_n5102_, new_n5103_, new_n5104_, new_n5105_,
    new_n5106_, new_n5107_, new_n5108_, new_n5109_, new_n5110_, new_n5111_,
    new_n5112_, new_n5113_, new_n5114_, new_n5115_, new_n5116_, new_n5117_,
    new_n5118_, new_n5119_, new_n5120_, new_n5121_, new_n5122_, new_n5123_,
    new_n5124_, new_n5125_, new_n5126_, new_n5127_, new_n5128_, new_n5129_,
    new_n5130_, new_n5131_, new_n5132_, new_n5133_, new_n5134_, new_n5135_,
    new_n5136_, new_n5137_, new_n5138_, new_n5139_, new_n5140_, new_n5141_,
    new_n5142_, new_n5143_, new_n5144_, new_n5145_, new_n5146_, new_n5147_,
    new_n5148_, new_n5149_, new_n5150_, new_n5151_, new_n5152_, new_n5153_,
    new_n5154_, new_n5155_, new_n5156_, new_n5157_, new_n5158_, new_n5159_,
    new_n5160_, new_n5161_, new_n5162_, new_n5163_, new_n5164_, new_n5165_,
    new_n5166_, new_n5167_, new_n5168_, new_n5169_, new_n5170_, new_n5171_,
    new_n5172_, new_n5173_, new_n5174_, new_n5175_, new_n5176_, new_n5177_,
    new_n5178_, new_n5179_, new_n5180_, new_n5181_, new_n5182_, new_n5183_,
    new_n5184_, new_n5185_, new_n5186_, new_n5187_, new_n5188_, new_n5189_,
    new_n5190_, new_n5191_, new_n5192_, new_n5193_, new_n5194_, new_n5195_,
    new_n5196_, new_n5197_, new_n5198_, new_n5199_, new_n5200_, new_n5201_,
    new_n5202_, new_n5203_, new_n5204_, new_n5205_, new_n5206_, new_n5207_,
    new_n5208_, new_n5209_, new_n5210_, new_n5211_, new_n5212_, new_n5213_,
    new_n5214_, new_n5215_, new_n5216_, new_n5217_, new_n5218_, new_n5219_,
    new_n5220_, new_n5221_, new_n5222_, new_n5223_, new_n5224_, new_n5225_,
    new_n5226_, new_n5227_, new_n5228_, new_n5229_, new_n5230_, new_n5231_,
    new_n5232_, new_n5233_, new_n5234_, new_n5235_, new_n5236_, new_n5237_,
    new_n5238_, new_n5239_, new_n5240_, new_n5241_, new_n5242_, new_n5243_,
    new_n5244_, new_n5245_, new_n5246_, new_n5247_, new_n5248_, new_n5249_,
    new_n5250_, new_n5251_, new_n5252_, new_n5253_, new_n5254_, new_n5255_,
    new_n5256_, new_n5257_, new_n5258_, new_n5259_, new_n5260_, new_n5261_,
    new_n5262_, new_n5263_, new_n5264_, new_n5265_, new_n5266_, new_n5267_,
    new_n5268_, new_n5269_, new_n5270_, new_n5271_, new_n5272_, new_n5273_,
    new_n5274_, new_n5275_, new_n5276_, new_n5277_, new_n5278_, new_n5279_,
    new_n5280_, new_n5281_, new_n5282_, new_n5283_, new_n5284_, new_n5285_,
    new_n5286_, new_n5287_, new_n5288_, new_n5289_, new_n5290_, new_n5291_,
    new_n5292_, new_n5293_, new_n5294_, new_n5295_, new_n5296_, new_n5297_,
    new_n5298_, new_n5299_, new_n5300_, new_n5301_, new_n5302_, new_n5303_,
    new_n5304_, new_n5305_, new_n5306_, new_n5307_, new_n5308_, new_n5309_,
    new_n5310_, new_n5311_, new_n5312_, new_n5313_, new_n5314_, new_n5315_,
    new_n5316_, new_n5317_, new_n5318_, new_n5319_, new_n5320_, new_n5321_,
    new_n5322_, new_n5323_, new_n5324_, new_n5325_, new_n5326_, new_n5327_,
    new_n5328_, new_n5329_, new_n5330_, new_n5331_, new_n5332_, new_n5333_,
    new_n5334_, new_n5335_, new_n5336_, new_n5337_, new_n5338_, new_n5339_,
    new_n5340_, new_n5341_, new_n5342_, new_n5343_, new_n5344_, new_n5345_,
    new_n5346_, new_n5347_, new_n5348_, new_n5349_, new_n5350_, new_n5351_,
    new_n5352_, new_n5353_, new_n5354_, new_n5355_, new_n5356_, new_n5357_,
    new_n5358_, new_n5359_, new_n5360_, new_n5361_, new_n5362_, new_n5363_,
    new_n5364_, new_n5365_, new_n5366_, new_n5367_, new_n5368_, new_n5369_,
    new_n5370_, new_n5371_, new_n5372_, new_n5373_, new_n5374_, new_n5375_,
    new_n5376_, new_n5377_, new_n5378_, new_n5379_, new_n5380_, new_n5381_,
    new_n5382_, new_n5383_, new_n5384_, new_n5385_, new_n5386_, new_n5387_,
    new_n5388_, new_n5389_, new_n5390_, new_n5391_, new_n5392_, new_n5393_,
    new_n5394_, new_n5395_, new_n5396_, new_n5397_, new_n5398_, new_n5399_,
    new_n5400_, new_n5401_, new_n5402_, new_n5403_, new_n5404_, new_n5405_,
    new_n5406_, new_n5407_, new_n5408_, new_n5409_, new_n5410_, new_n5411_,
    new_n5412_, new_n5413_, new_n5414_, new_n5415_, new_n5416_, new_n5417_,
    new_n5418_, new_n5419_, new_n5420_, new_n5421_, new_n5422_, new_n5423_,
    new_n5424_, new_n5425_, new_n5426_, new_n5427_, new_n5428_, new_n5429_,
    new_n5430_, new_n5431_, new_n5432_, new_n5433_, new_n5434_, new_n5435_,
    new_n5436_, new_n5437_, new_n5438_, new_n5439_, new_n5440_, new_n5441_,
    new_n5442_, new_n5443_, new_n5444_, new_n5445_, new_n5446_, new_n5447_,
    new_n5448_, new_n5449_, new_n5450_, new_n5451_, new_n5452_, new_n5453_,
    new_n5454_, new_n5455_, new_n5456_, new_n5457_, new_n5458_, new_n5459_,
    new_n5460_, new_n5461_, new_n5462_, new_n5463_, new_n5464_, new_n5465_,
    new_n5466_, new_n5467_, new_n5468_, new_n5469_, new_n5470_, new_n5471_,
    new_n5472_, new_n5473_, new_n5474_, new_n5475_, new_n5476_, new_n5477_,
    new_n5478_, new_n5479_, new_n5480_, new_n5481_, new_n5482_, new_n5483_,
    new_n5484_, new_n5485_, new_n5486_, new_n5487_, new_n5488_, new_n5489_,
    new_n5490_, new_n5491_, new_n5492_, new_n5493_, new_n5494_, new_n5495_,
    new_n5496_, new_n5497_, new_n5498_, new_n5499_, new_n5500_, new_n5501_,
    new_n5502_, new_n5503_, new_n5504_, new_n5505_, new_n5506_, new_n5507_,
    new_n5508_, new_n5509_, new_n5510_, new_n5511_, new_n5512_, new_n5513_,
    new_n5514_, new_n5515_, new_n5516_, new_n5517_, new_n5518_, new_n5519_,
    new_n5520_, new_n5521_, new_n5522_, new_n5523_, new_n5524_, new_n5525_,
    new_n5526_, new_n5527_, new_n5528_, new_n5529_, new_n5530_, new_n5531_,
    new_n5532_, new_n5533_, new_n5534_, new_n5535_, new_n5536_, new_n5537_,
    new_n5538_, new_n5539_, new_n5540_, new_n5541_, new_n5542_, new_n5543_,
    new_n5544_, new_n5545_, new_n5546_, new_n5547_, new_n5548_, new_n5549_,
    new_n5550_, new_n5551_, new_n5552_, new_n5553_, new_n5554_, new_n5555_,
    new_n5556_, new_n5557_, new_n5558_, new_n5559_, new_n5560_, new_n5561_,
    new_n5562_, new_n5563_, new_n5564_, new_n5565_, new_n5566_, new_n5567_,
    new_n5568_, new_n5569_, new_n5570_, new_n5571_, new_n5572_, new_n5573_,
    new_n5574_, new_n5575_, new_n5576_, new_n5577_, new_n5578_, new_n5579_,
    new_n5580_, new_n5581_, new_n5582_, new_n5583_, new_n5584_, new_n5585_,
    new_n5586_, new_n5587_, new_n5588_, new_n5589_, new_n5590_, new_n5591_,
    new_n5592_, new_n5593_, new_n5594_, new_n5595_, new_n5596_, new_n5597_,
    new_n5598_, new_n5599_, new_n5600_, new_n5601_, new_n5602_, new_n5603_,
    new_n5604_, new_n5605_, new_n5606_, new_n5607_, new_n5608_, new_n5609_,
    new_n5610_, new_n5611_, new_n5612_, new_n5613_, new_n5614_, new_n5615_,
    new_n5616_, new_n5617_, new_n5618_, new_n5619_, new_n5620_, new_n5621_,
    new_n5622_, new_n5623_, new_n5624_, new_n5625_, new_n5626_, new_n5627_,
    new_n5628_, new_n5629_, new_n5630_, new_n5631_, new_n5632_, new_n5633_,
    new_n5634_, new_n5635_, new_n5636_, new_n5637_, new_n5638_, new_n5639_,
    new_n5640_, new_n5641_, new_n5642_, new_n5643_, new_n5644_, new_n5645_,
    new_n5646_, new_n5647_, new_n5648_, new_n5649_, new_n5650_, new_n5651_,
    new_n5652_, new_n5653_, new_n5654_, new_n5655_, new_n5656_, new_n5657_,
    new_n5658_, new_n5659_, new_n5660_, new_n5661_, new_n5662_, new_n5663_,
    new_n5664_, new_n5665_, new_n5666_, new_n5667_, new_n5668_, new_n5669_,
    new_n5670_, new_n5671_, new_n5672_, new_n5673_, new_n5674_, new_n5675_,
    new_n5676_, new_n5677_, new_n5678_, new_n5679_, new_n5680_, new_n5681_,
    new_n5682_, new_n5683_, new_n5684_, new_n5685_, new_n5686_, new_n5687_,
    new_n5688_, new_n5689_, new_n5690_, new_n5691_, new_n5692_, new_n5693_,
    new_n5694_, new_n5695_, new_n5696_, new_n5697_, new_n5698_, new_n5699_,
    new_n5700_, new_n5701_, new_n5702_, new_n5703_, new_n5704_, new_n5705_,
    new_n5706_, new_n5707_, new_n5708_, new_n5709_, new_n5710_, new_n5711_,
    new_n5712_, new_n5713_, new_n5714_, new_n5715_, new_n5716_, new_n5717_,
    new_n5718_, new_n5719_, new_n5720_, new_n5721_, new_n5722_, new_n5723_,
    new_n5724_, new_n5725_, new_n5726_, new_n5727_, new_n5728_, new_n5729_,
    new_n5730_, new_n5731_, new_n5732_, new_n5733_, new_n5734_, new_n5735_,
    new_n5736_, new_n5737_, new_n5738_, new_n5739_, new_n5740_, new_n5741_,
    new_n5742_, new_n5743_, new_n5744_, new_n5745_, new_n5746_, new_n5747_,
    new_n5748_, new_n5749_, new_n5750_, new_n5751_, new_n5752_, new_n5753_,
    new_n5754_, new_n5755_, new_n5756_, new_n5757_, new_n5758_, new_n5759_,
    new_n5760_, new_n5761_, new_n5762_, new_n5763_, new_n5764_, new_n5765_,
    new_n5766_, new_n5767_, new_n5768_, new_n5769_, new_n5770_, new_n5771_,
    new_n5772_, new_n5773_, new_n5774_, new_n5775_, new_n5776_, new_n5777_,
    new_n5778_, new_n5779_, new_n5780_, new_n5781_, new_n5782_, new_n5783_,
    new_n5784_, new_n5785_, new_n5786_, new_n5787_, new_n5788_, new_n5789_,
    new_n5790_, new_n5791_, new_n5792_, new_n5793_, new_n5794_, new_n5795_,
    new_n5796_, new_n5797_, new_n5798_, new_n5799_, new_n5800_, new_n5801_,
    new_n5802_, new_n5803_, new_n5804_, new_n5805_, new_n5806_, new_n5807_,
    new_n5808_, new_n5809_, new_n5810_, new_n5811_, new_n5812_, new_n5813_,
    new_n5814_, new_n5815_, new_n5816_, new_n5817_, new_n5818_, new_n5819_,
    new_n5820_, new_n5821_, new_n5822_, new_n5823_, new_n5824_, new_n5825_,
    new_n5826_, new_n5827_, new_n5828_, new_n5829_, new_n5830_, new_n5831_,
    new_n5832_, new_n5833_, new_n5834_, new_n5835_, new_n5836_, new_n5837_,
    new_n5838_, new_n5839_, new_n5840_, new_n5841_, new_n5842_, new_n5843_,
    new_n5844_, new_n5845_, new_n5846_, new_n5847_, new_n5848_, new_n5849_,
    new_n5850_, new_n5851_, new_n5852_, new_n5853_, new_n5854_, new_n5855_,
    new_n5856_, new_n5857_, new_n5858_, new_n5859_, new_n5860_, new_n5861_,
    new_n5862_, new_n5863_, new_n5864_, new_n5865_, new_n5866_, new_n5867_,
    new_n5868_, new_n5869_, new_n5870_, new_n5871_, new_n5872_, new_n5873_,
    new_n5874_, new_n5875_, new_n5876_, new_n5877_, new_n5878_, new_n5879_,
    new_n5880_, new_n5881_, new_n5882_, new_n5883_, new_n5884_, new_n5885_,
    new_n5886_, new_n5887_, new_n5888_, new_n5889_, new_n5890_, new_n5891_,
    new_n5892_, new_n5893_, new_n5894_, new_n5895_, new_n5896_, new_n5897_,
    new_n5898_, new_n5899_, new_n5900_, new_n5901_, new_n5902_, new_n5903_,
    new_n5904_, new_n5905_, new_n5906_, new_n5907_, new_n5908_, new_n5909_,
    new_n5910_, new_n5911_, new_n5912_, new_n5913_, new_n5914_, new_n5915_,
    new_n5916_, new_n5917_, new_n5918_, new_n5919_, new_n5920_, new_n5921_,
    new_n5922_, new_n5923_, new_n5924_, new_n5925_, new_n5926_, new_n5927_,
    new_n5928_, new_n5929_, new_n5930_, new_n5931_, new_n5932_, new_n5933_,
    new_n5934_, new_n5935_, new_n5936_, new_n5937_, new_n5938_, new_n5939_,
    new_n5940_, new_n5941_, new_n5942_, new_n5943_, new_n5944_, new_n5945_,
    new_n5946_, new_n5947_, new_n5948_, new_n5949_, new_n5950_, new_n5951_,
    new_n5952_, new_n5953_, new_n5954_, new_n5955_, new_n5956_, new_n5957_,
    new_n5958_, new_n5959_, new_n5960_, new_n5961_, new_n5962_, new_n5963_,
    new_n5964_, new_n5965_, new_n5966_, new_n5967_, new_n5968_, new_n5969_,
    new_n5970_, new_n5971_, new_n5972_, new_n5973_, new_n5974_, new_n5975_,
    new_n5976_, new_n5977_, new_n5978_, new_n5979_, new_n5980_, new_n5981_,
    new_n5982_, new_n5983_, new_n5984_, new_n5985_, new_n5986_, new_n5987_,
    new_n5988_, new_n5989_, new_n5990_, new_n5991_, new_n5992_, new_n5993_,
    new_n5994_, new_n5995_, new_n5996_, new_n5997_, new_n5998_, new_n5999_,
    new_n6000_, new_n6001_, new_n6002_, new_n6003_, new_n6004_, new_n6005_,
    new_n6006_, new_n6007_, new_n6008_, new_n6009_, new_n6010_, new_n6011_,
    new_n6012_, new_n6013_, new_n6014_, new_n6015_, new_n6016_, new_n6017_,
    new_n6018_, new_n6019_, new_n6020_, new_n6021_, new_n6022_, new_n6023_,
    new_n6024_, new_n6025_, new_n6026_, new_n6027_, new_n6028_, new_n6029_,
    new_n6030_, new_n6031_, new_n6032_, new_n6033_, new_n6034_, new_n6035_,
    new_n6036_, new_n6037_, new_n6038_, new_n6039_, new_n6040_, new_n6041_,
    new_n6042_, new_n6043_, new_n6044_, new_n6045_, new_n6046_, new_n6047_,
    new_n6048_, new_n6049_, new_n6050_, new_n6051_, new_n6052_, new_n6053_,
    new_n6054_, new_n6055_, new_n6056_, new_n6057_, new_n6058_, new_n6059_,
    new_n6060_, new_n6061_, new_n6062_, new_n6063_, new_n6064_, new_n6065_,
    new_n6066_, new_n6067_, new_n6068_, new_n6069_, new_n6070_, new_n6071_,
    new_n6072_, new_n6073_, new_n6074_, new_n6075_, new_n6076_, new_n6077_,
    new_n6078_, new_n6079_, new_n6080_, new_n6081_, new_n6082_, new_n6083_,
    new_n6084_, new_n6085_, new_n6086_, new_n6087_, new_n6088_, new_n6089_,
    new_n6090_, new_n6091_, new_n6092_, new_n6093_, new_n6094_, new_n6095_,
    new_n6096_, new_n6097_, new_n6098_, new_n6099_, new_n6100_, new_n6101_,
    new_n6102_, new_n6103_, new_n6104_, new_n6105_, new_n6106_, new_n6107_,
    new_n6108_, new_n6109_, new_n6110_, new_n6111_, new_n6112_, new_n6113_,
    new_n6114_, new_n6115_, new_n6116_, new_n6117_, new_n6118_, new_n6119_,
    new_n6120_, new_n6121_, new_n6122_, new_n6123_, new_n6124_, new_n6125_,
    new_n6126_, new_n6127_, new_n6128_, new_n6129_, new_n6130_, new_n6131_,
    new_n6132_, new_n6133_, new_n6134_, new_n6135_, new_n6136_, new_n6137_,
    new_n6138_, new_n6139_, new_n6140_, new_n6141_, new_n6142_, new_n6143_,
    new_n6144_, new_n6145_, new_n6146_, new_n6147_, new_n6148_, new_n6149_,
    new_n6150_, new_n6151_, new_n6152_, new_n6153_, new_n6154_, new_n6155_,
    new_n6156_, new_n6157_, new_n6158_, new_n6159_, new_n6160_, new_n6161_,
    new_n6162_, new_n6163_, new_n6164_, new_n6165_, new_n6166_, new_n6167_,
    new_n6168_, new_n6169_, new_n6170_, new_n6171_, new_n6172_, new_n6173_,
    new_n6174_, new_n6175_, new_n6176_, new_n6177_, new_n6178_, new_n6179_,
    new_n6180_, new_n6181_, new_n6182_, new_n6183_, new_n6184_, new_n6185_,
    new_n6186_, new_n6187_, new_n6188_, new_n6189_, new_n6190_, new_n6191_,
    new_n6192_, new_n6193_, new_n6194_, new_n6195_, new_n6196_, new_n6197_,
    new_n6198_, new_n6199_, new_n6200_, new_n6201_, new_n6202_, new_n6203_,
    new_n6204_, new_n6205_, new_n6206_, new_n6207_, new_n6208_, new_n6209_,
    new_n6210_, new_n6211_, new_n6212_, new_n6213_, new_n6214_, new_n6215_,
    new_n6216_, new_n6217_, new_n6218_, new_n6219_, new_n6220_, new_n6221_,
    new_n6222_, new_n6223_, new_n6224_, new_n6225_, new_n6226_, new_n6227_,
    new_n6228_, new_n6229_, new_n6230_, new_n6231_, new_n6232_, new_n6233_,
    new_n6234_, new_n6235_, new_n6236_, new_n6237_, new_n6238_, new_n6239_,
    new_n6240_, new_n6241_, new_n6242_, new_n6243_, new_n6244_, new_n6245_,
    new_n6246_, new_n6247_, new_n6248_, new_n6249_, new_n6250_, new_n6251_,
    new_n6252_, new_n6253_, new_n6254_, new_n6255_, new_n6256_, new_n6257_,
    new_n6258_, new_n6259_, new_n6260_, new_n6261_, new_n6262_, new_n6263_,
    new_n6264_, new_n6265_, new_n6266_, new_n6267_, new_n6268_, new_n6269_,
    new_n6270_, new_n6271_, new_n6272_, new_n6273_, new_n6274_, new_n6275_,
    new_n6276_, new_n6277_, new_n6278_, new_n6279_, new_n6280_, new_n6281_,
    new_n6282_, new_n6283_, new_n6284_, new_n6285_, new_n6286_, new_n6287_,
    new_n6288_, new_n6289_, new_n6290_, new_n6291_, new_n6292_, new_n6293_,
    new_n6294_, new_n6295_, new_n6296_, new_n6297_, new_n6298_, new_n6299_,
    new_n6300_, new_n6301_, new_n6302_, new_n6303_, new_n6304_, new_n6305_,
    new_n6306_, new_n6307_, new_n6308_, new_n6309_, new_n6310_, new_n6311_,
    new_n6312_, new_n6313_, new_n6314_, new_n6315_, new_n6316_, new_n6317_,
    new_n6318_, new_n6319_, new_n6320_, new_n6321_, new_n6322_, new_n6323_,
    new_n6324_, new_n6325_, new_n6326_, new_n6327_, new_n6328_, new_n6329_,
    new_n6330_, new_n6331_, new_n6332_, new_n6333_, new_n6334_, new_n6335_,
    new_n6336_, new_n6337_, new_n6338_, new_n6339_, new_n6340_, new_n6341_,
    new_n6342_, new_n6343_, new_n6344_, new_n6345_, new_n6346_, new_n6347_,
    new_n6348_, new_n6349_, new_n6350_, new_n6351_, new_n6352_, new_n6353_,
    new_n6354_, new_n6355_, new_n6356_, new_n6357_, new_n6358_, new_n6359_,
    new_n6360_, new_n6361_, new_n6362_, new_n6363_, new_n6364_, new_n6365_,
    new_n6366_, new_n6367_, new_n6368_, new_n6369_, new_n6370_, new_n6371_,
    new_n6372_, new_n6373_, new_n6374_, new_n6375_, new_n6376_, new_n6377_,
    new_n6378_, new_n6379_, new_n6380_, new_n6381_, new_n6382_, new_n6383_,
    new_n6384_, new_n6385_, new_n6386_, new_n6387_, new_n6388_, new_n6389_,
    new_n6390_, new_n6391_, new_n6392_, new_n6393_, new_n6394_, new_n6395_,
    new_n6396_, new_n6397_, new_n6398_, new_n6399_, new_n6400_, new_n6401_,
    new_n6402_, new_n6403_, new_n6404_, new_n6405_, new_n6406_, new_n6407_,
    new_n6408_, new_n6409_, new_n6410_, new_n6411_, new_n6412_, new_n6413_,
    new_n6414_, new_n6415_, new_n6416_, new_n6417_, new_n6418_, new_n6419_,
    new_n6420_, new_n6421_, new_n6422_, new_n6423_, new_n6424_, new_n6425_,
    new_n6426_, new_n6427_, new_n6428_, new_n6429_, new_n6430_, new_n6431_,
    new_n6432_, new_n6433_, new_n6434_, new_n6435_, new_n6436_, new_n6437_,
    new_n6438_, new_n6439_, new_n6440_, new_n6441_, new_n6442_, new_n6443_,
    new_n6444_, new_n6445_, new_n6446_, new_n6447_, new_n6448_, new_n6449_,
    new_n6450_, new_n6451_, new_n6452_, new_n6453_, new_n6454_, new_n6455_,
    new_n6456_, new_n6457_, new_n6458_, new_n6459_, new_n6460_, new_n6461_,
    new_n6462_, new_n6463_, new_n6464_, new_n6465_, new_n6466_, new_n6467_,
    new_n6468_, new_n6469_, new_n6470_, new_n6471_, new_n6472_, new_n6473_,
    new_n6474_, new_n6475_, new_n6476_, new_n6477_, new_n6478_, new_n6479_,
    new_n6480_, new_n6481_, new_n6482_, new_n6483_, new_n6484_, new_n6485_,
    new_n6486_, new_n6487_, new_n6488_, new_n6489_, new_n6490_, new_n6491_,
    new_n6492_, new_n6493_, new_n6494_, new_n6495_, new_n6496_, new_n6497_,
    new_n6498_, new_n6499_, new_n6500_, new_n6501_, new_n6502_, new_n6503_,
    new_n6504_, new_n6505_, new_n6506_, new_n6507_, new_n6508_, new_n6509_,
    new_n6510_, new_n6511_, new_n6512_, new_n6513_, new_n6514_, new_n6515_,
    new_n6516_, new_n6517_, new_n6518_, new_n6519_, new_n6520_, new_n6521_,
    new_n6522_, new_n6523_, new_n6524_, new_n6525_, new_n6526_, new_n6527_,
    new_n6528_, new_n6529_, new_n6530_, new_n6531_, new_n6532_, new_n6533_,
    new_n6534_, new_n6535_, new_n6536_, new_n6537_, new_n6538_, new_n6539_,
    new_n6540_, new_n6541_, new_n6542_, new_n6543_, new_n6544_, new_n6545_,
    new_n6546_, new_n6547_, new_n6548_, new_n6549_, new_n6550_, new_n6551_,
    new_n6552_, new_n6553_, new_n6554_, new_n6555_, new_n6556_, new_n6557_,
    new_n6558_, new_n6559_, new_n6560_, new_n6561_, new_n6562_, new_n6563_,
    new_n6564_, new_n6565_, new_n6566_, new_n6567_, new_n6568_, new_n6569_,
    new_n6570_, new_n6571_, new_n6572_, new_n6573_, new_n6574_, new_n6575_,
    new_n6576_, new_n6577_, new_n6578_, new_n6579_, new_n6580_, new_n6581_,
    new_n6582_, new_n6583_, new_n6584_, new_n6585_, new_n6586_, new_n6587_,
    new_n6588_, new_n6589_, new_n6590_, new_n6591_, new_n6592_, new_n6593_,
    new_n6594_, new_n6595_, new_n6596_, new_n6597_, new_n6598_, new_n6599_,
    new_n6600_, new_n6601_, new_n6602_, new_n6603_, new_n6604_, new_n6605_,
    new_n6606_, new_n6607_, new_n6608_, new_n6609_, new_n6610_, new_n6611_,
    new_n6612_, new_n6613_, new_n6614_, new_n6615_, new_n6616_, new_n6617_,
    new_n6618_, new_n6619_, new_n6620_, new_n6621_, new_n6622_, new_n6623_,
    new_n6624_, new_n6625_, new_n6626_, new_n6627_, new_n6628_, new_n6629_,
    new_n6630_, new_n6631_, new_n6632_, new_n6633_, new_n6634_, new_n6635_,
    new_n6636_, new_n6637_, new_n6638_, new_n6639_, new_n6640_, new_n6641_,
    new_n6642_, new_n6643_, new_n6644_, new_n6645_, new_n6646_, new_n6647_,
    new_n6648_, new_n6649_, new_n6650_, new_n6651_, new_n6652_, new_n6653_,
    new_n6654_, new_n6655_, new_n6656_, new_n6657_, new_n6658_, new_n6659_,
    new_n6660_, new_n6661_, new_n6662_, new_n6663_, new_n6664_, new_n6665_,
    new_n6666_, new_n6667_, new_n6668_, new_n6669_, new_n6670_, new_n6671_,
    new_n6672_, new_n6673_, new_n6674_, new_n6675_, new_n6676_, new_n6677_,
    new_n6678_, new_n6679_, new_n6680_, new_n6681_, new_n6682_, new_n6683_,
    new_n6684_, new_n6685_, new_n6686_, new_n6687_, new_n6688_, new_n6689_,
    new_n6690_, new_n6691_, new_n6692_, new_n6693_, new_n6694_, new_n6695_,
    new_n6696_, new_n6697_, new_n6698_, new_n6699_, new_n6700_, new_n6701_,
    new_n6702_, new_n6703_, new_n6704_, new_n6705_, new_n6706_, new_n6707_,
    new_n6708_, new_n6709_, new_n6710_, new_n6711_, new_n6712_, new_n6713_,
    new_n6714_, new_n6715_, new_n6716_, new_n6717_, new_n6718_, new_n6719_,
    new_n6720_, new_n6721_, new_n6722_, new_n6723_, new_n6724_, new_n6725_,
    new_n6726_, new_n6727_, new_n6728_, new_n6729_, new_n6730_, new_n6731_,
    new_n6732_, new_n6733_, new_n6734_, new_n6735_, new_n6736_, new_n6737_,
    new_n6738_, new_n6739_, new_n6740_, new_n6741_, new_n6742_, new_n6743_,
    new_n6744_, new_n6745_, new_n6746_, new_n6747_, new_n6748_, new_n6749_,
    new_n6750_, new_n6751_, new_n6752_, new_n6753_, new_n6754_, new_n6755_,
    new_n6756_, new_n6757_, new_n6758_, new_n6759_, new_n6760_, new_n6761_,
    new_n6762_, new_n6763_, new_n6764_, new_n6765_, new_n6766_, new_n6767_,
    new_n6768_, new_n6769_, new_n6770_, new_n6771_, new_n6772_, new_n6773_,
    new_n6774_, new_n6775_, new_n6776_, new_n6777_, new_n6778_, new_n6779_,
    new_n6780_, new_n6781_, new_n6782_, new_n6783_, new_n6784_, new_n6785_,
    new_n6786_, new_n6787_, new_n6788_, new_n6789_, new_n6790_, new_n6791_,
    new_n6792_, new_n6793_, new_n6794_, new_n6795_, new_n6796_, new_n6797_,
    new_n6798_, new_n6799_, new_n6800_, new_n6801_, new_n6802_, new_n6803_,
    new_n6804_, new_n6805_, new_n6806_, new_n6807_, new_n6808_, new_n6809_,
    new_n6810_, new_n6811_, new_n6812_, new_n6813_, new_n6814_, new_n6815_,
    new_n6816_, new_n6817_, new_n6818_, new_n6819_, new_n6820_, new_n6821_,
    new_n6822_, new_n6823_, new_n6824_, new_n6825_, new_n6826_, new_n6827_,
    new_n6828_, new_n6829_, new_n6830_, new_n6831_, new_n6832_, new_n6833_,
    new_n6834_, new_n6835_, new_n6836_, new_n6837_, new_n6838_, new_n6839_,
    new_n6840_, new_n6841_, new_n6842_, new_n6843_, new_n6844_, new_n6845_,
    new_n6846_, new_n6847_, new_n6848_, new_n6849_, new_n6850_, new_n6851_,
    new_n6852_, new_n6853_, new_n6854_, new_n6855_, new_n6856_, new_n6857_,
    new_n6858_, new_n6859_, new_n6860_, new_n6861_, new_n6862_, new_n6863_,
    new_n6864_, new_n6865_, new_n6866_, new_n6867_, new_n6868_, new_n6869_,
    new_n6870_, new_n6871_, new_n6872_, new_n6873_, new_n6874_, new_n6875_,
    new_n6876_, new_n6877_, new_n6878_, new_n6879_, new_n6880_, new_n6881_,
    new_n6882_, new_n6883_, new_n6884_, new_n6885_, new_n6886_, new_n6887_,
    new_n6888_, new_n6889_, new_n6890_, new_n6891_, new_n6892_, new_n6893_,
    new_n6894_, new_n6895_, new_n6896_, new_n6897_, new_n6898_, new_n6899_,
    new_n6900_, new_n6901_, new_n6902_, new_n6903_, new_n6904_, new_n6905_,
    new_n6906_, new_n6907_, new_n6908_, new_n6909_, new_n6910_, new_n6911_,
    new_n6912_, new_n6913_, new_n6914_, new_n6915_, new_n6916_, new_n6917_,
    new_n6918_, new_n6919_, new_n6920_, new_n6921_, new_n6922_, new_n6923_,
    new_n6924_, new_n6925_, new_n6926_, new_n6927_, new_n6928_, new_n6929_,
    new_n6930_, new_n6931_, new_n6932_, new_n6933_, new_n6934_, new_n6935_,
    new_n6936_, new_n6937_, new_n6938_, new_n6939_, new_n6940_, new_n6941_,
    new_n6942_, new_n6943_, new_n6944_, new_n6945_, new_n6946_, new_n6947_,
    new_n6948_, new_n6949_, new_n6950_, new_n6951_, new_n6952_, new_n6953_,
    new_n6954_, new_n6955_, new_n6956_, new_n6957_, new_n6958_, new_n6959_,
    new_n6960_, new_n6961_, new_n6962_, new_n6963_, new_n6964_, new_n6965_,
    new_n6966_, new_n6967_, new_n6968_, new_n6969_, new_n6970_, new_n6971_,
    new_n6972_, new_n6973_, new_n6974_, new_n6975_, new_n6976_, new_n6977_,
    new_n6978_, new_n6979_, new_n6980_, new_n6981_, new_n6982_, new_n6983_,
    new_n6984_, new_n6985_, new_n6986_, new_n6987_, new_n6988_, new_n6989_,
    new_n6990_, new_n6991_, new_n6992_, new_n6993_, new_n6994_, new_n6995_,
    new_n6996_, new_n6997_, new_n6998_, new_n6999_, new_n7000_, new_n7001_,
    new_n7002_, new_n7003_, new_n7004_, new_n7005_, new_n7006_, new_n7007_,
    new_n7008_, new_n7009_, new_n7010_, new_n7011_, new_n7012_, new_n7013_,
    new_n7014_, new_n7015_, new_n7016_, new_n7017_, new_n7018_, new_n7019_,
    new_n7020_, new_n7021_, new_n7022_, new_n7023_, new_n7024_, new_n7025_,
    new_n7026_, new_n7027_, new_n7028_, new_n7029_, new_n7030_, new_n7031_,
    new_n7032_, new_n7033_, new_n7034_, new_n7035_, new_n7036_, new_n7037_,
    new_n7038_, new_n7039_, new_n7040_, new_n7041_, new_n7042_, new_n7043_,
    new_n7044_, new_n7045_, new_n7046_, new_n7047_, new_n7048_, new_n7049_,
    new_n7050_, new_n7051_, new_n7052_, new_n7053_, new_n7054_, new_n7055_,
    new_n7056_, new_n7057_, new_n7058_, new_n7059_, new_n7060_, new_n7061_,
    new_n7062_, new_n7063_, new_n7064_, new_n7065_, new_n7066_, new_n7067_,
    new_n7068_, new_n7069_, new_n7070_, new_n7071_, new_n7072_, new_n7073_,
    new_n7074_, new_n7075_, new_n7076_, new_n7077_, new_n7078_, new_n7079_,
    new_n7080_, new_n7081_, new_n7082_, new_n7083_, new_n7084_, new_n7085_,
    new_n7086_, new_n7087_, new_n7088_, new_n7089_, new_n7090_, new_n7091_,
    new_n7092_, new_n7093_, new_n7094_, new_n7095_, new_n7096_, new_n7097_,
    new_n7098_, new_n7099_, new_n7100_, new_n7101_, new_n7102_, new_n7103_,
    new_n7104_, new_n7105_, new_n7106_, new_n7107_, new_n7108_, new_n7109_,
    new_n7110_, new_n7111_, new_n7112_, new_n7113_, new_n7114_, new_n7115_,
    new_n7116_, new_n7117_, new_n7118_, new_n7119_, new_n7120_, new_n7121_,
    new_n7122_, new_n7123_, new_n7124_, new_n7125_, new_n7126_, new_n7127_,
    new_n7128_, new_n7129_, new_n7130_, new_n7131_, new_n7132_, new_n7133_,
    new_n7134_, new_n7135_, new_n7136_, new_n7137_, new_n7138_, new_n7139_,
    new_n7140_, new_n7141_, new_n7142_, new_n7143_, new_n7144_, new_n7145_,
    new_n7146_, new_n7147_, new_n7148_, new_n7149_, new_n7150_, new_n7151_,
    new_n7152_, new_n7153_, new_n7154_, new_n7155_, new_n7156_, new_n7157_,
    new_n7158_, new_n7159_, new_n7160_, new_n7161_, new_n7162_, new_n7163_,
    new_n7164_, new_n7165_, new_n7166_, new_n7167_, new_n7168_, new_n7169_,
    new_n7170_, new_n7171_, new_n7172_, new_n7173_, new_n7174_, new_n7175_,
    new_n7176_, new_n7177_, new_n7178_, new_n7179_, new_n7180_, new_n7181_,
    new_n7182_, new_n7183_, new_n7184_, new_n7185_, new_n7186_, new_n7187_,
    new_n7188_, new_n7189_, new_n7190_, new_n7191_, new_n7192_, new_n7193_,
    new_n7194_, new_n7195_, new_n7196_, new_n7197_, new_n7198_, new_n7199_,
    new_n7200_, new_n7201_, new_n7202_, new_n7203_, new_n7204_, new_n7205_,
    new_n7206_, new_n7207_, new_n7208_, new_n7209_, new_n7210_, new_n7211_,
    new_n7212_, new_n7213_, new_n7214_, new_n7215_, new_n7216_, new_n7217_,
    new_n7218_, new_n7219_, new_n7220_, new_n7221_, new_n7222_, new_n7223_,
    new_n7224_, new_n7225_, new_n7226_, new_n7227_, new_n7228_, new_n7229_,
    new_n7230_, new_n7231_, new_n7232_, new_n7233_, new_n7234_, new_n7235_,
    new_n7236_, new_n7237_, new_n7238_, new_n7239_, new_n7240_, new_n7241_,
    new_n7242_, new_n7243_, new_n7244_, new_n7245_, new_n7246_, new_n7247_,
    new_n7248_, new_n7249_, new_n7250_, new_n7251_, new_n7252_, new_n7253_,
    new_n7254_, new_n7255_, new_n7256_, new_n7257_, new_n7258_, new_n7259_,
    new_n7260_, new_n7261_, new_n7262_, new_n7263_, new_n7264_, new_n7265_,
    new_n7266_, new_n7267_, new_n7268_, new_n7269_, new_n7270_, new_n7271_,
    new_n7272_, new_n7273_, new_n7274_, new_n7275_, new_n7276_, new_n7277_,
    new_n7278_, new_n7279_, new_n7280_, new_n7281_, new_n7282_, new_n7283_,
    new_n7284_, new_n7285_, new_n7286_, new_n7287_, new_n7288_, new_n7289_,
    new_n7290_, new_n7291_, new_n7292_, new_n7293_, new_n7294_, new_n7295_,
    new_n7296_, new_n7297_, new_n7298_, new_n7299_, new_n7300_, new_n7301_,
    new_n7302_, new_n7303_, new_n7304_, new_n7305_, new_n7306_, new_n7307_,
    new_n7308_, new_n7309_, new_n7310_, new_n7311_, new_n7312_, new_n7313_,
    new_n7314_, new_n7315_, new_n7316_, new_n7317_, new_n7318_, new_n7319_,
    new_n7320_, new_n7321_, new_n7322_, new_n7323_, new_n7324_, new_n7325_,
    new_n7326_, new_n7327_, new_n7328_, new_n7329_, new_n7330_, new_n7331_,
    new_n7332_, new_n7333_, new_n7334_, new_n7335_, new_n7336_, new_n7337_,
    new_n7338_, new_n7339_, new_n7340_, new_n7341_, new_n7342_, new_n7343_,
    new_n7344_, new_n7345_, new_n7346_, new_n7347_, new_n7348_, new_n7349_,
    new_n7350_, new_n7351_, new_n7352_, new_n7353_, new_n7354_, new_n7355_,
    new_n7356_, new_n7357_, new_n7358_, new_n7359_, new_n7360_, new_n7361_,
    new_n7362_, new_n7363_, new_n7364_, new_n7365_, new_n7366_, new_n7367_,
    new_n7368_, new_n7369_, new_n7370_, new_n7371_, new_n7372_, new_n7373_,
    new_n7374_, new_n7375_, new_n7376_, new_n7377_, new_n7378_, new_n7379_,
    new_n7380_, new_n7381_, new_n7382_, new_n7383_, new_n7384_, new_n7385_,
    new_n7386_, new_n7387_, new_n7388_, new_n7389_, new_n7390_, new_n7391_,
    new_n7392_, new_n7393_, new_n7394_, new_n7395_, new_n7396_, new_n7397_,
    new_n7398_, new_n7399_, new_n7400_, new_n7401_, new_n7402_, new_n7403_,
    new_n7404_, new_n7405_, new_n7406_, new_n7407_, new_n7408_, new_n7409_,
    new_n7410_, new_n7411_, new_n7412_, new_n7413_, new_n7414_, new_n7415_,
    new_n7416_, new_n7417_, new_n7418_, new_n7419_, new_n7420_, new_n7421_,
    new_n7422_, new_n7423_, new_n7424_, new_n7425_, new_n7426_, new_n7427_,
    new_n7428_, new_n7429_, new_n7430_, new_n7431_, new_n7432_, new_n7433_,
    new_n7434_, new_n7435_, new_n7436_, new_n7437_, new_n7438_, new_n7439_,
    new_n7440_, new_n7441_, new_n7442_, new_n7443_, new_n7444_, new_n7445_,
    new_n7446_, new_n7447_, new_n7448_, new_n7449_, new_n7450_, new_n7451_,
    new_n7452_, new_n7453_, new_n7454_, new_n7455_, new_n7456_, new_n7457_,
    new_n7458_, new_n7459_, new_n7460_, new_n7461_, new_n7462_, new_n7463_,
    new_n7464_, new_n7465_, new_n7466_, new_n7467_, new_n7468_, new_n7469_,
    new_n7470_, new_n7471_, new_n7472_, new_n7473_, new_n7474_, new_n7475_,
    new_n7476_, new_n7477_, new_n7478_, new_n7479_, new_n7480_, new_n7481_,
    new_n7482_, new_n7483_, new_n7484_, new_n7485_, new_n7486_, new_n7487_,
    new_n7488_, new_n7489_, new_n7490_, new_n7491_, new_n7492_, new_n7493_,
    new_n7494_, new_n7495_, new_n7496_, new_n7497_, new_n7498_, new_n7499_,
    new_n7500_, new_n7501_, new_n7502_, new_n7503_, new_n7504_, new_n7505_,
    new_n7506_, new_n7507_, new_n7508_, new_n7509_, new_n7510_, new_n7511_,
    new_n7512_, new_n7513_, new_n7514_, new_n7515_, new_n7516_, new_n7517_,
    new_n7518_, new_n7519_, new_n7520_, new_n7521_, new_n7522_, new_n7523_,
    new_n7524_, new_n7525_, new_n7526_, new_n7527_, new_n7528_, new_n7529_,
    new_n7530_, new_n7531_, new_n7532_, new_n7533_, new_n7534_, new_n7535_,
    new_n7536_, new_n7537_, new_n7538_, new_n7539_, new_n7540_, new_n7541_,
    new_n7542_, new_n7543_, new_n7544_, new_n7545_, new_n7546_, new_n7547_,
    new_n7548_, new_n7549_, new_n7550_, new_n7551_, new_n7552_, new_n7553_,
    new_n7554_, new_n7555_, new_n7556_, new_n7557_, new_n7558_, new_n7559_,
    new_n7560_, new_n7561_, new_n7562_, new_n7563_, new_n7564_, new_n7565_,
    new_n7566_, new_n7567_, new_n7568_, new_n7569_, new_n7570_, new_n7571_,
    new_n7572_, new_n7573_, new_n7574_, new_n7575_, new_n7576_, new_n7577_,
    new_n7578_, new_n7579_, new_n7580_, new_n7581_, new_n7582_, new_n7583_,
    new_n7584_, new_n7585_, new_n7586_, new_n7587_, new_n7588_, new_n7589_,
    new_n7590_, new_n7591_, new_n7592_, new_n7593_, new_n7594_, new_n7595_,
    new_n7596_, new_n7597_, new_n7598_, new_n7599_, new_n7600_, new_n7601_,
    new_n7602_, new_n7603_, new_n7604_, new_n7605_, new_n7606_, new_n7607_,
    new_n7608_, new_n7609_, new_n7610_, new_n7611_, new_n7612_, new_n7613_,
    new_n7614_, new_n7615_, new_n7616_, new_n7617_, new_n7618_, new_n7619_,
    new_n7620_, new_n7621_, new_n7622_, new_n7623_, new_n7624_, new_n7625_,
    new_n7626_, new_n7627_, new_n7628_, new_n7629_, new_n7630_, new_n7631_,
    new_n7632_, new_n7633_, new_n7634_, new_n7635_, new_n7636_, new_n7637_,
    new_n7638_, new_n7639_, new_n7640_, new_n7641_, new_n7642_, new_n7643_,
    new_n7644_, new_n7645_, new_n7646_, new_n7647_, new_n7648_, new_n7649_,
    new_n7650_, new_n7651_, new_n7652_, new_n7653_, new_n7654_, new_n7655_,
    new_n7656_, new_n7657_, new_n7658_, new_n7659_, new_n7660_, new_n7661_,
    new_n7662_, new_n7663_, new_n7664_, new_n7665_, new_n7666_, new_n7667_,
    new_n7668_, new_n7669_, new_n7670_, new_n7671_, new_n7672_, new_n7673_,
    new_n7674_, new_n7675_, new_n7676_, new_n7677_, new_n7678_, new_n7679_,
    new_n7680_, new_n7681_, new_n7682_, new_n7683_, new_n7684_, new_n7685_,
    new_n7686_, new_n7687_, new_n7688_, new_n7689_, new_n7690_, new_n7691_,
    new_n7692_, new_n7693_, new_n7694_, new_n7695_, new_n7696_, new_n7697_,
    new_n7698_, new_n7699_, new_n7700_, new_n7701_, new_n7702_, new_n7703_,
    new_n7704_, new_n7705_, new_n7706_, new_n7707_, new_n7708_, new_n7709_,
    new_n7710_, new_n7711_, new_n7712_, new_n7713_, new_n7714_, new_n7715_,
    new_n7716_, new_n7717_, new_n7718_, new_n7719_, new_n7720_, new_n7721_,
    new_n7722_, new_n7723_, new_n7724_, new_n7725_, new_n7726_, new_n7727_,
    new_n7728_, new_n7729_, new_n7730_, new_n7731_, new_n7732_, new_n7733_,
    new_n7734_, new_n7735_, new_n7736_, new_n7737_, new_n7738_, new_n7739_,
    new_n7740_, new_n7741_, new_n7742_, new_n7743_, new_n7744_, new_n7745_,
    new_n7746_, new_n7747_, new_n7748_, new_n7749_, new_n7750_, new_n7751_,
    new_n7752_, new_n7753_, new_n7754_, new_n7755_, new_n7756_, new_n7757_,
    new_n7758_, new_n7759_, new_n7760_, new_n7761_, new_n7762_, new_n7763_,
    new_n7764_, new_n7765_, new_n7766_, new_n7767_, new_n7768_, new_n7769_,
    new_n7770_, new_n7771_, new_n7772_, new_n7773_, new_n7774_, new_n7775_,
    new_n7776_, new_n7777_, new_n7778_, new_n7779_, new_n7780_, new_n7781_,
    new_n7782_, new_n7783_, new_n7784_, new_n7785_, new_n7786_, new_n7787_,
    new_n7788_, new_n7789_, new_n7790_, new_n7791_, new_n7792_, new_n7793_,
    new_n7794_, new_n7795_, new_n7796_, new_n7797_, new_n7798_, new_n7799_,
    new_n7800_, new_n7801_, new_n7802_, new_n7803_, new_n7804_, new_n7805_,
    new_n7806_, new_n7807_, new_n7808_, new_n7809_, new_n7810_, new_n7811_,
    new_n7812_, new_n7813_, new_n7814_, new_n7815_, new_n7816_, new_n7817_,
    new_n7818_, new_n7819_, new_n7820_, new_n7821_, new_n7822_, new_n7823_,
    new_n7824_, new_n7825_, new_n7826_, new_n7827_, new_n7828_, new_n7829_,
    new_n7830_, new_n7831_, new_n7832_, new_n7833_, new_n7834_, new_n7835_,
    new_n7836_, new_n7837_, new_n7838_, new_n7839_, new_n7840_, new_n7841_,
    new_n7842_, new_n7843_, new_n7844_, new_n7845_, new_n7846_, new_n7847_,
    new_n7848_, new_n7849_, new_n7850_, new_n7851_, new_n7852_, new_n7853_,
    new_n7854_, new_n7855_, new_n7856_, new_n7857_, new_n7858_, new_n7859_,
    new_n7860_, new_n7861_, new_n7862_, new_n7863_, new_n7864_, new_n7865_,
    new_n7866_, new_n7867_, new_n7868_, new_n7869_, new_n7870_, new_n7871_,
    new_n7872_, new_n7873_, new_n7874_, new_n7875_, new_n7876_, new_n7877_,
    new_n7878_, new_n7879_, new_n7880_, new_n7881_, new_n7882_, new_n7883_,
    new_n7884_, new_n7885_, new_n7886_, new_n7887_, new_n7888_, new_n7889_,
    new_n7890_, new_n7891_, new_n7892_, new_n7893_, new_n7894_, new_n7895_,
    new_n7896_, new_n7897_, new_n7898_, new_n7899_, new_n7900_, new_n7901_,
    new_n7902_, new_n7903_, new_n7904_, new_n7905_, new_n7906_, new_n7907_,
    new_n7908_, new_n7909_, new_n7910_, new_n7911_, new_n7912_, new_n7913_,
    new_n7914_, new_n7915_, new_n7916_, new_n7917_, new_n7918_, new_n7919_,
    new_n7920_, new_n7921_, new_n7922_, new_n7923_, new_n7924_, new_n7925_,
    new_n7926_, new_n7927_, new_n7928_, new_n7929_, new_n7930_, new_n7931_,
    new_n7932_, new_n7933_, new_n7934_, new_n7935_, new_n7936_, new_n7937_,
    new_n7938_, new_n7939_, new_n7940_, new_n7941_, new_n7942_, new_n7943_,
    new_n7944_, new_n7945_, new_n7946_, new_n7947_, new_n7948_, new_n7949_,
    new_n7950_, new_n7951_, new_n7952_, new_n7953_, new_n7954_, new_n7955_,
    new_n7956_, new_n7957_, new_n7958_, new_n7959_, new_n7960_, new_n7961_,
    new_n7962_, new_n7963_, new_n7964_, new_n7965_, new_n7966_, new_n7967_,
    new_n7968_, new_n7969_, new_n7970_, new_n7971_, new_n7972_, new_n7973_,
    new_n7974_, new_n7975_, new_n7976_, new_n7977_, new_n7978_, new_n7979_,
    new_n7980_, new_n7981_, new_n7982_, new_n7983_, new_n7984_, new_n7985_,
    new_n7986_, new_n7987_, new_n7988_, new_n7989_, new_n7990_, new_n7991_,
    new_n7992_, new_n7993_, new_n7994_, new_n7995_, new_n7996_, new_n7997_,
    new_n7998_, new_n7999_, new_n8000_, new_n8001_, new_n8002_, new_n8003_,
    new_n8004_, new_n8005_, new_n8006_, new_n8007_, new_n8008_, new_n8009_,
    new_n8010_, new_n8011_, new_n8012_, new_n8013_, new_n8014_, new_n8015_,
    new_n8016_, new_n8017_, new_n8018_, new_n8019_, new_n8020_, new_n8021_,
    new_n8022_, new_n8023_, new_n8024_, new_n8025_, new_n8026_, new_n8027_,
    new_n8028_, new_n8029_, new_n8030_, new_n8031_, new_n8032_, new_n8033_,
    new_n8034_, new_n8035_, new_n8036_, new_n8037_, new_n8038_, new_n8039_,
    new_n8040_, new_n8041_, new_n8042_, new_n8043_, new_n8044_, new_n8045_,
    new_n8046_, new_n8047_, new_n8048_, new_n8049_, new_n8050_, new_n8051_,
    new_n8052_, new_n8053_, new_n8054_, new_n8055_, new_n8056_, new_n8057_,
    new_n8058_, new_n8059_, new_n8060_, new_n8061_, new_n8062_, new_n8063_,
    new_n8064_, new_n8065_, new_n8066_, new_n8067_, new_n8068_, new_n8069_,
    new_n8070_, new_n8071_, new_n8072_, new_n8073_, new_n8074_, new_n8075_,
    new_n8076_, new_n8077_, new_n8078_, new_n8079_, new_n8080_, new_n8081_,
    new_n8082_, new_n8083_, new_n8084_, new_n8085_, new_n8086_, new_n8087_,
    new_n8088_, new_n8089_, new_n8090_, new_n8091_, new_n8092_, new_n8093_,
    new_n8094_, new_n8095_, new_n8096_, new_n8097_, new_n8098_, new_n8099_,
    new_n8100_, new_n8101_, new_n8102_, new_n8103_, new_n8104_, new_n8105_,
    new_n8106_, new_n8107_, new_n8108_, new_n8109_, new_n8110_, new_n8111_,
    new_n8112_, new_n8113_, new_n8114_, new_n8115_, new_n8116_, new_n8117_,
    new_n8118_, new_n8119_, new_n8120_, new_n8121_, new_n8122_, new_n8123_,
    new_n8124_, new_n8125_, new_n8126_, new_n8127_, new_n8128_, new_n8129_,
    new_n8130_, new_n8131_, new_n8132_, new_n8133_, new_n8134_, new_n8135_,
    new_n8136_, new_n8137_, new_n8138_, new_n8139_, new_n8140_, new_n8141_,
    new_n8142_, new_n8143_, new_n8144_, new_n8145_, new_n8146_, new_n8147_,
    new_n8148_, new_n8149_, new_n8150_, new_n8151_, new_n8152_, new_n8153_,
    new_n8154_, new_n8155_, new_n8156_, new_n8157_, new_n8158_, new_n8159_,
    new_n8160_, new_n8161_, new_n8162_, new_n8163_, new_n8164_, new_n8165_,
    new_n8166_, new_n8167_, new_n8168_, new_n8169_, new_n8170_, new_n8171_,
    new_n8172_, new_n8173_, new_n8174_, new_n8175_, new_n8176_, new_n8177_,
    new_n8178_, new_n8179_, new_n8180_, new_n8181_, new_n8182_, new_n8183_,
    new_n8184_, new_n8185_, new_n8186_, new_n8187_, new_n8188_, new_n8189_,
    new_n8190_, new_n8191_, new_n8192_, new_n8193_, new_n8194_, new_n8195_,
    new_n8196_, new_n8197_, new_n8198_, new_n8199_, new_n8200_, new_n8201_,
    new_n8202_, new_n8203_, new_n8204_, new_n8205_, new_n8206_, new_n8207_,
    new_n8208_, new_n8209_, new_n8210_, new_n8211_, new_n8212_, new_n8213_,
    new_n8214_, new_n8215_, new_n8216_, new_n8217_, new_n8218_, new_n8219_,
    new_n8220_, new_n8221_, new_n8222_, new_n8223_, new_n8224_, new_n8225_,
    new_n8226_, new_n8227_, new_n8228_, new_n8229_, new_n8230_, new_n8231_,
    new_n8232_, new_n8233_, new_n8234_, new_n8235_, new_n8236_, new_n8237_,
    new_n8238_, new_n8239_, new_n8240_, new_n8241_, new_n8242_, new_n8243_,
    new_n8244_, new_n8245_, new_n8246_, new_n8247_, new_n8248_, new_n8249_,
    new_n8250_, new_n8251_, new_n8252_, new_n8253_, new_n8254_, new_n8255_,
    new_n8256_, new_n8257_, new_n8258_, new_n8259_, new_n8260_, new_n8261_,
    new_n8262_, new_n8263_, new_n8264_, new_n8265_, new_n8266_, new_n8267_,
    new_n8268_, new_n8269_, new_n8270_, new_n8271_, new_n8272_, new_n8273_,
    new_n8274_, new_n8275_, new_n8276_, new_n8277_, new_n8278_, new_n8279_,
    new_n8280_, new_n8281_, new_n8282_, new_n8283_, new_n8284_, new_n8285_,
    new_n8286_, new_n8287_, new_n8288_, new_n8289_, new_n8290_, new_n8291_,
    new_n8292_, new_n8293_, new_n8294_, new_n8295_, new_n8296_, new_n8297_,
    new_n8298_, new_n8299_, new_n8300_, new_n8301_, new_n8302_, new_n8303_,
    new_n8304_, new_n8305_, new_n8306_, new_n8307_, new_n8308_, new_n8309_,
    new_n8310_, new_n8311_, new_n8312_, new_n8313_, new_n8314_, new_n8315_,
    new_n8316_, new_n8317_, new_n8318_, new_n8319_, new_n8320_, new_n8321_,
    new_n8322_, new_n8323_, new_n8324_, new_n8325_, new_n8326_, new_n8327_,
    new_n8328_, new_n8329_, new_n8330_, new_n8331_, new_n8332_, new_n8333_,
    new_n8334_, new_n8335_, new_n8336_, new_n8337_, new_n8338_, new_n8339_,
    new_n8340_, new_n8341_, new_n8342_, new_n8343_, new_n8344_, new_n8345_,
    new_n8346_, new_n8347_, new_n8348_, new_n8349_, new_n8350_, new_n8351_,
    new_n8352_, new_n8353_, new_n8354_, new_n8355_, new_n8356_, new_n8357_,
    new_n8358_, new_n8359_, new_n8360_, new_n8361_, new_n8362_, new_n8363_,
    new_n8364_, new_n8365_, new_n8366_, new_n8367_, new_n8368_, new_n8369_,
    new_n8370_, new_n8371_, new_n8372_, new_n8373_, new_n8374_, new_n8375_,
    new_n8376_, new_n8377_, new_n8378_, new_n8379_, new_n8380_, new_n8381_,
    new_n8382_, new_n8383_, new_n8384_, new_n8385_, new_n8386_, new_n8387_,
    new_n8388_, new_n8389_, new_n8390_, new_n8391_, new_n8392_, new_n8393_,
    new_n8394_, new_n8395_, new_n8396_, new_n8397_, new_n8398_, new_n8399_,
    new_n8400_, new_n8401_, new_n8402_, new_n8403_, new_n8404_, new_n8405_,
    new_n8406_, new_n8407_, new_n8408_, new_n8409_, new_n8410_, new_n8411_,
    new_n8412_, new_n8413_, new_n8414_, new_n8415_, new_n8416_, new_n8417_,
    new_n8418_, new_n8419_, new_n8420_, new_n8421_, new_n8422_, new_n8423_,
    new_n8424_, new_n8425_, new_n8426_, new_n8427_, new_n8428_, new_n8429_,
    new_n8430_, new_n8431_, new_n8432_, new_n8433_, new_n8434_, new_n8435_,
    new_n8436_, new_n8437_, new_n8438_, new_n8439_, new_n8440_, new_n8441_,
    new_n8442_, new_n8443_, new_n8444_, new_n8445_, new_n8446_, new_n8447_,
    new_n8448_, new_n8449_, new_n8450_, new_n8451_, new_n8452_, new_n8453_,
    new_n8454_, new_n8455_, new_n8456_, new_n8457_, new_n8458_, new_n8459_,
    new_n8460_, new_n8461_, new_n8462_, new_n8463_, new_n8464_, new_n8465_,
    new_n8466_, new_n8467_, new_n8468_, new_n8469_, new_n8470_, new_n8471_,
    new_n8472_, new_n8473_, new_n8474_, new_n8475_, new_n8476_, new_n8477_,
    new_n8478_, new_n8479_, new_n8480_, new_n8481_, new_n8482_, new_n8483_,
    new_n8484_, new_n8485_, new_n8486_, new_n8487_, new_n8488_, new_n8489_,
    new_n8490_, new_n8491_, new_n8492_, new_n8493_, new_n8494_, new_n8495_,
    new_n8496_, new_n8497_, new_n8498_, new_n8499_, new_n8500_, new_n8501_,
    new_n8502_, new_n8503_, new_n8504_, new_n8505_, new_n8506_, new_n8507_,
    new_n8508_, new_n8509_, new_n8510_, new_n8511_, new_n8512_, new_n8513_,
    new_n8514_, new_n8515_, new_n8516_, new_n8517_, new_n8518_, new_n8519_,
    new_n8520_, new_n8521_, new_n8522_, new_n8523_, new_n8524_, new_n8525_,
    new_n8526_, new_n8527_, new_n8528_, new_n8529_, new_n8530_, new_n8531_,
    new_n8532_, new_n8533_, new_n8534_, new_n8535_, new_n8536_, new_n8537_,
    new_n8538_, new_n8539_, new_n8540_, new_n8541_, new_n8542_, new_n8543_,
    new_n8544_, new_n8545_, new_n8546_, new_n8547_, new_n8548_, new_n8549_,
    new_n8550_, new_n8551_, new_n8552_, new_n8553_, new_n8554_, new_n8555_,
    new_n8556_, new_n8557_, new_n8558_, new_n8559_, new_n8560_, new_n8561_,
    new_n8562_, new_n8563_, new_n8564_, new_n8565_, new_n8566_, new_n8567_,
    new_n8568_, new_n8569_, new_n8570_, new_n8571_, new_n8572_, new_n8573_,
    new_n8574_, new_n8575_, new_n8576_, new_n8577_, new_n8578_, new_n8579_,
    new_n8580_, new_n8581_, new_n8582_, new_n8583_, new_n8584_, new_n8585_,
    new_n8586_, new_n8587_, new_n8588_, new_n8589_, new_n8590_, new_n8591_,
    new_n8592_, new_n8593_, new_n8594_, new_n8595_, new_n8596_, new_n8597_,
    new_n8598_, new_n8599_, new_n8600_, new_n8601_, new_n8602_, new_n8603_,
    new_n8604_, new_n8605_, new_n8606_, new_n8607_, new_n8608_, new_n8609_,
    new_n8610_, new_n8611_, new_n8612_, new_n8613_, new_n8614_, new_n8615_,
    new_n8616_, new_n8617_, new_n8618_, new_n8619_, new_n8620_, new_n8621_,
    new_n8622_, new_n8623_, new_n8624_, new_n8625_, new_n8626_, new_n8627_,
    new_n8628_, new_n8629_, new_n8630_, new_n8631_, new_n8632_, new_n8633_,
    new_n8634_, new_n8635_, new_n8636_, new_n8637_, new_n8638_, new_n8639_,
    new_n8640_, new_n8641_, new_n8642_, new_n8643_, new_n8644_, new_n8645_,
    new_n8646_, new_n8647_, new_n8648_, new_n8649_, new_n8650_, new_n8651_,
    new_n8652_, new_n8653_, new_n8654_, new_n8655_, new_n8656_, new_n8657_,
    new_n8658_, new_n8659_, new_n8660_, new_n8661_, new_n8662_, new_n8663_,
    new_n8664_, new_n8665_, new_n8666_, new_n8667_, new_n8668_, new_n8669_,
    new_n8670_, new_n8671_, new_n8672_, new_n8673_, new_n8674_, new_n8675_,
    new_n8676_, new_n8677_, new_n8678_, new_n8679_, new_n8680_, new_n8681_,
    new_n8682_, new_n8683_, new_n8684_, new_n8685_, new_n8686_, new_n8687_,
    new_n8688_, new_n8689_, new_n8690_, new_n8691_, new_n8692_, new_n8693_,
    new_n8694_, new_n8695_, new_n8696_, new_n8697_, new_n8698_, new_n8699_,
    new_n8700_, new_n8701_, new_n8702_, new_n8703_, new_n8704_, new_n8705_,
    new_n8706_, new_n8707_, new_n8708_, new_n8709_, new_n8710_, new_n8711_,
    new_n8712_, new_n8713_, new_n8714_, new_n8715_, new_n8716_, new_n8717_,
    new_n8718_, new_n8719_, new_n8720_, new_n8721_, new_n8722_, new_n8723_,
    new_n8724_, new_n8725_, new_n8726_, new_n8727_, new_n8728_, new_n8729_,
    new_n8730_, new_n8731_, new_n8732_, new_n8733_, new_n8734_, new_n8735_,
    new_n8736_, new_n8737_, new_n8738_, new_n8739_, new_n8740_, new_n8741_,
    new_n8742_, new_n8743_, new_n8744_, new_n8745_, new_n8746_, new_n8747_,
    new_n8748_, new_n8749_, new_n8750_, new_n8751_, new_n8752_, new_n8753_,
    new_n8754_, new_n8755_, new_n8756_, new_n8757_, new_n8758_, new_n8759_,
    new_n8760_, new_n8761_, new_n8762_, new_n8763_, new_n8764_, new_n8765_,
    new_n8766_, new_n8767_, new_n8768_, new_n8769_, new_n8770_, new_n8771_,
    new_n8772_, new_n8773_, new_n8774_, new_n8775_, new_n8776_, new_n8777_,
    new_n8778_, new_n8779_, new_n8780_, new_n8781_, new_n8782_, new_n8783_,
    new_n8784_, new_n8785_, new_n8786_, new_n8787_, new_n8788_, new_n8789_,
    new_n8790_, new_n8791_, new_n8792_, new_n8793_, new_n8794_, new_n8795_,
    new_n8796_, new_n8797_, new_n8798_, new_n8799_, new_n8800_, new_n8801_,
    new_n8802_, new_n8803_, new_n8804_, new_n8805_, new_n8806_, new_n8807_,
    new_n8808_, new_n8809_, new_n8810_, new_n8811_, new_n8812_, new_n8813_,
    new_n8814_, new_n8815_, new_n8816_, new_n8817_, new_n8818_, new_n8819_,
    new_n8820_, new_n8821_, new_n8822_, new_n8823_, new_n8824_, new_n8825_,
    new_n8826_, new_n8827_, new_n8828_, new_n8829_, new_n8830_, new_n8831_,
    new_n8832_, new_n8833_, new_n8834_, new_n8835_, new_n8836_, new_n8837_,
    new_n8838_, new_n8839_, new_n8840_, new_n8841_, new_n8842_, new_n8843_,
    new_n8844_, new_n8845_, new_n8846_, new_n8847_, new_n8848_, new_n8849_,
    new_n8850_, new_n8851_, new_n8852_, new_n8853_, new_n8854_, new_n8855_,
    new_n8856_, new_n8857_, new_n8858_, new_n8859_, new_n8860_, new_n8861_,
    new_n8862_, new_n8863_, new_n8864_, new_n8865_, new_n8866_, new_n8867_,
    new_n8868_, new_n8869_, new_n8870_, new_n8871_, new_n8872_, new_n8873_,
    new_n8874_, new_n8875_, new_n8876_, new_n8877_, new_n8878_, new_n8879_,
    new_n8880_, new_n8881_, new_n8882_, new_n8883_, new_n8884_, new_n8885_,
    new_n8886_, new_n8887_, new_n8888_, new_n8889_, new_n8890_, new_n8891_,
    new_n8892_, new_n8893_, new_n8894_, new_n8895_, new_n8896_, new_n8897_,
    new_n8898_, new_n8899_, new_n8900_, new_n8901_, new_n8902_, new_n8903_,
    new_n8904_, new_n8905_, new_n8906_, new_n8907_, new_n8908_, new_n8909_,
    new_n8910_, new_n8911_, new_n8912_, new_n8913_, new_n8914_, new_n8915_,
    new_n8916_, new_n8917_, new_n8918_, new_n8919_, new_n8920_, new_n8921_,
    new_n8922_, new_n8923_, new_n8924_, new_n8925_, new_n8926_, new_n8927_,
    new_n8928_, new_n8929_, new_n8930_, new_n8931_, new_n8932_, new_n8933_,
    new_n8934_, new_n8935_, new_n8936_, new_n8937_, new_n8938_, new_n8939_,
    new_n8940_, new_n8941_, new_n8942_, new_n8943_, new_n8944_, new_n8945_,
    new_n8946_, new_n8947_, new_n8948_, new_n8949_, new_n8950_, new_n8951_,
    new_n8952_, new_n8953_, new_n8954_, new_n8955_, new_n8956_, new_n8957_,
    new_n8958_, new_n8959_, new_n8960_, new_n8961_, new_n8962_, new_n8963_,
    new_n8964_, new_n8965_, new_n8966_, new_n8967_, new_n8968_, new_n8969_,
    new_n8970_, new_n8971_, new_n8972_, new_n8973_, new_n8974_, new_n8975_,
    new_n8976_, new_n8977_, new_n8978_, new_n8979_, new_n8980_, new_n8981_,
    new_n8982_, new_n8983_, new_n8984_, new_n8985_, new_n8986_, new_n8987_,
    new_n8988_, new_n8989_, new_n8990_, new_n8991_, new_n8992_, new_n8993_,
    new_n8994_, new_n8995_, new_n8996_, new_n8997_, new_n8998_, new_n8999_,
    new_n9000_, new_n9001_, new_n9002_, new_n9003_, new_n9004_, new_n9005_,
    new_n9006_, new_n9007_, new_n9008_, new_n9009_, new_n9010_, new_n9011_,
    new_n9012_, new_n9013_, new_n9014_, new_n9015_, new_n9016_, new_n9017_,
    new_n9018_, new_n9019_, new_n9020_, new_n9021_, new_n9022_, new_n9023_,
    new_n9024_, new_n9025_, new_n9026_, new_n9027_, new_n9028_, new_n9029_,
    new_n9030_, new_n9031_, new_n9032_, new_n9033_, new_n9034_, new_n9035_,
    new_n9036_, new_n9037_, new_n9038_, new_n9039_, new_n9040_, new_n9041_,
    new_n9042_, new_n9043_, new_n9044_, new_n9045_, new_n9046_, new_n9047_,
    new_n9048_, new_n9049_, new_n9050_, new_n9051_, new_n9052_, new_n9053_,
    new_n9054_, new_n9055_, new_n9056_, new_n9057_, new_n9058_, new_n9059_,
    new_n9060_, new_n9061_, new_n9062_, new_n9063_, new_n9064_, new_n9065_,
    new_n9066_, new_n9067_, new_n9068_, new_n9069_, new_n9070_, new_n9071_,
    new_n9072_, new_n9073_, new_n9074_, new_n9075_, new_n9076_, new_n9077_,
    new_n9078_, new_n9079_, new_n9080_, new_n9081_, new_n9082_, new_n9083_,
    new_n9084_, new_n9085_, new_n9086_, new_n9087_, new_n9088_, new_n9089_,
    new_n9090_, new_n9091_, new_n9092_, new_n9093_, new_n9094_, new_n9095_,
    new_n9096_, new_n9097_, new_n9098_, new_n9099_, new_n9100_, new_n9101_,
    new_n9102_, new_n9103_, new_n9104_, new_n9105_, new_n9106_, new_n9107_,
    new_n9108_, new_n9109_, new_n9110_, new_n9111_, new_n9112_, new_n9113_,
    new_n9114_, new_n9115_, new_n9116_, new_n9117_, new_n9118_, new_n9119_,
    new_n9120_, new_n9121_, new_n9122_, new_n9123_, new_n9124_, new_n9125_,
    new_n9126_, new_n9127_, new_n9128_, new_n9129_, new_n9130_, new_n9131_,
    new_n9132_, new_n9133_, new_n9134_, new_n9135_, new_n9136_, new_n9137_,
    new_n9138_, new_n9139_, new_n9140_, new_n9141_, new_n9142_, new_n9143_,
    new_n9144_, new_n9145_, new_n9146_, new_n9147_, new_n9148_, new_n9149_,
    new_n9150_, new_n9151_, new_n9152_, new_n9153_, new_n9154_, new_n9155_,
    new_n9156_, new_n9157_, new_n9158_, new_n9159_, new_n9160_, new_n9161_,
    new_n9162_, new_n9163_, new_n9164_, new_n9165_, new_n9166_, new_n9167_,
    new_n9168_, new_n9169_, new_n9170_, new_n9171_, new_n9172_, new_n9173_,
    new_n9174_, new_n9175_, new_n9176_, new_n9177_, new_n9178_, new_n9179_,
    new_n9180_, new_n9181_, new_n9182_, new_n9183_, new_n9184_, new_n9185_,
    new_n9186_, new_n9187_, new_n9188_, new_n9189_, new_n9190_, new_n9191_,
    new_n9192_, new_n9193_, new_n9194_, new_n9195_, new_n9196_, new_n9197_,
    new_n9198_, new_n9199_, new_n9200_, new_n9201_, new_n9202_, new_n9203_,
    new_n9204_, new_n9205_, new_n9206_, new_n9207_, new_n9208_, new_n9209_,
    new_n9210_, new_n9211_, new_n9212_, new_n9213_, new_n9214_, new_n9215_,
    new_n9216_, new_n9217_, new_n9218_, new_n9219_, new_n9220_, new_n9221_,
    new_n9222_, new_n9223_, new_n9224_, new_n9225_, new_n9226_, new_n9227_,
    new_n9228_, new_n9229_, new_n9230_, new_n9231_, new_n9232_, new_n9233_,
    new_n9234_, new_n9235_, new_n9236_, new_n9237_, new_n9238_, new_n9239_,
    new_n9240_, new_n9241_, new_n9242_, new_n9243_, new_n9244_, new_n9245_,
    new_n9246_, new_n9247_, new_n9248_, new_n9249_, new_n9250_, new_n9251_,
    new_n9252_, new_n9253_, new_n9254_, new_n9255_, new_n9256_, new_n9257_,
    new_n9258_, new_n9259_, new_n9260_, new_n9261_, new_n9262_, new_n9263_,
    new_n9264_, new_n9265_, new_n9266_, new_n9267_, new_n9268_, new_n9269_,
    new_n9270_, new_n9271_, new_n9272_, new_n9273_, new_n9274_, new_n9275_,
    new_n9276_, new_n9277_, new_n9278_, new_n9279_, new_n9280_, new_n9281_,
    new_n9282_, new_n9283_, new_n9284_, new_n9285_, new_n9286_, new_n9287_,
    new_n9288_, new_n9289_, new_n9290_, new_n9291_, new_n9292_, new_n9293_,
    new_n9294_, new_n9295_, new_n9296_, new_n9297_, new_n9298_, new_n9299_,
    new_n9300_, new_n9301_, new_n9302_, new_n9303_, new_n9304_, new_n9305_,
    new_n9306_, new_n9307_, new_n9308_, new_n9309_, new_n9310_, new_n9311_,
    new_n9312_, new_n9313_, new_n9314_, new_n9315_, new_n9316_, new_n9317_,
    new_n9318_, new_n9319_, new_n9320_, new_n9321_, new_n9322_, new_n9323_,
    new_n9324_, new_n9325_, new_n9326_, new_n9327_, new_n9328_, new_n9329_,
    new_n9330_, new_n9331_, new_n9332_, new_n9333_, new_n9334_, new_n9335_,
    new_n9336_, new_n9337_, new_n9338_, new_n9339_, new_n9340_, new_n9341_,
    new_n9342_, new_n9343_, new_n9344_, new_n9345_, new_n9346_, new_n9347_,
    new_n9348_, new_n9349_, new_n9350_, new_n9351_, new_n9352_, new_n9353_,
    new_n9354_, new_n9355_, new_n9356_, new_n9357_, new_n9358_, new_n9359_,
    new_n9360_, new_n9361_, new_n9362_, new_n9363_, new_n9364_, new_n9365_,
    new_n9366_, new_n9367_, new_n9368_, new_n9369_, new_n9370_, new_n9371_,
    new_n9372_, new_n9373_, new_n9374_, new_n9375_, new_n9376_, new_n9377_,
    new_n9378_, new_n9379_, new_n9380_, new_n9381_, new_n9382_, new_n9383_,
    new_n9384_, new_n9385_, new_n9386_, new_n9387_, new_n9388_, new_n9389_,
    new_n9390_, new_n9391_, new_n9392_, new_n9393_, new_n9394_, new_n9395_,
    new_n9396_, new_n9397_, new_n9398_, new_n9399_, new_n9400_, new_n9401_,
    new_n9402_, new_n9403_, new_n9404_, new_n9405_, new_n9406_, new_n9407_,
    new_n9408_, new_n9409_, new_n9410_, new_n9411_, new_n9412_, new_n9413_,
    new_n9414_, new_n9415_, new_n9416_, new_n9417_, new_n9418_, new_n9419_,
    new_n9420_, new_n9421_, new_n9422_, new_n9423_, new_n9424_, new_n9425_,
    new_n9426_, new_n9427_, new_n9428_, new_n9429_, new_n9430_, new_n9431_,
    new_n9432_, new_n9433_, new_n9434_, new_n9435_, new_n9436_, new_n9437_,
    new_n9438_, new_n9439_, new_n9440_, new_n9441_, new_n9442_, new_n9443_,
    new_n9444_, new_n9445_, new_n9446_, new_n9447_, new_n9448_, new_n9449_,
    new_n9450_, new_n9451_, new_n9452_, new_n9453_, new_n9454_, new_n9455_,
    new_n9456_, new_n9457_, new_n9458_, new_n9459_, new_n9460_, new_n9461_,
    new_n9462_, new_n9463_, new_n9464_, new_n9465_, new_n9466_, new_n9467_,
    new_n9468_, new_n9469_, new_n9470_, new_n9471_, new_n9472_, new_n9473_,
    new_n9474_, new_n9475_, new_n9476_, new_n9477_, new_n9478_, new_n9479_,
    new_n9480_, new_n9481_, new_n9482_, new_n9483_, new_n9484_, new_n9485_,
    new_n9486_, new_n9487_, new_n9488_, new_n9489_, new_n9490_, new_n9491_,
    new_n9492_, new_n9493_, new_n9494_, new_n9495_, new_n9496_, new_n9497_,
    new_n9498_, new_n9499_, new_n9500_, new_n9501_, new_n9502_, new_n9503_,
    new_n9504_, new_n9505_, new_n9506_, new_n9507_, new_n9508_, new_n9509_,
    new_n9510_, new_n9511_, new_n9512_, new_n9513_, new_n9514_, new_n9515_,
    new_n9516_, new_n9517_, new_n9518_, new_n9519_, new_n9520_, new_n9521_,
    new_n9522_, new_n9523_, new_n9524_, new_n9525_, new_n9526_, new_n9527_,
    new_n9528_, new_n9529_, new_n9530_, new_n9531_, new_n9532_, new_n9533_,
    new_n9534_, new_n9535_, new_n9536_, new_n9537_, new_n9538_, new_n9539_,
    new_n9540_, new_n9541_, new_n9542_, new_n9543_, new_n9544_, new_n9545_,
    new_n9546_, new_n9547_, new_n9548_, new_n9549_, new_n9550_, new_n9551_,
    new_n9552_, new_n9553_, new_n9554_, new_n9555_, new_n9556_, new_n9557_,
    new_n9558_, new_n9559_, new_n9560_, new_n9561_, new_n9562_, new_n9563_,
    new_n9564_, new_n9565_, new_n9566_, new_n9567_, new_n9568_, new_n9569_,
    new_n9570_, new_n9571_, new_n9572_, new_n9573_, new_n9574_, new_n9575_,
    new_n9576_, new_n9577_, new_n9578_, new_n9579_, new_n9580_, new_n9581_,
    new_n9582_, new_n9583_, new_n9584_, new_n9585_, new_n9586_, new_n9587_,
    new_n9588_, new_n9589_, new_n9590_, new_n9591_, new_n9592_, new_n9593_,
    new_n9594_, new_n9595_, new_n9596_, new_n9597_, new_n9598_, new_n9599_,
    new_n9600_, new_n9601_, new_n9602_, new_n9603_, new_n9604_, new_n9605_,
    new_n9606_, new_n9607_, new_n9608_, new_n9609_, new_n9610_, new_n9611_,
    new_n9612_, new_n9613_, new_n9614_, new_n9615_, new_n9616_, new_n9617_,
    new_n9618_, new_n9619_, new_n9620_, new_n9621_, new_n9622_, new_n9623_,
    new_n9624_, new_n9625_, new_n9626_, new_n9627_, new_n9628_, new_n9629_,
    new_n9630_, new_n9631_, new_n9632_, new_n9633_, new_n9634_, new_n9635_,
    new_n9636_, new_n9637_, new_n9638_, new_n9639_, new_n9640_, new_n9641_,
    new_n9642_, new_n9643_, new_n9644_, new_n9645_, new_n9646_, new_n9647_,
    new_n9648_, new_n9649_, new_n9650_, new_n9651_, new_n9652_, new_n9653_,
    new_n9654_, new_n9655_, new_n9656_, new_n9657_, new_n9658_, new_n9659_,
    new_n9660_, new_n9661_, new_n9662_, new_n9663_, new_n9664_, new_n9665_,
    new_n9666_, new_n9667_, new_n9668_, new_n9669_, new_n9670_, new_n9671_,
    new_n9672_, new_n9673_, new_n9674_, new_n9675_, new_n9676_, new_n9677_,
    new_n9678_, new_n9679_, new_n9680_, new_n9681_, new_n9682_, new_n9683_,
    new_n9684_, new_n9685_, new_n9686_, new_n9687_, new_n9688_, new_n9689_,
    new_n9690_, new_n9691_, new_n9692_, new_n9693_, new_n9694_, new_n9695_,
    new_n9696_, new_n9697_, new_n9698_, new_n9699_, new_n9700_, new_n9701_,
    new_n9702_, new_n9703_, new_n9704_, new_n9705_, new_n9706_, new_n9707_,
    new_n9708_, new_n9709_, new_n9710_, new_n9711_, new_n9712_, new_n9713_,
    new_n9714_, new_n9715_, new_n9716_, new_n9717_, new_n9718_, new_n9719_,
    new_n9720_, new_n9721_, new_n9722_, new_n9723_, new_n9724_, new_n9725_,
    new_n9726_, new_n9727_, new_n9728_, new_n9729_, new_n9730_, new_n9731_,
    new_n9732_, new_n9733_, new_n9734_, new_n9735_, new_n9736_, new_n9737_,
    new_n9738_, new_n9739_, new_n9740_, new_n9741_, new_n9742_, new_n9743_,
    new_n9744_, new_n9745_, new_n9746_, new_n9747_, new_n9748_, new_n9749_,
    new_n9750_, new_n9751_, new_n9752_, new_n9753_, new_n9754_, new_n9755_,
    new_n9756_, new_n9757_, new_n9758_, new_n9759_, new_n9760_, new_n9761_,
    new_n9762_, new_n9763_, new_n9764_, new_n9765_, new_n9766_, new_n9767_,
    new_n9768_, new_n9769_, new_n9770_, new_n9771_, new_n9772_, new_n9773_,
    new_n9774_, new_n9775_, new_n9776_, new_n9777_, new_n9778_, new_n9779_,
    new_n9780_, new_n9781_, new_n9782_, new_n9783_, new_n9784_, new_n9785_,
    new_n9786_, new_n9787_, new_n9788_, new_n9789_, new_n9790_, new_n9791_,
    new_n9792_, new_n9793_, new_n9794_, new_n9795_, new_n9796_, new_n9797_,
    new_n9798_, new_n9799_, new_n9800_, new_n9801_, new_n9802_, new_n9803_,
    new_n9804_, new_n9805_, new_n9806_, new_n9807_, new_n9808_, new_n9809_,
    new_n9810_, new_n9811_, new_n9812_, new_n9813_, new_n9814_, new_n9815_,
    new_n9816_, new_n9817_, new_n9818_, new_n9819_, new_n9820_, new_n9821_,
    new_n9822_, new_n9823_, new_n9824_, new_n9825_, new_n9826_, new_n9827_,
    new_n9828_, new_n9829_, new_n9830_, new_n9831_, new_n9832_, new_n9833_,
    new_n9834_, new_n9835_, new_n9836_, new_n9837_, new_n9838_, new_n9839_,
    new_n9840_, new_n9841_, new_n9842_, new_n9843_, new_n9844_, new_n9845_,
    new_n9846_, new_n9847_, new_n9848_, new_n9849_, new_n9850_, new_n9851_,
    new_n9852_, new_n9853_, new_n9854_, new_n9855_, new_n9856_, new_n9857_,
    new_n9858_, new_n9859_, new_n9860_, new_n9861_, new_n9862_, new_n9863_,
    new_n9864_, new_n9865_, new_n9866_, new_n9867_, new_n9868_, new_n9869_,
    new_n9870_, new_n9871_, new_n9872_, new_n9873_, new_n9874_, new_n9875_,
    new_n9876_, new_n9877_, new_n9878_, new_n9879_, new_n9880_, new_n9881_,
    new_n9882_, new_n9883_, new_n9884_, new_n9885_, new_n9886_, new_n9887_,
    new_n9888_, new_n9889_, new_n9890_, new_n9891_, new_n9892_, new_n9893_,
    new_n9894_, new_n9895_, new_n9896_, new_n9897_, new_n9898_, new_n9899_,
    new_n9900_, new_n9901_, new_n9902_, new_n9903_, new_n9904_, new_n9905_,
    new_n9906_, new_n9907_, new_n9908_, new_n9909_, new_n9910_, new_n9911_,
    new_n9912_, new_n9913_, new_n9914_, new_n9915_, new_n9916_, new_n9917_,
    new_n9918_, new_n9919_, new_n9920_, new_n9921_, new_n9922_, new_n9923_,
    new_n9924_, new_n9925_, new_n9926_, new_n9927_, new_n9928_, new_n9929_,
    new_n9930_, new_n9931_, new_n9932_, new_n9933_, new_n9934_, new_n9935_,
    new_n9936_, new_n9937_, new_n9938_, new_n9939_, new_n9940_, new_n9941_,
    new_n9942_, new_n9943_, new_n9944_, new_n9945_, new_n9946_, new_n9947_,
    new_n9948_, new_n9949_, new_n9950_, new_n9951_, new_n9952_, new_n9953_,
    new_n9954_, new_n9955_, new_n9956_, new_n9957_, new_n9958_, new_n9959_,
    new_n9960_, new_n9961_, new_n9962_, new_n9963_, new_n9964_, new_n9965_,
    new_n9966_, new_n9967_, new_n9968_, new_n9969_, new_n9970_, new_n9971_,
    new_n9972_, new_n9973_, new_n9974_, new_n9975_, new_n9976_, new_n9977_,
    new_n9978_, new_n9979_, new_n9980_, new_n9981_, new_n9982_, new_n9983_,
    new_n9984_, new_n9985_, new_n9986_, new_n9987_, new_n9988_, new_n9989_,
    new_n9990_, new_n9991_, new_n9992_, new_n9993_, new_n9994_, new_n9995_,
    new_n9996_, new_n9997_, new_n9998_, new_n9999_, new_n10000_,
    new_n10001_, new_n10002_, new_n10003_, new_n10004_, new_n10005_,
    new_n10006_, new_n10007_, new_n10008_, new_n10009_, new_n10010_,
    new_n10011_, new_n10012_, new_n10013_, new_n10014_, new_n10015_,
    new_n10016_, new_n10017_, new_n10018_, new_n10019_, new_n10020_,
    new_n10021_, new_n10022_, new_n10023_, new_n10024_, new_n10025_,
    new_n10026_, new_n10027_, new_n10028_, new_n10029_, new_n10030_,
    new_n10031_, new_n10032_, new_n10033_, new_n10034_, new_n10035_,
    new_n10036_, new_n10037_, new_n10038_, new_n10039_, new_n10040_,
    new_n10041_, new_n10042_, new_n10043_, new_n10044_, new_n10045_,
    new_n10046_, new_n10047_, new_n10048_, new_n10049_, new_n10050_,
    new_n10051_, new_n10052_, new_n10053_, new_n10054_, new_n10055_,
    new_n10056_, new_n10057_, new_n10058_, new_n10059_, new_n10060_,
    new_n10061_, new_n10062_, new_n10063_, new_n10064_, new_n10065_,
    new_n10066_, new_n10067_, new_n10068_, new_n10069_, new_n10070_,
    new_n10071_, new_n10072_, new_n10073_, new_n10074_, new_n10075_,
    new_n10076_, new_n10077_, new_n10078_, new_n10079_, new_n10080_,
    new_n10081_, new_n10082_, new_n10083_, new_n10084_, new_n10085_,
    new_n10086_, new_n10087_, new_n10088_, new_n10089_, new_n10090_,
    new_n10091_, new_n10092_, new_n10093_, new_n10094_, new_n10095_,
    new_n10096_, new_n10097_, new_n10098_, new_n10099_, new_n10100_,
    new_n10101_, new_n10102_, new_n10103_, new_n10104_, new_n10105_,
    new_n10106_, new_n10107_, new_n10108_, new_n10109_, new_n10110_,
    new_n10111_, new_n10112_, new_n10113_, new_n10114_, new_n10115_,
    new_n10116_, new_n10117_, new_n10118_, new_n10119_, new_n10120_,
    new_n10121_, new_n10122_, new_n10123_, new_n10124_, new_n10125_,
    new_n10126_, new_n10127_, new_n10128_, new_n10129_, new_n10130_,
    new_n10131_, new_n10132_, new_n10133_, new_n10134_, new_n10135_,
    new_n10136_, new_n10137_, new_n10138_, new_n10139_, new_n10140_,
    new_n10141_, new_n10142_, new_n10143_, new_n10144_, new_n10145_,
    new_n10146_, new_n10147_, new_n10148_, new_n10149_, new_n10150_,
    new_n10151_, new_n10152_, new_n10153_, new_n10154_, new_n10155_,
    new_n10156_, new_n10157_, new_n10158_, new_n10159_, new_n10160_,
    new_n10161_, new_n10162_, new_n10163_, new_n10164_, new_n10165_,
    new_n10166_, new_n10167_, new_n10168_, new_n10169_, new_n10170_,
    new_n10171_, new_n10172_, new_n10173_, new_n10174_, new_n10175_,
    new_n10176_, new_n10177_, new_n10178_, new_n10179_, new_n10180_,
    new_n10181_, new_n10182_, new_n10183_, new_n10184_, new_n10185_,
    new_n10186_, new_n10187_, new_n10188_, new_n10189_, new_n10190_,
    new_n10191_, new_n10192_, new_n10193_, new_n10194_, new_n10195_,
    new_n10196_, new_n10197_, new_n10198_, new_n10199_, new_n10200_,
    new_n10201_, new_n10202_, new_n10203_, new_n10204_, new_n10205_,
    new_n10206_, new_n10207_, new_n10208_, new_n10209_, new_n10210_,
    new_n10211_, new_n10212_, new_n10213_, new_n10214_, new_n10215_,
    new_n10216_, new_n10217_, new_n10218_, new_n10219_, new_n10220_,
    new_n10221_, new_n10222_, new_n10223_, new_n10224_, new_n10225_,
    new_n10226_, new_n10227_, new_n10228_, new_n10229_, new_n10230_,
    new_n10231_, new_n10232_, new_n10233_, new_n10234_, new_n10235_,
    new_n10236_, new_n10237_, new_n10238_, new_n10239_, new_n10240_,
    new_n10241_, new_n10242_, new_n10243_, new_n10244_, new_n10245_,
    new_n10246_, new_n10247_, new_n10248_, new_n10249_, new_n10250_,
    new_n10251_, new_n10252_, new_n10253_, new_n10254_, new_n10255_,
    new_n10256_, new_n10257_, new_n10258_, new_n10259_, new_n10260_,
    new_n10261_, new_n10262_, new_n10263_, new_n10264_, new_n10265_,
    new_n10266_, new_n10267_, new_n10268_, new_n10269_, new_n10270_,
    new_n10271_, new_n10272_, new_n10273_, new_n10274_, new_n10275_,
    new_n10276_, new_n10277_, new_n10278_, new_n10279_, new_n10280_,
    new_n10281_, new_n10282_, new_n10283_, new_n10284_, new_n10285_,
    new_n10286_, new_n10287_, new_n10288_, new_n10289_, new_n10290_,
    new_n10291_, new_n10292_, new_n10293_, new_n10294_, new_n10295_,
    new_n10296_, new_n10297_, new_n10298_, new_n10299_, new_n10300_,
    new_n10301_, new_n10302_, new_n10303_, new_n10304_, new_n10305_,
    new_n10306_, new_n10307_, new_n10308_, new_n10309_, new_n10310_,
    new_n10311_, new_n10312_, new_n10313_, new_n10314_, new_n10315_,
    new_n10316_, new_n10317_, new_n10318_, new_n10319_, new_n10320_,
    new_n10321_, new_n10322_, new_n10323_, new_n10324_, new_n10325_,
    new_n10326_, new_n10327_, new_n10328_, new_n10329_, new_n10330_,
    new_n10331_, new_n10332_, new_n10333_, new_n10334_, new_n10335_,
    new_n10336_, new_n10337_, new_n10338_, new_n10339_, new_n10340_,
    new_n10341_, new_n10342_, new_n10343_, new_n10344_, new_n10345_,
    new_n10346_, new_n10347_, new_n10348_, new_n10349_, new_n10350_,
    new_n10351_, new_n10352_, new_n10353_, new_n10354_, new_n10355_,
    new_n10356_, new_n10357_, new_n10358_, new_n10359_, new_n10360_,
    new_n10361_, new_n10362_, new_n10363_, new_n10364_, new_n10365_,
    new_n10366_, new_n10367_, new_n10368_, new_n10369_, new_n10370_,
    new_n10371_, new_n10372_, new_n10373_, new_n10374_, new_n10375_,
    new_n10376_, new_n10377_, new_n10378_, new_n10379_, new_n10380_,
    new_n10381_, new_n10382_, new_n10383_, new_n10384_, new_n10385_,
    new_n10386_, new_n10387_, new_n10388_, new_n10389_, new_n10390_,
    new_n10391_, new_n10392_, new_n10393_, new_n10394_, new_n10395_,
    new_n10396_, new_n10397_, new_n10398_, new_n10399_, new_n10400_,
    new_n10401_, new_n10402_, new_n10403_, new_n10404_, new_n10405_,
    new_n10406_, new_n10407_, new_n10408_, new_n10409_, new_n10410_,
    new_n10411_, new_n10412_, new_n10413_, new_n10414_, new_n10415_,
    new_n10416_, new_n10417_, new_n10418_, new_n10419_, new_n10420_,
    new_n10421_, new_n10422_, new_n10423_, new_n10424_, new_n10425_,
    new_n10426_, new_n10427_, new_n10428_, new_n10429_, new_n10430_,
    new_n10431_, new_n10432_, new_n10433_, new_n10434_, new_n10435_,
    new_n10436_, new_n10437_, new_n10438_, new_n10439_, new_n10440_,
    new_n10441_, new_n10442_, new_n10443_, new_n10444_, new_n10445_,
    new_n10446_, new_n10447_, new_n10448_, new_n10449_, new_n10450_,
    new_n10451_, new_n10452_, new_n10453_, new_n10454_, new_n10455_,
    new_n10456_, new_n10457_, new_n10458_, new_n10459_, new_n10460_,
    new_n10461_, new_n10462_, new_n10463_, new_n10464_, new_n10465_,
    new_n10466_, new_n10467_, new_n10468_, new_n10469_, new_n10470_,
    new_n10471_, new_n10472_, new_n10473_, new_n10474_, new_n10475_,
    new_n10476_, new_n10477_, new_n10478_, new_n10479_, new_n10480_,
    new_n10481_, new_n10482_, new_n10483_, new_n10484_, new_n10485_,
    new_n10486_, new_n10487_, new_n10488_, new_n10489_, new_n10490_,
    new_n10491_, new_n10492_, new_n10493_, new_n10494_, new_n10495_,
    new_n10496_, new_n10497_, new_n10498_, new_n10499_, new_n10500_,
    new_n10501_, new_n10502_, new_n10503_, new_n10504_, new_n10505_,
    new_n10506_, new_n10507_, new_n10508_, new_n10509_, new_n10510_,
    new_n10511_, new_n10512_, new_n10513_, new_n10514_, new_n10515_,
    new_n10516_, new_n10517_, new_n10518_, new_n10519_, new_n10520_,
    new_n10521_, new_n10522_, new_n10523_, new_n10524_, new_n10525_,
    new_n10526_, new_n10527_, new_n10528_, new_n10529_, new_n10530_,
    new_n10531_, new_n10532_, new_n10533_, new_n10534_, new_n10535_,
    new_n10536_, new_n10537_, new_n10538_, new_n10539_, new_n10540_,
    new_n10541_, new_n10542_, new_n10543_, new_n10544_, new_n10545_,
    new_n10546_, new_n10547_, new_n10548_, new_n10549_, new_n10550_,
    new_n10551_, new_n10552_, new_n10553_, new_n10554_, new_n10555_,
    new_n10556_, new_n10557_, new_n10558_, new_n10559_, new_n10560_,
    new_n10561_, new_n10562_, new_n10563_, new_n10564_, new_n10565_,
    new_n10566_, new_n10567_, new_n10568_, new_n10569_, new_n10570_,
    new_n10571_, new_n10572_, new_n10573_, new_n10574_, new_n10575_,
    new_n10576_, new_n10577_, new_n10578_, new_n10579_, new_n10580_,
    new_n10581_, new_n10582_, new_n10583_, new_n10584_, new_n10585_,
    new_n10586_, new_n10587_, new_n10588_, new_n10589_, new_n10590_,
    new_n10591_, new_n10592_, new_n10593_, new_n10594_, new_n10595_,
    new_n10596_, new_n10597_, new_n10598_, new_n10599_, new_n10600_,
    new_n10601_, new_n10602_, new_n10603_, new_n10604_, new_n10605_,
    new_n10606_, new_n10607_, new_n10608_, new_n10609_, new_n10610_,
    new_n10611_, new_n10612_, new_n10613_, new_n10614_, new_n10615_,
    new_n10616_, new_n10617_, new_n10618_, new_n10619_, new_n10620_,
    new_n10621_, new_n10622_, new_n10623_, new_n10624_, new_n10625_,
    new_n10626_, new_n10627_, new_n10628_, new_n10629_, new_n10630_,
    new_n10631_, new_n10632_, new_n10633_, new_n10634_, new_n10635_,
    new_n10636_, new_n10637_, new_n10638_, new_n10639_, new_n10640_,
    new_n10641_, new_n10642_, new_n10643_, new_n10644_, new_n10645_,
    new_n10646_, new_n10647_, new_n10648_, new_n10649_, new_n10650_,
    new_n10651_, new_n10652_, new_n10653_, new_n10654_, new_n10655_,
    new_n10656_, new_n10657_, new_n10658_, new_n10659_, new_n10660_,
    new_n10661_, new_n10662_, new_n10663_, new_n10664_, new_n10665_,
    new_n10666_, new_n10667_, new_n10668_, new_n10669_, new_n10670_,
    new_n10671_, new_n10672_, new_n10673_, new_n10674_, new_n10675_,
    new_n10676_, new_n10677_, new_n10678_, new_n10679_, new_n10680_,
    new_n10681_, new_n10682_, new_n10683_, new_n10684_, new_n10685_,
    new_n10686_, new_n10687_, new_n10688_, new_n10689_, new_n10690_,
    new_n10691_, new_n10692_, new_n10693_, new_n10694_, new_n10695_,
    new_n10696_, new_n10697_, new_n10698_, new_n10699_, new_n10700_,
    new_n10701_, new_n10702_, new_n10703_, new_n10704_, new_n10705_,
    new_n10706_, new_n10707_, new_n10708_, new_n10709_, new_n10710_,
    new_n10711_, new_n10712_, new_n10713_, new_n10714_, new_n10715_,
    new_n10716_, new_n10717_, new_n10718_, new_n10719_, new_n10720_,
    new_n10721_, new_n10722_, new_n10723_, new_n10724_, new_n10725_,
    new_n10726_, new_n10727_, new_n10728_, new_n10729_, new_n10730_,
    new_n10731_, new_n10732_, new_n10733_, new_n10734_, new_n10735_,
    new_n10736_, new_n10737_, new_n10738_, new_n10739_, new_n10740_,
    new_n10741_, new_n10742_, new_n10743_, new_n10744_, new_n10745_,
    new_n10746_, new_n10747_, new_n10748_, new_n10749_, new_n10750_,
    new_n10751_, new_n10752_, new_n10753_, new_n10754_, new_n10755_,
    new_n10756_, new_n10757_, new_n10758_, new_n10759_, new_n10760_,
    new_n10761_, new_n10762_, new_n10763_, new_n10764_, new_n10765_,
    new_n10766_, new_n10767_, new_n10768_, new_n10769_, new_n10770_,
    new_n10771_, new_n10772_, new_n10773_, new_n10774_, new_n10775_,
    new_n10776_, new_n10777_, new_n10778_, new_n10779_, new_n10780_,
    new_n10781_, new_n10782_, new_n10783_, new_n10784_, new_n10785_,
    new_n10786_, new_n10787_, new_n10788_, new_n10789_, new_n10790_,
    new_n10791_, new_n10792_, new_n10793_, new_n10794_, new_n10795_,
    new_n10796_, new_n10797_, new_n10798_, new_n10799_, new_n10800_,
    new_n10801_, new_n10802_, new_n10803_, new_n10804_, new_n10805_,
    new_n10806_, new_n10807_, new_n10808_, new_n10809_, new_n10810_,
    new_n10811_, new_n10812_, new_n10813_, new_n10814_, new_n10815_,
    new_n10816_, new_n10817_, new_n10818_, new_n10819_, new_n10820_,
    new_n10821_, new_n10822_, new_n10823_, new_n10824_, new_n10825_,
    new_n10826_, new_n10827_, new_n10828_, new_n10829_, new_n10830_,
    new_n10831_, new_n10832_, new_n10833_, new_n10834_, new_n10835_,
    new_n10836_, new_n10837_, new_n10838_, new_n10839_, new_n10840_,
    new_n10841_, new_n10842_, new_n10843_, new_n10844_, new_n10845_,
    new_n10846_, new_n10847_, new_n10848_, new_n10849_, new_n10850_,
    new_n10851_, new_n10852_, new_n10853_, new_n10854_, new_n10855_,
    new_n10856_, new_n10857_, new_n10858_, new_n10859_, new_n10860_,
    new_n10861_, new_n10862_, new_n10863_, new_n10864_, new_n10865_,
    new_n10866_, new_n10867_, new_n10868_, new_n10869_, new_n10870_,
    new_n10871_, new_n10872_, new_n10873_, new_n10874_, new_n10875_,
    new_n10876_, new_n10877_, new_n10878_, new_n10879_, new_n10880_,
    new_n10881_, new_n10882_, new_n10883_, new_n10884_, new_n10885_,
    new_n10886_, new_n10887_, new_n10888_, new_n10889_, new_n10890_,
    new_n10891_, new_n10892_, new_n10893_, new_n10894_, new_n10895_,
    new_n10896_, new_n10897_, new_n10898_, new_n10899_, new_n10900_,
    new_n10901_, new_n10902_, new_n10903_, new_n10904_, new_n10905_,
    new_n10906_, new_n10907_, new_n10908_, new_n10909_, new_n10910_,
    new_n10911_, new_n10912_, new_n10913_, new_n10914_, new_n10915_,
    new_n10916_, new_n10917_, new_n10918_, new_n10919_, new_n10920_,
    new_n10921_, new_n10922_, new_n10923_, new_n10924_, new_n10925_,
    new_n10926_, new_n10927_, new_n10928_, new_n10929_, new_n10930_,
    new_n10931_, new_n10932_, new_n10933_, new_n10934_, new_n10935_,
    new_n10936_, new_n10937_, new_n10938_, new_n10939_, new_n10940_,
    new_n10941_, new_n10942_, new_n10943_, new_n10944_, new_n10945_,
    new_n10946_, new_n10947_, new_n10948_, new_n10949_, new_n10950_,
    new_n10951_, new_n10952_, new_n10953_, new_n10954_, new_n10955_,
    new_n10956_, new_n10957_, new_n10958_, new_n10959_, new_n10960_,
    new_n10961_, new_n10962_, new_n10963_, new_n10964_, new_n10965_,
    new_n10966_, new_n10967_, new_n10968_, new_n10969_, new_n10970_,
    new_n10971_, new_n10972_, new_n10973_, new_n10974_, new_n10975_,
    new_n10976_, new_n10977_, new_n10978_, new_n10979_, new_n10980_,
    new_n10981_, new_n10982_, new_n10983_, new_n10984_, new_n10985_,
    new_n10986_, new_n10987_, new_n10988_, new_n10989_, new_n10990_,
    new_n10991_, new_n10992_, new_n10993_, new_n10994_, new_n10995_,
    new_n10996_, new_n10997_, new_n10998_, new_n10999_, new_n11000_,
    new_n11001_, new_n11002_, new_n11003_, new_n11004_, new_n11005_,
    new_n11006_, new_n11007_, new_n11008_, new_n11009_, new_n11010_,
    new_n11011_, new_n11012_, new_n11013_, new_n11014_, new_n11015_,
    new_n11016_, new_n11017_, new_n11018_, new_n11019_, new_n11020_,
    new_n11021_, new_n11022_, new_n11023_, new_n11024_, new_n11025_,
    new_n11026_, new_n11027_, new_n11028_, new_n11029_, new_n11030_,
    new_n11031_, new_n11032_, new_n11033_, new_n11034_, new_n11035_,
    new_n11036_, new_n11037_, new_n11038_, new_n11039_, new_n11040_,
    new_n11041_, new_n11042_, new_n11043_, new_n11044_, new_n11045_,
    new_n11046_, new_n11047_, new_n11048_, new_n11049_, new_n11050_,
    new_n11051_, new_n11052_, new_n11053_, new_n11054_, new_n11055_,
    new_n11056_, new_n11057_, new_n11058_, new_n11059_, new_n11060_,
    new_n11061_, new_n11062_, new_n11063_, new_n11064_, new_n11065_,
    new_n11066_, new_n11067_, new_n11068_, new_n11069_, new_n11070_,
    new_n11071_, new_n11072_, new_n11073_, new_n11074_, new_n11075_,
    new_n11076_, new_n11077_, new_n11078_, new_n11079_, new_n11080_,
    new_n11081_, new_n11082_, new_n11083_, new_n11084_, new_n11085_,
    new_n11086_, new_n11087_, new_n11088_, new_n11089_, new_n11090_,
    new_n11091_, new_n11092_, new_n11093_, new_n11094_, new_n11095_,
    new_n11096_, new_n11097_, new_n11098_, new_n11099_, new_n11100_,
    new_n11101_, new_n11102_, new_n11103_, new_n11104_, new_n11105_,
    new_n11106_, new_n11107_, new_n11108_, new_n11109_, new_n11110_,
    new_n11111_, new_n11112_, new_n11113_, new_n11114_, new_n11115_,
    new_n11116_, new_n11117_, new_n11118_, new_n11119_, new_n11120_,
    new_n11121_, new_n11122_, new_n11123_, new_n11124_, new_n11125_,
    new_n11126_, new_n11127_, new_n11128_, new_n11129_, new_n11130_,
    new_n11131_, new_n11132_, new_n11133_, new_n11134_, new_n11135_,
    new_n11136_, new_n11137_, new_n11138_, new_n11139_, new_n11140_,
    new_n11141_, new_n11142_, new_n11143_, new_n11144_, new_n11145_,
    new_n11146_, new_n11147_, new_n11148_, new_n11149_, new_n11150_,
    new_n11151_, new_n11152_, new_n11153_, new_n11154_, new_n11155_,
    new_n11156_, new_n11157_, new_n11158_, new_n11159_, new_n11160_,
    new_n11161_, new_n11162_, new_n11163_, new_n11164_, new_n11165_,
    new_n11166_, new_n11167_, new_n11168_, new_n11169_, new_n11170_,
    new_n11171_, new_n11172_, new_n11173_, new_n11174_, new_n11175_,
    new_n11176_, new_n11177_, new_n11178_, new_n11179_, new_n11180_,
    new_n11181_, new_n11182_, new_n11183_, new_n11184_, new_n11185_,
    new_n11186_, new_n11187_, new_n11188_, new_n11189_, new_n11190_,
    new_n11191_, new_n11192_, new_n11193_, new_n11194_, new_n11195_,
    new_n11196_, new_n11197_, new_n11198_, new_n11199_, new_n11200_,
    new_n11201_, new_n11202_, new_n11203_, new_n11204_, new_n11205_,
    new_n11206_, new_n11207_, new_n11208_, new_n11209_, new_n11210_,
    new_n11211_, new_n11212_, new_n11213_, new_n11214_, new_n11215_,
    new_n11216_, new_n11217_, new_n11218_, new_n11219_, new_n11220_,
    new_n11221_, new_n11222_, new_n11223_, new_n11224_, new_n11225_,
    new_n11226_, new_n11227_, new_n11228_, new_n11229_, new_n11230_,
    new_n11231_, new_n11232_, new_n11233_, new_n11234_, new_n11235_,
    new_n11236_, new_n11237_, new_n11238_, new_n11239_, new_n11240_,
    new_n11241_, new_n11242_, new_n11243_, new_n11244_, new_n11245_,
    new_n11246_, new_n11247_, new_n11248_, new_n11249_, new_n11250_,
    new_n11251_, new_n11252_, new_n11253_, new_n11254_, new_n11255_,
    new_n11256_, new_n11257_, new_n11258_, new_n11259_, new_n11260_,
    new_n11261_, new_n11262_, new_n11263_, new_n11264_, new_n11265_,
    new_n11266_, new_n11267_, new_n11268_, new_n11269_, new_n11270_,
    new_n11271_, new_n11272_, new_n11273_, new_n11274_, new_n11275_,
    new_n11276_, new_n11277_, new_n11278_, new_n11279_, new_n11280_,
    new_n11281_, new_n11282_, new_n11283_, new_n11284_, new_n11285_,
    new_n11286_, new_n11287_, new_n11288_, new_n11289_, new_n11290_,
    new_n11291_, new_n11292_, new_n11293_, new_n11294_, new_n11295_,
    new_n11296_, new_n11297_, new_n11298_, new_n11299_, new_n11300_,
    new_n11301_, new_n11302_, new_n11303_, new_n11304_, new_n11305_,
    new_n11306_, new_n11307_, new_n11308_, new_n11309_, new_n11310_,
    new_n11311_, new_n11312_, new_n11313_, new_n11314_, new_n11315_,
    new_n11316_, new_n11317_, new_n11318_, new_n11319_, new_n11320_,
    new_n11321_, new_n11322_, new_n11323_, new_n11324_, new_n11325_,
    new_n11326_, new_n11327_, new_n11328_, new_n11329_, new_n11330_,
    new_n11331_, new_n11332_, new_n11333_, new_n11334_, new_n11335_,
    new_n11336_, new_n11337_, new_n11338_, new_n11339_, new_n11340_,
    new_n11341_, new_n11342_, new_n11343_, new_n11344_, new_n11345_,
    new_n11346_, new_n11347_, new_n11348_, new_n11349_, new_n11350_,
    new_n11351_, new_n11352_, new_n11353_, new_n11354_, new_n11355_,
    new_n11356_, new_n11357_, new_n11358_, new_n11359_, new_n11360_,
    new_n11361_, new_n11362_, new_n11363_, new_n11364_, new_n11365_,
    new_n11366_, new_n11367_, new_n11368_, new_n11369_, new_n11370_,
    new_n11371_, new_n11372_, new_n11373_, new_n11374_, new_n11375_,
    new_n11376_, new_n11377_, new_n11378_, new_n11379_, new_n11380_,
    new_n11381_, new_n11382_, new_n11383_, new_n11384_, new_n11385_,
    new_n11386_, new_n11387_, new_n11388_, new_n11389_, new_n11390_,
    new_n11391_, new_n11392_, new_n11393_, new_n11394_, new_n11395_,
    new_n11396_, new_n11397_, new_n11398_, new_n11399_, new_n11400_,
    new_n11401_, new_n11402_, new_n11403_, new_n11404_, new_n11405_,
    new_n11406_, new_n11407_, new_n11408_, new_n11409_, new_n11410_,
    new_n11411_, new_n11412_, new_n11413_, new_n11414_, new_n11415_,
    new_n11416_, new_n11417_, new_n11418_, new_n11419_, new_n11420_,
    new_n11421_, new_n11422_, new_n11423_, new_n11424_, new_n11425_,
    new_n11426_, new_n11427_, new_n11428_, new_n11429_, new_n11430_,
    new_n11431_, new_n11432_, new_n11433_, new_n11434_, new_n11435_,
    new_n11436_, new_n11437_, new_n11438_, new_n11439_, new_n11440_,
    new_n11441_, new_n11442_, new_n11443_, new_n11444_, new_n11445_,
    new_n11446_, new_n11447_, new_n11448_, new_n11449_, new_n11450_,
    new_n11451_, new_n11452_, new_n11453_, new_n11454_, new_n11455_,
    new_n11456_, new_n11457_, new_n11458_, new_n11459_, new_n11460_,
    new_n11461_, new_n11462_, new_n11463_, new_n11464_, new_n11465_,
    new_n11466_, new_n11467_, new_n11468_, new_n11469_, new_n11470_,
    new_n11471_, new_n11472_, new_n11473_, new_n11474_, new_n11475_,
    new_n11476_, new_n11477_, new_n11478_, new_n11479_, new_n11480_,
    new_n11481_, new_n11482_, new_n11483_, new_n11484_, new_n11485_,
    new_n11486_, new_n11487_, new_n11488_, new_n11489_, new_n11490_,
    new_n11491_, new_n11492_, new_n11493_, new_n11494_, new_n11495_,
    new_n11496_, new_n11497_, new_n11498_, new_n11499_, new_n11500_,
    new_n11501_, new_n11502_, new_n11503_, new_n11504_, new_n11505_,
    new_n11506_, new_n11507_, new_n11508_, new_n11509_, new_n11510_,
    new_n11511_, new_n11512_, new_n11513_, new_n11514_, new_n11515_,
    new_n11516_, new_n11517_, new_n11518_, new_n11519_, new_n11520_,
    new_n11521_, new_n11522_, new_n11523_, new_n11524_, new_n11525_,
    new_n11526_, new_n11527_, new_n11528_, new_n11529_, new_n11530_,
    new_n11531_, new_n11532_, new_n11533_, new_n11534_, new_n11535_,
    new_n11536_, new_n11537_, new_n11538_, new_n11539_, new_n11540_,
    new_n11541_, new_n11542_, new_n11543_, new_n11544_, new_n11545_,
    new_n11546_, new_n11547_, new_n11548_, new_n11549_, new_n11550_,
    new_n11551_, new_n11552_, new_n11553_, new_n11554_, new_n11555_,
    new_n11556_, new_n11557_, new_n11558_, new_n11559_, new_n11560_,
    new_n11561_, new_n11562_, new_n11563_, new_n11564_, new_n11565_,
    new_n11566_, new_n11567_, new_n11568_, new_n11569_, new_n11570_,
    new_n11571_, new_n11572_, new_n11573_, new_n11574_, new_n11575_,
    new_n11576_, new_n11577_, new_n11578_, new_n11579_, new_n11580_,
    new_n11581_, new_n11582_, new_n11583_, new_n11584_, new_n11585_,
    new_n11586_, new_n11587_, new_n11588_, new_n11589_, new_n11590_,
    new_n11591_, new_n11592_, new_n11593_, new_n11594_, new_n11595_,
    new_n11596_, new_n11597_, new_n11598_, new_n11599_, new_n11600_,
    new_n11601_, new_n11602_, new_n11603_, new_n11604_, new_n11605_,
    new_n11606_, new_n11607_, new_n11608_, new_n11609_, new_n11610_,
    new_n11611_, new_n11612_, new_n11613_, new_n11614_, new_n11615_,
    new_n11616_, new_n11617_, new_n11618_, new_n11619_, new_n11620_,
    new_n11621_, new_n11622_, new_n11623_, new_n11624_, new_n11625_,
    new_n11626_, new_n11627_, new_n11628_, new_n11629_, new_n11630_,
    new_n11631_, new_n11632_, new_n11633_, new_n11634_, new_n11635_,
    new_n11636_, new_n11637_, new_n11638_, new_n11639_, new_n11640_,
    new_n11641_, new_n11642_, new_n11643_, new_n11644_, new_n11645_,
    new_n11646_, new_n11647_, new_n11648_, new_n11649_, new_n11650_,
    new_n11651_, new_n11652_, new_n11653_, new_n11654_, new_n11655_,
    new_n11656_, new_n11657_, new_n11658_, new_n11659_, new_n11660_,
    new_n11661_, new_n11662_, new_n11663_, new_n11664_, new_n11665_,
    new_n11666_, new_n11667_, new_n11668_, new_n11669_, new_n11670_,
    new_n11671_, new_n11672_, new_n11673_, new_n11674_, new_n11675_,
    new_n11676_, new_n11677_, new_n11678_, new_n11679_, new_n11680_,
    new_n11681_, new_n11682_, new_n11683_, new_n11684_, new_n11685_,
    new_n11686_, new_n11687_, new_n11688_, new_n11689_, new_n11690_,
    new_n11691_, new_n11692_, new_n11693_, new_n11694_, new_n11695_,
    new_n11696_, new_n11697_, new_n11698_, new_n11699_, new_n11700_,
    new_n11701_, new_n11702_, new_n11703_, new_n11704_, new_n11705_,
    new_n11706_, new_n11707_, new_n11708_, new_n11709_, new_n11710_,
    new_n11711_, new_n11712_, new_n11713_, new_n11714_, new_n11715_,
    new_n11716_, new_n11717_, new_n11718_, new_n11719_, new_n11720_,
    new_n11721_, new_n11722_, new_n11723_, new_n11724_, new_n11725_,
    new_n11726_, new_n11727_, new_n11728_, new_n11729_, new_n11730_,
    new_n11731_, new_n11732_, new_n11733_, new_n11734_, new_n11735_,
    new_n11736_, new_n11737_, new_n11738_, new_n11739_, new_n11740_,
    new_n11741_, new_n11742_, new_n11743_, new_n11744_, new_n11745_,
    new_n11746_, new_n11747_, new_n11748_, new_n11749_, new_n11750_,
    new_n11751_, new_n11752_, new_n11753_, new_n11754_, new_n11755_,
    new_n11756_, new_n11757_, new_n11758_, new_n11759_, new_n11760_,
    new_n11761_, new_n11762_, new_n11763_, new_n11764_, new_n11765_,
    new_n11766_, new_n11767_, new_n11768_, new_n11769_, new_n11770_,
    new_n11771_, new_n11772_, new_n11773_, new_n11774_, new_n11775_,
    new_n11776_, new_n11777_, new_n11778_, new_n11779_, new_n11780_,
    new_n11781_, new_n11782_, new_n11783_, new_n11784_, new_n11785_,
    new_n11786_, new_n11787_, new_n11788_, new_n11789_, new_n11790_,
    new_n11791_, new_n11792_, new_n11793_, new_n11794_, new_n11795_,
    new_n11796_, new_n11797_, new_n11798_, new_n11799_, new_n11800_,
    new_n11801_, new_n11802_, new_n11803_, new_n11804_, new_n11805_,
    new_n11806_, new_n11807_, new_n11808_, new_n11809_, new_n11810_,
    new_n11811_, new_n11812_, new_n11813_, new_n11814_, new_n11815_,
    new_n11816_, new_n11817_, new_n11818_, new_n11819_, new_n11820_,
    new_n11821_, new_n11822_, new_n11823_, new_n11824_, new_n11825_,
    new_n11826_, new_n11827_, new_n11828_, new_n11829_, new_n11830_,
    new_n11831_, new_n11832_, new_n11833_, new_n11834_, new_n11835_,
    new_n11836_, new_n11837_, new_n11838_, new_n11839_, new_n11840_,
    new_n11841_, new_n11842_, new_n11843_, new_n11844_, new_n11845_,
    new_n11846_, new_n11847_, new_n11848_, new_n11849_, new_n11850_,
    new_n11851_, new_n11852_, new_n11853_, new_n11854_, new_n11855_,
    new_n11856_, new_n11857_, new_n11858_, new_n11859_, new_n11860_,
    new_n11861_, new_n11862_, new_n11863_, new_n11864_, new_n11865_,
    new_n11866_, new_n11867_, new_n11868_, new_n11869_, new_n11870_,
    new_n11871_, new_n11872_, new_n11873_, new_n11874_, new_n11875_,
    new_n11876_, new_n11877_, new_n11878_, new_n11879_, new_n11880_,
    new_n11881_, new_n11882_, new_n11883_, new_n11884_, new_n11885_,
    new_n11886_, new_n11887_, new_n11888_, new_n11889_, new_n11890_,
    new_n11891_, new_n11892_, new_n11893_, new_n11894_, new_n11895_,
    new_n11896_, new_n11897_, new_n11898_, new_n11899_, new_n11900_,
    new_n11901_, new_n11902_, new_n11903_, new_n11904_, new_n11905_,
    new_n11906_, new_n11907_, new_n11908_, new_n11909_, new_n11910_,
    new_n11911_, new_n11912_, new_n11913_, new_n11914_, new_n11915_,
    new_n11916_, new_n11917_, new_n11918_, new_n11919_, new_n11920_,
    new_n11921_, new_n11922_, new_n11923_, new_n11924_, new_n11925_,
    new_n11926_, new_n11927_, new_n11928_, new_n11929_, new_n11930_,
    new_n11931_, new_n11932_, new_n11933_, new_n11934_, new_n11935_,
    new_n11936_, new_n11937_, new_n11938_, new_n11939_, new_n11940_,
    new_n11941_, new_n11942_, new_n11943_, new_n11944_, new_n11945_,
    new_n11946_, new_n11947_, new_n11948_, new_n11949_, new_n11950_,
    new_n11951_, new_n11952_, new_n11953_, new_n11954_, new_n11955_,
    new_n11956_, new_n11957_, new_n11958_, new_n11959_, new_n11960_,
    new_n11961_, new_n11962_, new_n11963_, new_n11964_, new_n11965_,
    new_n11966_, new_n11967_, new_n11968_, new_n11969_, new_n11970_,
    new_n11971_, new_n11972_, new_n11973_, new_n11974_, new_n11975_,
    new_n11976_, new_n11977_, new_n11978_, new_n11979_, new_n11980_,
    new_n11981_, new_n11982_, new_n11983_, new_n11984_, new_n11985_,
    new_n11986_, new_n11987_, new_n11988_, new_n11989_, new_n11990_,
    new_n11991_, new_n11992_, new_n11993_, new_n11994_, new_n11995_,
    new_n11996_, new_n11997_, new_n11998_, new_n11999_, new_n12000_,
    new_n12001_, new_n12002_, new_n12003_, new_n12004_, new_n12005_,
    new_n12006_, new_n12007_, new_n12008_, new_n12009_, new_n12010_,
    new_n12011_, new_n12012_, new_n12013_, new_n12014_, new_n12015_,
    new_n12016_, new_n12017_, new_n12018_, new_n12019_, new_n12020_,
    new_n12021_, new_n12022_, new_n12023_, new_n12024_, new_n12025_,
    new_n12026_, new_n12027_, new_n12028_, new_n12029_, new_n12030_,
    new_n12031_, new_n12032_, new_n12033_, new_n12034_, new_n12035_,
    new_n12036_, new_n12037_, new_n12038_, new_n12039_, new_n12040_,
    new_n12041_, new_n12042_, new_n12043_, new_n12044_, new_n12045_,
    new_n12046_, new_n12047_, new_n12048_, new_n12049_, new_n12050_,
    new_n12051_, new_n12052_, new_n12053_, new_n12054_, new_n12055_,
    new_n12056_, new_n12057_, new_n12058_, new_n12059_, new_n12060_,
    new_n12061_, new_n12062_, new_n12063_, new_n12064_, new_n12065_,
    new_n12066_, new_n12067_, new_n12068_, new_n12069_, new_n12070_,
    new_n12071_, new_n12072_, new_n12073_, new_n12074_, new_n12075_,
    new_n12076_, new_n12077_, new_n12078_, new_n12079_, new_n12080_,
    new_n12081_, new_n12082_, new_n12083_, new_n12084_, new_n12085_,
    new_n12086_, new_n12087_, new_n12088_, new_n12089_, new_n12090_,
    new_n12091_, new_n12092_, new_n12093_, new_n12094_, new_n12095_,
    new_n12096_, new_n12097_, new_n12098_, new_n12099_, new_n12100_,
    new_n12101_, new_n12102_, new_n12103_, new_n12104_, new_n12105_,
    new_n12106_, new_n12107_, new_n12108_, new_n12109_, new_n12110_,
    new_n12111_, new_n12112_, new_n12113_, new_n12114_, new_n12115_,
    new_n12116_, new_n12117_, new_n12118_, new_n12119_, new_n12120_,
    new_n12121_, new_n12122_, new_n12123_, new_n12124_, new_n12125_,
    new_n12126_, new_n12127_, new_n12128_, new_n12129_, new_n12130_,
    new_n12131_, new_n12132_, new_n12133_, new_n12134_, new_n12135_,
    new_n12136_, new_n12137_, new_n12138_, new_n12139_, new_n12140_,
    new_n12141_, new_n12142_, new_n12143_, new_n12144_, new_n12145_,
    new_n12146_, new_n12147_, new_n12148_, new_n12149_, new_n12150_,
    new_n12151_, new_n12152_, new_n12153_, new_n12154_, new_n12155_,
    new_n12156_, new_n12157_, new_n12158_, new_n12159_, new_n12160_,
    new_n12161_, new_n12162_, new_n12163_, new_n12164_, new_n12165_,
    new_n12166_, new_n12167_, new_n12168_, new_n12169_, new_n12170_,
    new_n12171_, new_n12172_, new_n12173_, new_n12174_, new_n12175_,
    new_n12176_, new_n12177_, new_n12178_, new_n12179_, new_n12180_,
    new_n12181_, new_n12182_, new_n12183_, new_n12184_, new_n12185_,
    new_n12186_, new_n12187_, new_n12188_, new_n12189_, new_n12190_,
    new_n12191_, new_n12192_, new_n12193_, new_n12194_, new_n12195_,
    new_n12196_, new_n12197_, new_n12198_, new_n12199_, new_n12200_,
    new_n12201_, new_n12202_, new_n12203_, new_n12204_, new_n12205_,
    new_n12206_, new_n12207_, new_n12208_, new_n12209_, new_n12210_,
    new_n12211_, new_n12212_, new_n12213_, new_n12214_, new_n12215_,
    new_n12216_, new_n12217_, new_n12218_, new_n12219_, new_n12220_,
    new_n12221_, new_n12222_, new_n12223_, new_n12224_, new_n12225_,
    new_n12226_, new_n12227_, new_n12228_, new_n12229_, new_n12230_,
    new_n12231_, new_n12232_, new_n12233_, new_n12234_, new_n12235_,
    new_n12236_, new_n12237_, new_n12238_, new_n12239_, new_n12240_,
    new_n12241_, new_n12242_, new_n12243_, new_n12244_, new_n12245_,
    new_n12246_, new_n12247_, new_n12248_, new_n12249_, new_n12250_,
    new_n12251_, new_n12252_, new_n12253_, new_n12254_, new_n12255_,
    new_n12256_, new_n12257_, new_n12258_, new_n12259_, new_n12260_,
    new_n12261_, new_n12262_, new_n12263_, new_n12264_, new_n12265_,
    new_n12266_, new_n12267_, new_n12268_, new_n12269_, new_n12270_,
    new_n12271_, new_n12272_, new_n12273_, new_n12274_, new_n12275_,
    new_n12276_, new_n12277_, new_n12278_, new_n12279_, new_n12280_,
    new_n12281_, new_n12282_, new_n12283_, new_n12284_, new_n12285_,
    new_n12286_, new_n12287_, new_n12288_, new_n12289_, new_n12290_,
    new_n12291_, new_n12292_, new_n12293_, new_n12294_, new_n12295_,
    new_n12296_, new_n12297_, new_n12298_, new_n12299_, new_n12300_,
    new_n12301_, new_n12302_, new_n12303_, new_n12304_, new_n12305_,
    new_n12306_, new_n12307_, new_n12308_, new_n12309_, new_n12310_,
    new_n12311_, new_n12312_, new_n12313_, new_n12314_, new_n12315_,
    new_n12316_, new_n12317_, new_n12318_, new_n12319_, new_n12320_,
    new_n12321_, new_n12322_, new_n12323_, new_n12324_, new_n12325_,
    new_n12326_, new_n12327_, new_n12328_, new_n12329_, new_n12330_,
    new_n12331_, new_n12332_, new_n12333_, new_n12334_, new_n12335_,
    new_n12336_, new_n12337_, new_n12338_, new_n12339_, new_n12340_,
    new_n12341_, new_n12342_, new_n12343_, new_n12344_, new_n12345_,
    new_n12346_, new_n12347_, new_n12348_, new_n12349_, new_n12350_,
    new_n12351_, new_n12352_, new_n12353_, new_n12354_, new_n12355_,
    new_n12356_, new_n12357_, new_n12358_, new_n12359_, new_n12360_,
    new_n12361_, new_n12362_, new_n12363_, new_n12364_, new_n12365_,
    new_n12366_, new_n12367_, new_n12368_, new_n12369_, new_n12370_,
    new_n12371_, new_n12372_, new_n12373_, new_n12374_, new_n12375_,
    new_n12376_, new_n12377_, new_n12378_, new_n12379_, new_n12380_,
    new_n12381_, new_n12382_, new_n12383_, new_n12384_, new_n12385_,
    new_n12386_, new_n12387_, new_n12388_, new_n12389_, new_n12390_,
    new_n12391_, new_n12392_, new_n12393_, new_n12394_, new_n12395_,
    new_n12396_, new_n12397_, new_n12398_, new_n12399_, new_n12400_,
    new_n12401_, new_n12402_, new_n12403_, new_n12404_, new_n12405_,
    new_n12406_, new_n12407_, new_n12408_, new_n12409_, new_n12410_,
    new_n12411_, new_n12412_, new_n12413_, new_n12414_, new_n12415_,
    new_n12416_, new_n12417_, new_n12418_, new_n12419_, new_n12420_,
    new_n12421_, new_n12422_, new_n12423_, new_n12424_, new_n12425_,
    new_n12426_, new_n12427_, new_n12428_, new_n12429_, new_n12430_,
    new_n12431_, new_n12432_, new_n12433_, new_n12434_, new_n12435_,
    new_n12436_, new_n12437_, new_n12438_, new_n12439_, new_n12440_,
    new_n12441_, new_n12442_, new_n12443_, new_n12444_, new_n12445_,
    new_n12446_, new_n12447_, new_n12448_, new_n12449_, new_n12450_,
    new_n12451_, new_n12452_, new_n12453_, new_n12454_, new_n12455_,
    new_n12456_, new_n12457_, new_n12458_, new_n12459_, new_n12460_,
    new_n12461_, new_n12462_, new_n12463_, new_n12464_, new_n12465_,
    new_n12466_, new_n12467_, new_n12468_, new_n12469_, new_n12470_,
    new_n12471_, new_n12472_, new_n12473_, new_n12474_, new_n12475_,
    new_n12476_, new_n12477_, new_n12478_, new_n12479_, new_n12480_,
    new_n12481_, new_n12482_, new_n12483_, new_n12484_, new_n12485_,
    new_n12486_, new_n12487_, new_n12488_, new_n12489_, new_n12490_,
    new_n12491_, new_n12492_, new_n12493_, new_n12494_, new_n12495_,
    new_n12496_, new_n12497_, new_n12498_, new_n12499_, new_n12500_,
    new_n12501_, new_n12502_, new_n12503_, new_n12504_, new_n12505_,
    new_n12506_, new_n12507_, new_n12508_, new_n12509_, new_n12510_,
    new_n12511_, new_n12512_, new_n12513_, new_n12514_, new_n12515_,
    new_n12516_, new_n12517_, new_n12518_, new_n12519_, new_n12520_,
    new_n12521_, new_n12522_, new_n12523_, new_n12524_, new_n12525_,
    new_n12526_, new_n12527_, new_n12528_, new_n12529_, new_n12530_,
    new_n12531_, new_n12532_, new_n12533_, new_n12534_, new_n12535_,
    new_n12536_, new_n12537_, new_n12538_, new_n12539_, new_n12540_,
    new_n12541_, new_n12542_, new_n12543_, new_n12544_, new_n12545_,
    new_n12546_, new_n12547_, new_n12548_, new_n12549_, new_n12550_,
    new_n12551_, new_n12552_, new_n12553_, new_n12554_, new_n12555_,
    new_n12556_, new_n12557_, new_n12558_, new_n12559_, new_n12560_,
    new_n12561_, new_n12562_, new_n12563_, new_n12564_, new_n12565_,
    new_n12566_, new_n12567_, new_n12568_, new_n12569_, new_n12570_,
    new_n12571_, new_n12572_, new_n12573_, new_n12574_, new_n12575_,
    new_n12576_, new_n12577_, new_n12578_, new_n12579_, new_n12580_,
    new_n12581_, new_n12582_, new_n12583_, new_n12584_, new_n12585_,
    new_n12586_, new_n12587_, new_n12588_, new_n12589_, new_n12590_,
    new_n12591_, new_n12592_, new_n12593_, new_n12594_, new_n12595_,
    new_n12596_, new_n12597_, new_n12598_, new_n12599_, new_n12600_,
    new_n12601_, new_n12602_, new_n12603_, new_n12604_, new_n12605_,
    new_n12606_, new_n12607_, new_n12608_, new_n12609_, new_n12610_,
    new_n12611_, new_n12612_, new_n12613_, new_n12614_, new_n12615_,
    new_n12616_, new_n12617_, new_n12618_, new_n12619_, new_n12620_,
    new_n12621_, new_n12622_, new_n12623_, new_n12624_, new_n12625_,
    new_n12626_, new_n12627_, new_n12628_, new_n12629_, new_n12630_,
    new_n12631_, new_n12632_, new_n12633_, new_n12634_, new_n12635_,
    new_n12636_, new_n12637_, new_n12638_, new_n12639_, new_n12640_,
    new_n12641_, new_n12642_, new_n12643_, new_n12644_, new_n12645_,
    new_n12646_, new_n12647_, new_n12648_, new_n12649_, new_n12650_,
    new_n12651_, new_n12652_, new_n12653_, new_n12654_, new_n12655_,
    new_n12656_, new_n12657_, new_n12658_, new_n12659_, new_n12660_,
    new_n12661_, new_n12662_, new_n12663_, new_n12664_, new_n12665_,
    new_n12666_, new_n12667_, new_n12668_, new_n12669_, new_n12670_,
    new_n12671_, new_n12672_, new_n12673_, new_n12674_, new_n12675_,
    new_n12676_, new_n12677_, new_n12678_, new_n12679_, new_n12680_,
    new_n12681_, new_n12682_, new_n12683_, new_n12684_, new_n12685_,
    new_n12686_, new_n12687_, new_n12688_, new_n12689_, new_n12690_,
    new_n12691_, new_n12692_, new_n12693_, new_n12694_, new_n12695_,
    new_n12696_, new_n12697_, new_n12698_, new_n12699_, new_n12700_,
    new_n12701_, new_n12702_, new_n12703_, new_n12704_, new_n12705_,
    new_n12706_, new_n12707_, new_n12708_, new_n12709_, new_n12710_,
    new_n12711_, new_n12712_, new_n12713_, new_n12714_, new_n12715_,
    new_n12716_, new_n12717_, new_n12718_, new_n12719_, new_n12720_,
    new_n12721_, new_n12722_, new_n12723_, new_n12724_, new_n12725_,
    new_n12726_, new_n12727_, new_n12728_, new_n12729_, new_n12730_,
    new_n12731_, new_n12732_, new_n12733_, new_n12734_, new_n12735_,
    new_n12736_, new_n12737_, new_n12738_, new_n12739_, new_n12740_,
    new_n12741_, new_n12742_, new_n12743_, new_n12744_, new_n12745_,
    new_n12746_, new_n12747_, new_n12748_, new_n12749_, new_n12750_,
    new_n12751_, new_n12752_, new_n12753_, new_n12754_, new_n12755_,
    new_n12756_, new_n12757_, new_n12758_, new_n12759_, new_n12760_,
    new_n12761_, new_n12762_, new_n12763_, new_n12764_, new_n12765_,
    new_n12766_, new_n12767_, new_n12768_, new_n12769_, new_n12770_,
    new_n12771_, new_n12772_, new_n12773_, new_n12774_, new_n12775_,
    new_n12776_, new_n12777_, new_n12778_, new_n12779_, new_n12780_,
    new_n12781_, new_n12782_, new_n12783_, new_n12784_, new_n12785_,
    new_n12786_, new_n12787_, new_n12788_, new_n12789_, new_n12790_,
    new_n12791_, new_n12792_, new_n12793_, new_n12794_, new_n12795_,
    new_n12796_, new_n12797_, new_n12798_, new_n12799_, new_n12800_,
    new_n12801_, new_n12802_, new_n12803_, new_n12804_, new_n12805_,
    new_n12806_, new_n12807_, new_n12808_, new_n12809_, new_n12810_,
    new_n12811_, new_n12812_, new_n12813_, new_n12814_, new_n12815_,
    new_n12816_, new_n12817_, new_n12818_, new_n12819_, new_n12820_,
    new_n12821_, new_n12822_, new_n12823_, new_n12824_, new_n12825_,
    new_n12826_, new_n12827_, new_n12828_, new_n12829_, new_n12830_,
    new_n12831_, new_n12832_, new_n12833_, new_n12834_, new_n12835_,
    new_n12836_, new_n12837_, new_n12838_, new_n12839_, new_n12840_,
    new_n12841_, new_n12842_, new_n12843_, new_n12844_, new_n12845_,
    new_n12846_, new_n12847_, new_n12848_, new_n12849_, new_n12850_,
    new_n12851_, new_n12852_, new_n12853_, new_n12854_, new_n12855_,
    new_n12856_, new_n12857_, new_n12858_, new_n12859_, new_n12860_,
    new_n12861_, new_n12862_, new_n12863_, new_n12864_, new_n12865_,
    new_n12866_, new_n12867_, new_n12868_, new_n12869_, new_n12870_,
    new_n12871_, new_n12872_, new_n12873_, new_n12874_, new_n12875_,
    new_n12876_, new_n12877_, new_n12878_, new_n12879_, new_n12880_,
    new_n12881_, new_n12882_, new_n12883_, new_n12884_, new_n12885_,
    new_n12886_, new_n12887_, new_n12888_, new_n12889_, new_n12890_,
    new_n12891_, new_n12892_, new_n12893_, new_n12894_, new_n12895_,
    new_n12896_, new_n12897_, new_n12898_, new_n12899_, new_n12900_,
    new_n12901_, new_n12902_, new_n12903_, new_n12904_, new_n12905_,
    new_n12906_, new_n12907_, new_n12908_, new_n12909_, new_n12910_,
    new_n12911_, new_n12912_, new_n12913_, new_n12914_, new_n12915_,
    new_n12916_, new_n12917_, new_n12918_, new_n12919_, new_n12920_,
    new_n12921_, new_n12922_, new_n12923_, new_n12924_, new_n12925_,
    new_n12926_, new_n12927_, new_n12928_, new_n12929_, new_n12930_,
    new_n12931_, new_n12932_, new_n12933_, new_n12934_, new_n12935_,
    new_n12936_, new_n12937_, new_n12938_, new_n12939_, new_n12940_,
    new_n12941_, new_n12942_, new_n12943_, new_n12944_, new_n12945_,
    new_n12946_, new_n12947_, new_n12948_, new_n12949_, new_n12950_,
    new_n12951_, new_n12952_, new_n12953_, new_n12954_, new_n12955_,
    new_n12956_, new_n12957_, new_n12958_, new_n12959_, new_n12960_,
    new_n12961_, new_n12962_, new_n12963_, new_n12964_, new_n12965_,
    new_n12966_, new_n12967_, new_n12968_, new_n12969_, new_n12970_,
    new_n12971_, new_n12972_, new_n12973_, new_n12974_, new_n12975_,
    new_n12976_, new_n12977_, new_n12978_, new_n12979_, new_n12980_,
    new_n12981_, new_n12982_, new_n12983_, new_n12984_, new_n12985_,
    new_n12986_, new_n12987_, new_n12988_, new_n12989_, new_n12990_,
    new_n12991_, new_n12992_, new_n12993_, new_n12994_, new_n12995_,
    new_n12996_, new_n12997_, new_n12998_, new_n12999_, new_n13000_,
    new_n13001_, new_n13002_, new_n13003_, new_n13004_, new_n13005_,
    new_n13006_, new_n13007_, new_n13008_, new_n13009_, new_n13010_,
    new_n13011_, new_n13012_, new_n13013_, new_n13014_, new_n13015_,
    new_n13016_, new_n13017_, new_n13018_, new_n13019_, new_n13020_,
    new_n13021_, new_n13022_, new_n13023_, new_n13024_, new_n13025_,
    new_n13026_, new_n13027_, new_n13028_, new_n13029_, new_n13030_,
    new_n13031_, new_n13032_, new_n13033_, new_n13034_, new_n13035_,
    new_n13036_, new_n13037_, new_n13038_, new_n13039_, new_n13040_,
    new_n13041_, new_n13042_, new_n13043_, new_n13044_, new_n13045_,
    new_n13046_, new_n13047_, new_n13048_, new_n13049_, new_n13050_,
    new_n13051_, new_n13052_, new_n13053_, new_n13054_, new_n13055_,
    new_n13056_, new_n13057_, new_n13058_, new_n13059_, new_n13060_,
    new_n13061_, new_n13062_, new_n13063_, new_n13064_, new_n13065_,
    new_n13066_, new_n13067_, new_n13068_, new_n13069_, new_n13070_,
    new_n13071_, new_n13072_, new_n13073_, new_n13074_, new_n13075_,
    new_n13076_, new_n13077_, new_n13078_, new_n13079_, new_n13080_,
    new_n13081_, new_n13082_, new_n13083_, new_n13084_, new_n13085_,
    new_n13086_, new_n13087_, new_n13088_, new_n13089_, new_n13090_,
    new_n13091_, new_n13092_, new_n13093_, new_n13094_, new_n13095_,
    new_n13096_, new_n13097_, new_n13098_, new_n13099_, new_n13100_,
    new_n13101_, new_n13102_, new_n13103_, new_n13104_, new_n13105_,
    new_n13106_, new_n13107_, new_n13108_, new_n13109_, new_n13110_,
    new_n13111_, new_n13112_, new_n13113_, new_n13114_, new_n13115_,
    new_n13116_, new_n13117_, new_n13118_, new_n13119_, new_n13120_,
    new_n13121_, new_n13122_, new_n13123_, new_n13124_, new_n13125_,
    new_n13126_, new_n13127_, new_n13128_, new_n13129_, new_n13130_,
    new_n13131_, new_n13132_, new_n13133_, new_n13134_, new_n13135_,
    new_n13136_, new_n13137_, new_n13138_, new_n13139_, new_n13140_,
    new_n13141_, new_n13142_, new_n13143_, new_n13144_, new_n13145_,
    new_n13146_, new_n13147_, new_n13148_, new_n13149_, new_n13150_,
    new_n13151_, new_n13152_, new_n13153_, new_n13154_, new_n13155_,
    new_n13156_, new_n13157_, new_n13158_, new_n13159_, new_n13160_,
    new_n13161_, new_n13162_, new_n13163_, new_n13164_, new_n13165_,
    new_n13166_, new_n13167_, new_n13168_, new_n13169_, new_n13170_,
    new_n13171_, new_n13172_, new_n13173_, new_n13174_, new_n13175_,
    new_n13176_, new_n13177_, new_n13178_, new_n13179_, new_n13180_,
    new_n13181_, new_n13182_, new_n13183_, new_n13184_, new_n13185_,
    new_n13186_, new_n13187_, new_n13188_, new_n13189_, new_n13190_,
    new_n13191_, new_n13192_, new_n13193_, new_n13194_, new_n13195_,
    new_n13196_, new_n13197_, new_n13198_, new_n13199_, new_n13200_,
    new_n13201_, new_n13202_, new_n13203_, new_n13204_, new_n13205_,
    new_n13206_, new_n13207_, new_n13208_, new_n13209_, new_n13210_,
    new_n13211_, new_n13212_, new_n13213_, new_n13214_, new_n13215_,
    new_n13216_, new_n13217_, new_n13218_, new_n13219_, new_n13220_,
    new_n13221_, new_n13222_, new_n13223_, new_n13224_, new_n13225_,
    new_n13226_, new_n13227_, new_n13228_, new_n13229_, new_n13230_,
    new_n13231_, new_n13232_, new_n13233_, new_n13234_, new_n13235_,
    new_n13236_, new_n13237_, new_n13238_, new_n13239_, new_n13240_,
    new_n13241_, new_n13242_, new_n13243_, new_n13244_, new_n13245_,
    new_n13246_, new_n13247_, new_n13248_, new_n13249_, new_n13250_,
    new_n13251_, new_n13252_, new_n13253_, new_n13254_, new_n13255_,
    new_n13256_, new_n13257_, new_n13258_, new_n13259_, new_n13260_,
    new_n13261_, new_n13262_, new_n13263_, new_n13264_, new_n13265_,
    new_n13266_, new_n13267_, new_n13268_, new_n13269_, new_n13270_,
    new_n13271_, new_n13272_, new_n13273_, new_n13274_, new_n13275_,
    new_n13276_, new_n13277_, new_n13278_, new_n13279_, new_n13280_,
    new_n13281_, new_n13282_, new_n13283_, new_n13284_, new_n13285_,
    new_n13286_, new_n13287_, new_n13288_, new_n13289_, new_n13290_,
    new_n13291_, new_n13292_, new_n13293_, new_n13294_, new_n13295_,
    new_n13296_, new_n13297_, new_n13298_, new_n13299_, new_n13300_,
    new_n13301_, new_n13302_, new_n13303_, new_n13304_, new_n13305_,
    new_n13306_, new_n13307_, new_n13308_, new_n13309_, new_n13310_,
    new_n13311_, new_n13312_, new_n13313_, new_n13314_, new_n13315_,
    new_n13316_, new_n13317_, new_n13318_, new_n13319_, new_n13320_,
    new_n13321_, new_n13322_, new_n13323_, new_n13324_, new_n13325_,
    new_n13326_, new_n13327_, new_n13328_, new_n13329_, new_n13330_,
    new_n13331_, new_n13332_, new_n13333_, new_n13334_, new_n13335_,
    new_n13336_, new_n13337_, new_n13338_, new_n13339_, new_n13340_,
    new_n13341_, new_n13342_, new_n13343_, new_n13344_, new_n13345_,
    new_n13346_, new_n13347_, new_n13348_, new_n13349_, new_n13350_,
    new_n13351_, new_n13352_, new_n13353_, new_n13354_, new_n13355_,
    new_n13356_, new_n13357_, new_n13358_, new_n13359_, new_n13360_,
    new_n13361_, new_n13362_, new_n13363_, new_n13364_, new_n13365_,
    new_n13366_, new_n13367_, new_n13368_, new_n13369_, new_n13370_,
    new_n13371_, new_n13372_, new_n13373_, new_n13374_, new_n13375_,
    new_n13376_, new_n13377_, new_n13378_, new_n13379_, new_n13380_,
    new_n13381_, new_n13382_, new_n13383_, new_n13384_, new_n13385_,
    new_n13386_, new_n13387_, new_n13388_, new_n13389_, new_n13390_,
    new_n13391_, new_n13392_, new_n13393_, new_n13394_, new_n13395_,
    new_n13396_, new_n13397_, new_n13398_, new_n13399_, new_n13400_,
    new_n13401_, new_n13402_, new_n13403_, new_n13404_, new_n13405_,
    new_n13406_, new_n13407_, new_n13408_, new_n13409_, new_n13410_,
    new_n13411_, new_n13412_, new_n13413_, new_n13414_, new_n13415_,
    new_n13416_, new_n13417_, new_n13418_, new_n13419_, new_n13420_,
    new_n13421_, new_n13422_, new_n13423_, new_n13424_, new_n13425_,
    new_n13426_, new_n13427_, new_n13428_, new_n13429_, new_n13430_,
    new_n13431_, new_n13432_, new_n13433_, new_n13434_, new_n13435_,
    new_n13436_, new_n13437_, new_n13438_, new_n13439_, new_n13440_,
    new_n13441_, new_n13442_, new_n13443_, new_n13444_, new_n13445_,
    new_n13446_, new_n13447_, new_n13448_, new_n13449_, new_n13450_,
    new_n13451_, new_n13452_, new_n13453_, new_n13454_, new_n13455_,
    new_n13456_, new_n13457_, new_n13458_, new_n13459_, new_n13460_,
    new_n13461_, new_n13462_, new_n13463_, new_n13464_, new_n13465_,
    new_n13466_, new_n13467_, new_n13468_, new_n13469_, new_n13470_,
    new_n13471_, new_n13472_, new_n13473_, new_n13474_, new_n13475_,
    new_n13476_, new_n13477_, new_n13478_, new_n13479_, new_n13480_,
    new_n13481_, new_n13482_, new_n13483_, new_n13484_, new_n13485_,
    new_n13486_, new_n13487_, new_n13488_, new_n13489_, new_n13490_,
    new_n13491_, new_n13492_, new_n13493_, new_n13494_, new_n13495_,
    new_n13496_, new_n13497_, new_n13498_, new_n13499_, new_n13500_,
    new_n13501_, new_n13502_, new_n13503_, new_n13504_, new_n13505_,
    new_n13506_, new_n13507_, new_n13508_, new_n13509_, new_n13510_,
    new_n13511_, new_n13512_, new_n13513_, new_n13514_, new_n13515_,
    new_n13516_, new_n13517_, new_n13518_, new_n13519_, new_n13520_,
    new_n13521_, new_n13522_, new_n13523_, new_n13524_, new_n13525_,
    new_n13526_, new_n13527_, new_n13528_, new_n13529_, new_n13530_,
    new_n13531_, new_n13532_, new_n13533_, new_n13534_, new_n13535_,
    new_n13536_, new_n13537_, new_n13538_, new_n13539_, new_n13540_,
    new_n13541_, new_n13542_, new_n13543_, new_n13544_, new_n13545_,
    new_n13546_, new_n13547_, new_n13548_, new_n13549_, new_n13550_,
    new_n13551_, new_n13552_, new_n13553_, new_n13554_, new_n13555_,
    new_n13556_, new_n13557_, new_n13558_, new_n13559_, new_n13560_,
    new_n13561_, new_n13562_, new_n13563_, new_n13564_, new_n13565_,
    new_n13566_, new_n13567_, new_n13568_, new_n13569_, new_n13570_,
    new_n13571_, new_n13572_, new_n13573_, new_n13574_, new_n13575_,
    new_n13576_, new_n13577_, new_n13578_, new_n13579_, new_n13580_,
    new_n13581_, new_n13582_, new_n13583_, new_n13584_, new_n13585_,
    new_n13586_, new_n13587_, new_n13588_, new_n13589_, new_n13590_,
    new_n13591_, new_n13592_, new_n13593_, new_n13594_, new_n13595_,
    new_n13596_, new_n13597_, new_n13598_, new_n13599_, new_n13600_,
    new_n13601_, new_n13602_, new_n13603_, new_n13604_, new_n13605_,
    new_n13606_, new_n13607_, new_n13608_, new_n13609_, new_n13610_,
    new_n13611_, new_n13612_, new_n13613_, new_n13614_, new_n13615_,
    new_n13616_, new_n13617_, new_n13618_, new_n13619_, new_n13620_,
    new_n13621_, new_n13622_, new_n13623_, new_n13624_, new_n13625_,
    new_n13626_, new_n13627_, new_n13628_, new_n13629_, new_n13630_,
    new_n13631_, new_n13632_, new_n13633_, new_n13634_, new_n13635_,
    new_n13636_, new_n13637_, new_n13638_, new_n13639_, new_n13640_,
    new_n13641_, new_n13642_, new_n13643_, new_n13644_, new_n13645_,
    new_n13646_, new_n13647_, new_n13648_, new_n13649_, new_n13650_,
    new_n13651_, new_n13652_, new_n13653_, new_n13654_, new_n13655_,
    new_n13656_, new_n13657_, new_n13658_, new_n13659_, new_n13660_,
    new_n13661_, new_n13662_, new_n13663_, new_n13664_, new_n13665_,
    new_n13666_, new_n13667_, new_n13668_, new_n13669_, new_n13670_,
    new_n13671_, new_n13672_, new_n13673_, new_n13674_, new_n13675_,
    new_n13676_, new_n13677_, new_n13678_, new_n13679_, new_n13680_,
    new_n13681_, new_n13682_, new_n13683_, new_n13684_, new_n13685_,
    new_n13686_, new_n13687_, new_n13688_, new_n13689_, new_n13690_,
    new_n13691_, new_n13692_, new_n13693_, new_n13694_, new_n13695_,
    new_n13696_, new_n13697_, new_n13698_, new_n13699_, new_n13700_,
    new_n13701_, new_n13702_, new_n13703_, new_n13704_, new_n13705_,
    new_n13706_, new_n13707_, new_n13708_, new_n13709_, new_n13710_,
    new_n13711_, new_n13712_, new_n13713_, new_n13714_, new_n13715_,
    new_n13716_, new_n13717_, new_n13718_, new_n13719_, new_n13720_,
    new_n13721_, new_n13722_, new_n13723_, new_n13724_, new_n13725_,
    new_n13726_, new_n13727_, new_n13728_, new_n13729_, new_n13730_,
    new_n13731_, new_n13732_, new_n13733_, new_n13734_, new_n13735_,
    new_n13736_, new_n13737_, new_n13738_, new_n13739_, new_n13740_,
    new_n13741_, new_n13742_, new_n13743_, new_n13744_, new_n13745_,
    new_n13746_, new_n13747_, new_n13748_, new_n13749_, new_n13750_,
    new_n13751_, new_n13752_, new_n13753_, new_n13754_, new_n13755_,
    new_n13756_, new_n13757_, new_n13758_, new_n13759_, new_n13760_,
    new_n13761_, new_n13762_, new_n13763_, new_n13764_, new_n13765_,
    new_n13766_, new_n13767_, new_n13768_, new_n13769_, new_n13770_,
    new_n13771_, new_n13772_, new_n13773_, new_n13774_, new_n13775_,
    new_n13776_, new_n13777_, new_n13778_, new_n13779_, new_n13780_,
    new_n13781_, new_n13782_, new_n13783_, new_n13784_, new_n13785_,
    new_n13786_, new_n13787_, new_n13788_, new_n13789_, new_n13790_,
    new_n13791_, new_n13792_, new_n13793_, new_n13794_, new_n13795_,
    new_n13796_, new_n13797_, new_n13798_, new_n13799_, new_n13800_,
    new_n13801_, new_n13802_, new_n13803_, new_n13804_, new_n13805_,
    new_n13806_, new_n13807_, new_n13808_, new_n13809_, new_n13810_,
    new_n13811_, new_n13812_, new_n13813_, new_n13814_, new_n13815_,
    new_n13816_, new_n13817_, new_n13818_, new_n13819_, new_n13820_,
    new_n13821_, new_n13822_, new_n13823_, new_n13824_, new_n13825_,
    new_n13826_, new_n13827_, new_n13828_, new_n13829_, new_n13830_,
    new_n13831_, new_n13832_, new_n13833_, new_n13834_, new_n13835_,
    new_n13836_, new_n13837_, new_n13838_, new_n13839_, new_n13840_,
    new_n13841_, new_n13842_, new_n13843_, new_n13844_, new_n13845_,
    new_n13846_, new_n13847_, new_n13848_, new_n13849_, new_n13850_,
    new_n13851_, new_n13852_, new_n13853_, new_n13854_, new_n13855_,
    new_n13856_, new_n13857_, new_n13858_, new_n13859_, new_n13860_,
    new_n13861_, new_n13862_, new_n13863_, new_n13864_, new_n13865_,
    new_n13866_, new_n13867_, new_n13868_, new_n13869_, new_n13870_,
    new_n13871_, new_n13872_, new_n13873_, new_n13874_, new_n13875_,
    new_n13876_, new_n13877_, new_n13878_, new_n13879_, new_n13880_,
    new_n13881_, new_n13882_, new_n13883_, new_n13884_, new_n13885_,
    new_n13886_, new_n13887_, new_n13888_, new_n13889_, new_n13890_,
    new_n13891_, new_n13892_, new_n13893_, new_n13894_, new_n13895_,
    new_n13896_, new_n13897_, new_n13898_, new_n13899_, new_n13900_,
    new_n13901_, new_n13902_, new_n13903_, new_n13904_, new_n13905_,
    new_n13906_, new_n13907_, new_n13908_, new_n13909_, new_n13910_,
    new_n13911_, new_n13912_, new_n13913_, new_n13914_, new_n13915_,
    new_n13916_, new_n13917_, new_n13918_, new_n13919_, new_n13920_,
    new_n13921_, new_n13922_, new_n13923_, new_n13924_, new_n13925_,
    new_n13926_, new_n13927_, new_n13928_, new_n13929_, new_n13930_,
    new_n13931_, new_n13932_, new_n13933_, new_n13934_, new_n13935_,
    new_n13936_, new_n13937_, new_n13938_, new_n13939_, new_n13940_,
    new_n13941_, new_n13942_, new_n13943_, new_n13944_, new_n13945_,
    new_n13946_, new_n13947_, new_n13948_, new_n13949_, new_n13950_,
    new_n13951_, new_n13952_, new_n13953_, new_n13954_, new_n13955_,
    new_n13956_, new_n13957_, new_n13958_, new_n13959_, new_n13960_,
    new_n13961_, new_n13962_, new_n13963_, new_n13964_, new_n13965_,
    new_n13966_, new_n13967_, new_n13968_, new_n13969_, new_n13970_,
    new_n13971_, new_n13972_, new_n13973_, new_n13974_, new_n13975_,
    new_n13976_, new_n13977_, new_n13978_, new_n13979_, new_n13980_,
    new_n13981_, new_n13982_, new_n13983_, new_n13984_, new_n13985_,
    new_n13986_, new_n13987_, new_n13988_, new_n13989_, new_n13990_,
    new_n13991_, new_n13992_, new_n13993_, new_n13994_, new_n13995_,
    new_n13996_, new_n13997_, new_n13998_, new_n13999_, new_n14000_,
    new_n14001_, new_n14002_, new_n14003_, new_n14004_, new_n14005_,
    new_n14006_, new_n14007_, new_n14008_, new_n14009_, new_n14010_,
    new_n14011_, new_n14012_, new_n14013_, new_n14014_, new_n14015_,
    new_n14016_, new_n14017_, new_n14018_, new_n14019_, new_n14020_,
    new_n14021_, new_n14022_, new_n14023_, new_n14024_, new_n14025_,
    new_n14026_, new_n14027_, new_n14028_, new_n14029_, new_n14030_,
    new_n14031_, new_n14032_, new_n14033_, new_n14034_, new_n14035_,
    new_n14036_, new_n14037_, new_n14038_, new_n14039_, new_n14040_,
    new_n14041_, new_n14042_, new_n14043_, new_n14044_, new_n14045_,
    new_n14046_, new_n14047_, new_n14048_, new_n14049_, new_n14050_,
    new_n14051_, new_n14052_, new_n14053_, new_n14054_, new_n14055_,
    new_n14056_, new_n14057_, new_n14058_, new_n14059_, new_n14060_,
    new_n14061_, new_n14062_, new_n14063_, new_n14064_, new_n14065_,
    new_n14066_, new_n14067_, new_n14068_, new_n14069_, new_n14070_,
    new_n14071_, new_n14072_, new_n14073_, new_n14074_, new_n14075_,
    new_n14076_, new_n14077_, new_n14078_, new_n14079_, new_n14080_,
    new_n14081_, new_n14082_, new_n14083_, new_n14084_, new_n14085_,
    new_n14086_, new_n14087_, new_n14088_, new_n14089_, new_n14090_,
    new_n14091_, new_n14092_, new_n14093_, new_n14094_, new_n14095_,
    new_n14096_, new_n14097_, new_n14098_, new_n14099_, new_n14100_,
    new_n14101_, new_n14102_, new_n14103_, new_n14104_, new_n14105_,
    new_n14106_, new_n14107_, new_n14108_, new_n14109_, new_n14110_,
    new_n14111_, new_n14112_, new_n14113_, new_n14114_, new_n14115_,
    new_n14116_, new_n14117_, new_n14118_, new_n14119_, new_n14120_,
    new_n14121_, new_n14122_, new_n14123_, new_n14124_, new_n14125_,
    new_n14126_, new_n14127_, new_n14128_, new_n14129_, new_n14130_,
    new_n14131_, new_n14132_, new_n14133_, new_n14134_, new_n14135_,
    new_n14136_, new_n14137_, new_n14138_, new_n14139_, new_n14140_,
    new_n14141_, new_n14142_, new_n14143_, new_n14144_, new_n14145_,
    new_n14146_, new_n14147_, new_n14148_, new_n14149_, new_n14150_,
    new_n14151_, new_n14152_, new_n14153_, new_n14154_, new_n14155_,
    new_n14156_, new_n14157_, new_n14158_, new_n14159_, new_n14160_,
    new_n14161_, new_n14162_, new_n14163_, new_n14164_, new_n14165_,
    new_n14166_, new_n14167_, new_n14168_, new_n14169_, new_n14170_,
    new_n14171_, new_n14172_, new_n14173_, new_n14174_, new_n14175_,
    new_n14176_, new_n14177_, new_n14178_, new_n14179_, new_n14180_,
    new_n14181_, new_n14182_, new_n14183_, new_n14184_, new_n14185_,
    new_n14186_, new_n14187_, new_n14188_, new_n14189_, new_n14190_,
    new_n14191_, new_n14192_, new_n14193_, new_n14194_, new_n14195_,
    new_n14196_, new_n14197_, new_n14198_, new_n14199_, new_n14200_,
    new_n14201_, new_n14202_, new_n14203_, new_n14204_, new_n14205_,
    new_n14206_, new_n14207_, new_n14208_, new_n14209_, new_n14210_,
    new_n14211_, new_n14212_, new_n14213_, new_n14214_, new_n14215_,
    new_n14216_, new_n14217_, new_n14218_, new_n14219_, new_n14220_,
    new_n14221_, new_n14222_, new_n14223_, new_n14224_, new_n14225_,
    new_n14226_, new_n14227_, new_n14228_, new_n14229_, new_n14230_,
    new_n14231_, new_n14232_, new_n14233_, new_n14234_, new_n14235_,
    new_n14236_, new_n14237_, new_n14238_, new_n14239_, new_n14240_,
    new_n14241_, new_n14242_, new_n14243_, new_n14244_, new_n14245_,
    new_n14246_, new_n14247_, new_n14248_, new_n14249_, new_n14250_,
    new_n14251_, new_n14252_, new_n14253_, new_n14254_, new_n14255_,
    new_n14256_, new_n14257_, new_n14258_, new_n14259_, new_n14260_,
    new_n14261_, new_n14262_, new_n14263_, new_n14264_, new_n14265_,
    new_n14266_, new_n14267_, new_n14268_, new_n14269_, new_n14270_,
    new_n14271_, new_n14272_, new_n14273_, new_n14274_, new_n14275_,
    new_n14276_, new_n14277_, new_n14278_, new_n14279_, new_n14280_,
    new_n14281_, new_n14282_, new_n14283_, new_n14284_, new_n14285_,
    new_n14286_, new_n14287_, new_n14288_, new_n14289_, new_n14290_,
    new_n14291_, new_n14292_, new_n14293_, new_n14294_, new_n14295_,
    new_n14296_, new_n14297_, new_n14298_, new_n14299_, new_n14300_,
    new_n14301_, new_n14302_, new_n14303_, new_n14304_, new_n14305_,
    new_n14306_, new_n14307_, new_n14308_, new_n14309_, new_n14310_,
    new_n14311_, new_n14312_, new_n14313_, new_n14314_, new_n14315_,
    new_n14316_, new_n14317_, new_n14318_, new_n14319_, new_n14320_,
    new_n14321_, new_n14322_, new_n14323_, new_n14324_, new_n14325_,
    new_n14326_, new_n14327_, new_n14328_, new_n14329_, new_n14330_,
    new_n14331_, new_n14332_, new_n14333_, new_n14334_, new_n14335_,
    new_n14336_, new_n14337_, new_n14338_, new_n14339_, new_n14340_,
    new_n14341_, new_n14342_, new_n14343_, new_n14344_, new_n14345_,
    new_n14346_, new_n14347_, new_n14348_, new_n14349_, new_n14350_,
    new_n14351_, new_n14352_, new_n14353_, new_n14354_, new_n14355_,
    new_n14356_, new_n14357_, new_n14358_, new_n14359_, new_n14360_,
    new_n14361_, new_n14362_, new_n14363_, new_n14364_, new_n14365_,
    new_n14366_, new_n14367_, new_n14368_, new_n14369_, new_n14370_,
    new_n14371_, new_n14372_, new_n14373_, new_n14374_, new_n14375_,
    new_n14376_, new_n14377_, new_n14378_, new_n14379_, new_n14380_,
    new_n14381_, new_n14382_, new_n14383_, new_n14384_, new_n14385_,
    new_n14386_, new_n14387_, new_n14388_, new_n14389_, new_n14390_,
    new_n14391_, new_n14392_, new_n14393_, new_n14394_, new_n14395_,
    new_n14396_, new_n14397_, new_n14398_, new_n14399_, new_n14400_,
    new_n14401_, new_n14402_, new_n14403_, new_n14404_, new_n14405_,
    new_n14406_, new_n14407_, new_n14408_, new_n14409_, new_n14410_,
    new_n14411_, new_n14412_, new_n14413_, new_n14414_, new_n14415_,
    new_n14416_, new_n14417_, new_n14418_, new_n14419_, new_n14420_,
    new_n14421_, new_n14422_, new_n14423_, new_n14424_, new_n14425_,
    new_n14426_, new_n14427_, new_n14428_, new_n14429_, new_n14430_,
    new_n14431_, new_n14432_, new_n14433_, new_n14434_, new_n14435_,
    new_n14436_, new_n14437_, new_n14438_, new_n14439_, new_n14440_,
    new_n14441_, new_n14442_, new_n14443_, new_n14444_, new_n14445_,
    new_n14446_, new_n14447_, new_n14448_, new_n14449_, new_n14450_,
    new_n14451_, new_n14452_, new_n14453_, new_n14454_, new_n14455_,
    new_n14456_, new_n14457_, new_n14458_, new_n14459_, new_n14460_,
    new_n14461_, new_n14462_, new_n14463_, new_n14464_, new_n14465_,
    new_n14466_, new_n14467_, new_n14468_, new_n14469_, new_n14470_,
    new_n14471_, new_n14472_, new_n14473_, new_n14474_, new_n14475_,
    new_n14476_, new_n14477_, new_n14478_, new_n14479_, new_n14480_,
    new_n14481_, new_n14482_, new_n14483_, new_n14484_, new_n14485_,
    new_n14486_, new_n14487_, new_n14488_, new_n14489_, new_n14490_,
    new_n14491_, new_n14492_, new_n14493_, new_n14494_, new_n14495_,
    new_n14496_, new_n14497_, new_n14498_, new_n14499_, new_n14500_,
    new_n14501_, new_n14502_, new_n14503_, new_n14504_, new_n14505_,
    new_n14506_, new_n14507_, new_n14508_, new_n14509_, new_n14510_,
    new_n14511_, new_n14512_, new_n14513_, new_n14514_, new_n14515_,
    new_n14516_, new_n14517_, new_n14518_, new_n14519_, new_n14520_,
    new_n14521_, new_n14522_, new_n14523_, new_n14524_, new_n14525_,
    new_n14526_, new_n14527_, new_n14528_, new_n14529_, new_n14530_,
    new_n14531_, new_n14532_, new_n14533_, new_n14534_, new_n14535_,
    new_n14536_, new_n14537_, new_n14538_, new_n14539_, new_n14540_,
    new_n14541_, new_n14542_, new_n14543_, new_n14544_, new_n14545_,
    new_n14546_, new_n14547_, new_n14548_, new_n14549_, new_n14550_,
    new_n14551_, new_n14552_, new_n14553_, new_n14554_, new_n14555_,
    new_n14556_, new_n14557_, new_n14558_, new_n14559_, new_n14560_,
    new_n14561_, new_n14562_, new_n14563_, new_n14564_, new_n14565_,
    new_n14566_, new_n14567_, new_n14568_, new_n14569_, new_n14570_,
    new_n14571_, new_n14572_, new_n14573_, new_n14574_, new_n14575_,
    new_n14576_, new_n14577_, new_n14578_, new_n14579_, new_n14580_,
    new_n14581_, new_n14582_, new_n14583_, new_n14584_, new_n14585_,
    new_n14586_, new_n14587_, new_n14588_, new_n14589_, new_n14590_,
    new_n14591_, new_n14592_, new_n14593_, new_n14594_, new_n14595_,
    new_n14596_, new_n14597_, new_n14598_, new_n14599_, new_n14600_,
    new_n14601_, new_n14602_, new_n14603_, new_n14604_, new_n14605_,
    new_n14606_, new_n14607_, new_n14608_, new_n14609_, new_n14610_,
    new_n14611_, new_n14612_, new_n14613_, new_n14614_, new_n14615_,
    new_n14616_, new_n14617_, new_n14618_, new_n14619_, new_n14620_,
    new_n14621_, new_n14622_, new_n14623_, new_n14624_, new_n14625_,
    new_n14626_, new_n14627_, new_n14628_, new_n14629_, new_n14630_,
    new_n14631_, new_n14632_, new_n14633_, new_n14634_, new_n14635_,
    new_n14636_, new_n14637_, new_n14638_, new_n14639_, new_n14640_,
    new_n14641_, new_n14642_, new_n14643_, new_n14644_, new_n14645_,
    new_n14646_, new_n14647_, new_n14648_, new_n14649_, new_n14650_,
    new_n14651_, new_n14652_, new_n14653_, new_n14654_, new_n14655_,
    new_n14656_, new_n14657_, new_n14658_, new_n14659_, new_n14660_,
    new_n14661_, new_n14662_, new_n14663_, new_n14664_, new_n14665_,
    new_n14666_, new_n14667_, new_n14668_, new_n14669_, new_n14670_,
    new_n14671_, new_n14672_, new_n14673_, new_n14674_, new_n14675_,
    new_n14676_, new_n14677_, new_n14678_, new_n14679_, new_n14680_,
    new_n14681_, new_n14682_, new_n14683_, new_n14684_, new_n14685_,
    new_n14686_, new_n14687_, new_n14688_, new_n14689_, new_n14690_,
    new_n14691_, new_n14692_, new_n14693_, new_n14694_, new_n14695_,
    new_n14696_, new_n14697_, new_n14698_, new_n14699_, new_n14700_,
    new_n14701_, new_n14702_, new_n14703_, new_n14704_, new_n14705_,
    new_n14706_, new_n14707_, new_n14708_, new_n14709_, new_n14710_,
    new_n14711_, new_n14712_, new_n14713_, new_n14714_, new_n14715_,
    new_n14716_, new_n14717_, new_n14718_, new_n14719_, new_n14720_,
    new_n14721_, new_n14722_, new_n14723_, new_n14724_, new_n14725_,
    new_n14726_, new_n14727_, new_n14728_, new_n14729_, new_n14730_,
    new_n14731_, new_n14732_, new_n14733_, new_n14734_, new_n14735_,
    new_n14736_, new_n14737_, new_n14738_, new_n14739_, new_n14740_,
    new_n14741_, new_n14742_, new_n14743_, new_n14744_, new_n14745_,
    new_n14746_, new_n14747_, new_n14748_, new_n14749_, new_n14750_,
    new_n14751_, new_n14752_, new_n14753_, new_n14754_, new_n14755_,
    new_n14756_, new_n14757_, new_n14758_, new_n14759_, new_n14760_,
    new_n14761_, new_n14762_, new_n14763_, new_n14764_, new_n14765_,
    new_n14766_, new_n14767_, new_n14768_, new_n14769_, new_n14770_,
    new_n14771_, new_n14772_, new_n14773_, new_n14774_, new_n14775_,
    new_n14776_, new_n14777_, new_n14778_, new_n14779_, new_n14780_,
    new_n14781_, new_n14782_, new_n14783_, new_n14784_, new_n14785_,
    new_n14786_, new_n14787_, new_n14788_, new_n14789_, new_n14790_,
    new_n14791_, new_n14792_, new_n14793_, new_n14794_, new_n14795_,
    new_n14796_, new_n14797_, new_n14798_, new_n14799_, new_n14800_,
    new_n14801_, new_n14802_, new_n14803_, new_n14804_, new_n14805_,
    new_n14806_, new_n14807_, new_n14808_, new_n14809_, new_n14810_,
    new_n14811_, new_n14812_, new_n14813_, new_n14814_, new_n14815_,
    new_n14816_, new_n14817_, new_n14818_, new_n14819_, new_n14820_,
    new_n14821_, new_n14822_, new_n14823_, new_n14824_, new_n14825_,
    new_n14826_, new_n14827_, new_n14828_, new_n14829_, new_n14830_,
    new_n14831_, new_n14832_, new_n14833_, new_n14834_, new_n14835_,
    new_n14836_, new_n14837_, new_n14838_, new_n14839_, new_n14840_,
    new_n14841_, new_n14842_, new_n14843_, new_n14844_, new_n14845_,
    new_n14846_, new_n14847_, new_n14848_, new_n14849_, new_n14850_,
    new_n14851_, new_n14852_, new_n14853_, new_n14854_, new_n14855_,
    new_n14856_, new_n14857_, new_n14858_, new_n14859_, new_n14860_,
    new_n14861_, new_n14862_, new_n14863_, new_n14864_, new_n14865_,
    new_n14866_, new_n14867_, new_n14868_, new_n14869_, new_n14870_,
    new_n14871_, new_n14872_, new_n14873_, new_n14874_, new_n14875_,
    new_n14876_, new_n14877_, new_n14878_, new_n14879_, new_n14880_,
    new_n14881_, new_n14882_, new_n14883_, new_n14884_, new_n14885_,
    new_n14886_, new_n14887_, new_n14888_, new_n14889_, new_n14890_,
    new_n14891_, new_n14892_, new_n14893_, new_n14894_, new_n14895_,
    new_n14896_, new_n14897_, new_n14898_, new_n14899_, new_n14900_,
    new_n14901_, new_n14902_, new_n14903_, new_n14904_, new_n14905_,
    new_n14906_, new_n14907_, new_n14908_, new_n14909_, new_n14910_,
    new_n14911_, new_n14912_, new_n14913_, new_n14914_, new_n14915_,
    new_n14916_, new_n14917_, new_n14918_, new_n14919_, new_n14920_,
    new_n14921_, new_n14922_, new_n14923_, new_n14924_, new_n14925_,
    new_n14926_, new_n14927_, new_n14928_, new_n14929_, new_n14930_,
    new_n14931_, new_n14932_, new_n14933_, new_n14934_, new_n14935_,
    new_n14936_, new_n14937_, new_n14938_, new_n14939_, new_n14940_,
    new_n14941_, new_n14942_, new_n14943_, new_n14944_, new_n14945_,
    new_n14946_, new_n14947_, new_n14948_, new_n14949_, new_n14950_,
    new_n14951_, new_n14952_, new_n14953_, new_n14954_, new_n14955_,
    new_n14956_, new_n14957_, new_n14958_, new_n14959_, new_n14960_,
    new_n14961_, new_n14962_, new_n14963_, new_n14964_, new_n14965_,
    new_n14966_, new_n14967_, new_n14968_, new_n14969_, new_n14970_,
    new_n14971_, new_n14972_, new_n14973_, new_n14974_, new_n14975_,
    new_n14976_, new_n14977_, new_n14978_, new_n14979_, new_n14980_,
    new_n14981_, new_n14982_, new_n14983_, new_n14984_, new_n14985_,
    new_n14986_, new_n14987_, new_n14988_, new_n14989_, new_n14990_,
    new_n14991_, new_n14992_, new_n14993_, new_n14994_, new_n14995_,
    new_n14996_, new_n14997_, new_n14998_, new_n14999_, new_n15000_,
    new_n15001_, new_n15002_, new_n15003_, new_n15004_, new_n15005_,
    new_n15006_, new_n15007_, new_n15008_, new_n15009_, new_n15010_,
    new_n15011_, new_n15012_, new_n15013_, new_n15014_, new_n15015_,
    new_n15016_, new_n15017_, new_n15018_, new_n15019_, new_n15020_,
    new_n15021_, new_n15022_, new_n15023_, new_n15024_, new_n15025_,
    new_n15026_, new_n15027_, new_n15028_, new_n15029_, new_n15030_,
    new_n15031_, new_n15032_, new_n15033_, new_n15034_, new_n15035_,
    new_n15036_, new_n15037_, new_n15038_, new_n15039_, new_n15040_,
    new_n15041_, new_n15042_, new_n15043_, new_n15044_, new_n15045_,
    new_n15046_, new_n15047_, new_n15048_, new_n15049_, new_n15050_,
    new_n15051_, new_n15052_, new_n15053_, new_n15054_, new_n15055_,
    new_n15056_, new_n15057_, new_n15058_, new_n15059_, new_n15060_,
    new_n15061_, new_n15062_, new_n15063_, new_n15064_, new_n15065_,
    new_n15066_, new_n15067_, new_n15068_, new_n15069_, new_n15070_,
    new_n15071_, new_n15072_, new_n15073_, new_n15074_, new_n15075_,
    new_n15076_, new_n15077_, new_n15078_, new_n15079_, new_n15080_,
    new_n15081_, new_n15082_, new_n15083_, new_n15084_, new_n15085_,
    new_n15086_, new_n15087_, new_n15088_, new_n15089_, new_n15090_,
    new_n15091_, new_n15092_, new_n15093_, new_n15094_, new_n15095_,
    new_n15096_, new_n15097_, new_n15098_, new_n15099_, new_n15100_,
    new_n15101_, new_n15102_, new_n15103_, new_n15104_, new_n15105_,
    new_n15106_, new_n15107_, new_n15108_, new_n15109_, new_n15110_,
    new_n15111_, new_n15112_, new_n15113_, new_n15114_, new_n15115_,
    new_n15116_, new_n15117_, new_n15118_, new_n15119_, new_n15120_,
    new_n15121_, new_n15122_, new_n15123_, new_n15124_, new_n15125_,
    new_n15126_, new_n15127_, new_n15128_, new_n15129_, new_n15130_,
    new_n15131_, new_n15132_, new_n15133_, new_n15134_, new_n15135_,
    new_n15136_, new_n15137_, new_n15138_, new_n15139_, new_n15140_,
    new_n15141_, new_n15142_, new_n15143_, new_n15144_, new_n15145_,
    new_n15146_, new_n15147_, new_n15148_, new_n15149_, new_n15150_,
    new_n15151_, new_n15152_, new_n15153_, new_n15154_, new_n15155_,
    new_n15156_, new_n15157_, new_n15158_, new_n15159_, new_n15160_,
    new_n15161_, new_n15162_, new_n15163_, new_n15164_, new_n15165_,
    new_n15166_, new_n15167_, new_n15168_, new_n15169_, new_n15170_,
    new_n15171_, new_n15172_, new_n15173_, new_n15174_, new_n15175_,
    new_n15176_, new_n15177_, new_n15178_, new_n15179_, new_n15180_,
    new_n15181_, new_n15182_, new_n15183_, new_n15184_, new_n15185_,
    new_n15186_, new_n15187_, new_n15188_, new_n15189_, new_n15190_,
    new_n15191_, new_n15192_, new_n15193_, new_n15194_, new_n15195_,
    new_n15196_, new_n15197_, new_n15198_, new_n15199_, new_n15200_,
    new_n15201_, new_n15202_, new_n15203_, new_n15204_, new_n15205_,
    new_n15206_, new_n15207_, new_n15208_, new_n15209_, new_n15210_,
    new_n15211_, new_n15212_, new_n15213_, new_n15214_, new_n15215_,
    new_n15216_, new_n15217_, new_n15218_, new_n15219_, new_n15220_,
    new_n15221_, new_n15222_, new_n15223_, new_n15224_, new_n15225_,
    new_n15226_, new_n15227_, new_n15228_, new_n15229_, new_n15230_,
    new_n15231_, new_n15232_, new_n15233_, new_n15234_, new_n15235_,
    new_n15236_, new_n15237_, new_n15238_, new_n15239_, new_n15240_,
    new_n15241_, new_n15242_, new_n15243_, new_n15244_, new_n15245_,
    new_n15246_, new_n15247_, new_n15248_, new_n15249_, new_n15250_,
    new_n15251_, new_n15252_, new_n15253_, new_n15254_, new_n15255_,
    new_n15256_, new_n15257_, new_n15258_, new_n15259_, new_n15260_,
    new_n15261_, new_n15262_, new_n15263_, new_n15264_, new_n15265_,
    new_n15266_, new_n15267_, new_n15268_, new_n15269_, new_n15270_,
    new_n15271_, new_n15272_, new_n15273_, new_n15274_, new_n15275_,
    new_n15276_, new_n15277_, new_n15278_, new_n15279_, new_n15280_,
    new_n15281_, new_n15282_, new_n15283_, new_n15284_, new_n15285_,
    new_n15286_, new_n15287_, new_n15288_, new_n15289_, new_n15290_,
    new_n15291_, new_n15292_, new_n15293_, new_n15294_, new_n15295_,
    new_n15296_, new_n15297_, new_n15298_, new_n15299_, new_n15300_,
    new_n15301_, new_n15302_, new_n15303_, new_n15304_, new_n15305_,
    new_n15306_, new_n15307_, new_n15308_, new_n15309_, new_n15310_,
    new_n15311_, new_n15312_, new_n15313_, new_n15314_, new_n15315_,
    new_n15316_, new_n15317_, new_n15318_, new_n15319_, new_n15320_,
    new_n15321_, new_n15322_, new_n15323_, new_n15324_, new_n15325_,
    new_n15326_, new_n15327_, new_n15328_, new_n15329_, new_n15330_,
    new_n15331_, new_n15332_, new_n15333_, new_n15334_, new_n15335_,
    new_n15336_, new_n15337_, new_n15338_, new_n15339_, new_n15340_,
    new_n15341_, new_n15342_, new_n15343_, new_n15344_, new_n15345_,
    new_n15346_, new_n15347_, new_n15348_, new_n15349_, new_n15350_,
    new_n15351_, new_n15352_, new_n15353_, new_n15354_, new_n15355_,
    new_n15356_, new_n15357_, new_n15358_, new_n15359_, new_n15360_,
    new_n15361_, new_n15362_, new_n15363_, new_n15364_, new_n15365_,
    new_n15366_, new_n15367_, new_n15368_, new_n15369_, new_n15370_,
    new_n15371_, new_n15372_, new_n15373_, new_n15374_, new_n15375_,
    new_n15376_, new_n15377_, new_n15378_, new_n15379_, new_n15380_,
    new_n15381_, new_n15382_, new_n15383_, new_n15384_, new_n15385_,
    new_n15386_, new_n15387_, new_n15388_, new_n15389_, new_n15390_,
    new_n15391_, new_n15392_, new_n15393_, new_n15394_, new_n15395_,
    new_n15396_, new_n15397_, new_n15398_, new_n15399_, new_n15400_,
    new_n15401_, new_n15402_, new_n15403_, new_n15404_, new_n15405_,
    new_n15406_, new_n15407_, new_n15408_, new_n15409_, new_n15410_,
    new_n15411_, new_n15412_, new_n15413_, new_n15414_, new_n15415_,
    new_n15416_, new_n15417_, new_n15418_, new_n15419_, new_n15420_,
    new_n15421_, new_n15422_, new_n15423_, new_n15424_, new_n15425_,
    new_n15426_, new_n15427_, new_n15428_, new_n15429_, new_n15430_,
    new_n15431_, new_n15432_, new_n15433_, new_n15434_, new_n15435_,
    new_n15436_, new_n15437_, new_n15438_, new_n15439_, new_n15440_,
    new_n15441_, new_n15442_, new_n15443_, new_n15444_, new_n15445_,
    new_n15446_, new_n15447_, new_n15448_, new_n15449_, new_n15450_,
    new_n15451_, new_n15452_, new_n15453_, new_n15454_, new_n15455_,
    new_n15456_, new_n15457_, new_n15458_, new_n15459_, new_n15460_,
    new_n15461_, new_n15462_, new_n15463_, new_n15464_, new_n15465_,
    new_n15466_, new_n15467_, new_n15468_, new_n15469_, new_n15470_,
    new_n15471_, new_n15472_, new_n15473_, new_n15474_, new_n15475_,
    new_n15476_, new_n15477_, new_n15478_, new_n15479_, new_n15480_,
    new_n15481_, new_n15482_, new_n15483_, new_n15484_, new_n15485_,
    new_n15486_, new_n15487_, new_n15488_, new_n15489_, new_n15490_,
    new_n15491_, new_n15492_, new_n15493_, new_n15494_, new_n15495_,
    new_n15496_, new_n15497_, new_n15498_, new_n15499_, new_n15500_,
    new_n15501_, new_n15502_, new_n15503_, new_n15504_, new_n15505_,
    new_n15506_, new_n15507_, new_n15508_, new_n15509_, new_n15510_,
    new_n15511_, new_n15512_, new_n15513_, new_n15514_, new_n15515_,
    new_n15516_, new_n15517_, new_n15518_, new_n15519_, new_n15520_,
    new_n15521_, new_n15522_, new_n15523_, new_n15524_, new_n15525_,
    new_n15526_, new_n15527_, new_n15528_, new_n15529_, new_n15530_,
    new_n15531_, new_n15532_, new_n15533_, new_n15534_, new_n15535_,
    new_n15536_, new_n15537_, new_n15538_, new_n15539_, new_n15540_,
    new_n15541_, new_n15542_, new_n15543_, new_n15544_, new_n15545_,
    new_n15546_, new_n15547_, new_n15548_, new_n15549_, new_n15550_,
    new_n15551_, new_n15552_, new_n15553_, new_n15554_, new_n15555_,
    new_n15556_, new_n15557_, new_n15558_, new_n15559_, new_n15560_,
    new_n15561_, new_n15562_, new_n15563_, new_n15564_, new_n15565_,
    new_n15566_, new_n15567_, new_n15568_, new_n15569_, new_n15570_,
    new_n15571_, new_n15572_, new_n15573_, new_n15574_, new_n15575_,
    new_n15576_, new_n15577_, new_n15578_, new_n15579_, new_n15580_,
    new_n15581_, new_n15582_, new_n15583_, new_n15584_, new_n15585_,
    new_n15586_, new_n15587_, new_n15588_, new_n15589_, new_n15590_,
    new_n15591_, new_n15592_, new_n15593_, new_n15594_, new_n15595_,
    new_n15596_, new_n15597_, new_n15598_, new_n15599_, new_n15600_,
    new_n15601_, new_n15602_, new_n15603_, new_n15604_, new_n15605_,
    new_n15606_, new_n15607_, new_n15608_, new_n15609_, new_n15610_,
    new_n15611_, new_n15612_, new_n15613_, new_n15614_, new_n15615_,
    new_n15616_, new_n15617_, new_n15618_, new_n15619_, new_n15620_,
    new_n15621_, new_n15622_, new_n15623_, new_n15624_, new_n15625_,
    new_n15626_, new_n15627_, new_n15628_, new_n15629_, new_n15630_,
    new_n15631_, new_n15632_, new_n15633_, new_n15634_, new_n15635_,
    new_n15636_, new_n15637_, new_n15638_, new_n15639_, new_n15640_,
    new_n15641_, new_n15642_, new_n15643_, new_n15644_, new_n15645_,
    new_n15646_, new_n15647_, new_n15648_, new_n15649_, new_n15650_,
    new_n15651_, new_n15652_, new_n15653_, new_n15654_, new_n15655_,
    new_n15656_, new_n15657_, new_n15658_, new_n15659_, new_n15660_,
    new_n15661_, new_n15662_, new_n15663_, new_n15664_, new_n15665_,
    new_n15666_, new_n15667_, new_n15668_, new_n15669_, new_n15670_,
    new_n15671_, new_n15672_, new_n15673_, new_n15674_, new_n15675_,
    new_n15676_, new_n15677_, new_n15678_, new_n15679_, new_n15680_,
    new_n15681_, new_n15682_, new_n15683_, new_n15684_, new_n15685_,
    new_n15686_, new_n15687_, new_n15688_, new_n15689_, new_n15690_,
    new_n15691_, new_n15692_, new_n15693_, new_n15694_, new_n15695_,
    new_n15696_, new_n15697_, new_n15698_, new_n15699_, new_n15700_,
    new_n15701_, new_n15702_, new_n15703_, new_n15704_, new_n15705_,
    new_n15706_, new_n15707_, new_n15708_, new_n15709_, new_n15710_,
    new_n15711_, new_n15712_, new_n15713_, new_n15714_, new_n15715_,
    new_n15716_, new_n15717_, new_n15718_, new_n15719_, new_n15720_,
    new_n15721_, new_n15722_, new_n15723_, new_n15724_, new_n15725_,
    new_n15726_, new_n15727_, new_n15728_, new_n15729_, new_n15730_,
    new_n15731_, new_n15732_, new_n15733_, new_n15734_, new_n15735_,
    new_n15736_, new_n15737_, new_n15738_, new_n15739_, new_n15740_,
    new_n15741_, new_n15742_, new_n15743_, new_n15744_, new_n15745_,
    new_n15746_, new_n15747_, new_n15748_, new_n15749_, new_n15750_,
    new_n15751_, new_n15752_, new_n15753_, new_n15754_, new_n15755_,
    new_n15756_, new_n15757_, new_n15758_, new_n15759_, new_n15760_,
    new_n15761_, new_n15762_, new_n15763_, new_n15764_, new_n15765_,
    new_n15766_, new_n15767_, new_n15768_, new_n15769_, new_n15770_,
    new_n15771_, new_n15772_, new_n15773_, new_n15774_, new_n15775_,
    new_n15776_, new_n15777_, new_n15778_, new_n15779_, new_n15780_,
    new_n15781_, new_n15782_, new_n15783_, new_n15784_, new_n15785_,
    new_n15786_, new_n15787_, new_n15788_, new_n15789_, new_n15790_,
    new_n15791_, new_n15792_, new_n15793_, new_n15794_, new_n15795_,
    new_n15796_, new_n15797_, new_n15798_, new_n15799_, new_n15800_,
    new_n15801_, new_n15802_, new_n15803_, new_n15804_, new_n15805_,
    new_n15806_, new_n15807_, new_n15808_, new_n15809_, new_n15810_,
    new_n15811_, new_n15812_, new_n15813_, new_n15814_, new_n15815_,
    new_n15816_, new_n15817_, new_n15818_, new_n15819_, new_n15820_,
    new_n15821_, new_n15822_, new_n15823_, new_n15824_, new_n15825_,
    new_n15826_, new_n15827_, new_n15828_, new_n15829_, new_n15830_,
    new_n15831_, new_n15832_, new_n15833_, new_n15834_, new_n15835_,
    new_n15836_, new_n15837_, new_n15838_, new_n15839_, new_n15840_,
    new_n15841_, new_n15842_, new_n15843_, new_n15844_, new_n15845_,
    new_n15846_, new_n15847_, new_n15848_, new_n15849_, new_n15850_,
    new_n15851_, new_n15852_, new_n15853_, new_n15854_, new_n15855_,
    new_n15856_, new_n15857_, new_n15858_, new_n15859_, new_n15860_,
    new_n15861_, new_n15862_, new_n15863_, new_n15864_, new_n15865_,
    new_n15866_, new_n15867_, new_n15868_, new_n15869_, new_n15870_,
    new_n15871_, new_n15872_, new_n15873_, new_n15874_, new_n15875_,
    new_n15876_, new_n15877_, new_n15878_, new_n15879_, new_n15880_,
    new_n15881_, new_n15882_, new_n15883_, new_n15884_, new_n15885_,
    new_n15886_, new_n15887_, new_n15888_, new_n15889_, new_n15890_,
    new_n15891_, new_n15892_, new_n15893_, new_n15894_, new_n15895_,
    new_n15896_, new_n15897_, new_n15898_, new_n15899_, new_n15900_,
    new_n15901_, new_n15902_, new_n15903_, new_n15904_, new_n15905_,
    new_n15906_, new_n15907_, new_n15908_, new_n15909_, new_n15910_,
    new_n15911_, new_n15912_, new_n15913_, new_n15914_, new_n15915_,
    new_n15916_, new_n15917_, new_n15918_, new_n15919_, new_n15920_,
    new_n15921_, new_n15922_, new_n15923_, new_n15924_, new_n15925_,
    new_n15926_, new_n15927_, new_n15928_, new_n15929_, new_n15930_,
    new_n15931_, new_n15932_, new_n15933_, new_n15934_, new_n15935_,
    new_n15936_, new_n15937_, new_n15938_, new_n15939_, new_n15940_,
    new_n15941_, new_n15942_, new_n15943_, new_n15944_, new_n15945_,
    new_n15946_, new_n15947_, new_n15948_, new_n15949_, new_n15950_,
    new_n15951_, new_n15952_, new_n15953_, new_n15954_, new_n15955_,
    new_n15956_, new_n15957_, new_n15958_, new_n15959_, new_n15960_,
    new_n15961_, new_n15962_, new_n15963_, new_n15964_, new_n15965_,
    new_n15966_, new_n15967_, new_n15968_, new_n15969_, new_n15970_,
    new_n15971_, new_n15972_, new_n15973_, new_n15974_, new_n15975_,
    new_n15976_, new_n15977_, new_n15978_, new_n15979_, new_n15980_,
    new_n15981_, new_n15982_, new_n15983_, new_n15984_, new_n15985_,
    new_n15986_, new_n15987_, new_n15988_, new_n15989_, new_n15990_,
    new_n15991_, new_n15992_, new_n15993_, new_n15994_, new_n15995_,
    new_n15996_, new_n15997_, new_n15998_, new_n15999_, new_n16000_,
    new_n16001_, new_n16002_, new_n16003_, new_n16004_, new_n16005_,
    new_n16006_, new_n16007_, new_n16008_, new_n16009_, new_n16010_,
    new_n16011_, new_n16012_, new_n16013_, new_n16014_, new_n16015_,
    new_n16016_, new_n16017_, new_n16018_, new_n16019_, new_n16020_,
    new_n16021_, new_n16022_, new_n16023_, new_n16024_, new_n16025_,
    new_n16026_, new_n16027_, new_n16028_, new_n16029_, new_n16030_,
    new_n16031_, new_n16032_, new_n16033_, new_n16034_, new_n16035_,
    new_n16036_, new_n16037_, new_n16038_, new_n16039_, new_n16040_,
    new_n16041_, new_n16042_, new_n16043_, new_n16044_, new_n16045_,
    new_n16046_, new_n16047_, new_n16048_, new_n16049_, new_n16050_,
    new_n16051_, new_n16052_, new_n16053_, new_n16054_, new_n16055_,
    new_n16056_, new_n16057_, new_n16058_, new_n16059_, new_n16060_,
    new_n16061_, new_n16062_, new_n16063_, new_n16064_, new_n16065_,
    new_n16066_, new_n16067_, new_n16068_, new_n16069_, new_n16070_,
    new_n16071_, new_n16072_, new_n16073_, new_n16074_, new_n16075_,
    new_n16076_, new_n16077_, new_n16078_, new_n16079_, new_n16080_,
    new_n16081_, new_n16082_, new_n16083_, new_n16084_, new_n16085_,
    new_n16086_, new_n16087_, new_n16088_, new_n16089_, new_n16090_,
    new_n16091_, new_n16092_, new_n16093_, new_n16094_, new_n16095_,
    new_n16096_, new_n16097_, new_n16098_, new_n16099_, new_n16100_,
    new_n16101_, new_n16102_, new_n16103_, new_n16104_, new_n16105_,
    new_n16106_, new_n16107_, new_n16108_, new_n16109_, new_n16110_,
    new_n16111_, new_n16112_, new_n16113_, new_n16114_, new_n16115_,
    new_n16116_, new_n16117_, new_n16118_, new_n16119_, new_n16120_,
    new_n16121_, new_n16122_, new_n16123_, new_n16124_, new_n16125_,
    new_n16126_, new_n16127_, new_n16128_, new_n16129_, new_n16130_,
    new_n16131_, new_n16132_, new_n16133_, new_n16134_, new_n16135_,
    new_n16136_, new_n16137_, new_n16138_, new_n16139_, new_n16140_,
    new_n16141_, new_n16142_, new_n16143_, new_n16144_, new_n16145_,
    new_n16146_, new_n16147_, new_n16148_, new_n16149_, new_n16150_,
    new_n16151_, new_n16152_, new_n16153_, new_n16154_, new_n16155_,
    new_n16156_, new_n16157_, new_n16158_, new_n16159_, new_n16160_,
    new_n16161_, new_n16162_, new_n16163_, new_n16164_, new_n16165_,
    new_n16166_, new_n16167_, new_n16168_, new_n16169_, new_n16170_,
    new_n16171_, new_n16172_, new_n16173_, new_n16174_, new_n16175_,
    new_n16176_, new_n16177_, new_n16178_, new_n16179_, new_n16180_,
    new_n16181_, new_n16182_, new_n16183_, new_n16184_, new_n16185_,
    new_n16186_, new_n16187_, new_n16188_, new_n16189_, new_n16190_,
    new_n16191_, new_n16192_, new_n16193_, new_n16194_, new_n16195_,
    new_n16196_, new_n16197_, new_n16198_, new_n16199_, new_n16200_,
    new_n16201_, new_n16202_, new_n16203_, new_n16204_, new_n16205_,
    new_n16206_, new_n16207_, new_n16208_, new_n16209_, new_n16210_,
    new_n16211_, new_n16212_, new_n16213_, new_n16214_, new_n16215_,
    new_n16216_, new_n16217_, new_n16218_, new_n16219_, new_n16220_,
    new_n16221_, new_n16222_, new_n16223_, new_n16224_, new_n16225_,
    new_n16226_, new_n16227_, new_n16228_, new_n16229_, new_n16230_,
    new_n16231_, new_n16232_, new_n16233_, new_n16234_, new_n16235_,
    new_n16236_, new_n16237_, new_n16238_, new_n16239_, new_n16240_,
    new_n16241_, new_n16242_, new_n16243_, new_n16244_, new_n16245_,
    new_n16246_, new_n16247_, new_n16248_, new_n16249_, new_n16250_,
    new_n16251_, new_n16252_, new_n16253_, new_n16254_, new_n16255_,
    new_n16256_, new_n16257_, new_n16258_, new_n16259_, new_n16260_,
    new_n16261_, new_n16262_, new_n16263_, new_n16264_, new_n16265_,
    new_n16266_, new_n16267_, new_n16268_, new_n16269_, new_n16270_,
    new_n16271_, new_n16272_, new_n16273_, new_n16274_, new_n16275_,
    new_n16276_, new_n16277_, new_n16278_, new_n16279_, new_n16280_,
    new_n16281_, new_n16282_, new_n16283_, new_n16284_, new_n16285_,
    new_n16286_, new_n16287_, new_n16288_, new_n16289_, new_n16290_,
    new_n16291_, new_n16292_, new_n16293_, new_n16294_, new_n16295_,
    new_n16296_, new_n16297_, new_n16298_, new_n16299_, new_n16300_,
    new_n16301_, new_n16302_, new_n16303_, new_n16304_, new_n16305_,
    new_n16306_, new_n16307_, new_n16308_, new_n16309_, new_n16310_,
    new_n16311_, new_n16312_, new_n16313_, new_n16314_, new_n16315_,
    new_n16316_, new_n16317_, new_n16318_, new_n16319_, new_n16320_,
    new_n16321_, new_n16322_, new_n16323_, new_n16324_, new_n16325_,
    new_n16326_, new_n16327_, new_n16328_, new_n16329_, new_n16330_,
    new_n16331_, new_n16332_, new_n16333_, new_n16334_, new_n16335_,
    new_n16336_, new_n16337_, new_n16338_, new_n16339_, new_n16340_,
    new_n16341_, new_n16342_, new_n16343_, new_n16344_, new_n16345_,
    new_n16346_, new_n16347_, new_n16348_, new_n16349_, new_n16350_,
    new_n16351_, new_n16352_, new_n16353_, new_n16354_, new_n16355_,
    new_n16356_, new_n16357_, new_n16358_, new_n16359_, new_n16360_,
    new_n16361_, new_n16362_, new_n16363_, new_n16364_, new_n16365_,
    new_n16366_, new_n16367_, new_n16368_, new_n16369_, new_n16370_,
    new_n16371_, new_n16372_, new_n16373_, new_n16374_, new_n16375_,
    new_n16376_, new_n16377_, new_n16378_, new_n16379_, new_n16380_,
    new_n16381_, new_n16382_, new_n16383_, new_n16384_, new_n16385_,
    new_n16386_, new_n16387_, new_n16388_, new_n16389_, new_n16390_,
    new_n16391_, new_n16392_, new_n16393_, new_n16394_, new_n16395_,
    new_n16396_, new_n16397_, new_n16398_, new_n16399_, new_n16400_,
    new_n16401_, new_n16402_, new_n16403_, new_n16404_, new_n16405_,
    new_n16406_, new_n16407_, new_n16408_, new_n16409_, new_n16410_,
    new_n16411_, new_n16412_, new_n16413_, new_n16414_, new_n16415_,
    new_n16416_, new_n16417_, new_n16418_, new_n16419_, new_n16420_,
    new_n16421_, new_n16422_, new_n16423_, new_n16424_, new_n16425_,
    new_n16426_, new_n16427_, new_n16428_, new_n16429_, new_n16430_,
    new_n16431_, new_n16432_, new_n16433_, new_n16434_, new_n16435_,
    new_n16436_, new_n16437_, new_n16438_, new_n16439_, new_n16440_,
    new_n16441_, new_n16442_, new_n16443_, new_n16444_, new_n16445_,
    new_n16446_, new_n16447_, new_n16448_, new_n16449_, new_n16450_,
    new_n16451_, new_n16452_, new_n16453_, new_n16454_, new_n16455_,
    new_n16456_, new_n16457_, new_n16458_, new_n16459_, new_n16460_,
    new_n16461_, new_n16462_, new_n16463_, new_n16464_, new_n16465_,
    new_n16466_, new_n16467_, new_n16468_, new_n16469_, new_n16470_,
    new_n16471_, new_n16472_, new_n16473_, new_n16474_, new_n16475_,
    new_n16476_, new_n16477_, new_n16478_, new_n16479_, new_n16480_,
    new_n16481_, new_n16482_, new_n16483_, new_n16484_, new_n16485_,
    new_n16486_, new_n16487_, new_n16488_, new_n16489_, new_n16490_,
    new_n16491_, new_n16492_, new_n16493_, new_n16494_, new_n16495_,
    new_n16496_, new_n16497_, new_n16498_, new_n16499_, new_n16500_,
    new_n16501_, new_n16502_, new_n16503_, new_n16504_, new_n16505_,
    new_n16506_, new_n16507_, new_n16508_, new_n16509_, new_n16510_,
    new_n16511_, new_n16512_, new_n16513_, new_n16514_, new_n16515_,
    new_n16516_, new_n16517_, new_n16518_, new_n16519_, new_n16520_,
    new_n16521_, new_n16522_, new_n16523_, new_n16524_, new_n16525_,
    new_n16526_, new_n16527_, new_n16528_, new_n16529_, new_n16530_,
    new_n16531_, new_n16532_, new_n16533_, new_n16534_, new_n16535_,
    new_n16536_, new_n16537_, new_n16538_, new_n16539_, new_n16540_,
    new_n16541_, new_n16542_, new_n16543_, new_n16544_, new_n16545_,
    new_n16546_, new_n16547_, new_n16548_, new_n16549_, new_n16550_,
    new_n16551_, new_n16552_, new_n16553_, new_n16554_, new_n16555_,
    new_n16556_, new_n16557_, new_n16558_, new_n16559_, new_n16560_,
    new_n16561_, new_n16562_, new_n16563_, new_n16564_, new_n16565_,
    new_n16566_, new_n16567_, new_n16568_, new_n16569_, new_n16570_,
    new_n16571_, new_n16572_, new_n16573_, new_n16574_, new_n16575_,
    new_n16576_, new_n16577_, new_n16578_, new_n16579_, new_n16580_,
    new_n16581_, new_n16582_, new_n16583_, new_n16584_, new_n16585_,
    new_n16586_, new_n16587_, new_n16588_, new_n16589_, new_n16590_,
    new_n16591_, new_n16592_, new_n16593_, new_n16594_, new_n16595_,
    new_n16596_, new_n16597_, new_n16598_, new_n16599_, new_n16600_,
    new_n16601_, new_n16602_, new_n16603_, new_n16604_, new_n16605_,
    new_n16606_, new_n16607_, new_n16608_, new_n16609_, new_n16610_,
    new_n16611_, new_n16612_, new_n16613_, new_n16614_, new_n16615_,
    new_n16616_, new_n16617_, new_n16618_, new_n16619_, new_n16620_,
    new_n16621_, new_n16622_, new_n16623_, new_n16624_, new_n16625_,
    new_n16626_, new_n16627_, new_n16628_, new_n16629_, new_n16630_,
    new_n16631_, new_n16632_, new_n16633_, new_n16634_, new_n16635_,
    new_n16636_, new_n16637_, new_n16638_, new_n16639_, new_n16640_,
    new_n16641_, new_n16642_, new_n16643_, new_n16644_, new_n16645_,
    new_n16646_, new_n16647_, new_n16648_, new_n16649_, new_n16650_,
    new_n16651_, new_n16652_, new_n16653_, new_n16654_, new_n16655_,
    new_n16656_, new_n16657_, new_n16658_, new_n16659_, new_n16660_,
    new_n16661_, new_n16662_, new_n16663_, new_n16664_, new_n16665_,
    new_n16666_, new_n16667_, new_n16668_, new_n16669_, new_n16670_,
    new_n16671_, new_n16672_, new_n16673_, new_n16674_, new_n16675_,
    new_n16676_, new_n16677_, new_n16678_, new_n16679_, new_n16680_,
    new_n16681_, new_n16682_, new_n16683_, new_n16684_, new_n16685_,
    new_n16686_, new_n16687_, new_n16688_, new_n16689_, new_n16690_,
    new_n16691_, new_n16692_, new_n16693_, new_n16694_, new_n16695_,
    new_n16696_, new_n16697_, new_n16698_, new_n16699_, new_n16700_,
    new_n16701_, new_n16702_, new_n16703_, new_n16704_, new_n16705_,
    new_n16706_, new_n16707_, new_n16708_, new_n16709_, new_n16710_,
    new_n16711_, new_n16712_, new_n16713_, new_n16714_, new_n16715_,
    new_n16716_, new_n16717_, new_n16718_, new_n16719_, new_n16720_,
    new_n16721_, new_n16722_, new_n16723_, new_n16724_, new_n16725_,
    new_n16726_, new_n16727_, new_n16728_, new_n16729_, new_n16730_,
    new_n16731_, new_n16732_, new_n16733_, new_n16734_, new_n16735_,
    new_n16736_, new_n16737_, new_n16738_, new_n16739_, new_n16740_,
    new_n16741_, new_n16742_, new_n16743_, new_n16744_, new_n16745_,
    new_n16746_, new_n16747_, new_n16748_, new_n16749_, new_n16750_,
    new_n16751_, new_n16752_, new_n16753_, new_n16754_, new_n16755_,
    new_n16756_, new_n16757_, new_n16758_, new_n16759_, new_n16760_,
    new_n16761_, new_n16762_, new_n16763_, new_n16764_, new_n16765_,
    new_n16766_, new_n16767_, new_n16768_, new_n16769_, new_n16770_,
    new_n16771_, new_n16772_, new_n16773_, new_n16774_, new_n16775_,
    new_n16776_, new_n16777_, new_n16778_, new_n16779_, new_n16780_,
    new_n16781_, new_n16782_, new_n16783_, new_n16784_, new_n16785_,
    new_n16786_, new_n16787_, new_n16788_, new_n16789_, new_n16790_,
    new_n16791_, new_n16792_, new_n16793_, new_n16794_, new_n16795_,
    new_n16796_, new_n16797_, new_n16798_, new_n16799_, new_n16800_,
    new_n16801_, new_n16802_, new_n16803_, new_n16804_, new_n16805_,
    new_n16806_, new_n16807_, new_n16808_, new_n16809_, new_n16810_,
    new_n16811_, new_n16812_, new_n16813_, new_n16814_, new_n16815_,
    new_n16816_, new_n16817_, new_n16818_, new_n16819_, new_n16820_,
    new_n16821_, new_n16822_, new_n16823_, new_n16824_, new_n16825_,
    new_n16826_, new_n16827_, new_n16828_, new_n16829_, new_n16830_,
    new_n16831_, new_n16832_, new_n16833_, new_n16834_, new_n16835_,
    new_n16836_, new_n16837_, new_n16838_, new_n16839_, new_n16840_,
    new_n16841_, new_n16842_, new_n16843_, new_n16844_, new_n16845_,
    new_n16846_, new_n16847_, new_n16848_, new_n16849_, new_n16850_,
    new_n16851_, new_n16852_, new_n16853_, new_n16854_, new_n16855_,
    new_n16856_, new_n16857_, new_n16858_, new_n16859_, new_n16860_,
    new_n16861_, new_n16862_, new_n16863_, new_n16864_, new_n16865_,
    new_n16866_, new_n16867_, new_n16868_, new_n16869_, new_n16870_,
    new_n16871_, new_n16872_, new_n16873_, new_n16874_, new_n16875_,
    new_n16876_, new_n16877_, new_n16878_, new_n16879_, new_n16880_,
    new_n16881_, new_n16882_, new_n16883_, new_n16884_, new_n16885_,
    new_n16886_, new_n16887_, new_n16888_, new_n16889_, new_n16890_,
    new_n16891_, new_n16892_, new_n16893_, new_n16894_, new_n16895_,
    new_n16896_, new_n16897_, new_n16898_, new_n16899_, new_n16900_,
    new_n16901_, new_n16902_, new_n16903_, new_n16904_, new_n16905_,
    new_n16906_, new_n16907_, new_n16908_, new_n16909_, new_n16910_,
    new_n16911_, new_n16912_, new_n16913_, new_n16914_, new_n16915_,
    new_n16916_, new_n16917_, new_n16918_, new_n16919_, new_n16920_,
    new_n16921_, new_n16922_, new_n16923_, new_n16924_, new_n16925_,
    new_n16926_, new_n16927_, new_n16928_, new_n16929_, new_n16930_,
    new_n16931_, new_n16932_, new_n16933_, new_n16934_, new_n16935_,
    new_n16936_, new_n16937_, new_n16938_, new_n16939_, new_n16940_,
    new_n16941_, new_n16942_, new_n16943_, new_n16944_, new_n16945_,
    new_n16946_, new_n16947_, new_n16948_, new_n16949_, new_n16950_,
    new_n16951_, new_n16952_, new_n16953_, new_n16954_, new_n16955_,
    new_n16956_, new_n16957_, new_n16958_, new_n16959_, new_n16960_,
    new_n16961_, new_n16962_, new_n16963_, new_n16964_, new_n16965_,
    new_n16966_, new_n16967_, new_n16968_, new_n16969_, new_n16970_,
    new_n16971_, new_n16972_, new_n16973_, new_n16974_, new_n16975_,
    new_n16976_, new_n16977_, new_n16978_, new_n16979_, new_n16980_,
    new_n16981_, new_n16982_, new_n16983_, new_n16984_, new_n16985_,
    new_n16986_, new_n16987_, new_n16988_, new_n16989_, new_n16990_,
    new_n16991_, new_n16992_, new_n16993_, new_n16994_, new_n16995_,
    new_n16996_, new_n16997_, new_n16998_, new_n16999_, new_n17000_,
    new_n17001_, new_n17002_, new_n17003_, new_n17004_, new_n17005_,
    new_n17006_, new_n17007_, new_n17008_, new_n17009_, new_n17010_,
    new_n17011_, new_n17012_, new_n17013_, new_n17014_, new_n17015_,
    new_n17016_, new_n17017_, new_n17018_, new_n17019_, new_n17020_,
    new_n17021_, new_n17022_, new_n17023_, new_n17024_, new_n17025_,
    new_n17026_, new_n17027_, new_n17028_, new_n17029_, new_n17030_,
    new_n17031_, new_n17032_, new_n17033_, new_n17034_, new_n17035_,
    new_n17036_, new_n17037_, new_n17038_, new_n17039_, new_n17040_,
    new_n17041_, new_n17042_, new_n17043_, new_n17044_, new_n17045_,
    new_n17046_, new_n17047_, new_n17048_, new_n17049_, new_n17050_,
    new_n17051_, new_n17052_, new_n17053_, new_n17054_, new_n17055_,
    new_n17056_, new_n17057_, new_n17058_, new_n17059_, new_n17060_,
    new_n17061_, new_n17062_, new_n17063_, new_n17064_, new_n17065_,
    new_n17066_, new_n17067_, new_n17068_, new_n17069_, new_n17070_,
    new_n17071_, new_n17072_, new_n17073_, new_n17074_, new_n17075_,
    new_n17076_, new_n17077_, new_n17078_, new_n17079_, new_n17080_,
    new_n17081_, new_n17082_, new_n17083_, new_n17084_, new_n17085_,
    new_n17086_, new_n17087_, new_n17088_, new_n17089_, new_n17090_,
    new_n17091_, new_n17092_, new_n17093_, new_n17094_, new_n17095_,
    new_n17096_, new_n17097_, new_n17098_, new_n17099_, new_n17100_,
    new_n17101_, new_n17102_, new_n17103_, new_n17104_, new_n17105_,
    new_n17106_, new_n17107_, new_n17108_, new_n17109_, new_n17110_,
    new_n17111_, new_n17112_, new_n17113_, new_n17114_, new_n17115_,
    new_n17116_, new_n17117_, new_n17118_, new_n17119_, new_n17120_,
    new_n17121_, new_n17122_, new_n17123_, new_n17124_, new_n17125_,
    new_n17126_, new_n17127_, new_n17128_, new_n17129_, new_n17130_,
    new_n17131_, new_n17132_, new_n17133_, new_n17134_, new_n17135_,
    new_n17136_, new_n17137_, new_n17138_, new_n17139_, new_n17140_,
    new_n17141_, new_n17142_, new_n17143_, new_n17144_, new_n17145_,
    new_n17146_, new_n17147_, new_n17148_, new_n17149_, new_n17150_,
    new_n17151_, new_n17152_, new_n17153_, new_n17154_, new_n17155_,
    new_n17156_, new_n17157_, new_n17158_, new_n17159_, new_n17160_,
    new_n17161_, new_n17162_, new_n17163_, new_n17164_, new_n17165_,
    new_n17166_, new_n17167_, new_n17168_, new_n17169_, new_n17170_,
    new_n17171_, new_n17172_, new_n17173_, new_n17174_, new_n17175_,
    new_n17176_, new_n17177_, new_n17178_, new_n17179_, new_n17180_,
    new_n17181_, new_n17182_, new_n17183_, new_n17184_, new_n17185_,
    new_n17186_, new_n17187_, new_n17188_, new_n17189_, new_n17190_,
    new_n17191_, new_n17192_, new_n17193_, new_n17194_, new_n17195_,
    new_n17196_, new_n17197_, new_n17198_, new_n17199_, new_n17200_,
    new_n17201_, new_n17202_, new_n17203_, new_n17204_, new_n17205_,
    new_n17206_, new_n17207_, new_n17208_, new_n17209_, new_n17210_,
    new_n17211_, new_n17212_, new_n17213_, new_n17214_, new_n17215_,
    new_n17216_, new_n17217_, new_n17218_, new_n17219_, new_n17220_,
    new_n17221_, new_n17222_, new_n17223_, new_n17224_, new_n17225_,
    new_n17226_, new_n17227_, new_n17228_, new_n17229_, new_n17230_,
    new_n17231_, new_n17232_, new_n17233_, new_n17234_, new_n17235_,
    new_n17236_, new_n17237_, new_n17238_, new_n17239_, new_n17240_,
    new_n17241_, new_n17242_, new_n17243_, new_n17244_, new_n17245_,
    new_n17246_, new_n17247_, new_n17248_, new_n17249_, new_n17250_,
    new_n17251_, new_n17252_, new_n17253_, new_n17254_, new_n17255_,
    new_n17256_, new_n17257_, new_n17258_, new_n17259_, new_n17260_,
    new_n17261_, new_n17262_, new_n17263_, new_n17264_, new_n17265_,
    new_n17266_, new_n17267_, new_n17268_, new_n17269_, new_n17270_,
    new_n17271_, new_n17272_, new_n17273_, new_n17274_, new_n17275_,
    new_n17276_, new_n17277_, new_n17278_, new_n17279_, new_n17280_,
    new_n17281_, new_n17282_, new_n17283_, new_n17284_, new_n17285_,
    new_n17286_, new_n17287_, new_n17288_, new_n17289_, new_n17290_,
    new_n17291_, new_n17292_, new_n17293_, new_n17294_, new_n17295_,
    new_n17296_, new_n17297_, new_n17298_, new_n17299_, new_n17300_,
    new_n17301_, new_n17302_, new_n17303_, new_n17304_, new_n17305_,
    new_n17306_, new_n17307_, new_n17308_, new_n17309_, new_n17310_,
    new_n17311_, new_n17312_, new_n17313_, new_n17314_, new_n17315_,
    new_n17316_, new_n17317_, new_n17318_, new_n17319_, new_n17320_,
    new_n17321_, new_n17322_, new_n17323_, new_n17324_, new_n17325_,
    new_n17326_, new_n17327_, new_n17328_, new_n17329_, new_n17330_,
    new_n17331_, new_n17332_, new_n17333_, new_n17334_, new_n17335_,
    new_n17336_, new_n17337_, new_n17338_, new_n17339_, new_n17340_,
    new_n17341_, new_n17342_, new_n17343_, new_n17344_, new_n17345_,
    new_n17346_, new_n17347_, new_n17348_, new_n17349_, new_n17350_,
    new_n17351_, new_n17352_, new_n17353_, new_n17354_, new_n17355_,
    new_n17356_, new_n17357_, new_n17358_, new_n17359_, new_n17360_,
    new_n17361_, new_n17362_, new_n17363_, new_n17364_, new_n17365_,
    new_n17366_, new_n17367_, new_n17368_, new_n17369_, new_n17370_,
    new_n17371_, new_n17372_, new_n17373_, new_n17374_, new_n17375_,
    new_n17376_, new_n17377_, new_n17378_, new_n17379_, new_n17380_,
    new_n17381_, new_n17382_, new_n17383_, new_n17384_, new_n17385_,
    new_n17386_, new_n17387_, new_n17388_, new_n17389_, new_n17390_,
    new_n17391_, new_n17392_, new_n17393_, new_n17394_, new_n17395_,
    new_n17396_, new_n17397_, new_n17398_, new_n17399_, new_n17400_,
    new_n17401_, new_n17402_, new_n17403_, new_n17404_, new_n17405_,
    new_n17406_, new_n17407_, new_n17408_, new_n17409_, new_n17410_,
    new_n17411_, new_n17412_, new_n17413_, new_n17414_, new_n17415_,
    new_n17416_, new_n17417_, new_n17418_, new_n17419_, new_n17420_,
    new_n17421_, new_n17422_, new_n17423_, new_n17424_, new_n17425_,
    new_n17426_, new_n17427_, new_n17428_, new_n17429_, new_n17430_,
    new_n17431_, new_n17432_, new_n17433_, new_n17434_, new_n17435_,
    new_n17436_, new_n17437_, new_n17438_, new_n17439_, new_n17440_,
    new_n17441_, new_n17442_, new_n17443_, new_n17444_, new_n17445_,
    new_n17446_, new_n17447_, new_n17448_, new_n17449_, new_n17450_,
    new_n17451_, new_n17452_, new_n17453_, new_n17454_, new_n17455_,
    new_n17456_, new_n17457_, new_n17458_, new_n17459_, new_n17460_,
    new_n17461_, new_n17462_, new_n17463_, new_n17464_, new_n17465_,
    new_n17466_, new_n17467_, new_n17468_, new_n17469_, new_n17470_,
    new_n17471_, new_n17472_, new_n17473_, new_n17474_, new_n17475_,
    new_n17476_, new_n17477_, new_n17478_, new_n17479_, new_n17480_,
    new_n17481_, new_n17482_, new_n17483_, new_n17484_, new_n17485_,
    new_n17486_, new_n17487_, new_n17488_, new_n17489_, new_n17490_,
    new_n17491_, new_n17492_, new_n17493_, new_n17494_, new_n17495_,
    new_n17496_, new_n17497_, new_n17498_, new_n17499_, new_n17500_,
    new_n17501_, new_n17502_, new_n17503_, new_n17504_, new_n17505_,
    new_n17506_, new_n17507_, new_n17508_, new_n17509_, new_n17510_,
    new_n17511_, new_n17512_, new_n17513_, new_n17514_, new_n17515_,
    new_n17516_, new_n17517_, new_n17518_, new_n17519_, new_n17520_,
    new_n17521_, new_n17522_, new_n17523_, new_n17524_, new_n17525_,
    new_n17526_, new_n17527_, new_n17528_, new_n17529_, new_n17530_,
    new_n17531_, new_n17532_, new_n17533_, new_n17534_, new_n17535_,
    new_n17536_, new_n17537_, new_n17538_, new_n17539_, new_n17540_,
    new_n17541_, new_n17542_, new_n17543_, new_n17544_, new_n17545_,
    new_n17546_, new_n17547_, new_n17548_, new_n17549_, new_n17550_,
    new_n17551_, new_n17552_, new_n17553_, new_n17554_, new_n17555_,
    new_n17556_, new_n17557_, new_n17558_, new_n17559_, new_n17560_,
    new_n17561_, new_n17562_, new_n17563_, new_n17564_, new_n17565_,
    new_n17566_, new_n17567_, new_n17568_, new_n17569_, new_n17570_,
    new_n17571_, new_n17572_, new_n17573_, new_n17574_, new_n17575_,
    new_n17576_, new_n17577_, new_n17578_, new_n17579_, new_n17580_,
    new_n17581_, new_n17582_, new_n17583_, new_n17584_, new_n17585_,
    new_n17586_, new_n17587_, new_n17588_, new_n17589_, new_n17590_,
    new_n17591_, new_n17592_, new_n17593_, new_n17594_, new_n17595_,
    new_n17596_, new_n17597_, new_n17598_, new_n17599_, new_n17600_,
    new_n17601_, new_n17602_, new_n17603_, new_n17604_, new_n17605_,
    new_n17606_, new_n17607_, new_n17608_, new_n17609_, new_n17610_,
    new_n17611_, new_n17612_, new_n17613_, new_n17614_, new_n17615_,
    new_n17616_, new_n17617_, new_n17618_, new_n17619_, new_n17620_,
    new_n17621_, new_n17622_, new_n17623_, new_n17624_, new_n17625_,
    new_n17626_, new_n17627_, new_n17628_, new_n17629_, new_n17630_,
    new_n17631_, new_n17632_, new_n17633_, new_n17634_, new_n17635_,
    new_n17636_, new_n17637_, new_n17638_, new_n17639_, new_n17640_,
    new_n17641_, new_n17642_, new_n17643_, new_n17644_, new_n17645_,
    new_n17646_, new_n17647_, new_n17648_, new_n17649_, new_n17650_,
    new_n17651_, new_n17652_, new_n17653_, new_n17654_, new_n17655_,
    new_n17656_, new_n17657_, new_n17658_, new_n17659_, new_n17660_,
    new_n17661_, new_n17662_, new_n17663_, new_n17664_, new_n17665_,
    new_n17666_, new_n17667_, new_n17668_, new_n17669_, new_n17670_,
    new_n17671_, new_n17672_, new_n17673_, new_n17674_, new_n17675_,
    new_n17676_, new_n17677_, new_n17678_, new_n17679_, new_n17680_,
    new_n17681_, new_n17682_, new_n17683_, new_n17684_, new_n17685_,
    new_n17686_, new_n17687_, new_n17688_, new_n17689_, new_n17690_,
    new_n17691_, new_n17692_, new_n17693_, new_n17694_, new_n17695_,
    new_n17696_, new_n17697_, new_n17698_, new_n17699_, new_n17700_,
    new_n17701_, new_n17702_, new_n17703_, new_n17704_, new_n17705_,
    new_n17706_, new_n17707_, new_n17708_, new_n17709_, new_n17710_,
    new_n17711_, new_n17712_, new_n17713_, new_n17714_, new_n17715_,
    new_n17716_, new_n17717_, new_n17718_, new_n17719_, new_n17720_,
    new_n17721_, new_n17722_, new_n17723_, new_n17724_, new_n17725_,
    new_n17726_, new_n17727_, new_n17728_, new_n17729_, new_n17730_,
    new_n17731_, new_n17732_, new_n17733_, new_n17734_, new_n17735_,
    new_n17736_, new_n17737_, new_n17738_, new_n17739_, new_n17740_,
    new_n17741_, new_n17742_, new_n17743_, new_n17744_, new_n17745_,
    new_n17746_, new_n17747_, new_n17748_, new_n17749_, new_n17750_,
    new_n17751_, new_n17752_, new_n17753_, new_n17754_, new_n17755_,
    new_n17756_, new_n17757_, new_n17758_, new_n17759_, new_n17760_,
    new_n17761_, new_n17762_, new_n17763_, new_n17764_, new_n17765_,
    new_n17766_, new_n17767_, new_n17768_, new_n17769_, new_n17770_,
    new_n17771_, new_n17772_, new_n17773_, new_n17774_, new_n17775_,
    new_n17776_, new_n17777_, new_n17778_, new_n17779_, new_n17780_,
    new_n17781_, new_n17782_, new_n17783_, new_n17784_, new_n17785_,
    new_n17786_, new_n17787_, new_n17788_, new_n17789_, new_n17790_,
    new_n17791_, new_n17792_, new_n17793_, new_n17794_, new_n17795_,
    new_n17796_, new_n17797_, new_n17798_, new_n17799_, new_n17800_,
    new_n17801_, new_n17802_, new_n17803_, new_n17804_, new_n17805_,
    new_n17806_, new_n17807_, new_n17808_, new_n17809_, new_n17810_,
    new_n17811_, new_n17812_, new_n17813_, new_n17814_, new_n17815_,
    new_n17816_, new_n17817_, new_n17818_, new_n17819_, new_n17820_,
    new_n17821_, new_n17822_, new_n17823_, new_n17824_, new_n17825_,
    new_n17826_, new_n17827_, new_n17828_, new_n17829_, new_n17830_,
    new_n17831_, new_n17832_, new_n17833_, new_n17834_, new_n17835_,
    new_n17836_, new_n17837_, new_n17838_, new_n17839_, new_n17840_,
    new_n17841_, new_n17842_, new_n17843_, new_n17844_, new_n17845_,
    new_n17846_, new_n17847_, new_n17848_, new_n17849_, new_n17850_,
    new_n17851_, new_n17852_, new_n17853_, new_n17854_, new_n17855_,
    new_n17856_, new_n17857_, new_n17858_, new_n17859_, new_n17860_,
    new_n17861_, new_n17862_, new_n17863_, new_n17864_, new_n17865_,
    new_n17866_, new_n17867_, new_n17868_, new_n17869_, new_n17870_,
    new_n17871_, new_n17872_, new_n17873_, new_n17874_, new_n17875_,
    new_n17876_, new_n17877_, new_n17878_, new_n17879_, new_n17880_,
    new_n17881_, new_n17882_, new_n17883_, new_n17884_, new_n17885_,
    new_n17886_, new_n17887_, new_n17888_, new_n17889_, new_n17890_,
    new_n17891_, new_n17892_, new_n17893_, new_n17894_, new_n17895_,
    new_n17896_, new_n17897_, new_n17898_, new_n17899_, new_n17900_,
    new_n17901_, new_n17902_, new_n17903_, new_n17904_, new_n17905_,
    new_n17906_, new_n17907_, new_n17908_, new_n17909_, new_n17910_,
    new_n17911_, new_n17912_, new_n17913_, new_n17914_, new_n17915_,
    new_n17916_, new_n17917_, new_n17918_, new_n17919_, new_n17920_,
    new_n17921_, new_n17922_, new_n17923_, new_n17924_, new_n17925_,
    new_n17926_, new_n17927_, new_n17928_, new_n17929_, new_n17930_,
    new_n17931_, new_n17932_, new_n17933_, new_n17934_, new_n17935_,
    new_n17936_, new_n17937_, new_n17938_, new_n17939_, new_n17940_,
    new_n17941_, new_n17942_, new_n17943_, new_n17944_, new_n17945_,
    new_n17946_, new_n17947_, new_n17948_, new_n17949_, new_n17950_,
    new_n17951_, new_n17952_, new_n17953_, new_n17954_, new_n17955_,
    new_n17956_, new_n17957_, new_n17958_, new_n17959_, new_n17960_,
    new_n17961_, new_n17962_, new_n17963_, new_n17964_, new_n17965_,
    new_n17966_, new_n17967_, new_n17968_, new_n17969_, new_n17970_,
    new_n17971_, new_n17972_, new_n17973_, new_n17974_, new_n17975_,
    new_n17976_, new_n17977_, new_n17978_, new_n17979_, new_n17980_,
    new_n17981_, new_n17982_, new_n17983_, new_n17984_, new_n17985_,
    new_n17986_, new_n17987_, new_n17988_, new_n17989_, new_n17990_,
    new_n17991_, new_n17992_, new_n17993_, new_n17994_, new_n17995_,
    new_n17996_, new_n17997_, new_n17998_, new_n17999_, new_n18000_,
    new_n18001_, new_n18002_, new_n18003_, new_n18004_, new_n18005_,
    new_n18006_, new_n18007_, new_n18008_, new_n18009_, new_n18010_,
    new_n18011_, new_n18012_, new_n18013_, new_n18014_, new_n18015_,
    new_n18016_, new_n18017_, new_n18018_, new_n18019_, new_n18020_,
    new_n18021_, new_n18022_, new_n18023_, new_n18024_, new_n18025_,
    new_n18026_, new_n18027_, new_n18028_, new_n18029_, new_n18030_,
    new_n18031_, new_n18032_, new_n18033_, new_n18034_, new_n18035_,
    new_n18036_, new_n18037_, new_n18038_, new_n18039_, new_n18040_,
    new_n18041_, new_n18042_, new_n18043_, new_n18044_, new_n18045_,
    new_n18046_, new_n18047_, new_n18048_, new_n18049_, new_n18050_,
    new_n18051_, new_n18052_, new_n18053_, new_n18054_, new_n18055_,
    new_n18056_, new_n18057_, new_n18058_, new_n18059_, new_n18060_,
    new_n18061_, new_n18062_, new_n18063_, new_n18064_, new_n18065_,
    new_n18066_, new_n18067_, new_n18068_, new_n18069_, new_n18070_,
    new_n18071_, new_n18072_, new_n18073_, new_n18074_, new_n18075_,
    new_n18076_, new_n18077_, new_n18078_, new_n18079_, new_n18080_,
    new_n18081_, new_n18082_, new_n18083_, new_n18084_, new_n18085_,
    new_n18086_, new_n18087_, new_n18088_, new_n18089_, new_n18090_,
    new_n18091_, new_n18092_, new_n18093_, new_n18094_, new_n18095_,
    new_n18096_, new_n18097_, new_n18098_, new_n18099_, new_n18100_,
    new_n18101_, new_n18102_, new_n18103_, new_n18104_, new_n18105_,
    new_n18106_, new_n18107_, new_n18108_, new_n18109_, new_n18110_,
    new_n18111_, new_n18112_, new_n18113_, new_n18114_, new_n18115_,
    new_n18116_, new_n18117_, new_n18118_, new_n18119_, new_n18120_,
    new_n18121_, new_n18122_, new_n18123_, new_n18124_, new_n18125_,
    new_n18126_, new_n18127_, new_n18128_, new_n18129_, new_n18130_,
    new_n18131_, new_n18132_, new_n18133_, new_n18134_, new_n18135_,
    new_n18136_, new_n18137_, new_n18138_, new_n18139_, new_n18140_,
    new_n18141_, new_n18142_, new_n18143_, new_n18144_, new_n18145_,
    new_n18146_, new_n18147_, new_n18148_, new_n18149_, new_n18150_,
    new_n18151_, new_n18152_, new_n18153_, new_n18154_, new_n18155_,
    new_n18156_, new_n18157_, new_n18158_, new_n18159_, new_n18160_,
    new_n18161_, new_n18162_, new_n18163_, new_n18164_, new_n18165_,
    new_n18166_, new_n18167_, new_n18168_, new_n18169_, new_n18170_,
    new_n18171_, new_n18172_, new_n18173_, new_n18174_, new_n18175_,
    new_n18176_, new_n18177_, new_n18178_, new_n18179_, new_n18180_,
    new_n18181_, new_n18182_, new_n18183_, new_n18184_, new_n18185_,
    new_n18186_, new_n18187_, new_n18188_, new_n18189_, new_n18190_,
    new_n18191_, new_n18192_, new_n18193_, new_n18194_, new_n18195_,
    new_n18196_, new_n18197_, new_n18198_, new_n18199_, new_n18200_,
    new_n18201_, new_n18202_, new_n18203_, new_n18204_, new_n18205_,
    new_n18206_, new_n18207_, new_n18208_, new_n18209_, new_n18210_,
    new_n18211_, new_n18212_, new_n18213_, new_n18214_, new_n18215_,
    new_n18216_, new_n18217_, new_n18218_, new_n18219_, new_n18220_,
    new_n18221_, new_n18222_, new_n18223_, new_n18224_, new_n18225_,
    new_n18226_, new_n18227_, new_n18228_, new_n18229_, new_n18230_,
    new_n18231_, new_n18232_, new_n18233_, new_n18234_, new_n18235_,
    new_n18236_, new_n18237_, new_n18238_, new_n18239_, new_n18240_,
    new_n18241_, new_n18242_, new_n18243_, new_n18244_, new_n18245_,
    new_n18246_, new_n18247_, new_n18248_, new_n18249_, new_n18250_,
    new_n18251_, new_n18252_, new_n18253_, new_n18254_, new_n18255_,
    new_n18256_, new_n18257_, new_n18258_, new_n18259_, new_n18260_,
    new_n18261_, new_n18262_, new_n18263_, new_n18264_, new_n18265_,
    new_n18266_, new_n18267_, new_n18268_, new_n18269_, new_n18270_,
    new_n18271_, new_n18272_, new_n18273_, new_n18274_, new_n18275_,
    new_n18276_, new_n18277_, new_n18278_, new_n18279_, new_n18280_,
    new_n18281_, new_n18282_, new_n18283_, new_n18284_, new_n18285_,
    new_n18286_, new_n18287_, new_n18288_, new_n18289_, new_n18290_,
    new_n18291_, new_n18292_, new_n18293_, new_n18294_, new_n18295_,
    new_n18296_, new_n18297_, new_n18298_, new_n18299_, new_n18300_,
    new_n18301_, new_n18302_, new_n18303_, new_n18304_, new_n18305_,
    new_n18306_, new_n18307_, new_n18308_, new_n18309_, new_n18310_,
    new_n18311_, new_n18312_, new_n18313_, new_n18314_, new_n18315_,
    new_n18316_, new_n18317_, new_n18318_, new_n18319_, new_n18320_,
    new_n18321_, new_n18322_, new_n18323_, new_n18324_, new_n18325_,
    new_n18326_, new_n18327_, new_n18328_, new_n18329_, new_n18330_,
    new_n18331_, new_n18332_, new_n18333_, new_n18334_, new_n18335_,
    new_n18336_, new_n18337_, new_n18338_, new_n18339_, new_n18340_,
    new_n18341_, new_n18342_, new_n18343_, new_n18344_, new_n18345_,
    new_n18346_, new_n18347_, new_n18348_, new_n18349_, new_n18350_,
    new_n18351_, new_n18352_, new_n18353_, new_n18354_, new_n18355_,
    new_n18356_, new_n18357_, new_n18358_, new_n18359_, new_n18360_,
    new_n18361_, new_n18362_, new_n18363_, new_n18364_, new_n18365_,
    new_n18366_, new_n18367_, new_n18368_, new_n18369_, new_n18370_,
    new_n18371_, new_n18372_, new_n18373_, new_n18374_, new_n18375_,
    new_n18376_, new_n18377_, new_n18378_, new_n18379_, new_n18380_,
    new_n18381_, new_n18382_, new_n18383_, new_n18384_, new_n18385_,
    new_n18386_, new_n18387_, new_n18388_, new_n18389_, new_n18390_,
    new_n18391_, new_n18392_, new_n18393_, new_n18394_, new_n18395_,
    new_n18396_, new_n18397_, new_n18398_, new_n18399_, new_n18400_,
    new_n18401_, new_n18402_, new_n18403_, new_n18404_, new_n18405_,
    new_n18406_, new_n18407_, new_n18408_, new_n18409_, new_n18410_,
    new_n18411_, new_n18412_, new_n18413_, new_n18414_, new_n18415_,
    new_n18416_, new_n18417_, new_n18418_, new_n18419_, new_n18420_,
    new_n18421_, new_n18422_, new_n18423_, new_n18424_, new_n18425_,
    new_n18426_, new_n18427_, new_n18428_, new_n18429_, new_n18430_,
    new_n18431_, new_n18432_, new_n18433_, new_n18434_, new_n18435_,
    new_n18436_, new_n18437_, new_n18438_, new_n18439_, new_n18440_,
    new_n18441_, new_n18442_, new_n18443_, new_n18444_, new_n18445_,
    new_n18446_, new_n18447_, new_n18448_, new_n18449_, new_n18450_,
    new_n18451_, new_n18452_, new_n18453_, new_n18454_, new_n18455_,
    new_n18456_, new_n18457_, new_n18458_, new_n18459_, new_n18460_,
    new_n18461_, new_n18462_, new_n18463_, new_n18464_, new_n18465_,
    new_n18466_, new_n18467_, new_n18468_, new_n18469_, new_n18470_,
    new_n18471_, new_n18472_, new_n18473_, new_n18474_, new_n18475_,
    new_n18476_, new_n18477_, new_n18478_, new_n18479_, new_n18480_,
    new_n18481_, new_n18482_, new_n18483_, new_n18484_, new_n18485_,
    new_n18486_, new_n18487_, new_n18488_, new_n18489_, new_n18490_,
    new_n18491_, new_n18492_, new_n18493_, new_n18494_, new_n18495_,
    new_n18496_, new_n18497_, new_n18498_, new_n18499_, new_n18500_,
    new_n18501_, new_n18502_, new_n18503_, new_n18504_, new_n18505_,
    new_n18506_, new_n18507_, new_n18508_, new_n18509_, new_n18510_,
    new_n18511_, new_n18512_, new_n18513_, new_n18514_, new_n18515_,
    new_n18516_, new_n18517_, new_n18518_, new_n18519_, new_n18520_,
    new_n18521_, new_n18522_, new_n18523_, new_n18524_, new_n18525_,
    new_n18526_, new_n18527_, new_n18528_, new_n18529_, new_n18530_,
    new_n18531_, new_n18532_, new_n18533_, new_n18534_, new_n18535_,
    new_n18536_, new_n18537_, new_n18538_, new_n18539_, new_n18540_,
    new_n18541_, new_n18542_, new_n18543_, new_n18544_, new_n18545_,
    new_n18546_, new_n18547_, new_n18548_, new_n18549_, new_n18550_,
    new_n18551_, new_n18552_, new_n18553_, new_n18554_, new_n18555_,
    new_n18556_, new_n18557_, new_n18558_, new_n18559_, new_n18560_,
    new_n18561_, new_n18562_, new_n18563_, new_n18564_, new_n18565_,
    new_n18566_, new_n18567_, new_n18568_, new_n18569_, new_n18570_,
    new_n18571_, new_n18572_, new_n18573_, new_n18574_, new_n18575_,
    new_n18576_, new_n18577_, new_n18578_, new_n18579_, new_n18580_,
    new_n18581_, new_n18582_, new_n18583_, new_n18584_, new_n18585_,
    new_n18586_, new_n18587_, new_n18588_, new_n18589_, new_n18590_,
    new_n18591_, new_n18592_, new_n18593_, new_n18594_, new_n18595_,
    new_n18596_, new_n18597_, new_n18598_, new_n18599_, new_n18600_,
    new_n18601_, new_n18602_, new_n18603_, new_n18604_, new_n18605_,
    new_n18606_, new_n18607_, new_n18608_, new_n18609_, new_n18610_,
    new_n18611_, new_n18612_, new_n18613_, new_n18614_, new_n18615_,
    new_n18616_, new_n18617_, new_n18618_, new_n18619_, new_n18620_,
    new_n18621_, new_n18622_, new_n18623_, new_n18624_, new_n18625_,
    new_n18626_, new_n18627_, new_n18628_, new_n18629_, new_n18630_,
    new_n18631_, new_n18632_, new_n18633_, new_n18634_, new_n18635_,
    new_n18636_, new_n18637_, new_n18638_, new_n18639_, new_n18640_,
    new_n18641_, new_n18642_, new_n18643_, new_n18644_, new_n18645_,
    new_n18646_, new_n18647_, new_n18648_, new_n18649_, new_n18650_,
    new_n18651_, new_n18652_, new_n18653_, new_n18654_, new_n18655_,
    new_n18656_, new_n18657_, new_n18658_, new_n18659_, new_n18660_,
    new_n18661_, new_n18662_, new_n18663_, new_n18664_, new_n18665_,
    new_n18666_, new_n18667_, new_n18668_, new_n18669_, new_n18670_,
    new_n18671_, new_n18672_, new_n18673_, new_n18674_, new_n18675_,
    new_n18676_, new_n18677_, new_n18678_, new_n18679_, new_n18680_,
    new_n18681_, new_n18682_, new_n18683_, new_n18684_, new_n18685_,
    new_n18686_, new_n18687_, new_n18688_, new_n18689_, new_n18690_,
    new_n18691_, new_n18692_, new_n18693_, new_n18694_, new_n18695_,
    new_n18696_, new_n18697_, new_n18698_, new_n18699_, new_n18700_,
    new_n18701_, new_n18702_, new_n18703_, new_n18704_, new_n18705_,
    new_n18706_, new_n18707_, new_n18708_, new_n18709_, new_n18710_,
    new_n18711_, new_n18712_, new_n18713_, new_n18714_, new_n18715_,
    new_n18716_, new_n18717_, new_n18718_, new_n18719_, new_n18720_,
    new_n18721_, new_n18722_, new_n18723_, new_n18724_, new_n18725_,
    new_n18726_, new_n18727_, new_n18728_, new_n18729_, new_n18730_,
    new_n18731_, new_n18732_, new_n18733_, new_n18734_, new_n18735_,
    new_n18736_, new_n18737_, new_n18738_, new_n18739_, new_n18740_,
    new_n18741_, new_n18742_, new_n18743_, new_n18744_, new_n18745_,
    new_n18746_, new_n18747_, new_n18748_, new_n18749_, new_n18750_,
    new_n18751_, new_n18752_, new_n18753_, new_n18754_, new_n18755_,
    new_n18756_, new_n18757_, new_n18758_, new_n18759_, new_n18760_,
    new_n18761_, new_n18762_, new_n18763_, new_n18764_, new_n18765_,
    new_n18766_, new_n18767_, new_n18768_, new_n18769_, new_n18770_,
    new_n18771_, new_n18772_, new_n18773_, new_n18774_, new_n18775_,
    new_n18776_, new_n18777_, new_n18778_, new_n18779_, new_n18780_,
    new_n18781_, new_n18782_, new_n18783_, new_n18784_, new_n18785_,
    new_n18786_, new_n18787_, new_n18788_, new_n18789_, new_n18790_,
    new_n18791_, new_n18792_, new_n18793_, new_n18794_, new_n18795_,
    new_n18796_, new_n18797_, new_n18798_, new_n18799_, new_n18800_,
    new_n18801_, new_n18802_, new_n18803_, new_n18804_, new_n18805_,
    new_n18806_, new_n18807_, new_n18808_, new_n18809_, new_n18810_,
    new_n18811_, new_n18812_, new_n18813_, new_n18814_, new_n18815_,
    new_n18816_, new_n18817_, new_n18818_, new_n18819_, new_n18820_,
    new_n18821_, new_n18822_, new_n18823_, new_n18824_, new_n18825_,
    new_n18826_, new_n18827_, new_n18828_, new_n18829_, new_n18830_,
    new_n18831_, new_n18832_, new_n18833_, new_n18834_, new_n18835_,
    new_n18836_, new_n18837_, new_n18838_, new_n18839_, new_n18840_,
    new_n18841_, new_n18842_, new_n18843_, new_n18844_, new_n18845_,
    new_n18846_, new_n18847_, new_n18848_, new_n18849_, new_n18850_,
    new_n18851_, new_n18852_, new_n18853_, new_n18854_, new_n18855_,
    new_n18856_, new_n18857_, new_n18858_, new_n18859_, new_n18860_,
    new_n18861_, new_n18862_, new_n18863_, new_n18864_, new_n18865_,
    new_n18866_, new_n18867_, new_n18868_, new_n18869_, new_n18870_,
    new_n18871_, new_n18872_, new_n18873_, new_n18874_, new_n18875_,
    new_n18876_, new_n18877_, new_n18878_, new_n18879_, new_n18880_,
    new_n18881_, new_n18882_, new_n18883_, new_n18884_, new_n18885_,
    new_n18886_, new_n18887_, new_n18888_, new_n18889_, new_n18890_,
    new_n18891_, new_n18892_, new_n18893_, new_n18894_, new_n18895_,
    new_n18896_, new_n18897_, new_n18898_, new_n18899_, new_n18900_,
    new_n18901_, new_n18902_, new_n18903_, new_n18904_, new_n18905_,
    new_n18906_, new_n18907_, new_n18908_, new_n18909_, new_n18910_,
    new_n18911_, new_n18912_, new_n18913_, new_n18914_, new_n18915_,
    new_n18916_, new_n18917_, new_n18918_, new_n18919_, new_n18920_,
    new_n18921_, new_n18922_, new_n18923_, new_n18924_, new_n18925_,
    new_n18926_, new_n18927_, new_n18928_, new_n18929_, new_n18930_,
    new_n18931_, new_n18932_, new_n18933_, new_n18934_, new_n18935_,
    new_n18936_, new_n18937_, new_n18938_, new_n18939_, new_n18940_,
    new_n18941_, new_n18942_, new_n18943_, new_n18944_, new_n18945_,
    new_n18946_, new_n18947_, new_n18948_, new_n18949_, new_n18950_,
    new_n18951_, new_n18952_, new_n18953_, new_n18954_, new_n18955_,
    new_n18956_, new_n18957_, new_n18958_, new_n18959_, new_n18960_,
    new_n18961_, new_n18962_, new_n18963_, new_n18964_, new_n18965_,
    new_n18966_, new_n18967_, new_n18968_, new_n18969_, new_n18970_,
    new_n18971_, new_n18972_, new_n18973_, new_n18974_, new_n18975_,
    new_n18976_, new_n18977_, new_n18978_, new_n18979_, new_n18980_,
    new_n18981_, new_n18982_, new_n18983_, new_n18984_, new_n18985_,
    new_n18986_, new_n18987_, new_n18988_, new_n18989_, new_n18990_,
    new_n18991_, new_n18992_, new_n18993_, new_n18994_, new_n18995_,
    new_n18996_, new_n18997_, new_n18998_, new_n18999_, new_n19000_,
    new_n19001_, new_n19002_, new_n19003_, new_n19004_, new_n19005_,
    new_n19006_, new_n19007_, new_n19008_, new_n19009_, new_n19010_,
    new_n19011_, new_n19012_, new_n19013_, new_n19014_, new_n19015_,
    new_n19016_, new_n19017_, new_n19018_, new_n19019_, new_n19020_,
    new_n19021_, new_n19022_, new_n19023_, new_n19024_, new_n19025_,
    new_n19026_, new_n19027_, new_n19028_, new_n19029_, new_n19030_,
    new_n19031_, new_n19032_, new_n19033_, new_n19034_, new_n19035_,
    new_n19036_, new_n19037_, new_n19038_, new_n19039_, new_n19040_,
    new_n19041_, new_n19042_, new_n19043_, new_n19044_, new_n19045_,
    new_n19046_, new_n19047_, new_n19048_, new_n19049_, new_n19050_,
    new_n19051_, new_n19052_, new_n19053_, new_n19054_, new_n19055_,
    new_n19056_, new_n19057_, new_n19058_, new_n19059_, new_n19060_,
    new_n19061_, new_n19062_, new_n19063_, new_n19064_, new_n19065_,
    new_n19066_, new_n19067_, new_n19068_, new_n19069_, new_n19070_,
    new_n19071_, new_n19072_, new_n19073_, new_n19074_, new_n19075_,
    new_n19076_, new_n19077_, new_n19078_, new_n19079_, new_n19080_,
    new_n19081_, new_n19082_, new_n19083_, new_n19084_, new_n19085_,
    new_n19086_, new_n19087_, new_n19088_, new_n19089_, new_n19090_,
    new_n19091_, new_n19092_, new_n19093_, new_n19094_, new_n19095_,
    new_n19096_, new_n19097_, new_n19098_, new_n19099_, new_n19100_,
    new_n19101_, new_n19102_, new_n19103_, new_n19104_, new_n19105_,
    new_n19106_, new_n19107_, new_n19108_, new_n19109_, new_n19110_,
    new_n19111_, new_n19112_, new_n19113_, new_n19114_, new_n19115_,
    new_n19116_, new_n19117_, new_n19118_, new_n19119_, new_n19120_,
    new_n19121_, new_n19122_, new_n19123_, new_n19124_, new_n19125_,
    new_n19126_, new_n19127_, new_n19128_, new_n19129_, new_n19130_,
    new_n19131_, new_n19132_, new_n19133_, new_n19134_, new_n19135_,
    new_n19136_, new_n19137_, new_n19138_, new_n19139_, new_n19140_,
    new_n19141_, new_n19142_, new_n19143_, new_n19144_, new_n19145_,
    new_n19146_, new_n19147_, new_n19148_, new_n19149_, new_n19150_,
    new_n19151_, new_n19152_, new_n19153_, new_n19154_, new_n19155_,
    new_n19156_, new_n19157_, new_n19158_, new_n19159_, new_n19160_,
    new_n19161_, new_n19162_, new_n19163_, new_n19164_, new_n19165_,
    new_n19166_, new_n19167_, new_n19168_, new_n19169_, new_n19170_,
    new_n19171_, new_n19172_, new_n19173_, new_n19174_, new_n19175_,
    new_n19176_, new_n19177_, new_n19178_, new_n19179_, new_n19180_,
    new_n19181_, new_n19182_, new_n19183_, new_n19184_, new_n19185_,
    new_n19186_, new_n19187_, new_n19188_, new_n19189_, new_n19190_,
    new_n19191_, new_n19192_, new_n19193_, new_n19194_, new_n19195_,
    new_n19196_, new_n19197_, new_n19198_, new_n19199_, new_n19200_,
    new_n19201_, new_n19202_, new_n19203_, new_n19204_, new_n19205_,
    new_n19206_, new_n19207_, new_n19208_, new_n19209_, new_n19210_,
    new_n19211_, new_n19212_, new_n19213_, new_n19214_, new_n19215_,
    new_n19216_, new_n19217_, new_n19218_, new_n19219_, new_n19220_,
    new_n19221_, new_n19222_, new_n19223_, new_n19224_, new_n19225_,
    new_n19226_, new_n19227_, new_n19228_, new_n19229_, new_n19230_,
    new_n19231_, new_n19232_, new_n19233_, new_n19234_, new_n19235_,
    new_n19236_, new_n19237_, new_n19238_, new_n19239_, new_n19240_,
    new_n19241_, new_n19242_, new_n19243_, new_n19244_, new_n19245_,
    new_n19246_, new_n19247_, new_n19248_, new_n19249_, new_n19250_,
    new_n19251_, new_n19252_, new_n19253_, new_n19254_, new_n19255_,
    new_n19256_, new_n19257_, new_n19258_, new_n19259_, new_n19260_,
    new_n19261_, new_n19262_, new_n19263_, new_n19264_, new_n19265_,
    new_n19266_, new_n19267_, new_n19268_, new_n19269_, new_n19270_,
    new_n19271_, new_n19272_, new_n19273_, new_n19274_, new_n19275_,
    new_n19276_, new_n19277_, new_n19278_, new_n19279_, new_n19280_,
    new_n19281_, new_n19282_, new_n19283_, new_n19284_, new_n19285_,
    new_n19286_, new_n19287_, new_n19288_, new_n19289_, new_n19290_,
    new_n19291_, new_n19292_, new_n19293_, new_n19294_, new_n19295_,
    new_n19296_, new_n19297_, new_n19298_, new_n19299_, new_n19300_,
    new_n19301_, new_n19302_, new_n19303_, new_n19304_, new_n19305_,
    new_n19306_, new_n19307_, new_n19308_, new_n19309_, new_n19310_,
    new_n19311_, new_n19312_, new_n19313_, new_n19314_, new_n19315_,
    new_n19316_, new_n19317_, new_n19318_, new_n19319_, new_n19320_,
    new_n19321_, new_n19322_, new_n19323_, new_n19324_, new_n19325_,
    new_n19326_, new_n19327_, new_n19328_, new_n19329_, new_n19330_,
    new_n19331_, new_n19332_, new_n19333_, new_n19334_, new_n19335_,
    new_n19336_, new_n19337_, new_n19338_, new_n19339_, new_n19340_,
    new_n19341_, new_n19342_, new_n19343_, new_n19344_, new_n19345_,
    new_n19346_, new_n19347_, new_n19348_, new_n19349_, new_n19350_,
    new_n19351_, new_n19352_, new_n19353_, new_n19354_, new_n19355_,
    new_n19356_, new_n19357_, new_n19358_, new_n19359_, new_n19360_,
    new_n19361_, new_n19362_, new_n19363_, new_n19364_, new_n19365_,
    new_n19366_, new_n19367_, new_n19368_, new_n19369_, new_n19370_,
    new_n19371_, new_n19372_, new_n19373_, new_n19374_, new_n19375_,
    new_n19376_, new_n19377_, new_n19378_, new_n19379_, new_n19380_,
    new_n19381_, new_n19382_, new_n19383_, new_n19384_, new_n19385_,
    new_n19386_, new_n19387_, new_n19388_, new_n19389_, new_n19390_,
    new_n19391_, new_n19392_, new_n19393_, new_n19394_, new_n19395_,
    new_n19396_, new_n19397_, new_n19398_, new_n19399_, new_n19400_,
    new_n19401_, new_n19402_, new_n19403_, new_n19404_, new_n19405_,
    new_n19406_, new_n19407_, new_n19408_, new_n19409_, new_n19410_,
    new_n19411_, new_n19412_, new_n19413_, new_n19414_, new_n19415_,
    new_n19416_, new_n19417_, new_n19418_, new_n19419_, new_n19420_,
    new_n19421_, new_n19422_, new_n19423_, new_n19424_, new_n19425_,
    new_n19426_, new_n19427_, new_n19428_, new_n19429_, new_n19430_,
    new_n19431_, new_n19432_, new_n19433_, new_n19434_, new_n19435_,
    new_n19436_, new_n19437_, new_n19438_, new_n19439_, new_n19440_,
    new_n19441_, new_n19442_, new_n19443_, new_n19444_, new_n19445_,
    new_n19446_, new_n19447_, new_n19448_, new_n19449_, new_n19450_,
    new_n19451_, new_n19452_, new_n19453_, new_n19454_, new_n19455_,
    new_n19456_, new_n19457_, new_n19458_, new_n19459_, new_n19460_,
    new_n19461_, new_n19462_, new_n19463_, new_n19464_, new_n19465_,
    new_n19466_, new_n19467_, new_n19468_, new_n19469_, new_n19470_,
    new_n19471_, new_n19472_, new_n19473_, new_n19474_, new_n19475_,
    new_n19476_, new_n19477_, new_n19478_, new_n19479_, new_n19480_,
    new_n19481_, new_n19482_, new_n19483_, new_n19484_, new_n19485_,
    new_n19486_, new_n19487_, new_n19488_, new_n19489_, new_n19490_,
    new_n19491_, new_n19492_, new_n19493_, new_n19494_, new_n19495_,
    new_n19496_, new_n19497_, new_n19498_, new_n19499_, new_n19500_,
    new_n19501_, new_n19502_, new_n19503_, new_n19504_, new_n19505_,
    new_n19506_, new_n19507_, new_n19508_, new_n19509_, new_n19510_,
    new_n19511_, new_n19512_, new_n19513_, new_n19514_, new_n19515_,
    new_n19516_, new_n19517_, new_n19518_, new_n19519_, new_n19520_,
    new_n19521_, new_n19522_, new_n19523_, new_n19524_, new_n19525_,
    new_n19526_, new_n19527_, new_n19528_, new_n19529_, new_n19530_,
    new_n19531_, new_n19532_, new_n19533_, new_n19534_, new_n19535_,
    new_n19536_, new_n19537_, new_n19538_, new_n19539_, new_n19540_,
    new_n19541_, new_n19542_, new_n19543_, new_n19544_, new_n19545_,
    new_n19546_, new_n19547_, new_n19548_, new_n19549_, new_n19550_,
    new_n19551_, new_n19552_, new_n19553_, new_n19554_, new_n19555_,
    new_n19556_, new_n19557_, new_n19558_, new_n19559_, new_n19560_,
    new_n19561_, new_n19562_, new_n19563_, new_n19564_, new_n19565_,
    new_n19566_, new_n19567_, new_n19568_, new_n19569_, new_n19570_,
    new_n19571_, new_n19572_, new_n19573_, new_n19574_, new_n19575_,
    new_n19576_, new_n19577_, new_n19578_, new_n19579_, new_n19580_,
    new_n19581_, new_n19582_, new_n19583_, new_n19584_, new_n19585_,
    new_n19586_, new_n19587_, new_n19588_, new_n19589_, new_n19590_,
    new_n19591_, new_n19592_, new_n19593_, new_n19594_, new_n19595_,
    new_n19596_, new_n19597_, new_n19598_, new_n19599_, new_n19600_,
    new_n19601_, new_n19602_, new_n19603_, new_n19604_, new_n19605_,
    new_n19606_, new_n19607_, new_n19608_, new_n19609_, new_n19610_,
    new_n19611_, new_n19612_, new_n19613_, new_n19614_, new_n19615_,
    new_n19616_, new_n19617_, new_n19618_, new_n19619_, new_n19620_,
    new_n19621_, new_n19622_, new_n19623_, new_n19624_, new_n19625_,
    new_n19626_, new_n19627_, new_n19628_, new_n19629_, new_n19630_,
    new_n19631_, new_n19632_, new_n19633_, new_n19634_, new_n19635_,
    new_n19636_, new_n19637_, new_n19638_, new_n19639_, new_n19640_,
    new_n19641_, new_n19642_, new_n19643_, new_n19644_, new_n19645_,
    new_n19646_, new_n19647_, new_n19648_, new_n19649_, new_n19650_,
    new_n19651_, new_n19652_, new_n19653_, new_n19654_, new_n19655_,
    new_n19656_, new_n19657_, new_n19658_, new_n19659_, new_n19660_,
    new_n19661_, new_n19662_, new_n19663_, new_n19664_, new_n19665_,
    new_n19666_, new_n19667_, new_n19668_, new_n19669_, new_n19670_,
    new_n19671_, new_n19672_, new_n19673_, new_n19674_, new_n19675_,
    new_n19676_, new_n19677_, new_n19678_, new_n19679_, new_n19680_,
    new_n19681_, new_n19682_, new_n19683_, new_n19684_, new_n19685_,
    new_n19686_, new_n19687_, new_n19688_, new_n19689_, new_n19690_,
    new_n19691_, new_n19692_, new_n19693_, new_n19694_, new_n19695_,
    new_n19696_, new_n19697_, new_n19698_, new_n19699_, new_n19700_,
    new_n19701_, new_n19702_, new_n19703_, new_n19704_, new_n19705_,
    new_n19706_, new_n19707_, new_n19708_, new_n19709_, new_n19710_,
    new_n19711_, new_n19712_, new_n19713_, new_n19714_, new_n19715_,
    new_n19716_, new_n19717_, new_n19718_, new_n19719_, new_n19720_,
    new_n19721_, new_n19722_, new_n19723_, new_n19724_, new_n19725_,
    new_n19726_, new_n19727_, new_n19728_, new_n19729_, new_n19730_,
    new_n19731_, new_n19732_, new_n19733_, new_n19734_, new_n19735_,
    new_n19736_, new_n19737_, new_n19738_, new_n19739_, new_n19740_,
    new_n19741_, new_n19742_, new_n19743_, new_n19744_, new_n19745_,
    new_n19746_, new_n19747_, new_n19748_, new_n19749_, new_n19750_,
    new_n19751_, new_n19752_, new_n19753_, new_n19754_, new_n19755_,
    new_n19756_, new_n19757_, new_n19758_, new_n19759_, new_n19760_,
    new_n19761_, new_n19762_, new_n19763_, new_n19764_, new_n19765_,
    new_n19766_, new_n19767_, new_n19768_, new_n19769_, new_n19770_,
    new_n19771_, new_n19772_, new_n19773_, new_n19774_, new_n19775_,
    new_n19776_, new_n19777_, new_n19778_, new_n19779_, new_n19780_,
    new_n19781_, new_n19782_, new_n19783_, new_n19784_, new_n19785_,
    new_n19786_, new_n19787_, new_n19788_, new_n19789_, new_n19790_,
    new_n19791_, new_n19792_, new_n19793_, new_n19794_, new_n19795_,
    new_n19796_, new_n19797_, new_n19798_, new_n19799_, new_n19800_,
    new_n19801_, new_n19802_, new_n19803_, new_n19804_, new_n19805_,
    new_n19806_, new_n19807_, new_n19808_, new_n19809_, new_n19810_,
    new_n19811_, new_n19812_, new_n19813_, new_n19814_, new_n19815_,
    new_n19816_, new_n19817_, new_n19818_, new_n19819_, new_n19820_,
    new_n19821_, new_n19822_, new_n19823_, new_n19824_, new_n19825_,
    new_n19826_, new_n19827_, new_n19828_, new_n19829_, new_n19830_,
    new_n19831_, new_n19832_, new_n19833_, new_n19834_, new_n19835_,
    new_n19836_, new_n19837_, new_n19838_, new_n19839_, new_n19840_,
    new_n19841_, new_n19842_, new_n19843_, new_n19844_, new_n19845_,
    new_n19846_, new_n19847_, new_n19848_, new_n19849_, new_n19850_,
    new_n19851_, new_n19852_, new_n19853_, new_n19854_, new_n19855_,
    new_n19856_, new_n19857_, new_n19858_, new_n19859_, new_n19860_,
    new_n19861_, new_n19862_, new_n19863_, new_n19864_, new_n19865_,
    new_n19866_, new_n19867_, new_n19868_, new_n19869_, new_n19870_,
    new_n19871_, new_n19872_, new_n19873_, new_n19874_, new_n19875_,
    new_n19876_, new_n19877_, new_n19878_, new_n19879_, new_n19880_,
    new_n19881_, new_n19882_, new_n19883_, new_n19884_, new_n19885_,
    new_n19886_, new_n19887_, new_n19888_, new_n19889_, new_n19890_,
    new_n19891_, new_n19892_, new_n19893_, new_n19894_, new_n19895_,
    new_n19896_, new_n19897_, new_n19898_, new_n19899_, new_n19900_,
    new_n19901_, new_n19902_, new_n19903_, new_n19904_, new_n19905_,
    new_n19906_, new_n19907_, new_n19908_, new_n19909_, new_n19910_,
    new_n19911_, new_n19912_, new_n19913_, new_n19914_, new_n19915_,
    new_n19916_, new_n19917_, new_n19918_, new_n19919_, new_n19920_,
    new_n19921_, new_n19922_, new_n19923_, new_n19924_, new_n19925_,
    new_n19926_, new_n19927_, new_n19928_, new_n19929_, new_n19930_,
    new_n19931_, new_n19932_, new_n19933_, new_n19934_, new_n19935_,
    new_n19936_, new_n19937_, new_n19938_, new_n19939_, new_n19940_,
    new_n19941_, new_n19942_, new_n19943_, new_n19944_, new_n19945_,
    new_n19946_, new_n19947_, new_n19948_, new_n19949_, new_n19950_,
    new_n19951_, new_n19952_, new_n19953_, new_n19954_, new_n19955_,
    new_n19956_, new_n19957_, new_n19958_, new_n19959_, new_n19960_,
    new_n19961_, new_n19962_, new_n19963_, new_n19964_, new_n19965_,
    new_n19966_, new_n19967_, new_n19968_, new_n19969_, new_n19970_,
    new_n19971_, new_n19972_, new_n19973_, new_n19974_, new_n19975_,
    new_n19976_, new_n19977_, new_n19978_, new_n19979_, new_n19980_,
    new_n19981_, new_n19982_, new_n19983_, new_n19984_, new_n19985_,
    new_n19986_, new_n19987_, new_n19988_, new_n19989_, new_n19990_,
    new_n19991_, new_n19992_, new_n19993_, new_n19994_, new_n19995_,
    new_n19996_, new_n19997_, new_n19998_, new_n19999_, new_n20000_,
    new_n20001_, new_n20002_, new_n20003_, new_n20004_, new_n20005_,
    new_n20006_, new_n20007_, new_n20008_, new_n20009_, new_n20010_,
    new_n20011_, new_n20012_, new_n20013_, new_n20014_, new_n20015_,
    new_n20016_, new_n20017_, new_n20018_, new_n20019_, new_n20020_,
    new_n20021_, new_n20022_, new_n20023_, new_n20024_, new_n20025_,
    new_n20026_, new_n20027_, new_n20028_, new_n20029_, new_n20030_,
    new_n20031_, new_n20032_, new_n20033_, new_n20034_, new_n20035_,
    new_n20036_, new_n20037_, new_n20038_, new_n20039_, new_n20040_,
    new_n20041_, new_n20042_, new_n20043_, new_n20044_, new_n20045_,
    new_n20046_, new_n20047_, new_n20048_, new_n20049_, new_n20050_,
    new_n20051_, new_n20052_, new_n20053_, new_n20054_, new_n20055_,
    new_n20056_, new_n20057_, new_n20058_, new_n20059_, new_n20060_,
    new_n20061_, new_n20062_, new_n20063_, new_n20064_, new_n20065_,
    new_n20066_, new_n20067_, new_n20068_, new_n20069_, new_n20070_,
    new_n20071_, new_n20072_, new_n20073_, new_n20074_, new_n20075_,
    new_n20076_, new_n20077_, new_n20078_, new_n20079_, new_n20080_,
    new_n20081_, new_n20082_, new_n20083_, new_n20084_, new_n20085_,
    new_n20086_, new_n20087_, new_n20088_, new_n20089_, new_n20090_,
    new_n20091_, new_n20092_, new_n20093_, new_n20094_, new_n20095_,
    new_n20096_, new_n20097_, new_n20098_, new_n20099_, new_n20100_,
    new_n20101_, new_n20102_, new_n20103_, new_n20104_, new_n20105_,
    new_n20106_, new_n20107_, new_n20108_, new_n20109_, new_n20110_,
    new_n20111_, new_n20112_, new_n20113_, new_n20114_, new_n20115_,
    new_n20116_, new_n20117_, new_n20118_, new_n20119_, new_n20120_,
    new_n20121_, new_n20122_, new_n20123_, new_n20124_, new_n20125_,
    new_n20126_, new_n20127_, new_n20128_, new_n20129_, new_n20130_,
    new_n20131_, new_n20132_, new_n20133_, new_n20134_, new_n20135_,
    new_n20136_, new_n20137_, new_n20138_, new_n20139_, new_n20140_,
    new_n20141_, new_n20142_, new_n20143_, new_n20144_, new_n20145_,
    new_n20146_, new_n20147_, new_n20148_, new_n20149_, new_n20150_,
    new_n20151_, new_n20152_, new_n20153_, new_n20154_, new_n20155_,
    new_n20156_, new_n20157_, new_n20158_, new_n20159_, new_n20160_,
    new_n20161_, new_n20162_, new_n20163_, new_n20164_, new_n20165_,
    new_n20166_, new_n20167_, new_n20168_, new_n20169_, new_n20170_,
    new_n20171_, new_n20172_, new_n20173_, new_n20174_, new_n20175_,
    new_n20176_, new_n20177_, new_n20178_, new_n20179_, new_n20180_,
    new_n20181_, new_n20182_, new_n20183_, new_n20184_, new_n20185_,
    new_n20186_, new_n20187_, new_n20188_, new_n20189_, new_n20190_,
    new_n20191_, new_n20192_, new_n20193_, new_n20194_, new_n20195_,
    new_n20196_, new_n20197_, new_n20198_, new_n20199_, new_n20200_,
    new_n20201_, new_n20202_, new_n20203_, new_n20204_, new_n20205_,
    new_n20206_, new_n20207_, new_n20208_, new_n20209_, new_n20210_,
    new_n20211_, new_n20212_, new_n20213_, new_n20214_, new_n20215_,
    new_n20216_, new_n20217_, new_n20218_, new_n20219_, new_n20220_,
    new_n20221_, new_n20222_, new_n20223_, new_n20224_, new_n20225_,
    new_n20226_, new_n20227_, new_n20228_, new_n20229_, new_n20230_,
    new_n20231_, new_n20232_, new_n20233_, new_n20234_, new_n20235_,
    new_n20236_, new_n20237_, new_n20238_, new_n20239_, new_n20240_,
    new_n20241_, new_n20242_, new_n20243_, new_n20244_, new_n20245_,
    new_n20246_, new_n20247_, new_n20248_, new_n20249_, new_n20250_,
    new_n20251_, new_n20252_, new_n20253_, new_n20254_, new_n20255_,
    new_n20256_, new_n20257_, new_n20258_, new_n20259_, new_n20260_,
    new_n20261_, new_n20262_, new_n20263_, new_n20264_, new_n20265_,
    new_n20266_, new_n20267_, new_n20268_, new_n20269_, new_n20270_,
    new_n20271_, new_n20272_, new_n20273_, new_n20274_, new_n20275_,
    new_n20276_, new_n20277_, new_n20278_, new_n20279_, new_n20280_,
    new_n20281_, new_n20282_, new_n20283_, new_n20284_, new_n20285_,
    new_n20286_, new_n20287_, new_n20288_, new_n20289_, new_n20290_,
    new_n20291_, new_n20292_, new_n20293_, new_n20294_, new_n20295_,
    new_n20296_, new_n20297_, new_n20298_, new_n20299_, new_n20300_,
    new_n20301_, new_n20302_, new_n20303_, new_n20304_, new_n20305_,
    new_n20306_, new_n20307_, new_n20308_, new_n20309_, new_n20310_,
    new_n20311_, new_n20312_, new_n20313_, new_n20314_, new_n20315_,
    new_n20316_, new_n20317_, new_n20318_, new_n20319_, new_n20320_,
    new_n20321_, new_n20322_, new_n20323_, new_n20324_, new_n20325_,
    new_n20326_, new_n20327_, new_n20328_, new_n20329_, new_n20330_,
    new_n20331_, new_n20332_, new_n20333_, new_n20334_, new_n20335_,
    new_n20336_, new_n20337_, new_n20338_, new_n20339_, new_n20340_,
    new_n20341_, new_n20342_, new_n20343_, new_n20344_, new_n20345_,
    new_n20346_, new_n20347_, new_n20348_, new_n20349_, new_n20350_,
    new_n20351_, new_n20352_, new_n20353_, new_n20354_, new_n20355_,
    new_n20356_, new_n20357_, new_n20358_, new_n20359_, new_n20360_,
    new_n20361_, new_n20362_, new_n20363_, new_n20364_, new_n20365_,
    new_n20366_, new_n20367_, new_n20368_, new_n20369_, new_n20370_,
    new_n20371_, new_n20372_, new_n20373_, new_n20374_, new_n20375_,
    new_n20376_, new_n20377_, new_n20378_, new_n20379_, new_n20380_,
    new_n20381_, new_n20382_, new_n20383_, new_n20384_, new_n20385_,
    new_n20386_, new_n20387_, new_n20388_, new_n20389_, new_n20390_,
    new_n20391_, new_n20392_, new_n20393_, new_n20394_, new_n20395_,
    new_n20396_, new_n20397_, new_n20398_, new_n20399_, new_n20400_,
    new_n20401_, new_n20402_, new_n20403_, new_n20404_, new_n20405_,
    new_n20406_, new_n20407_, new_n20408_, new_n20409_, new_n20410_,
    new_n20411_, new_n20412_, new_n20413_, new_n20414_, new_n20415_,
    new_n20416_, new_n20417_, new_n20418_, new_n20419_, new_n20420_,
    new_n20421_, new_n20422_, new_n20423_, new_n20424_, new_n20425_,
    new_n20426_, new_n20427_, new_n20428_, new_n20429_, new_n20430_,
    new_n20431_, new_n20432_, new_n20433_, new_n20434_, new_n20435_,
    new_n20436_, new_n20437_, new_n20438_, new_n20439_, new_n20440_,
    new_n20441_, new_n20442_, new_n20443_, new_n20444_, new_n20445_,
    new_n20446_, new_n20447_, new_n20448_, new_n20449_, new_n20450_,
    new_n20451_, new_n20452_, new_n20453_, new_n20454_, new_n20455_,
    new_n20456_, new_n20457_, new_n20458_, new_n20459_, new_n20460_,
    new_n20461_, new_n20462_, new_n20463_, new_n20464_, new_n20465_,
    new_n20466_, new_n20467_, new_n20468_, new_n20469_, new_n20470_,
    new_n20471_, new_n20472_, new_n20473_, new_n20474_, new_n20475_,
    new_n20476_, new_n20477_, new_n20478_, new_n20479_, new_n20480_,
    new_n20481_, new_n20482_, new_n20483_, new_n20484_, new_n20485_,
    new_n20486_, new_n20487_, new_n20488_, new_n20489_, new_n20490_,
    new_n20491_, new_n20492_, new_n20493_, new_n20494_, new_n20495_,
    new_n20496_, new_n20497_, new_n20498_, new_n20499_, new_n20500_,
    new_n20501_, new_n20502_, new_n20503_, new_n20504_, new_n20505_,
    new_n20506_, new_n20507_, new_n20508_, new_n20509_, new_n20510_,
    new_n20511_, new_n20512_, new_n20513_, new_n20514_, new_n20515_,
    new_n20516_, new_n20517_, new_n20518_, new_n20519_, new_n20520_,
    new_n20521_, new_n20522_, new_n20523_, new_n20524_, new_n20525_,
    new_n20526_, new_n20527_, new_n20528_, new_n20529_, new_n20530_,
    new_n20531_, new_n20532_, new_n20533_, new_n20534_, new_n20535_,
    new_n20536_, new_n20537_, new_n20538_, new_n20539_, new_n20540_,
    new_n20541_, new_n20542_, new_n20543_, new_n20544_, new_n20545_,
    new_n20546_, new_n20547_, new_n20548_, new_n20549_, new_n20550_,
    new_n20551_, new_n20552_, new_n20553_, new_n20554_, new_n20555_,
    new_n20556_, new_n20557_, new_n20558_, new_n20559_, new_n20560_,
    new_n20561_, new_n20562_, new_n20563_, new_n20564_, new_n20565_,
    new_n20566_, new_n20567_, new_n20568_, new_n20569_, new_n20570_,
    new_n20571_, new_n20572_, new_n20573_, new_n20574_, new_n20575_,
    new_n20576_, new_n20577_, new_n20578_, new_n20579_, new_n20580_,
    new_n20581_, new_n20582_, new_n20583_, new_n20584_, new_n20585_,
    new_n20586_, new_n20587_, new_n20588_, new_n20589_, new_n20590_,
    new_n20591_, new_n20592_, new_n20593_, new_n20594_, new_n20595_,
    new_n20596_, new_n20597_, new_n20598_, new_n20599_, new_n20600_,
    new_n20601_, new_n20602_, new_n20603_, new_n20604_, new_n20605_,
    new_n20606_, new_n20607_, new_n20608_, new_n20609_, new_n20610_,
    new_n20611_, new_n20612_, new_n20613_, new_n20614_, new_n20615_,
    new_n20616_, new_n20617_, new_n20618_, new_n20619_, new_n20620_,
    new_n20621_, new_n20622_, new_n20623_, new_n20624_, new_n20625_,
    new_n20626_, new_n20627_, new_n20628_, new_n20629_, new_n20630_,
    new_n20631_, new_n20632_, new_n20633_, new_n20634_, new_n20635_,
    new_n20636_, new_n20637_, new_n20638_, new_n20639_, new_n20640_,
    new_n20641_, new_n20642_, new_n20643_, new_n20644_, new_n20645_,
    new_n20646_, new_n20647_, new_n20648_, new_n20649_, new_n20650_,
    new_n20651_, new_n20652_, new_n20653_, new_n20654_, new_n20655_,
    new_n20656_, new_n20657_, new_n20658_, new_n20659_, new_n20660_,
    new_n20661_, new_n20662_, new_n20663_, new_n20664_, new_n20665_,
    new_n20666_, new_n20667_, new_n20668_, new_n20669_, new_n20670_,
    new_n20671_, new_n20672_, new_n20673_, new_n20674_, new_n20675_,
    new_n20676_, new_n20677_, new_n20678_, new_n20679_, new_n20680_,
    new_n20681_, new_n20682_, new_n20683_, new_n20684_, new_n20685_,
    new_n20686_, new_n20687_, new_n20688_, new_n20689_, new_n20690_,
    new_n20691_, new_n20692_, new_n20693_, new_n20694_, new_n20695_,
    new_n20696_, new_n20697_, new_n20698_, new_n20699_, new_n20700_,
    new_n20701_, new_n20702_, new_n20703_, new_n20704_, new_n20705_,
    new_n20706_, new_n20707_, new_n20708_, new_n20709_, new_n20710_,
    new_n20711_, new_n20712_, new_n20713_, new_n20714_, new_n20715_,
    new_n20716_, new_n20717_, new_n20718_, new_n20719_, new_n20720_,
    new_n20721_, new_n20722_, new_n20723_, new_n20724_, new_n20725_,
    new_n20726_, new_n20727_, new_n20728_, new_n20729_, new_n20730_,
    new_n20731_, new_n20732_, new_n20733_, new_n20734_, new_n20735_,
    new_n20736_, new_n20737_, new_n20738_, new_n20739_, new_n20740_,
    new_n20741_, new_n20742_, new_n20743_, new_n20744_, new_n20745_,
    new_n20746_, new_n20747_, new_n20748_, new_n20749_, new_n20750_,
    new_n20751_, new_n20752_, new_n20753_, new_n20754_, new_n20755_,
    new_n20756_, new_n20757_, new_n20758_, new_n20759_, new_n20760_,
    new_n20761_, new_n20762_, new_n20763_, new_n20764_, new_n20765_,
    new_n20766_, new_n20767_, new_n20768_, new_n20769_, new_n20770_,
    new_n20771_, new_n20772_, new_n20773_, new_n20774_, new_n20775_,
    new_n20776_, new_n20777_, new_n20778_, new_n20779_, new_n20780_,
    new_n20781_, new_n20782_, new_n20783_, new_n20784_, new_n20785_,
    new_n20786_, new_n20787_, new_n20788_, new_n20789_, new_n20790_,
    new_n20791_, new_n20792_, new_n20793_, new_n20794_, new_n20795_,
    new_n20796_, new_n20797_, new_n20798_, new_n20799_, new_n20800_,
    new_n20801_, new_n20802_, new_n20803_, new_n20804_, new_n20805_,
    new_n20806_, new_n20807_, new_n20808_, new_n20809_, new_n20810_,
    new_n20811_, new_n20812_, new_n20813_, new_n20814_, new_n20815_,
    new_n20816_, new_n20817_, new_n20818_, new_n20819_, new_n20820_,
    new_n20821_, new_n20822_, new_n20823_, new_n20824_, new_n20825_,
    new_n20826_, new_n20827_, new_n20828_, new_n20829_, new_n20830_,
    new_n20831_, new_n20832_, new_n20833_, new_n20834_, new_n20835_,
    new_n20836_, new_n20837_, new_n20838_, new_n20839_, new_n20840_,
    new_n20841_, new_n20842_, new_n20843_, new_n20844_, new_n20845_,
    new_n20846_, new_n20847_, new_n20848_, new_n20849_, new_n20850_,
    new_n20851_, new_n20852_, new_n20853_, new_n20854_, new_n20855_,
    new_n20856_, new_n20857_, new_n20858_, new_n20859_, new_n20860_,
    new_n20861_, new_n20862_, new_n20863_, new_n20864_, new_n20865_,
    new_n20866_, new_n20867_, new_n20868_, new_n20869_, new_n20870_,
    new_n20871_, new_n20872_, new_n20873_, new_n20874_, new_n20875_,
    new_n20876_, new_n20877_, new_n20878_, new_n20879_, new_n20880_,
    new_n20881_, new_n20882_, new_n20883_, new_n20884_, new_n20885_,
    new_n20886_, new_n20887_, new_n20888_, new_n20889_, new_n20890_,
    new_n20891_, new_n20892_, new_n20893_, new_n20894_, new_n20895_,
    new_n20896_, new_n20897_, new_n20898_, new_n20899_, new_n20900_,
    new_n20901_, new_n20902_, new_n20903_, new_n20904_, new_n20905_,
    new_n20906_, new_n20907_, new_n20908_, new_n20909_, new_n20910_,
    new_n20911_, new_n20912_, new_n20913_, new_n20914_, new_n20915_,
    new_n20916_, new_n20917_, new_n20918_, new_n20919_, new_n20920_,
    new_n20921_, new_n20922_, new_n20923_, new_n20924_, new_n20925_,
    new_n20926_, new_n20927_, new_n20928_, new_n20929_, new_n20930_,
    new_n20931_, new_n20932_, new_n20933_, new_n20934_, new_n20935_,
    new_n20936_, new_n20937_, new_n20938_, new_n20939_, new_n20940_,
    new_n20941_, new_n20942_, new_n20943_, new_n20944_, new_n20945_,
    new_n20946_, new_n20947_, new_n20948_, new_n20949_, new_n20950_,
    new_n20951_, new_n20952_, new_n20953_, new_n20954_, new_n20955_,
    new_n20956_, new_n20957_, new_n20958_, new_n20959_, new_n20960_,
    new_n20961_, new_n20962_, new_n20963_, new_n20964_, new_n20965_,
    new_n20966_, new_n20967_, new_n20968_, new_n20969_, new_n20970_,
    new_n20971_, new_n20972_, new_n20973_, new_n20974_, new_n20975_,
    new_n20976_, new_n20977_, new_n20978_, new_n20979_, new_n20980_,
    new_n20981_, new_n20982_, new_n20983_, new_n20984_, new_n20985_,
    new_n20986_, new_n20987_, new_n20988_, new_n20989_, new_n20990_,
    new_n20991_, new_n20992_, new_n20993_, new_n20994_, new_n20995_,
    new_n20996_, new_n20997_, new_n20998_, new_n20999_, new_n21000_,
    new_n21001_, new_n21002_, new_n21003_, new_n21004_, new_n21005_,
    new_n21006_, new_n21007_, new_n21008_, new_n21009_, new_n21010_,
    new_n21011_, new_n21012_, new_n21013_, new_n21014_, new_n21015_,
    new_n21016_, new_n21017_, new_n21018_, new_n21019_, new_n21020_,
    new_n21021_, new_n21022_, new_n21023_, new_n21024_, new_n21025_,
    new_n21026_, new_n21027_, new_n21028_, new_n21029_, new_n21030_,
    new_n21031_, new_n21032_, new_n21033_, new_n21034_, new_n21035_,
    new_n21036_, new_n21037_, new_n21038_, new_n21039_, new_n21040_,
    new_n21041_, new_n21042_, new_n21043_, new_n21044_, new_n21045_,
    new_n21046_, new_n21047_, new_n21048_, new_n21049_, new_n21050_,
    new_n21051_, new_n21052_, new_n21053_, new_n21054_, new_n21055_,
    new_n21056_, new_n21057_, new_n21058_, new_n21059_, new_n21060_,
    new_n21061_, new_n21062_, new_n21063_, new_n21064_, new_n21065_,
    new_n21066_, new_n21067_, new_n21068_, new_n21069_, new_n21070_,
    new_n21071_, new_n21072_, new_n21073_, new_n21074_, new_n21075_,
    new_n21076_, new_n21077_, new_n21078_, new_n21079_, new_n21080_,
    new_n21081_, new_n21082_, new_n21083_, new_n21084_, new_n21085_,
    new_n21086_, new_n21087_, new_n21088_, new_n21089_, new_n21090_,
    new_n21091_, new_n21092_, new_n21093_, new_n21094_, new_n21095_,
    new_n21096_, new_n21097_, new_n21098_, new_n21099_, new_n21100_,
    new_n21101_, new_n21102_, new_n21103_, new_n21104_, new_n21105_,
    new_n21106_, new_n21107_, new_n21108_, new_n21109_, new_n21110_,
    new_n21111_, new_n21112_, new_n21113_, new_n21114_, new_n21115_,
    new_n21116_, new_n21117_, new_n21118_, new_n21119_, new_n21120_,
    new_n21121_, new_n21122_, new_n21123_, new_n21124_, new_n21125_,
    new_n21126_, new_n21127_, new_n21128_, new_n21129_, new_n21130_,
    new_n21131_, new_n21132_, new_n21133_, new_n21134_, new_n21135_,
    new_n21136_, new_n21137_, new_n21138_, new_n21139_, new_n21140_,
    new_n21141_, new_n21142_, new_n21143_, new_n21144_, new_n21145_,
    new_n21146_, new_n21147_, new_n21148_, new_n21149_, new_n21150_,
    new_n21151_, new_n21152_, new_n21153_, new_n21154_, new_n21155_,
    new_n21156_, new_n21157_, new_n21158_, new_n21159_, new_n21160_,
    new_n21161_, new_n21162_, new_n21163_, new_n21164_, new_n21165_,
    new_n21166_, new_n21167_, new_n21168_, new_n21169_, new_n21170_,
    new_n21171_, new_n21172_, new_n21173_, new_n21174_, new_n21175_,
    new_n21176_, new_n21177_, new_n21178_, new_n21179_, new_n21180_,
    new_n21181_, new_n21182_, new_n21183_, new_n21184_, new_n21185_,
    new_n21186_, new_n21187_, new_n21188_, new_n21189_, new_n21190_,
    new_n21191_, new_n21192_, new_n21193_, new_n21194_, new_n21195_,
    new_n21196_, new_n21197_, new_n21198_, new_n21199_, new_n21200_,
    new_n21201_, new_n21202_, new_n21203_, new_n21204_, new_n21205_,
    new_n21206_, new_n21207_, new_n21208_, new_n21209_, new_n21210_,
    new_n21211_, new_n21212_, new_n21213_, new_n21214_, new_n21215_,
    new_n21216_, new_n21217_, new_n21218_, new_n21219_, new_n21220_,
    new_n21221_, new_n21222_, new_n21223_, new_n21224_, new_n21225_,
    new_n21226_, new_n21227_, new_n21228_, new_n21229_, new_n21230_,
    new_n21231_, new_n21232_, new_n21233_, new_n21234_, new_n21235_,
    new_n21236_, new_n21237_, new_n21238_, new_n21239_, new_n21240_,
    new_n21241_, new_n21242_, new_n21243_, new_n21244_, new_n21245_,
    new_n21246_, new_n21247_, new_n21248_, new_n21249_, new_n21250_,
    new_n21251_, new_n21252_, new_n21253_, new_n21254_, new_n21255_,
    new_n21256_, new_n21257_, new_n21258_, new_n21259_, new_n21260_,
    new_n21261_, new_n21262_, new_n21263_, new_n21264_, new_n21265_,
    new_n21266_, new_n21267_, new_n21268_, new_n21269_, new_n21270_,
    new_n21271_, new_n21272_, new_n21273_, new_n21274_, new_n21275_,
    new_n21276_, new_n21277_, new_n21278_, new_n21279_, new_n21280_,
    new_n21281_, new_n21282_, new_n21283_, new_n21284_, new_n21285_,
    new_n21286_, new_n21287_, new_n21288_, new_n21289_, new_n21290_,
    new_n21291_, new_n21292_, new_n21293_, new_n21294_, new_n21295_,
    new_n21296_, new_n21297_, new_n21298_, new_n21299_, new_n21300_,
    new_n21301_, new_n21302_, new_n21303_, new_n21304_, new_n21305_,
    new_n21306_, new_n21307_, new_n21308_, new_n21309_, new_n21310_,
    new_n21311_, new_n21312_, new_n21313_, new_n21314_, new_n21315_,
    new_n21316_, new_n21317_, new_n21318_, new_n21319_, new_n21320_,
    new_n21321_, new_n21322_, new_n21323_, new_n21324_, new_n21325_,
    new_n21326_, new_n21327_, new_n21328_, new_n21329_, new_n21330_,
    new_n21331_, new_n21332_, new_n21333_, new_n21334_, new_n21335_,
    new_n21336_, new_n21337_, new_n21338_, new_n21339_, new_n21340_,
    new_n21341_, new_n21342_, new_n21343_, new_n21344_, new_n21345_,
    new_n21346_, new_n21347_, new_n21348_, new_n21349_, new_n21350_,
    new_n21351_, new_n21352_, new_n21353_, new_n21354_, new_n21355_,
    new_n21356_, new_n21357_, new_n21358_, new_n21359_, new_n21360_,
    new_n21361_, new_n21362_, new_n21363_, new_n21364_, new_n21365_,
    new_n21366_, new_n21367_, new_n21368_, new_n21369_, new_n21370_,
    new_n21371_, new_n21372_, new_n21373_, new_n21374_, new_n21375_,
    new_n21376_, new_n21377_, new_n21378_, new_n21379_, new_n21380_,
    new_n21381_, new_n21382_, new_n21383_, new_n21384_, new_n21385_,
    new_n21386_, new_n21387_, new_n21388_, new_n21389_, new_n21390_,
    new_n21391_, new_n21392_, new_n21393_, new_n21394_, new_n21395_,
    new_n21396_, new_n21397_, new_n21398_, new_n21399_, new_n21400_,
    new_n21401_, new_n21402_, new_n21403_, new_n21404_, new_n21405_,
    new_n21406_, new_n21407_, new_n21408_, new_n21409_, new_n21410_,
    new_n21411_, new_n21412_, new_n21413_, new_n21414_, new_n21415_,
    new_n21416_, new_n21417_, new_n21418_, new_n21419_, new_n21420_,
    new_n21421_, new_n21422_, new_n21423_, new_n21424_, new_n21425_,
    new_n21426_, new_n21427_, new_n21428_, new_n21429_, new_n21430_,
    new_n21431_, new_n21432_, new_n21433_, new_n21434_, new_n21435_,
    new_n21436_, new_n21437_, new_n21438_, new_n21439_, new_n21440_,
    new_n21441_, new_n21442_, new_n21443_, new_n21444_, new_n21445_,
    new_n21446_, new_n21447_, new_n21448_, new_n21449_, new_n21450_,
    new_n21451_, new_n21452_, new_n21453_, new_n21454_, new_n21455_,
    new_n21456_, new_n21457_, new_n21458_, new_n21459_, new_n21460_,
    new_n21461_, new_n21462_, new_n21463_, new_n21464_, new_n21465_,
    new_n21466_, new_n21467_, new_n21468_, new_n21469_, new_n21470_,
    new_n21471_, new_n21472_, new_n21473_, new_n21474_, new_n21475_,
    new_n21476_, new_n21477_, new_n21478_, new_n21479_, new_n21480_,
    new_n21481_, new_n21482_, new_n21483_, new_n21484_, new_n21485_,
    new_n21486_, new_n21487_, new_n21488_, new_n21489_, new_n21490_,
    new_n21491_, new_n21492_, new_n21493_, new_n21494_, new_n21495_,
    new_n21496_, new_n21497_, new_n21498_, new_n21499_, new_n21500_,
    new_n21501_, new_n21502_, new_n21503_, new_n21504_, new_n21505_,
    new_n21506_, new_n21507_, new_n21508_, new_n21509_, new_n21510_,
    new_n21511_, new_n21512_, new_n21513_, new_n21514_, new_n21515_,
    new_n21516_, new_n21517_, new_n21518_, new_n21519_, new_n21520_,
    new_n21521_, new_n21522_, new_n21523_, new_n21524_, new_n21525_,
    new_n21526_, new_n21527_, new_n21528_, new_n21529_, new_n21530_,
    new_n21531_, new_n21532_, new_n21533_, new_n21534_, new_n21535_,
    new_n21536_, new_n21537_, new_n21538_, new_n21539_, new_n21540_,
    new_n21541_, new_n21542_, new_n21543_, new_n21544_, new_n21545_,
    new_n21546_, new_n21547_, new_n21548_, new_n21549_, new_n21550_,
    new_n21551_, new_n21552_, new_n21553_, new_n21554_, new_n21555_,
    new_n21556_, new_n21557_, new_n21558_, new_n21559_, new_n21560_,
    new_n21561_, new_n21562_, new_n21563_, new_n21564_, new_n21565_,
    new_n21566_, new_n21567_, new_n21568_, new_n21569_, new_n21570_,
    new_n21571_, new_n21572_, new_n21573_, new_n21574_, new_n21575_,
    new_n21576_, new_n21577_, new_n21578_, new_n21579_, new_n21580_,
    new_n21581_, new_n21582_, new_n21583_, new_n21584_, new_n21585_,
    new_n21586_, new_n21587_, new_n21588_, new_n21589_, new_n21590_,
    new_n21591_, new_n21592_, new_n21593_, new_n21594_, new_n21595_,
    new_n21596_, new_n21597_, new_n21598_, new_n21599_, new_n21600_,
    new_n21601_, new_n21602_, new_n21603_, new_n21604_, new_n21605_,
    new_n21606_, new_n21607_, new_n21608_, new_n21609_, new_n21610_,
    new_n21611_, new_n21612_, new_n21613_, new_n21614_, new_n21615_,
    new_n21616_, new_n21617_, new_n21618_, new_n21619_, new_n21620_,
    new_n21621_, new_n21622_, new_n21623_, new_n21624_, new_n21625_,
    new_n21626_, new_n21627_, new_n21628_, new_n21629_, new_n21630_,
    new_n21631_, new_n21632_, new_n21633_, new_n21634_, new_n21635_,
    new_n21636_, new_n21637_, new_n21638_, new_n21639_, new_n21640_,
    new_n21641_, new_n21642_, new_n21643_, new_n21644_, new_n21645_,
    new_n21646_, new_n21647_, new_n21648_, new_n21649_, new_n21650_,
    new_n21651_, new_n21652_, new_n21653_, new_n21654_, new_n21655_,
    new_n21656_, new_n21657_, new_n21658_, new_n21659_, new_n21660_,
    new_n21661_, new_n21662_, new_n21663_, new_n21664_, new_n21665_,
    new_n21666_, new_n21667_, new_n21668_, new_n21669_, new_n21670_,
    new_n21671_, new_n21672_, new_n21673_, new_n21674_, new_n21675_,
    new_n21676_, new_n21677_, new_n21678_, new_n21679_, new_n21680_,
    new_n21681_, new_n21682_, new_n21683_, new_n21684_, new_n21685_,
    new_n21686_, new_n21687_, new_n21688_, new_n21689_, new_n21690_,
    new_n21691_, new_n21692_, new_n21693_, new_n21694_, new_n21695_,
    new_n21696_, new_n21697_, new_n21698_, new_n21699_, new_n21700_,
    new_n21701_, new_n21702_, new_n21703_, new_n21704_, new_n21705_,
    new_n21706_, new_n21707_, new_n21708_, new_n21709_, new_n21710_,
    new_n21711_, new_n21712_, new_n21713_, new_n21714_, new_n21715_,
    new_n21716_, new_n21717_, new_n21718_, new_n21719_, new_n21720_,
    new_n21721_, new_n21722_, new_n21723_, new_n21724_, new_n21725_,
    new_n21726_, new_n21727_, new_n21728_, new_n21729_, new_n21730_,
    new_n21731_, new_n21732_, new_n21733_, new_n21734_, new_n21735_,
    new_n21736_, new_n21737_, new_n21738_, new_n21739_, new_n21740_,
    new_n21741_, new_n21742_, new_n21743_, new_n21744_, new_n21745_,
    new_n21746_, new_n21747_, new_n21748_, new_n21749_, new_n21750_,
    new_n21751_, new_n21752_, new_n21753_, new_n21754_, new_n21755_,
    new_n21756_, new_n21757_, new_n21758_, new_n21759_, new_n21760_,
    new_n21761_, new_n21762_, new_n21763_, new_n21764_, new_n21765_,
    new_n21766_, new_n21767_, new_n21768_, new_n21769_, new_n21770_,
    new_n21771_, new_n21772_, new_n21773_, new_n21774_, new_n21775_,
    new_n21776_, new_n21777_, new_n21778_, new_n21779_, new_n21780_,
    new_n21781_, new_n21782_, new_n21783_, new_n21784_, new_n21785_,
    new_n21786_, new_n21787_, new_n21788_, new_n21789_, new_n21790_,
    new_n21791_, new_n21792_, new_n21793_, new_n21794_, new_n21795_,
    new_n21796_, new_n21797_, new_n21798_, new_n21799_, new_n21800_,
    new_n21801_, new_n21802_, new_n21803_, new_n21804_, new_n21805_,
    new_n21806_, new_n21807_, new_n21808_, new_n21809_, new_n21810_,
    new_n21811_, new_n21812_, new_n21813_, new_n21814_, new_n21815_,
    new_n21816_, new_n21817_, new_n21818_, new_n21819_, new_n21820_,
    new_n21821_, new_n21822_, new_n21823_, new_n21824_, new_n21825_,
    new_n21826_, new_n21827_, new_n21828_, new_n21829_, new_n21830_,
    new_n21831_, new_n21832_, new_n21833_, new_n21834_, new_n21835_,
    new_n21836_, new_n21837_, new_n21838_, new_n21839_, new_n21840_,
    new_n21841_, new_n21842_, new_n21843_, new_n21844_, new_n21845_,
    new_n21846_, new_n21847_, new_n21848_, new_n21849_, new_n21850_,
    new_n21851_, new_n21852_, new_n21853_, new_n21854_, new_n21855_,
    new_n21856_, new_n21857_, new_n21858_, new_n21859_, new_n21860_,
    new_n21861_, new_n21862_, new_n21863_, new_n21864_, new_n21865_,
    new_n21866_, new_n21867_, new_n21868_, new_n21869_, new_n21870_,
    new_n21871_, new_n21872_, new_n21873_, new_n21874_, new_n21875_,
    new_n21876_, new_n21877_, new_n21878_, new_n21879_, new_n21880_,
    new_n21881_, new_n21882_, new_n21883_, new_n21884_, new_n21885_,
    new_n21886_, new_n21887_, new_n21888_, new_n21889_, new_n21890_,
    new_n21891_, new_n21892_, new_n21893_, new_n21894_, new_n21895_,
    new_n21896_, new_n21897_, new_n21898_, new_n21899_, new_n21900_,
    new_n21901_, new_n21902_, new_n21903_, new_n21904_, new_n21905_,
    new_n21906_, new_n21907_, new_n21908_, new_n21909_, new_n21910_,
    new_n21911_, new_n21912_, new_n21913_, new_n21914_, new_n21915_,
    new_n21916_, new_n21917_, new_n21918_, new_n21919_, new_n21920_,
    new_n21921_, new_n21922_, new_n21923_, new_n21924_, new_n21925_,
    new_n21926_, new_n21927_, new_n21928_, new_n21929_, new_n21930_,
    new_n21931_, new_n21932_, new_n21933_, new_n21934_, new_n21935_,
    new_n21936_, new_n21937_, new_n21938_, new_n21939_, new_n21940_,
    new_n21941_, new_n21942_, new_n21943_, new_n21944_, new_n21945_,
    new_n21946_, new_n21947_, new_n21948_, new_n21949_, new_n21950_,
    new_n21951_, new_n21952_, new_n21953_, new_n21954_, new_n21955_,
    new_n21956_, new_n21957_, new_n21958_, new_n21959_, new_n21960_,
    new_n21961_, new_n21962_, new_n21963_, new_n21964_, new_n21965_,
    new_n21966_, new_n21967_, new_n21968_, new_n21969_, new_n21970_,
    new_n21971_, new_n21972_, new_n21973_, new_n21974_, new_n21975_,
    new_n21976_, new_n21977_, new_n21978_, new_n21979_, new_n21980_,
    new_n21981_, new_n21982_, new_n21983_, new_n21984_, new_n21985_,
    new_n21986_, new_n21987_, new_n21988_, new_n21989_, new_n21990_,
    new_n21991_, new_n21992_, new_n21993_, new_n21994_, new_n21995_,
    new_n21996_, new_n21997_, new_n21998_, new_n21999_, new_n22000_,
    new_n22001_, new_n22002_, new_n22003_, new_n22004_, new_n22005_,
    new_n22006_, new_n22007_, new_n22008_, new_n22009_, new_n22010_,
    new_n22011_, new_n22012_, new_n22013_, new_n22014_, new_n22015_,
    new_n22016_, new_n22017_, new_n22018_, new_n22019_, new_n22020_,
    new_n22021_, new_n22022_, new_n22023_, new_n22024_, new_n22025_,
    new_n22026_, new_n22027_, new_n22028_, new_n22029_, new_n22030_,
    new_n22031_, new_n22032_, new_n22033_, new_n22034_, new_n22035_,
    new_n22036_, new_n22037_, new_n22038_, new_n22039_, new_n22040_,
    new_n22041_, new_n22042_, new_n22043_, new_n22044_, new_n22045_,
    new_n22046_, new_n22047_, new_n22048_, new_n22049_, new_n22050_,
    new_n22051_, new_n22052_, new_n22053_, new_n22054_, new_n22055_,
    new_n22056_, new_n22057_, new_n22058_, new_n22059_, new_n22060_,
    new_n22061_, new_n22062_, new_n22063_, new_n22064_, new_n22065_,
    new_n22066_, new_n22067_, new_n22068_, new_n22069_, new_n22070_,
    new_n22071_, new_n22072_, new_n22073_, new_n22074_, new_n22075_,
    new_n22076_, new_n22077_, new_n22078_, new_n22079_, new_n22080_,
    new_n22081_, new_n22082_, new_n22083_, new_n22084_, new_n22085_,
    new_n22086_, new_n22087_, new_n22088_, new_n22089_, new_n22090_,
    new_n22091_, new_n22092_, new_n22093_, new_n22094_, new_n22095_,
    new_n22096_, new_n22097_, new_n22098_, new_n22099_, new_n22100_,
    new_n22101_, new_n22102_, new_n22103_, new_n22104_, new_n22105_,
    new_n22106_, new_n22107_, new_n22108_, new_n22109_, new_n22110_,
    new_n22111_, new_n22112_, new_n22113_, new_n22114_, new_n22115_,
    new_n22116_, new_n22117_, new_n22118_, new_n22119_, new_n22120_,
    new_n22121_, new_n22122_, new_n22123_, new_n22124_, new_n22125_,
    new_n22126_, new_n22127_, new_n22128_, new_n22129_, new_n22130_,
    new_n22131_, new_n22132_, new_n22133_, new_n22134_, new_n22135_,
    new_n22136_, new_n22137_, new_n22138_, new_n22139_, new_n22140_,
    new_n22141_, new_n22142_, new_n22143_, new_n22144_, new_n22145_,
    new_n22146_, new_n22147_, new_n22148_, new_n22149_, new_n22150_,
    new_n22151_, new_n22152_, new_n22153_, new_n22154_, new_n22155_,
    new_n22156_, new_n22157_, new_n22158_, new_n22159_, new_n22160_,
    new_n22161_, new_n22162_, new_n22163_, new_n22164_, new_n22165_,
    new_n22166_, new_n22167_, new_n22168_, new_n22169_, new_n22170_,
    new_n22171_, new_n22172_, new_n22173_, new_n22174_, new_n22175_,
    new_n22176_, new_n22177_, new_n22178_, new_n22179_, new_n22180_,
    new_n22181_, new_n22182_, new_n22183_, new_n22184_, new_n22185_,
    new_n22186_, new_n22187_, new_n22188_, new_n22189_, new_n22190_,
    new_n22191_, new_n22192_, new_n22193_, new_n22194_, new_n22195_,
    new_n22196_, new_n22197_, new_n22198_, new_n22199_, new_n22200_,
    new_n22201_, new_n22202_, new_n22203_, new_n22204_, new_n22205_,
    new_n22206_, new_n22207_, new_n22208_, new_n22209_, new_n22210_,
    new_n22211_, new_n22212_, new_n22213_, new_n22214_, new_n22215_,
    new_n22216_, new_n22217_, new_n22218_, new_n22219_, new_n22220_,
    new_n22221_, new_n22222_, new_n22223_, new_n22224_, new_n22225_,
    new_n22226_, new_n22227_, new_n22228_, new_n22229_, new_n22230_,
    new_n22231_, new_n22232_, new_n22233_, new_n22234_, new_n22235_,
    new_n22236_, new_n22237_, new_n22238_, new_n22239_, new_n22240_,
    new_n22241_, new_n22242_, new_n22243_, new_n22244_, new_n22245_,
    new_n22246_, new_n22247_, new_n22248_, new_n22249_, new_n22250_,
    new_n22251_, new_n22252_, new_n22253_, new_n22254_, new_n22255_,
    new_n22256_, new_n22257_, new_n22258_, new_n22259_, new_n22260_,
    new_n22261_, new_n22262_, new_n22263_, new_n22264_, new_n22265_,
    new_n22266_, new_n22267_, new_n22268_, new_n22269_, new_n22270_,
    new_n22271_, new_n22272_, new_n22273_, new_n22274_, new_n22275_,
    new_n22276_, new_n22277_, new_n22278_, new_n22279_, new_n22280_,
    new_n22281_, new_n22282_, new_n22283_, new_n22284_, new_n22285_,
    new_n22286_, new_n22287_, new_n22288_, new_n22289_, new_n22290_,
    new_n22291_, new_n22292_, new_n22293_, new_n22294_, new_n22295_,
    new_n22296_, new_n22297_, new_n22298_, new_n22299_, new_n22300_,
    new_n22301_, new_n22302_, new_n22303_, new_n22304_, new_n22305_,
    new_n22306_, new_n22307_, new_n22308_, new_n22309_, new_n22310_,
    new_n22311_, new_n22312_, new_n22313_, new_n22314_, new_n22315_,
    new_n22316_, new_n22317_, new_n22318_, new_n22319_, new_n22320_,
    new_n22321_, new_n22322_, new_n22323_, new_n22324_, new_n22325_,
    new_n22326_, new_n22327_, new_n22328_, new_n22329_, new_n22330_,
    new_n22331_, new_n22332_, new_n22333_, new_n22334_, new_n22335_,
    new_n22336_, new_n22337_, new_n22338_, new_n22339_, new_n22340_,
    new_n22341_, new_n22342_, new_n22343_, new_n22344_, new_n22345_,
    new_n22346_, new_n22347_, new_n22348_, new_n22349_, new_n22350_,
    new_n22351_, new_n22352_, new_n22353_, new_n22354_, new_n22355_,
    new_n22356_, new_n22357_, new_n22358_, new_n22359_, new_n22360_,
    new_n22361_, new_n22362_, new_n22363_, new_n22364_, new_n22365_,
    new_n22366_, new_n22367_, new_n22368_, new_n22369_, new_n22370_,
    new_n22371_, new_n22372_, new_n22373_, new_n22374_, new_n22375_,
    new_n22376_, new_n22377_, new_n22378_, new_n22379_, new_n22380_,
    new_n22381_, new_n22382_, new_n22383_, new_n22384_, new_n22385_,
    new_n22386_, new_n22387_, new_n22388_, new_n22389_, new_n22390_,
    new_n22391_, new_n22392_, new_n22393_, new_n22394_, new_n22395_,
    new_n22396_, new_n22397_, new_n22398_, new_n22399_, new_n22400_,
    new_n22401_, new_n22402_, new_n22403_, new_n22404_, new_n22405_,
    new_n22406_, new_n22407_, new_n22408_, new_n22409_, new_n22410_,
    new_n22411_, new_n22412_, new_n22413_, new_n22414_, new_n22415_,
    new_n22416_, new_n22417_, new_n22418_, new_n22419_, new_n22420_,
    new_n22421_, new_n22422_, new_n22423_, new_n22424_, new_n22425_,
    new_n22426_, new_n22427_, new_n22428_, new_n22429_, new_n22430_,
    new_n22431_, new_n22432_, new_n22433_, new_n22434_, new_n22435_,
    new_n22436_, new_n22437_, new_n22438_, new_n22439_, new_n22440_,
    new_n22441_, new_n22442_, new_n22443_, new_n22444_, new_n22445_,
    new_n22446_, new_n22447_, new_n22448_, new_n22449_, new_n22450_,
    new_n22451_, new_n22452_, new_n22453_, new_n22454_, new_n22455_,
    new_n22456_, new_n22457_, new_n22458_, new_n22459_, new_n22460_,
    new_n22461_, new_n22462_, new_n22463_, new_n22464_, new_n22465_,
    new_n22466_, new_n22467_, new_n22468_, new_n22469_, new_n22470_,
    new_n22471_, new_n22472_, new_n22473_, new_n22474_, new_n22475_,
    new_n22476_, new_n22477_, new_n22478_, new_n22479_, new_n22480_,
    new_n22481_, new_n22482_, new_n22483_, new_n22484_, new_n22485_,
    new_n22486_, new_n22487_, new_n22488_, new_n22489_, new_n22490_,
    new_n22491_, new_n22492_, new_n22493_, new_n22494_, new_n22495_,
    new_n22496_, new_n22497_, new_n22498_, new_n22499_, new_n22500_,
    new_n22501_, new_n22502_, new_n22503_, new_n22504_, new_n22505_,
    new_n22506_, new_n22507_, new_n22508_, new_n22509_, new_n22510_,
    new_n22511_, new_n22512_, new_n22513_, new_n22514_, new_n22515_,
    new_n22516_, new_n22517_, new_n22518_, new_n22519_, new_n22520_,
    new_n22521_, new_n22522_, new_n22523_, new_n22524_, new_n22525_,
    new_n22526_, new_n22527_, new_n22528_, new_n22529_, new_n22530_,
    new_n22531_, new_n22532_, new_n22533_, new_n22534_, new_n22535_,
    new_n22536_, new_n22537_, new_n22538_, new_n22539_, new_n22540_,
    new_n22541_, new_n22542_, new_n22543_, new_n22544_, new_n22545_,
    new_n22546_, new_n22547_, new_n22548_, new_n22549_, new_n22550_,
    new_n22551_, new_n22552_, new_n22553_, new_n22554_, new_n22555_,
    new_n22556_, new_n22557_, new_n22558_, new_n22559_, new_n22560_,
    new_n22561_, new_n22562_, new_n22563_, new_n22564_, new_n22565_,
    new_n22566_, new_n22567_, new_n22568_, new_n22569_, new_n22570_,
    new_n22571_, new_n22572_, new_n22573_, new_n22574_, new_n22575_,
    new_n22576_, new_n22577_, new_n22578_, new_n22579_, new_n22580_,
    new_n22581_, new_n22582_, new_n22583_, new_n22584_, new_n22585_,
    new_n22586_, new_n22587_, new_n22588_, new_n22589_, new_n22590_,
    new_n22591_, new_n22592_, new_n22593_, new_n22594_, new_n22595_,
    new_n22596_, new_n22597_, new_n22598_, new_n22599_, new_n22600_,
    new_n22601_, new_n22602_, new_n22603_, new_n22604_, new_n22605_,
    new_n22606_, new_n22607_, new_n22608_, new_n22609_, new_n22610_,
    new_n22611_, new_n22612_, new_n22613_, new_n22614_, new_n22615_,
    new_n22616_, new_n22617_, new_n22618_, new_n22619_, new_n22620_,
    new_n22621_, new_n22622_, new_n22623_, new_n22624_, new_n22625_,
    new_n22626_, new_n22627_, new_n22628_, new_n22629_, new_n22630_,
    new_n22631_, new_n22632_, new_n22633_, new_n22634_, new_n22635_,
    new_n22636_, new_n22637_, new_n22638_, new_n22639_, new_n22640_,
    new_n22641_, new_n22642_, new_n22643_, new_n22644_, new_n22645_,
    new_n22646_, new_n22647_, new_n22648_, new_n22649_, new_n22650_,
    new_n22651_, new_n22652_, new_n22653_, new_n22654_, new_n22655_,
    new_n22656_, new_n22657_, new_n22658_, new_n22659_, new_n22660_,
    new_n22661_, new_n22662_, new_n22663_, new_n22664_, new_n22665_,
    new_n22666_, new_n22667_, new_n22668_, new_n22669_, new_n22670_,
    new_n22671_, new_n22672_, new_n22673_, new_n22674_, new_n22675_,
    new_n22676_, new_n22677_, new_n22678_, new_n22679_, new_n22680_,
    new_n22681_, new_n22682_, new_n22683_, new_n22684_, new_n22685_,
    new_n22686_, new_n22687_, new_n22688_, new_n22689_, new_n22690_,
    new_n22691_, new_n22692_, new_n22693_, new_n22694_, new_n22695_,
    new_n22696_, new_n22697_, new_n22698_, new_n22699_, new_n22700_,
    new_n22701_, new_n22702_, new_n22703_, new_n22704_, new_n22705_,
    new_n22706_, new_n22707_, new_n22708_, new_n22709_, new_n22710_,
    new_n22711_, new_n22712_, new_n22713_, new_n22714_, new_n22715_,
    new_n22716_, new_n22717_, new_n22718_, new_n22719_, new_n22720_,
    new_n22721_, new_n22722_, new_n22723_, new_n22724_, new_n22725_,
    new_n22726_, new_n22727_, new_n22728_, new_n22729_, new_n22730_,
    new_n22731_, new_n22732_, new_n22733_, new_n22734_, new_n22735_,
    new_n22736_, new_n22737_, new_n22738_, new_n22739_, new_n22740_,
    new_n22741_, new_n22742_, new_n22743_, new_n22744_, new_n22745_,
    new_n22746_, new_n22747_, new_n22748_, new_n22749_, new_n22750_,
    new_n22751_, new_n22752_, new_n22753_, new_n22754_, new_n22755_,
    new_n22756_, new_n22757_, new_n22758_, new_n22759_, new_n22760_,
    new_n22761_, new_n22762_, new_n22763_, new_n22764_, new_n22765_,
    new_n22766_, new_n22767_, new_n22768_, new_n22769_, new_n22770_,
    new_n22771_, new_n22772_, new_n22773_, new_n22774_, new_n22775_,
    new_n22776_, new_n22777_, new_n22778_, new_n22779_, new_n22780_,
    new_n22781_, new_n22782_, new_n22783_, new_n22784_, new_n22785_,
    new_n22786_, new_n22787_, new_n22788_, new_n22789_, new_n22790_,
    new_n22791_, new_n22792_, new_n22793_, new_n22794_, new_n22795_,
    new_n22796_, new_n22797_, new_n22798_, new_n22799_, new_n22800_,
    new_n22801_, new_n22802_, new_n22803_, new_n22804_, new_n22805_,
    new_n22806_, new_n22807_, new_n22808_, new_n22809_, new_n22810_,
    new_n22811_, new_n22812_, new_n22813_, new_n22814_, new_n22815_,
    new_n22816_, new_n22817_, new_n22818_, new_n22819_, new_n22820_,
    new_n22821_, new_n22822_, new_n22823_, new_n22824_, new_n22825_,
    new_n22826_, new_n22827_, new_n22828_, new_n22829_, new_n22830_,
    new_n22831_, new_n22832_, new_n22833_, new_n22834_, new_n22835_,
    new_n22836_, new_n22837_, new_n22838_, new_n22839_, new_n22840_,
    new_n22841_, new_n22842_, new_n22843_, new_n22844_, new_n22845_,
    new_n22846_, new_n22847_, new_n22848_, new_n22849_, new_n22850_,
    new_n22851_, new_n22852_, new_n22853_, new_n22854_, new_n22855_,
    new_n22856_, new_n22857_, new_n22858_, new_n22859_, new_n22860_,
    new_n22861_, new_n22862_, new_n22863_, new_n22864_, new_n22865_,
    new_n22866_, new_n22867_, new_n22868_, new_n22869_, new_n22870_,
    new_n22871_, new_n22872_, new_n22873_, new_n22874_, new_n22875_,
    new_n22876_, new_n22877_, new_n22878_, new_n22879_, new_n22880_,
    new_n22881_, new_n22882_, new_n22883_, new_n22884_, new_n22885_,
    new_n22886_, new_n22887_, new_n22888_, new_n22889_, new_n22890_,
    new_n22891_, new_n22892_, new_n22893_, new_n22894_, new_n22895_,
    new_n22896_, new_n22897_, new_n22898_, new_n22899_, new_n22900_,
    new_n22901_, new_n22902_, new_n22903_, new_n22904_, new_n22905_,
    new_n22906_, new_n22907_, new_n22908_, new_n22909_, new_n22910_,
    new_n22911_, new_n22912_, new_n22913_, new_n22914_, new_n22915_,
    new_n22916_, new_n22917_, new_n22918_, new_n22919_, new_n22920_,
    new_n22921_, new_n22922_, new_n22923_, new_n22924_, new_n22925_,
    new_n22926_, new_n22927_, new_n22928_, new_n22929_, new_n22930_,
    new_n22931_, new_n22932_, new_n22933_, new_n22934_, new_n22935_,
    new_n22936_, new_n22937_, new_n22938_, new_n22939_, new_n22940_,
    new_n22941_, new_n22942_, new_n22943_, new_n22944_, new_n22945_,
    new_n22946_, new_n22947_, new_n22948_, new_n22949_, new_n22950_,
    new_n22951_, new_n22952_, new_n22953_, new_n22954_, new_n22955_,
    new_n22956_, new_n22957_, new_n22958_, new_n22959_, new_n22960_,
    new_n22961_, new_n22962_, new_n22963_, new_n22964_, new_n22965_,
    new_n22966_, new_n22967_, new_n22968_, new_n22969_, new_n22970_,
    new_n22971_, new_n22972_, new_n22973_, new_n22974_, new_n22975_,
    new_n22976_, new_n22977_, new_n22978_, new_n22979_, new_n22980_,
    new_n22981_, new_n22982_, new_n22983_, new_n22984_, new_n22985_,
    new_n22986_, new_n22987_, new_n22988_, new_n22989_, new_n22990_,
    new_n22991_, new_n22992_, new_n22993_, new_n22994_, new_n22995_,
    new_n22996_, new_n22997_, new_n22998_, new_n22999_, new_n23000_,
    new_n23001_, new_n23002_, new_n23003_, new_n23004_, new_n23005_,
    new_n23006_, new_n23007_, new_n23008_, new_n23009_, new_n23010_,
    new_n23011_, new_n23012_, new_n23013_, new_n23014_, new_n23015_,
    new_n23016_, new_n23017_, new_n23018_, new_n23019_, new_n23020_,
    new_n23021_, new_n23022_, new_n23023_, new_n23024_, new_n23025_,
    new_n23026_, new_n23027_, new_n23028_, new_n23029_, new_n23030_,
    new_n23031_, new_n23032_, new_n23033_, new_n23034_, new_n23035_,
    new_n23036_, new_n23037_, new_n23038_, new_n23039_, new_n23040_,
    new_n23041_, new_n23042_, new_n23043_, new_n23044_, new_n23045_,
    new_n23046_, new_n23047_, new_n23048_, new_n23049_, new_n23050_,
    new_n23051_, new_n23052_, new_n23053_, new_n23054_, new_n23055_,
    new_n23056_, new_n23057_, new_n23058_, new_n23059_, new_n23060_,
    new_n23061_, new_n23062_, new_n23063_, new_n23064_, new_n23065_,
    new_n23066_, new_n23067_, new_n23068_, new_n23069_, new_n23070_,
    new_n23071_, new_n23072_, new_n23073_, new_n23074_, new_n23075_,
    new_n23076_, new_n23077_, new_n23078_, new_n23079_, new_n23080_,
    new_n23081_, new_n23082_, new_n23083_, new_n23084_, new_n23085_,
    new_n23086_, new_n23087_, new_n23088_, new_n23089_, new_n23090_,
    new_n23091_, new_n23092_, new_n23093_, new_n23094_, new_n23095_,
    new_n23096_, new_n23097_, new_n23098_, new_n23099_, new_n23100_,
    new_n23101_, new_n23102_, new_n23103_, new_n23104_, new_n23105_,
    new_n23106_, new_n23107_, new_n23108_, new_n23109_, new_n23110_,
    new_n23111_, new_n23112_, new_n23113_, new_n23114_, new_n23115_,
    new_n23116_, new_n23117_, new_n23118_, new_n23119_, new_n23120_,
    new_n23121_, new_n23122_, new_n23123_, new_n23124_, new_n23125_,
    new_n23126_, new_n23127_, new_n23128_, new_n23129_, new_n23130_,
    new_n23131_, new_n23132_, new_n23133_, new_n23134_, new_n23135_,
    new_n23136_, new_n23137_, new_n23138_, new_n23139_, new_n23140_,
    new_n23141_, new_n23142_, new_n23143_, new_n23144_, new_n23145_,
    new_n23146_, new_n23147_, new_n23148_, new_n23149_, new_n23150_,
    new_n23151_, new_n23152_, new_n23153_, new_n23154_, new_n23155_,
    new_n23156_, new_n23157_, new_n23158_, new_n23159_, new_n23160_,
    new_n23161_, new_n23162_, new_n23163_, new_n23164_, new_n23165_,
    new_n23166_, new_n23167_, new_n23168_, new_n23169_, new_n23170_,
    new_n23171_, new_n23172_, new_n23173_, new_n23174_, new_n23175_,
    new_n23176_, new_n23177_, new_n23178_, new_n23179_, new_n23180_,
    new_n23181_, new_n23182_, new_n23183_, new_n23184_, new_n23185_,
    new_n23186_, new_n23187_, new_n23188_, new_n23189_, new_n23190_,
    new_n23191_, new_n23192_, new_n23193_, new_n23194_, new_n23195_,
    new_n23196_, new_n23197_, new_n23198_, new_n23199_, new_n23200_,
    new_n23201_, new_n23202_, new_n23203_, new_n23204_, new_n23205_,
    new_n23206_, new_n23207_, new_n23208_, new_n23209_, new_n23210_,
    new_n23211_, new_n23212_, new_n23213_, new_n23214_, new_n23215_,
    new_n23216_, new_n23217_, new_n23218_, new_n23219_, new_n23220_,
    new_n23221_, new_n23222_, new_n23223_, new_n23224_, new_n23225_,
    new_n23226_, new_n23227_, new_n23228_, new_n23229_, new_n23230_,
    new_n23231_, new_n23232_, new_n23233_, new_n23234_, new_n23235_,
    new_n23236_, new_n23237_, new_n23238_, new_n23239_, new_n23240_,
    new_n23241_, new_n23242_, new_n23243_, new_n23244_, new_n23245_,
    new_n23246_, new_n23247_, new_n23248_, new_n23249_, new_n23250_,
    new_n23251_, new_n23252_, new_n23253_, new_n23254_, new_n23255_,
    new_n23256_, new_n23257_, new_n23258_, new_n23259_, new_n23260_,
    new_n23261_, new_n23262_, new_n23263_, new_n23264_, new_n23265_,
    new_n23266_, new_n23267_, new_n23268_, new_n23269_, new_n23270_,
    new_n23271_, new_n23272_, new_n23273_, new_n23274_, new_n23275_,
    new_n23276_, new_n23277_, new_n23278_, new_n23279_, new_n23280_,
    new_n23281_, new_n23282_, new_n23283_, new_n23284_, new_n23285_,
    new_n23286_, new_n23287_, new_n23288_, new_n23289_, new_n23290_,
    new_n23291_, new_n23292_, new_n23293_, new_n23294_, new_n23295_,
    new_n23296_, new_n23297_, new_n23298_, new_n23299_, new_n23300_,
    new_n23301_, new_n23302_, new_n23303_, new_n23304_, new_n23305_,
    new_n23306_, new_n23307_, new_n23308_, new_n23309_, new_n23310_,
    new_n23311_, new_n23312_, new_n23313_, new_n23314_, new_n23315_,
    new_n23316_, new_n23317_, new_n23318_, new_n23319_, new_n23320_,
    new_n23321_, new_n23322_, new_n23323_, new_n23324_, new_n23325_,
    new_n23326_, new_n23327_, new_n23328_, new_n23329_, new_n23330_,
    new_n23331_, new_n23332_, new_n23333_, new_n23334_, new_n23335_,
    new_n23336_, new_n23337_, new_n23338_, new_n23339_, new_n23340_,
    new_n23341_, new_n23342_, new_n23343_, new_n23344_, new_n23345_,
    new_n23346_, new_n23347_, new_n23348_, new_n23349_, new_n23350_,
    new_n23351_, new_n23352_, new_n23353_, new_n23354_, new_n23355_,
    new_n23356_, new_n23357_, new_n23358_, new_n23359_, new_n23360_,
    new_n23361_, new_n23362_, new_n23363_, new_n23364_, new_n23365_,
    new_n23366_, new_n23367_, new_n23368_, new_n23369_, new_n23370_,
    new_n23371_, new_n23372_, new_n23373_, new_n23374_, new_n23375_,
    new_n23376_, new_n23377_, new_n23378_, new_n23379_, new_n23380_,
    new_n23381_, new_n23382_, new_n23383_, new_n23384_, new_n23385_,
    new_n23386_, new_n23387_, new_n23388_, new_n23389_, new_n23390_,
    new_n23391_, new_n23392_, new_n23393_, new_n23394_, new_n23395_,
    new_n23396_, new_n23397_, new_n23398_, new_n23399_, new_n23400_,
    new_n23401_, new_n23402_, new_n23403_, new_n23404_, new_n23405_,
    new_n23406_, new_n23407_, new_n23408_, new_n23409_, new_n23410_,
    new_n23411_, new_n23412_, new_n23413_, new_n23414_, new_n23415_,
    new_n23416_, new_n23417_, new_n23418_, new_n23419_, new_n23420_,
    new_n23421_, new_n23422_, new_n23423_, new_n23424_, new_n23425_,
    new_n23426_, new_n23427_, new_n23428_, new_n23429_, new_n23430_,
    new_n23431_, new_n23432_, new_n23433_, new_n23434_, new_n23435_,
    new_n23436_, new_n23437_, new_n23438_, new_n23439_, new_n23440_,
    new_n23441_, new_n23442_, new_n23443_, new_n23444_, new_n23445_,
    new_n23446_, new_n23447_, new_n23448_, new_n23449_, new_n23450_,
    new_n23451_, new_n23452_, new_n23453_, new_n23454_, new_n23455_,
    new_n23456_, new_n23457_, new_n23458_, new_n23459_, new_n23460_,
    new_n23461_, new_n23462_, new_n23463_, new_n23464_, new_n23465_,
    new_n23466_, new_n23467_, new_n23468_, new_n23469_, new_n23470_,
    new_n23471_, new_n23472_, new_n23473_, new_n23474_, new_n23475_,
    new_n23476_, new_n23477_, new_n23478_, new_n23479_, new_n23480_,
    new_n23481_, new_n23482_, new_n23483_, new_n23484_, new_n23485_,
    new_n23486_, new_n23487_, new_n23488_, new_n23489_, new_n23490_,
    new_n23491_, new_n23492_, new_n23493_, new_n23494_, new_n23495_,
    new_n23496_, new_n23497_, new_n23498_, new_n23499_, new_n23500_,
    new_n23501_, new_n23502_, new_n23503_, new_n23504_, new_n23505_,
    new_n23506_, new_n23507_, new_n23508_, new_n23509_, new_n23510_,
    new_n23511_, new_n23512_, new_n23513_, new_n23514_, new_n23515_,
    new_n23516_, new_n23517_, new_n23518_, new_n23519_, new_n23520_,
    new_n23521_, new_n23522_, new_n23523_, new_n23524_, new_n23525_,
    new_n23526_, new_n23527_, new_n23528_, new_n23529_, new_n23530_,
    new_n23531_, new_n23532_, new_n23533_, new_n23534_, new_n23535_,
    new_n23536_, new_n23537_, new_n23538_, new_n23539_, new_n23540_,
    new_n23541_, new_n23542_, new_n23543_, new_n23544_, new_n23545_,
    new_n23546_, new_n23547_, new_n23548_, new_n23549_, new_n23550_,
    new_n23551_, new_n23552_, new_n23553_, new_n23554_, new_n23555_,
    new_n23556_, new_n23557_, new_n23558_, new_n23559_, new_n23560_,
    new_n23561_, new_n23562_, new_n23563_, new_n23564_, new_n23565_,
    new_n23566_, new_n23567_, new_n23568_, new_n23569_, new_n23570_,
    new_n23571_, new_n23572_, new_n23573_, new_n23574_, new_n23575_,
    new_n23576_, new_n23577_, new_n23578_, new_n23579_, new_n23580_,
    new_n23581_, new_n23582_, new_n23583_, new_n23584_, new_n23585_,
    new_n23586_, new_n23587_, new_n23588_, new_n23589_, new_n23590_,
    new_n23591_, new_n23592_, new_n23593_, new_n23594_, new_n23595_,
    new_n23596_, new_n23597_, new_n23598_, new_n23599_, new_n23600_,
    new_n23601_, new_n23602_, new_n23603_, new_n23604_, new_n23605_,
    new_n23606_, new_n23607_, new_n23608_, new_n23609_, new_n23610_,
    new_n23611_, new_n23612_, new_n23613_, new_n23614_, new_n23615_,
    new_n23616_, new_n23617_, new_n23618_, new_n23619_, new_n23620_,
    new_n23621_, new_n23622_, new_n23623_, new_n23624_, new_n23625_,
    new_n23626_, new_n23627_, new_n23628_, new_n23629_, new_n23630_,
    new_n23631_, new_n23632_, new_n23633_, new_n23634_, new_n23635_,
    new_n23636_, new_n23637_, new_n23638_, new_n23639_, new_n23640_,
    new_n23641_, new_n23642_, new_n23643_, new_n23644_, new_n23645_,
    new_n23646_, new_n23647_, new_n23648_, new_n23649_, new_n23650_,
    new_n23651_, new_n23652_, new_n23653_, new_n23654_, new_n23655_,
    new_n23656_, new_n23657_, new_n23658_, new_n23659_, new_n23660_,
    new_n23661_, new_n23662_, new_n23663_, new_n23664_, new_n23665_,
    new_n23666_, new_n23667_, new_n23668_, new_n23669_, new_n23670_,
    new_n23671_, new_n23672_, new_n23673_, new_n23674_, new_n23675_,
    new_n23676_, new_n23677_, new_n23678_, new_n23679_, new_n23680_,
    new_n23681_, new_n23682_, new_n23683_, new_n23684_, new_n23685_,
    new_n23686_, new_n23687_, new_n23688_, new_n23689_, new_n23690_,
    new_n23691_, new_n23692_, new_n23693_, new_n23694_, new_n23695_,
    new_n23696_, new_n23697_, new_n23698_, new_n23699_, new_n23700_,
    new_n23701_, new_n23702_, new_n23703_, new_n23704_, new_n23705_,
    new_n23706_, new_n23707_, new_n23708_, new_n23709_, new_n23710_,
    new_n23711_, new_n23712_, new_n23713_, new_n23714_, new_n23715_,
    new_n23716_, new_n23717_, new_n23718_, new_n23719_, new_n23720_,
    new_n23721_, new_n23722_, new_n23723_, new_n23724_, new_n23725_,
    new_n23726_, new_n23727_, new_n23728_, new_n23729_, new_n23730_,
    new_n23731_, new_n23732_, new_n23733_, new_n23734_, new_n23735_,
    new_n23736_, new_n23737_, new_n23738_, new_n23739_, new_n23740_,
    new_n23741_, new_n23742_, new_n23743_, new_n23744_, new_n23745_,
    new_n23746_, new_n23747_, new_n23748_, new_n23749_, new_n23750_,
    new_n23751_, new_n23752_, new_n23753_, new_n23754_, new_n23755_,
    new_n23756_, new_n23757_, new_n23758_, new_n23759_, new_n23760_,
    new_n23761_, new_n23762_, new_n23763_, new_n23764_, new_n23765_,
    new_n23766_, new_n23767_, new_n23768_, new_n23769_, new_n23770_,
    new_n23771_, new_n23772_, new_n23773_, new_n23774_, new_n23775_,
    new_n23776_, new_n23777_, new_n23778_, new_n23779_, new_n23780_,
    new_n23781_, new_n23782_, new_n23783_, new_n23784_, new_n23785_,
    new_n23786_, new_n23787_, new_n23788_, new_n23789_, new_n23790_,
    new_n23791_, new_n23792_, new_n23793_, new_n23794_, new_n23795_,
    new_n23796_, new_n23797_, new_n23798_, new_n23799_, new_n23800_,
    new_n23801_, new_n23802_, new_n23803_, new_n23804_, new_n23805_,
    new_n23806_, new_n23807_, new_n23808_, new_n23809_, new_n23810_,
    new_n23811_, new_n23812_, new_n23813_, new_n23814_, new_n23815_,
    new_n23816_, new_n23817_, new_n23818_, new_n23819_, new_n23820_,
    new_n23821_, new_n23822_, new_n23823_, new_n23824_, new_n23825_,
    new_n23826_, new_n23827_, new_n23828_, new_n23829_, new_n23830_,
    new_n23831_, new_n23832_, new_n23833_, new_n23834_, new_n23835_,
    new_n23836_, new_n23837_, new_n23838_, new_n23839_, new_n23840_,
    new_n23841_, new_n23842_, new_n23843_, new_n23844_, new_n23845_,
    new_n23846_, new_n23847_, new_n23848_, new_n23849_, new_n23850_,
    new_n23851_, new_n23852_, new_n23853_, new_n23854_, new_n23855_,
    new_n23856_, new_n23857_, new_n23858_, new_n23859_, new_n23860_,
    new_n23861_, new_n23862_, new_n23863_, new_n23864_, new_n23865_,
    new_n23866_, new_n23867_, new_n23868_, new_n23869_, new_n23870_,
    new_n23871_, new_n23872_, new_n23873_, new_n23874_, new_n23875_,
    new_n23876_, new_n23877_, new_n23878_, new_n23879_, new_n23880_,
    new_n23881_, new_n23882_, new_n23883_, new_n23884_, new_n23885_,
    new_n23886_, new_n23887_, new_n23888_, new_n23889_, new_n23890_,
    new_n23891_, new_n23892_, new_n23893_, new_n23894_, new_n23895_,
    new_n23896_, new_n23897_, new_n23898_, new_n23899_, new_n23900_,
    new_n23901_, new_n23902_, new_n23903_, new_n23904_, new_n23905_,
    new_n23906_, new_n23907_, new_n23908_, new_n23909_, new_n23910_,
    new_n23911_, new_n23912_, new_n23913_, new_n23914_, new_n23915_,
    new_n23916_, new_n23917_, new_n23918_, new_n23919_, new_n23920_,
    new_n23921_, new_n23922_, new_n23923_, new_n23924_, new_n23925_,
    new_n23926_, new_n23927_, new_n23928_, new_n23929_, new_n23930_,
    new_n23931_, new_n23932_, new_n23933_, new_n23934_, new_n23935_,
    new_n23936_, new_n23937_, new_n23938_, new_n23939_, new_n23940_,
    new_n23941_, new_n23942_, new_n23943_, new_n23944_, new_n23945_,
    new_n23946_, new_n23947_, new_n23948_, new_n23949_, new_n23950_,
    new_n23951_, new_n23952_, new_n23953_, new_n23954_, new_n23955_,
    new_n23956_, new_n23957_, new_n23958_, new_n23959_, new_n23960_,
    new_n23961_, new_n23962_, new_n23963_, new_n23964_, new_n23965_,
    new_n23966_, new_n23967_, new_n23968_, new_n23969_, new_n23970_,
    new_n23971_, new_n23972_, new_n23973_, new_n23974_, new_n23975_,
    new_n23976_, new_n23977_, new_n23978_, new_n23979_, new_n23980_,
    new_n23981_, new_n23982_, new_n23983_, new_n23984_, new_n23985_,
    new_n23986_, new_n23987_, new_n23988_, new_n23989_, new_n23990_,
    new_n23991_, new_n23992_, new_n23993_, new_n23994_, new_n23995_,
    new_n23996_, new_n23997_, new_n23998_, new_n23999_, new_n24000_,
    new_n24001_, new_n24002_, new_n24003_, new_n24004_, new_n24005_,
    new_n24006_, new_n24007_, new_n24008_, new_n24009_, new_n24010_,
    new_n24011_, new_n24012_, new_n24013_, new_n24014_, new_n24015_,
    new_n24016_, new_n24017_, new_n24018_, new_n24019_, new_n24020_,
    new_n24021_, new_n24022_, new_n24023_, new_n24024_, new_n24025_,
    new_n24026_, new_n24027_, new_n24028_, new_n24029_, new_n24030_,
    new_n24031_, new_n24032_, new_n24033_, new_n24034_, new_n24035_,
    new_n24036_, new_n24037_, new_n24038_, new_n24039_, new_n24040_,
    new_n24041_, new_n24042_, new_n24043_, new_n24044_, new_n24045_,
    new_n24046_, new_n24047_, new_n24048_, new_n24049_, new_n24050_,
    new_n24051_, new_n24052_, new_n24053_, new_n24054_, new_n24055_,
    new_n24056_, new_n24057_, new_n24058_, new_n24059_, new_n24060_,
    new_n24061_, new_n24062_, new_n24063_, new_n24064_, new_n24065_,
    new_n24066_, new_n24067_, new_n24068_, new_n24069_, new_n24070_,
    new_n24071_, new_n24072_, new_n24073_, new_n24074_, new_n24075_,
    new_n24076_, new_n24077_, new_n24078_, new_n24079_, new_n24080_,
    new_n24081_, new_n24082_, new_n24083_, new_n24084_, new_n24085_,
    new_n24086_, new_n24087_, new_n24088_, new_n24089_, new_n24090_,
    new_n24091_, new_n24092_, new_n24093_, new_n24094_, new_n24095_,
    new_n24096_, new_n24097_, new_n24098_, new_n24099_, new_n24100_,
    new_n24101_, new_n24102_, new_n24103_, new_n24104_, new_n24105_,
    new_n24106_, new_n24107_, new_n24108_, new_n24109_, new_n24110_,
    new_n24111_, new_n24112_, new_n24113_, new_n24114_, new_n24115_,
    new_n24116_, new_n24117_, new_n24118_, new_n24119_, new_n24120_,
    new_n24121_, new_n24122_, new_n24123_, new_n24124_, new_n24125_,
    new_n24126_, new_n24127_, new_n24128_, new_n24129_, new_n24130_,
    new_n24131_, new_n24132_, new_n24133_, new_n24134_, new_n24135_,
    new_n24136_, new_n24137_, new_n24138_, new_n24139_, new_n24140_,
    new_n24141_, new_n24142_, new_n24143_, new_n24144_, new_n24145_,
    new_n24146_, new_n24147_, new_n24148_, new_n24149_, new_n24150_,
    new_n24151_, new_n24152_, new_n24153_, new_n24154_, new_n24155_,
    new_n24156_, new_n24157_, new_n24158_, new_n24159_, new_n24160_,
    new_n24161_, new_n24162_, new_n24163_, new_n24164_, new_n24165_,
    new_n24166_, new_n24167_, new_n24168_, new_n24169_, new_n24170_,
    new_n24171_, new_n24172_, new_n24173_, new_n24174_, new_n24175_,
    new_n24176_, new_n24177_, new_n24178_, new_n24179_, new_n24180_,
    new_n24181_, new_n24182_, new_n24183_, new_n24184_, new_n24185_,
    new_n24186_, new_n24187_, new_n24188_, new_n24189_, new_n24190_,
    new_n24191_, new_n24192_, new_n24193_, new_n24194_, new_n24195_,
    new_n24196_, new_n24197_, new_n24198_, new_n24199_, new_n24200_,
    new_n24201_, new_n24202_, new_n24203_, new_n24204_, new_n24205_,
    new_n24206_, new_n24207_, new_n24208_, new_n24209_, new_n24210_,
    new_n24211_, new_n24212_, new_n24213_, new_n24214_, new_n24215_,
    new_n24216_, new_n24217_, new_n24218_, new_n24219_, new_n24220_,
    new_n24221_, new_n24222_, new_n24223_, new_n24224_, new_n24225_,
    new_n24226_, new_n24227_, new_n24228_, new_n24229_, new_n24230_,
    new_n24231_, new_n24232_, new_n24233_, new_n24234_, new_n24235_,
    new_n24236_, new_n24237_, new_n24238_, new_n24239_, new_n24240_,
    new_n24241_, new_n24242_, new_n24243_, new_n24244_, new_n24245_,
    new_n24246_, new_n24247_, new_n24248_, new_n24249_, new_n24250_,
    new_n24251_, new_n24252_, new_n24253_, new_n24254_, new_n24255_,
    new_n24256_, new_n24257_, new_n24258_, new_n24259_, new_n24260_,
    new_n24261_, new_n24262_, new_n24263_, new_n24264_, new_n24265_,
    new_n24266_, new_n24267_, new_n24268_, new_n24269_, new_n24270_,
    new_n24271_, new_n24272_, new_n24273_, new_n24274_, new_n24275_,
    new_n24276_, new_n24277_, new_n24278_, new_n24279_, new_n24280_,
    new_n24281_, new_n24282_, new_n24283_, new_n24284_, new_n24285_,
    new_n24286_, new_n24287_, new_n24288_, new_n24289_, new_n24290_,
    new_n24291_, new_n24292_, new_n24293_, new_n24294_, new_n24295_,
    new_n24296_, new_n24297_, new_n24298_, new_n24299_, new_n24300_,
    new_n24301_, new_n24302_, new_n24303_, new_n24304_, new_n24305_,
    new_n24306_, new_n24307_, new_n24308_, new_n24309_, new_n24310_,
    new_n24311_, new_n24312_, new_n24313_, new_n24314_, new_n24315_,
    new_n24316_, new_n24317_, new_n24318_, new_n24319_, new_n24320_,
    new_n24321_, new_n24322_, new_n24323_, new_n24324_, new_n24325_,
    new_n24326_, new_n24327_, new_n24328_, new_n24329_, new_n24330_,
    new_n24331_, new_n24332_, new_n24333_, new_n24334_, new_n24335_,
    new_n24336_, new_n24337_, new_n24338_, new_n24339_, new_n24340_,
    new_n24341_, new_n24342_, new_n24343_, new_n24344_, new_n24345_,
    new_n24346_, new_n24347_, new_n24348_, new_n24349_, new_n24350_,
    new_n24351_, new_n24352_, new_n24353_, new_n24354_, new_n24355_,
    new_n24356_, new_n24357_, new_n24358_, new_n24359_, new_n24360_,
    new_n24361_, new_n24362_, new_n24363_, new_n24364_, new_n24365_,
    new_n24366_, new_n24367_, new_n24368_, new_n24369_, new_n24370_,
    new_n24371_, new_n24372_, new_n24373_, new_n24374_, new_n24375_,
    new_n24376_, new_n24377_, new_n24378_, new_n24379_, new_n24380_,
    new_n24381_, new_n24382_, new_n24383_, new_n24384_, new_n24385_,
    new_n24386_, new_n24387_, new_n24388_, new_n24389_, new_n24390_,
    new_n24391_, new_n24392_, new_n24393_, new_n24394_, new_n24395_,
    new_n24396_, new_n24397_, new_n24398_, new_n24399_, new_n24400_,
    new_n24401_, new_n24402_, new_n24403_, new_n24404_, new_n24405_,
    new_n24406_, new_n24407_, new_n24408_, new_n24409_, new_n24410_,
    new_n24411_, new_n24412_, new_n24413_, new_n24414_, new_n24415_,
    new_n24416_, new_n24417_, new_n24418_, new_n24419_, new_n24420_,
    new_n24421_, new_n24422_, new_n24423_, new_n24424_, new_n24425_,
    new_n24426_, new_n24427_, new_n24428_, new_n24429_, new_n24430_,
    new_n24431_, new_n24432_, new_n24433_, new_n24434_, new_n24435_,
    new_n24436_, new_n24437_, new_n24438_, new_n24439_, new_n24440_,
    new_n24441_, new_n24442_, new_n24443_, new_n24444_, new_n24445_,
    new_n24446_, new_n24447_, new_n24448_, new_n24449_, new_n24450_,
    new_n24451_, new_n24452_, new_n24453_, new_n24454_, new_n24455_,
    new_n24456_, new_n24457_, new_n24458_, new_n24459_, new_n24460_,
    new_n24461_, new_n24462_, new_n24463_, new_n24464_, new_n24465_,
    new_n24466_, new_n24467_, new_n24468_, new_n24469_, new_n24470_,
    new_n24471_, new_n24472_, new_n24473_, new_n24474_, new_n24475_,
    new_n24476_, new_n24477_, new_n24478_, new_n24479_, new_n24480_,
    new_n24481_, new_n24482_, new_n24483_, new_n24484_, new_n24485_,
    new_n24486_, new_n24487_, new_n24488_, new_n24489_, new_n24490_,
    new_n24491_, new_n24492_, new_n24493_, new_n24494_, new_n24495_,
    new_n24496_, new_n24497_, new_n24498_, new_n24499_, new_n24500_,
    new_n24501_, new_n24502_, new_n24503_, new_n24504_, new_n24505_,
    new_n24506_, new_n24507_, new_n24508_, new_n24509_, new_n24510_,
    new_n24511_, new_n24512_, new_n24513_, new_n24514_, new_n24515_,
    new_n24516_, new_n24517_, new_n24518_, new_n24519_, new_n24520_,
    new_n24521_, new_n24522_, new_n24523_, new_n24524_, new_n24525_,
    new_n24526_, new_n24527_, new_n24528_, new_n24529_, new_n24530_,
    new_n24531_, new_n24532_, new_n24533_, new_n24534_, new_n24535_,
    new_n24536_, new_n24537_, new_n24538_, new_n24539_, new_n24540_,
    new_n24541_, new_n24542_, new_n24543_, new_n24544_, new_n24545_,
    new_n24546_, new_n24547_, new_n24548_, new_n24549_, new_n24550_,
    new_n24551_, new_n24552_, new_n24553_, new_n24554_, new_n24555_,
    new_n24556_, new_n24557_, new_n24558_, new_n24559_, new_n24560_,
    new_n24561_, new_n24562_, new_n24563_, new_n24564_, new_n24565_,
    new_n24566_, new_n24567_, new_n24568_, new_n24569_, new_n24570_,
    new_n24571_, new_n24572_, new_n24573_, new_n24574_, new_n24575_,
    new_n24576_, new_n24577_, new_n24578_, new_n24579_, new_n24580_,
    new_n24581_, new_n24582_, new_n24583_, new_n24584_, new_n24585_,
    new_n24586_, new_n24587_, new_n24588_, new_n24589_, new_n24590_,
    new_n24591_, new_n24592_, new_n24593_, new_n24594_, new_n24595_,
    new_n24596_, new_n24597_, new_n24598_, new_n24599_, new_n24600_,
    new_n24601_, new_n24602_, new_n24603_, new_n24604_, new_n24605_,
    new_n24606_, new_n24607_, new_n24608_, new_n24609_, new_n24610_,
    new_n24611_, new_n24612_, new_n24613_, new_n24614_, new_n24615_,
    new_n24616_, new_n24617_, new_n24618_, new_n24619_, new_n24620_,
    new_n24621_, new_n24622_, new_n24623_, new_n24624_, new_n24625_,
    new_n24626_, new_n24627_, new_n24628_, new_n24629_, new_n24630_,
    new_n24631_, new_n24632_, new_n24633_, new_n24634_, new_n24635_,
    new_n24636_, new_n24637_, new_n24638_, new_n24639_, new_n24640_,
    new_n24641_, new_n24642_, new_n24643_, new_n24644_, new_n24645_,
    new_n24646_, new_n24647_, new_n24648_, new_n24649_, new_n24650_,
    new_n24651_, new_n24652_, new_n24653_, new_n24654_, new_n24655_,
    new_n24656_, new_n24657_, new_n24658_, new_n24659_, new_n24660_,
    new_n24661_, new_n24662_, new_n24663_, new_n24664_, new_n24665_,
    new_n24666_, new_n24667_, new_n24668_, new_n24669_, new_n24670_,
    new_n24671_, new_n24672_, new_n24673_, new_n24674_, new_n24675_,
    new_n24676_, new_n24677_, new_n24678_, new_n24679_, new_n24680_,
    new_n24681_, new_n24682_, new_n24683_, new_n24684_, new_n24685_,
    new_n24686_, new_n24687_, new_n24688_, new_n24689_, new_n24690_,
    new_n24691_, new_n24692_, new_n24693_, new_n24694_, new_n24695_,
    new_n24696_, new_n24697_, new_n24698_, new_n24699_, new_n24700_,
    new_n24701_, new_n24702_, new_n24703_, new_n24704_, new_n24705_,
    new_n24706_, new_n24707_, new_n24708_, new_n24709_, new_n24710_,
    new_n24711_, new_n24712_, new_n24713_, new_n24714_, new_n24715_,
    new_n24716_, new_n24717_, new_n24718_, new_n24719_, new_n24720_,
    new_n24721_, new_n24722_, new_n24723_, new_n24724_, new_n24725_,
    new_n24726_, new_n24727_, new_n24728_, new_n24729_, new_n24730_,
    new_n24731_, new_n24732_, new_n24733_, new_n24734_, new_n24735_,
    new_n24736_, new_n24737_, new_n24738_, new_n24739_, new_n24740_,
    new_n24741_, new_n24742_, new_n24743_, new_n24744_, new_n24745_,
    new_n24746_, new_n24747_, new_n24748_, new_n24749_, new_n24750_,
    new_n24751_, new_n24752_, new_n24753_, new_n24754_, new_n24755_,
    new_n24756_, new_n24757_, new_n24758_, new_n24759_, new_n24760_,
    new_n24761_, new_n24762_, new_n24763_, new_n24764_, new_n24765_,
    new_n24766_, new_n24767_, new_n24768_, new_n24769_, new_n24770_,
    new_n24771_, new_n24772_, new_n24773_, new_n24774_, new_n24775_,
    new_n24776_, new_n24777_, new_n24778_, new_n24779_, new_n24780_,
    new_n24781_, new_n24782_, new_n24783_, new_n24784_, new_n24785_,
    new_n24786_, new_n24787_, new_n24788_, new_n24789_, new_n24790_,
    new_n24791_, new_n24792_, new_n24793_, new_n24794_, new_n24795_,
    new_n24796_, new_n24797_, new_n24798_, new_n24799_, new_n24800_,
    new_n24801_, new_n24802_, new_n24803_, new_n24804_, new_n24805_,
    new_n24806_, new_n24807_, new_n24808_, new_n24809_, new_n24810_,
    new_n24811_, new_n24812_, new_n24813_, new_n24814_, new_n24815_,
    new_n24816_, new_n24817_, new_n24818_, new_n24819_, new_n24820_,
    new_n24821_, new_n24822_, new_n24823_, new_n24824_, new_n24825_,
    new_n24826_, new_n24827_, new_n24828_, new_n24829_, new_n24830_,
    new_n24831_, new_n24832_, new_n24833_, new_n24834_, new_n24835_,
    new_n24836_, new_n24837_, new_n24838_, new_n24839_, new_n24840_,
    new_n24841_, new_n24842_, new_n24843_, new_n24844_, new_n24845_,
    new_n24846_, new_n24847_, new_n24848_, new_n24849_, new_n24850_,
    new_n24851_, new_n24852_, new_n24853_, new_n24854_, new_n24855_,
    new_n24856_, new_n24857_, new_n24858_, new_n24859_, new_n24860_,
    new_n24861_, new_n24862_, new_n24863_, new_n24864_, new_n24865_,
    new_n24866_, new_n24867_, new_n24868_, new_n24869_, new_n24870_,
    new_n24871_, new_n24872_, new_n24873_, new_n24874_, new_n24875_,
    new_n24876_, new_n24877_, new_n24878_, new_n24879_, new_n24880_,
    new_n24881_, new_n24882_, new_n24883_, new_n24884_, new_n24885_,
    new_n24886_, new_n24887_, new_n24888_, new_n24889_, new_n24890_,
    new_n24891_, new_n24892_, new_n24893_, new_n24894_, new_n24895_,
    new_n24896_, new_n24897_, new_n24898_, new_n24899_, new_n24900_,
    new_n24901_, new_n24902_, new_n24903_, new_n24904_, new_n24905_,
    new_n24906_, new_n24907_, new_n24908_, new_n24909_, new_n24910_,
    new_n24911_, new_n24912_, new_n24913_, new_n24914_, new_n24915_,
    new_n24916_, new_n24917_, new_n24918_, new_n24919_, new_n24920_,
    new_n24921_, new_n24922_, new_n24923_, new_n24924_, new_n24925_,
    new_n24926_, new_n24927_, new_n24928_, new_n24929_, new_n24930_,
    new_n24931_, new_n24932_, new_n24933_, new_n24934_, new_n24935_,
    new_n24936_, new_n24937_, new_n24938_, new_n24939_, new_n24940_,
    new_n24941_, new_n24942_, new_n24943_, new_n24944_, new_n24945_,
    new_n24946_, new_n24947_, new_n24948_, new_n24949_, new_n24950_,
    new_n24951_, new_n24952_, new_n24953_, new_n24954_, new_n24955_,
    new_n24956_, new_n24957_, new_n24958_, new_n24959_, new_n24960_,
    new_n24961_, new_n24962_, new_n24963_, new_n24964_, new_n24965_,
    new_n24966_, new_n24967_, new_n24968_, new_n24969_, new_n24970_,
    new_n24971_, new_n24972_, new_n24973_, new_n24974_, new_n24975_,
    new_n24976_, new_n24977_, new_n24978_, new_n24979_, new_n24980_,
    new_n24981_, new_n24982_, new_n24983_, new_n24984_, new_n24985_,
    new_n24986_, new_n24987_, new_n24988_, new_n24989_, new_n24990_,
    new_n24991_, new_n24992_, new_n24993_, new_n24994_, new_n24995_,
    new_n24996_, new_n24997_, new_n24998_, new_n24999_, new_n25000_,
    new_n25001_, new_n25002_, new_n25003_, new_n25004_, new_n25005_,
    new_n25006_, new_n25007_, new_n25008_, new_n25009_, new_n25010_,
    new_n25011_, new_n25012_, new_n25013_, new_n25014_, new_n25015_,
    new_n25016_, new_n25017_, new_n25018_, new_n25019_, new_n25020_,
    new_n25021_, new_n25022_, new_n25023_, new_n25024_, new_n25025_,
    new_n25026_, new_n25027_, new_n25028_, new_n25029_, new_n25030_,
    new_n25031_, new_n25032_, new_n25033_, new_n25034_, new_n25035_,
    new_n25036_, new_n25037_, new_n25038_, new_n25039_, new_n25040_,
    new_n25041_, new_n25042_, new_n25043_, new_n25044_, new_n25045_,
    new_n25046_, new_n25047_, new_n25048_, new_n25049_, new_n25050_,
    new_n25051_, new_n25052_, new_n25053_, new_n25054_, new_n25055_,
    new_n25056_, new_n25057_, new_n25058_, new_n25059_, new_n25060_,
    new_n25061_, new_n25062_, new_n25063_, new_n25064_, new_n25065_,
    new_n25066_, new_n25067_, new_n25068_, new_n25069_, new_n25070_,
    new_n25071_, new_n25072_, new_n25073_, new_n25074_, new_n25075_,
    new_n25076_, new_n25077_, new_n25078_, new_n25079_, new_n25080_,
    new_n25081_, new_n25082_, new_n25083_, new_n25084_, new_n25085_,
    new_n25086_, new_n25087_, new_n25088_, new_n25089_, new_n25090_,
    new_n25091_, new_n25092_, new_n25093_, new_n25094_, new_n25095_,
    new_n25096_, new_n25097_, new_n25098_, new_n25099_, new_n25100_,
    new_n25101_, new_n25102_, new_n25103_, new_n25104_, new_n25105_,
    new_n25106_, new_n25107_, new_n25108_, new_n25109_, new_n25110_,
    new_n25111_, new_n25112_, new_n25113_, new_n25114_, new_n25115_,
    new_n25116_, new_n25117_, new_n25118_, new_n25119_, new_n25120_,
    new_n25121_, new_n25122_, new_n25123_, new_n25124_, new_n25125_,
    new_n25126_, new_n25127_, new_n25128_, new_n25129_, new_n25130_,
    new_n25131_, new_n25132_, new_n25133_, new_n25134_, new_n25135_,
    new_n25136_, new_n25137_, new_n25138_, new_n25139_, new_n25140_,
    new_n25141_, new_n25142_, new_n25143_, new_n25144_, new_n25145_,
    new_n25146_, new_n25147_, new_n25148_, new_n25149_, new_n25150_,
    new_n25151_, new_n25152_, new_n25153_, new_n25154_, new_n25155_,
    new_n25156_, new_n25157_, new_n25158_, new_n25159_, new_n25160_,
    new_n25161_, new_n25162_, new_n25163_, new_n25164_, new_n25165_,
    new_n25166_, new_n25167_, new_n25168_, new_n25169_, new_n25170_,
    new_n25171_, new_n25172_, new_n25173_, new_n25174_, new_n25175_,
    new_n25176_, new_n25177_, new_n25178_, new_n25179_, new_n25180_,
    new_n25181_, new_n25182_, new_n25183_, new_n25184_, new_n25185_,
    new_n25186_, new_n25187_, new_n25188_, new_n25189_, new_n25190_,
    new_n25191_, new_n25192_, new_n25193_, new_n25194_, new_n25195_,
    new_n25196_, new_n25197_, new_n25198_, new_n25199_, new_n25200_,
    new_n25201_, new_n25202_, new_n25203_, new_n25204_, new_n25205_,
    new_n25206_, new_n25207_, new_n25208_, new_n25209_, new_n25210_,
    new_n25211_, new_n25212_, new_n25213_, new_n25214_, new_n25215_,
    new_n25216_, new_n25217_, new_n25218_, new_n25219_, new_n25220_,
    new_n25221_, new_n25222_, new_n25223_, new_n25224_, new_n25225_,
    new_n25226_, new_n25227_, new_n25228_, new_n25229_, new_n25230_,
    new_n25231_, new_n25232_, new_n25233_, new_n25234_, new_n25235_,
    new_n25236_, new_n25237_, new_n25238_, new_n25239_, new_n25240_,
    new_n25241_, new_n25242_, new_n25243_, new_n25244_, new_n25245_,
    new_n25246_, new_n25247_, new_n25248_, new_n25249_, new_n25250_,
    new_n25251_, new_n25252_, new_n25253_, new_n25254_, new_n25255_,
    new_n25256_, new_n25257_, new_n25258_, new_n25259_, new_n25260_,
    new_n25261_, new_n25262_, new_n25263_, new_n25264_, new_n25265_,
    new_n25266_, new_n25267_, new_n25268_, new_n25269_, new_n25270_,
    new_n25271_, new_n25272_, new_n25273_, new_n25274_, new_n25275_,
    new_n25276_, new_n25277_, new_n25278_, new_n25279_, new_n25280_,
    new_n25281_, new_n25282_, new_n25283_, new_n25284_, new_n25285_,
    new_n25286_, new_n25287_, new_n25288_, new_n25289_, new_n25290_,
    new_n25291_, new_n25292_, new_n25293_, new_n25294_, new_n25295_,
    new_n25296_, new_n25297_, new_n25298_, new_n25299_, new_n25300_,
    new_n25301_, new_n25302_, new_n25303_, new_n25304_, new_n25305_,
    new_n25306_, new_n25307_, new_n25308_, new_n25309_, new_n25310_,
    new_n25311_, new_n25312_, new_n25313_, new_n25314_, new_n25315_,
    new_n25316_, new_n25317_, new_n25318_, new_n25319_, new_n25320_,
    new_n25321_, new_n25322_, new_n25323_, new_n25324_, new_n25325_,
    new_n25326_, new_n25327_, new_n25328_, new_n25329_, new_n25330_,
    new_n25331_, new_n25332_, new_n25333_, new_n25334_, new_n25335_,
    new_n25336_, new_n25337_, new_n25338_, new_n25339_, new_n25340_,
    new_n25341_, new_n25342_, new_n25343_, new_n25344_, new_n25345_,
    new_n25346_, new_n25347_, new_n25348_, new_n25349_, new_n25350_,
    new_n25351_, new_n25352_, new_n25353_, new_n25354_, new_n25355_,
    new_n25356_, new_n25357_, new_n25358_, new_n25359_, new_n25360_,
    new_n25361_, new_n25362_, new_n25363_, new_n25364_, new_n25365_,
    new_n25366_, new_n25367_, new_n25368_, new_n25369_, new_n25370_,
    new_n25371_, new_n25372_, new_n25373_, new_n25374_, new_n25375_,
    new_n25376_, new_n25377_, new_n25378_, new_n25379_, new_n25380_,
    new_n25381_, new_n25382_, new_n25383_, new_n25384_, new_n25385_,
    new_n25386_, new_n25387_, new_n25388_, new_n25389_, new_n25390_,
    new_n25391_, new_n25392_, new_n25393_, new_n25394_, new_n25395_,
    new_n25396_, new_n25397_, new_n25398_, new_n25399_, new_n25400_,
    new_n25401_, new_n25402_, new_n25403_, new_n25404_, new_n25405_,
    new_n25406_, new_n25407_, new_n25408_, new_n25409_, new_n25410_,
    new_n25411_, new_n25412_, new_n25413_, new_n25414_, new_n25415_,
    new_n25416_, new_n25417_, new_n25418_, new_n25419_, new_n25420_,
    new_n25421_, new_n25422_, new_n25423_, new_n25424_, new_n25425_,
    new_n25426_, new_n25427_, new_n25428_, new_n25429_, new_n25430_,
    new_n25431_, new_n25432_, new_n25433_, new_n25434_, new_n25435_,
    new_n25436_, new_n25437_, new_n25438_, new_n25439_, new_n25440_,
    new_n25441_, new_n25442_, new_n25443_, new_n25444_, new_n25445_,
    new_n25446_, new_n25447_, new_n25448_, new_n25449_, new_n25450_,
    new_n25451_, new_n25452_, new_n25453_, new_n25454_, new_n25455_,
    new_n25456_, new_n25457_, new_n25458_, new_n25459_, new_n25460_,
    new_n25461_, new_n25462_, new_n25463_, new_n25464_, new_n25465_,
    new_n25466_, new_n25467_, new_n25468_, new_n25469_, new_n25470_,
    new_n25471_, new_n25472_, new_n25473_, new_n25474_, new_n25475_,
    new_n25476_, new_n25477_, new_n25478_, new_n25479_, new_n25480_,
    new_n25481_, new_n25482_, new_n25483_, new_n25484_, new_n25485_,
    new_n25486_, new_n25487_, new_n25488_, new_n25489_, new_n25490_,
    new_n25491_, new_n25492_, new_n25493_, new_n25494_, new_n25495_,
    new_n25496_, new_n25497_, new_n25498_, new_n25499_, new_n25500_,
    new_n25501_, new_n25502_, new_n25503_, new_n25504_, new_n25505_,
    new_n25506_, new_n25507_, new_n25508_, new_n25509_, new_n25510_,
    new_n25511_, new_n25512_, new_n25513_, new_n25514_, new_n25515_,
    new_n25516_, new_n25517_, new_n25518_, new_n25519_, new_n25520_,
    new_n25521_, new_n25522_, new_n25523_, new_n25524_, new_n25525_,
    new_n25526_, new_n25527_, new_n25528_, new_n25529_, new_n25530_,
    new_n25531_, new_n25532_, new_n25533_, new_n25534_, new_n25535_,
    new_n25536_, new_n25537_, new_n25538_, new_n25539_, new_n25540_,
    new_n25541_, new_n25542_, new_n25543_, new_n25544_, new_n25545_,
    new_n25546_, new_n25547_, new_n25548_, new_n25549_, new_n25550_,
    new_n25551_, new_n25552_, new_n25553_, new_n25554_, new_n25555_,
    new_n25556_, new_n25557_, new_n25558_, new_n25559_, new_n25560_,
    new_n25561_, new_n25562_, new_n25563_, new_n25564_, new_n25565_,
    new_n25566_, new_n25567_, new_n25568_, new_n25569_, new_n25570_,
    new_n25571_, new_n25572_, new_n25573_, new_n25574_, new_n25575_,
    new_n25576_, new_n25577_, new_n25578_, new_n25579_, new_n25580_,
    new_n25581_, new_n25582_, new_n25583_, new_n25584_, new_n25585_,
    new_n25586_, new_n25587_, new_n25588_, new_n25589_, new_n25590_,
    new_n25591_, new_n25592_, new_n25593_, new_n25594_, new_n25595_,
    new_n25596_, new_n25597_, new_n25598_, new_n25599_, new_n25600_,
    new_n25601_, new_n25602_, new_n25603_, new_n25604_, new_n25605_,
    new_n25606_, new_n25607_, new_n25608_, new_n25609_, new_n25610_,
    new_n25611_, new_n25612_, new_n25613_, new_n25614_, new_n25615_,
    new_n25616_, new_n25617_, new_n25618_, new_n25619_, new_n25620_,
    new_n25621_, new_n25622_, new_n25623_, new_n25624_, new_n25625_,
    new_n25626_, new_n25627_, new_n25628_, new_n25629_, new_n25630_,
    new_n25631_, new_n25632_, new_n25633_, new_n25634_, new_n25635_,
    new_n25636_, new_n25637_, new_n25638_, new_n25639_, new_n25640_,
    new_n25641_, new_n25642_, new_n25643_, new_n25644_, new_n25645_,
    new_n25646_, new_n25647_, new_n25648_, new_n25649_, new_n25650_,
    new_n25651_, new_n25652_, new_n25653_, new_n25654_, new_n25655_,
    new_n25656_, new_n25657_, new_n25658_, new_n25659_, new_n25660_,
    new_n25661_, new_n25662_, new_n25663_, new_n25664_, new_n25665_,
    new_n25666_, new_n25667_, new_n25668_, new_n25669_, new_n25670_,
    new_n25671_, new_n25672_, new_n25673_, new_n25674_, new_n25675_,
    new_n25676_, new_n25677_, new_n25678_, new_n25679_, new_n25680_,
    new_n25681_, new_n25682_, new_n25683_, new_n25684_, new_n25685_,
    new_n25686_, new_n25687_, new_n25688_, new_n25689_, new_n25690_,
    new_n25691_, new_n25692_, new_n25693_, new_n25694_, new_n25695_,
    new_n25696_, new_n25697_, new_n25698_, new_n25699_, new_n25700_,
    new_n25701_, new_n25702_, new_n25703_, new_n25704_, new_n25705_,
    new_n25706_, new_n25707_, new_n25708_, new_n25709_, new_n25710_,
    new_n25711_, new_n25712_, new_n25713_, new_n25714_, new_n25715_,
    new_n25716_, new_n25717_, new_n25718_, new_n25719_, new_n25720_,
    new_n25721_, new_n25722_, new_n25723_, new_n25724_, new_n25725_,
    new_n25726_, new_n25727_, new_n25728_, new_n25729_, new_n25730_,
    new_n25731_, new_n25732_, new_n25733_, new_n25734_, new_n25735_,
    new_n25736_, new_n25737_, new_n25738_, new_n25739_, new_n25740_,
    new_n25741_, new_n25742_, new_n25743_, new_n25744_, new_n25745_,
    new_n25746_, new_n25747_, new_n25748_, new_n25749_, new_n25750_,
    new_n25751_, new_n25752_, new_n25753_, new_n25754_, new_n25755_,
    new_n25756_, new_n25757_, new_n25758_, new_n25759_, new_n25760_,
    new_n25761_, new_n25762_, new_n25763_, new_n25764_, new_n25765_,
    new_n25766_, new_n25767_, new_n25768_, new_n25769_, new_n25770_,
    new_n25771_, new_n25772_, new_n25773_, new_n25774_, new_n25775_,
    new_n25776_, new_n25777_, new_n25778_, new_n25779_, new_n25780_,
    new_n25781_, new_n25782_, new_n25783_, new_n25784_, new_n25785_,
    new_n25786_, new_n25787_, new_n25788_, new_n25789_, new_n25790_,
    new_n25791_, new_n25792_, new_n25793_, new_n25794_, new_n25795_,
    new_n25796_, new_n25797_, new_n25798_, new_n25799_, new_n25800_,
    new_n25801_, new_n25802_, new_n25803_, new_n25804_, new_n25805_,
    new_n25806_, new_n25807_, new_n25808_, new_n25809_, new_n25810_,
    new_n25811_, new_n25812_, new_n25813_, new_n25814_, new_n25815_,
    new_n25816_, new_n25817_, new_n25818_, new_n25819_, new_n25820_,
    new_n25821_, new_n25822_, new_n25823_, new_n25824_, new_n25825_,
    new_n25826_, new_n25827_, new_n25828_, new_n25829_, new_n25830_,
    new_n25831_, new_n25832_, new_n25833_, new_n25834_, new_n25835_,
    new_n25836_, new_n25837_, new_n25838_, new_n25839_, new_n25840_,
    new_n25841_, new_n25842_, new_n25843_, new_n25844_, new_n25845_,
    new_n25846_, new_n25847_, new_n25848_, new_n25849_, new_n25850_,
    new_n25851_, new_n25852_, new_n25853_, new_n25854_, new_n25855_,
    new_n25856_, new_n25857_, new_n25858_, new_n25859_, new_n25860_,
    new_n25861_, new_n25862_, new_n25863_, new_n25864_, new_n25865_,
    new_n25866_, new_n25867_, new_n25868_, new_n25869_, new_n25870_,
    new_n25871_, new_n25872_, new_n25873_, new_n25874_, new_n25875_,
    new_n25876_, new_n25877_, new_n25878_, new_n25879_, new_n25880_,
    new_n25881_, new_n25882_, new_n25883_, new_n25884_, new_n25885_,
    new_n25886_, new_n25887_, new_n25888_, new_n25889_, new_n25890_,
    new_n25891_, new_n25892_, new_n25893_, new_n25894_, new_n25895_,
    new_n25896_, new_n25897_, new_n25898_, new_n25899_, new_n25900_,
    new_n25901_, new_n25902_, new_n25903_, new_n25904_, new_n25905_,
    new_n25906_, new_n25907_, new_n25908_, new_n25909_, new_n25910_,
    new_n25911_, new_n25912_, new_n25913_, new_n25914_, new_n25915_,
    new_n25916_, new_n25917_, new_n25918_, new_n25919_, new_n25920_,
    new_n25921_, new_n25922_, new_n25923_, new_n25924_, new_n25925_,
    new_n25926_, new_n25927_, new_n25928_, new_n25929_, new_n25930_,
    new_n25931_, new_n25932_, new_n25933_, new_n25934_, new_n25935_,
    new_n25936_, new_n25937_, new_n25938_, new_n25939_, new_n25940_,
    new_n25941_, new_n25942_, new_n25943_, new_n25944_, new_n25945_,
    new_n25946_, new_n25947_, new_n25948_, new_n25949_, new_n25950_,
    new_n25951_, new_n25952_, new_n25953_, new_n25954_, new_n25955_,
    new_n25956_, new_n25957_, new_n25958_, new_n25959_, new_n25960_,
    new_n25961_, new_n25962_, new_n25963_, new_n25964_, new_n25965_,
    new_n25966_, new_n25967_, new_n25968_, new_n25969_, new_n25970_,
    new_n25971_, new_n25972_, new_n25973_, new_n25974_, new_n25975_,
    new_n25976_, new_n25977_, new_n25978_, new_n25979_, new_n25980_,
    new_n25981_, new_n25982_, new_n25983_, new_n25984_, new_n25985_,
    new_n25986_, new_n25987_, new_n25988_, new_n25989_, new_n25990_,
    new_n25991_, new_n25992_, new_n25993_, new_n25994_, new_n25995_,
    new_n25996_, new_n25997_, new_n25998_, new_n25999_, new_n26000_,
    new_n26001_, new_n26002_, new_n26003_, new_n26004_, new_n26005_,
    new_n26006_, new_n26007_, new_n26008_, new_n26009_, new_n26010_,
    new_n26011_, new_n26012_, new_n26013_, new_n26014_, new_n26015_,
    new_n26016_, new_n26017_, new_n26018_, new_n26019_, new_n26020_,
    new_n26021_, new_n26022_, new_n26023_, new_n26024_, new_n26025_,
    new_n26026_, new_n26027_, new_n26028_, new_n26029_, new_n26030_,
    new_n26031_, new_n26032_, new_n26033_, new_n26034_, new_n26035_,
    new_n26036_, new_n26037_, new_n26038_, new_n26039_, new_n26040_,
    new_n26041_, new_n26042_, new_n26043_, new_n26044_, new_n26045_,
    new_n26046_, new_n26047_, new_n26048_, new_n26049_, new_n26050_,
    new_n26051_, new_n26052_, new_n26053_, new_n26054_, new_n26055_,
    new_n26056_, new_n26057_, new_n26058_, new_n26059_, new_n26060_,
    new_n26061_, new_n26062_, new_n26063_, new_n26064_, new_n26065_,
    new_n26066_, new_n26067_, new_n26068_, new_n26069_, new_n26070_,
    new_n26071_, new_n26072_, new_n26073_, new_n26074_, new_n26075_,
    new_n26076_, new_n26077_, new_n26078_, new_n26079_, new_n26080_,
    new_n26081_, new_n26082_, new_n26083_, new_n26084_, new_n26085_,
    new_n26086_, new_n26087_, new_n26088_, new_n26089_, new_n26090_,
    new_n26091_, new_n26092_, new_n26093_, new_n26094_, new_n26095_,
    new_n26096_, new_n26097_, new_n26098_, new_n26099_, new_n26100_,
    new_n26101_, new_n26102_, new_n26103_, new_n26104_, new_n26105_,
    new_n26106_, new_n26107_, new_n26108_, new_n26109_, new_n26110_,
    new_n26111_, new_n26112_, new_n26113_, new_n26114_, new_n26115_,
    new_n26116_, new_n26117_, new_n26118_, new_n26119_, new_n26120_,
    new_n26121_, new_n26122_, new_n26123_, new_n26124_, new_n26125_,
    new_n26126_, new_n26127_, new_n26128_, new_n26129_, new_n26130_,
    new_n26131_, new_n26132_, new_n26133_, new_n26134_, new_n26135_,
    new_n26136_, new_n26137_, new_n26138_, new_n26139_, new_n26140_,
    new_n26141_, new_n26142_, new_n26143_, new_n26144_, new_n26145_,
    new_n26146_, new_n26147_, new_n26148_, new_n26149_, new_n26150_,
    new_n26151_, new_n26152_, new_n26153_, new_n26154_, new_n26155_,
    new_n26156_, new_n26157_, new_n26158_, new_n26159_, new_n26160_,
    new_n26161_, new_n26162_, new_n26163_, new_n26164_, new_n26165_,
    new_n26166_, new_n26167_, new_n26168_, new_n26169_, new_n26170_,
    new_n26171_, new_n26172_, new_n26173_, new_n26174_, new_n26175_,
    new_n26176_, new_n26177_, new_n26178_, new_n26179_, new_n26180_,
    new_n26181_, new_n26182_, new_n26183_, new_n26184_, new_n26185_,
    new_n26186_, new_n26187_, new_n26188_, new_n26189_, new_n26190_,
    new_n26191_, new_n26192_, new_n26193_, new_n26194_, new_n26195_,
    new_n26196_, new_n26197_, new_n26198_, new_n26199_, new_n26200_,
    new_n26201_, new_n26202_, new_n26203_, new_n26204_, new_n26205_,
    new_n26206_, new_n26207_, new_n26208_, new_n26209_, new_n26210_,
    new_n26211_, new_n26212_, new_n26213_, new_n26214_, new_n26215_,
    new_n26216_, new_n26217_, new_n26218_, new_n26219_, new_n26220_,
    new_n26221_, new_n26222_, new_n26223_, new_n26224_, new_n26225_,
    new_n26226_, new_n26227_, new_n26228_, new_n26229_, new_n26230_,
    new_n26231_, new_n26232_, new_n26233_, new_n26234_, new_n26235_,
    new_n26236_, new_n26237_, new_n26238_, new_n26239_, new_n26240_,
    new_n26241_, new_n26242_, new_n26243_, new_n26244_, new_n26245_,
    new_n26246_, new_n26247_, new_n26248_, new_n26249_, new_n26250_,
    new_n26251_, new_n26252_, new_n26253_, new_n26254_, new_n26255_,
    new_n26256_, new_n26257_, new_n26258_, new_n26259_, new_n26260_,
    new_n26261_, new_n26262_, new_n26263_, new_n26264_, new_n26265_,
    new_n26266_, new_n26267_, new_n26268_, new_n26269_, new_n26270_,
    new_n26271_, new_n26272_, new_n26273_, new_n26274_, new_n26275_,
    new_n26276_, new_n26277_, new_n26278_, new_n26279_, new_n26280_,
    new_n26281_, new_n26282_, new_n26283_, new_n26284_, new_n26285_,
    new_n26286_, new_n26287_, new_n26288_, new_n26289_, new_n26290_,
    new_n26291_, new_n26292_, new_n26293_, new_n26294_, new_n26295_,
    new_n26296_, new_n26297_, new_n26298_, new_n26299_, new_n26300_,
    new_n26301_, new_n26302_, new_n26303_, new_n26304_, new_n26305_,
    new_n26306_, new_n26307_, new_n26308_, new_n26309_, new_n26310_,
    new_n26311_, new_n26312_, new_n26313_, new_n26314_, new_n26315_,
    new_n26316_, new_n26317_, new_n26318_, new_n26319_, new_n26320_,
    new_n26321_, new_n26322_, new_n26323_, new_n26324_, new_n26325_,
    new_n26326_, new_n26327_, new_n26328_, new_n26329_, new_n26330_,
    new_n26331_, new_n26332_, new_n26333_, new_n26334_, new_n26335_,
    new_n26336_, new_n26337_, new_n26338_, new_n26339_, new_n26340_,
    new_n26341_, new_n26342_, new_n26343_, new_n26344_, new_n26345_,
    new_n26346_, new_n26347_, new_n26348_, new_n26349_, new_n26350_,
    new_n26351_, new_n26352_, new_n26353_, new_n26354_, new_n26355_,
    new_n26356_, new_n26357_, new_n26358_, new_n26359_, new_n26360_,
    new_n26361_, new_n26362_, new_n26363_, new_n26364_, new_n26365_,
    new_n26366_, new_n26367_, new_n26368_, new_n26369_, new_n26370_,
    new_n26371_, new_n26372_, new_n26373_, new_n26374_, new_n26375_,
    new_n26376_, new_n26377_, new_n26378_, new_n26379_, new_n26380_,
    new_n26381_, new_n26382_, new_n26383_, new_n26384_, new_n26385_,
    new_n26386_, new_n26387_, new_n26388_, new_n26389_, new_n26390_,
    new_n26391_, new_n26392_, new_n26393_, new_n26394_, new_n26395_,
    new_n26396_, new_n26397_, new_n26398_, new_n26399_, new_n26400_,
    new_n26401_, new_n26402_, new_n26403_, new_n26404_, new_n26405_,
    new_n26406_, new_n26407_, new_n26408_, new_n26409_, new_n26410_,
    new_n26411_, new_n26412_, new_n26413_, new_n26414_, new_n26415_,
    new_n26416_, new_n26417_, new_n26418_, new_n26419_, new_n26420_,
    new_n26421_, new_n26422_, new_n26423_, new_n26424_, new_n26425_,
    new_n26426_, new_n26427_, new_n26428_, new_n26429_, new_n26430_,
    new_n26431_, new_n26432_, new_n26433_, new_n26434_, new_n26435_,
    new_n26436_, new_n26437_, new_n26438_, new_n26439_, new_n26440_,
    new_n26441_, new_n26442_, new_n26443_, new_n26444_, new_n26445_,
    new_n26446_, new_n26447_, new_n26448_, new_n26449_, new_n26450_,
    new_n26451_, new_n26452_, new_n26453_, new_n26454_, new_n26455_,
    new_n26456_, new_n26457_, new_n26458_, new_n26459_, new_n26460_,
    new_n26461_, new_n26462_, new_n26463_, new_n26464_, new_n26465_,
    new_n26466_, new_n26467_, new_n26468_, new_n26469_, new_n26470_,
    new_n26471_, new_n26472_, new_n26473_, new_n26474_, new_n26475_,
    new_n26476_, new_n26477_, new_n26478_, new_n26479_, new_n26480_,
    new_n26481_, new_n26482_, new_n26483_, new_n26484_, new_n26485_,
    new_n26486_, new_n26487_, new_n26488_, new_n26489_, new_n26490_,
    new_n26491_, new_n26492_, new_n26493_, new_n26494_, new_n26495_,
    new_n26496_, new_n26497_, new_n26498_, new_n26499_, new_n26500_,
    new_n26501_, new_n26502_, new_n26503_, new_n26504_, new_n26505_,
    new_n26506_, new_n26507_, new_n26508_, new_n26509_, new_n26510_,
    new_n26511_, new_n26512_, new_n26513_, new_n26514_, new_n26515_,
    new_n26516_, new_n26517_, new_n26518_, new_n26519_, new_n26520_,
    new_n26521_, new_n26522_, new_n26523_, new_n26524_, new_n26525_,
    new_n26526_, new_n26527_, new_n26528_, new_n26529_, new_n26530_,
    new_n26531_, new_n26532_, new_n26533_, new_n26534_, new_n26535_,
    new_n26536_, new_n26537_, new_n26538_, new_n26539_, new_n26540_,
    new_n26541_, new_n26542_, new_n26543_, new_n26544_, new_n26545_,
    new_n26546_, new_n26547_, new_n26548_, new_n26549_, new_n26550_,
    new_n26551_, new_n26552_, new_n26553_, new_n26554_, new_n26555_,
    new_n26556_, new_n26557_, new_n26558_, new_n26559_, new_n26560_,
    new_n26561_, new_n26562_, new_n26563_, new_n26564_, new_n26565_,
    new_n26566_, new_n26567_, new_n26568_, new_n26569_, new_n26570_,
    new_n26571_, new_n26572_, new_n26573_, new_n26574_, new_n26575_,
    new_n26576_, new_n26577_, new_n26578_, new_n26579_, new_n26580_,
    new_n26581_, new_n26582_, new_n26583_, new_n26584_, new_n26585_,
    new_n26586_, new_n26587_, new_n26588_, new_n26589_, new_n26590_,
    new_n26591_, new_n26592_, new_n26593_, new_n26594_, new_n26595_,
    new_n26596_, new_n26597_, new_n26598_, new_n26599_, new_n26600_,
    new_n26601_, new_n26602_, new_n26603_, new_n26604_, new_n26605_,
    new_n26606_, new_n26607_, new_n26608_, new_n26609_, new_n26610_,
    new_n26611_, new_n26612_, new_n26613_, new_n26614_, new_n26615_,
    new_n26616_, new_n26617_, new_n26618_, new_n26619_, new_n26620_,
    new_n26621_, new_n26622_, new_n26623_, new_n26624_, new_n26625_,
    new_n26626_, new_n26627_, new_n26628_, new_n26629_, new_n26630_,
    new_n26631_, new_n26632_, new_n26633_, new_n26634_, new_n26635_,
    new_n26636_, new_n26637_, new_n26638_, new_n26639_, new_n26640_,
    new_n26641_, new_n26642_, new_n26643_, new_n26644_, new_n26645_,
    new_n26646_, new_n26647_, new_n26648_, new_n26649_, new_n26650_,
    new_n26651_, new_n26652_, new_n26653_, new_n26654_, new_n26655_,
    new_n26656_, new_n26657_, new_n26658_, new_n26659_, new_n26660_,
    new_n26661_, new_n26662_, new_n26663_, new_n26664_, new_n26665_,
    new_n26666_, new_n26667_, new_n26668_, new_n26669_, new_n26670_,
    new_n26671_, new_n26672_, new_n26673_, new_n26674_, new_n26675_,
    new_n26676_, new_n26677_, new_n26678_, new_n26679_, new_n26680_,
    new_n26681_, new_n26682_, new_n26683_, new_n26684_, new_n26685_,
    new_n26686_, new_n26687_, new_n26688_, new_n26689_, new_n26690_,
    new_n26691_, new_n26692_, new_n26693_, new_n26694_, new_n26695_,
    new_n26696_, new_n26697_, new_n26698_, new_n26699_, new_n26700_,
    new_n26701_, new_n26702_, new_n26703_, new_n26704_, new_n26705_,
    new_n26706_, new_n26707_, new_n26708_, new_n26709_, new_n26710_,
    new_n26711_, new_n26712_, new_n26713_, new_n26714_, new_n26715_,
    new_n26716_, new_n26717_, new_n26718_, new_n26719_, new_n26720_,
    new_n26721_, new_n26722_, new_n26723_, new_n26724_, new_n26725_,
    new_n26726_, new_n26727_, new_n26728_, new_n26729_, new_n26730_,
    new_n26731_, new_n26732_, new_n26733_, new_n26734_, new_n26735_,
    new_n26736_, new_n26737_, new_n26738_, new_n26739_, new_n26740_,
    new_n26741_, new_n26742_, new_n26743_, new_n26744_, new_n26745_,
    new_n26746_, new_n26747_, new_n26748_, new_n26749_, new_n26750_,
    new_n26751_, new_n26752_, new_n26753_, new_n26754_, new_n26755_,
    new_n26756_, new_n26757_, new_n26758_, new_n26759_, new_n26760_,
    new_n26761_, new_n26762_, new_n26763_, new_n26764_, new_n26765_,
    new_n26766_, new_n26767_, new_n26768_, new_n26769_, new_n26770_,
    new_n26771_, new_n26772_, new_n26773_, new_n26774_, new_n26775_,
    new_n26776_, new_n26777_, new_n26778_, new_n26779_, new_n26780_,
    new_n26781_, new_n26782_, new_n26783_, new_n26784_, new_n26785_,
    new_n26786_, new_n26787_, new_n26788_, new_n26789_, new_n26790_,
    new_n26791_, new_n26792_, new_n26793_, new_n26794_, new_n26795_,
    new_n26796_, new_n26797_, new_n26798_, new_n26799_, new_n26800_,
    new_n26801_, new_n26802_, new_n26803_, new_n26804_, new_n26805_,
    new_n26806_, new_n26807_, new_n26808_, new_n26809_, new_n26810_,
    new_n26811_, new_n26812_, new_n26813_, new_n26814_, new_n26815_,
    new_n26816_, new_n26817_, new_n26818_, new_n26819_, new_n26820_,
    new_n26821_, new_n26822_, new_n26823_, new_n26824_, new_n26825_,
    new_n26826_, new_n26827_, new_n26828_, new_n26829_, new_n26830_,
    new_n26831_, new_n26832_, new_n26833_, new_n26834_, new_n26835_,
    new_n26836_, new_n26837_, new_n26838_, new_n26839_, new_n26840_,
    new_n26841_, new_n26842_, new_n26843_, new_n26844_, new_n26845_,
    new_n26846_, new_n26847_, new_n26848_, new_n26849_, new_n26850_,
    new_n26851_, new_n26852_, new_n26853_, new_n26854_, new_n26855_,
    new_n26856_, new_n26857_, new_n26858_, new_n26859_, new_n26860_,
    new_n26861_, new_n26862_, new_n26863_, new_n26864_, new_n26865_,
    new_n26866_, new_n26867_, new_n26868_, new_n26869_, new_n26870_,
    new_n26871_, new_n26872_, new_n26873_, new_n26874_, new_n26875_,
    new_n26876_, new_n26877_, new_n26878_, new_n26879_, new_n26880_,
    new_n26881_, new_n26882_, new_n26883_, new_n26884_, new_n26885_,
    new_n26886_, new_n26887_, new_n26888_, new_n26889_, new_n26890_,
    new_n26891_, new_n26892_, new_n26893_, new_n26894_, new_n26895_,
    new_n26896_, new_n26897_, new_n26898_, new_n26899_, new_n26900_,
    new_n26901_, new_n26902_, new_n26903_, new_n26904_, new_n26905_,
    new_n26906_, new_n26907_, new_n26908_, new_n26909_, new_n26910_,
    new_n26911_, new_n26912_, new_n26913_, new_n26914_, new_n26915_,
    new_n26916_, new_n26917_, new_n26918_, new_n26919_, new_n26920_,
    new_n26921_, new_n26922_, new_n26923_, new_n26924_, new_n26925_,
    new_n26926_, new_n26927_, new_n26928_, new_n26929_, new_n26930_,
    new_n26931_, new_n26932_, new_n26933_, new_n26934_, new_n26935_,
    new_n26936_, new_n26937_, new_n26938_, new_n26939_, new_n26940_,
    new_n26941_, new_n26942_, new_n26943_, new_n26944_, new_n26945_,
    new_n26946_, new_n26947_, new_n26948_, new_n26949_, new_n26950_,
    new_n26951_, new_n26952_, new_n26953_, new_n26954_, new_n26955_,
    new_n26956_, new_n26957_, new_n26958_, new_n26959_, new_n26960_,
    new_n26961_, new_n26962_, new_n26963_, new_n26964_, new_n26965_,
    new_n26966_, new_n26967_, new_n26968_, new_n26969_, new_n26970_,
    new_n26971_, new_n26972_, new_n26973_, new_n26974_, new_n26975_,
    new_n26976_, new_n26977_, new_n26978_, new_n26979_, new_n26980_,
    new_n26981_, new_n26982_, new_n26983_, new_n26984_, new_n26985_,
    new_n26986_, new_n26987_, new_n26988_, new_n26989_, new_n26990_,
    new_n26991_, new_n26992_, new_n26993_, new_n26994_, new_n26995_,
    new_n26996_, new_n26997_, new_n26998_, new_n26999_, new_n27000_,
    new_n27001_, new_n27002_, new_n27003_, new_n27004_, new_n27005_,
    new_n27006_, new_n27007_, new_n27008_, new_n27009_, new_n27010_,
    new_n27011_, new_n27012_, new_n27013_, new_n27014_, new_n27015_,
    new_n27016_, new_n27017_, new_n27018_, new_n27019_, new_n27020_,
    new_n27021_, new_n27022_, new_n27023_, new_n27024_, new_n27025_,
    new_n27026_, new_n27027_, new_n27028_, new_n27029_, new_n27030_,
    new_n27031_, new_n27032_, new_n27033_, new_n27034_, new_n27035_,
    new_n27036_, new_n27037_, new_n27038_, new_n27039_, new_n27040_,
    new_n27041_, new_n27042_, new_n27043_, new_n27044_, new_n27045_,
    new_n27046_, new_n27047_, new_n27048_, new_n27049_, new_n27050_,
    new_n27051_, new_n27052_, new_n27053_, new_n27054_, new_n27055_,
    new_n27056_, new_n27057_, new_n27058_, new_n27059_, new_n27060_,
    new_n27061_, new_n27062_, new_n27063_, new_n27064_, new_n27065_,
    new_n27066_, new_n27067_, new_n27068_, new_n27069_, new_n27070_,
    new_n27071_, new_n27072_, new_n27073_, new_n27074_, new_n27075_,
    new_n27076_, new_n27077_, new_n27078_, new_n27079_, new_n27080_,
    new_n27081_, new_n27082_, new_n27083_, new_n27084_, new_n27085_,
    new_n27086_, new_n27087_, new_n27088_, new_n27089_, new_n27090_,
    new_n27091_, new_n27092_, new_n27093_, new_n27094_, new_n27095_,
    new_n27096_, new_n27097_, new_n27098_, new_n27099_, new_n27100_,
    new_n27101_, new_n27102_, new_n27103_, new_n27104_, new_n27105_,
    new_n27106_, new_n27107_, new_n27108_, new_n27109_, new_n27110_,
    new_n27111_, new_n27112_, new_n27113_, new_n27114_, new_n27115_,
    new_n27116_, new_n27117_, new_n27118_, new_n27119_, new_n27120_,
    new_n27121_, new_n27122_, new_n27123_, new_n27124_, new_n27125_,
    new_n27126_, new_n27127_, new_n27128_, new_n27129_, new_n27130_,
    new_n27131_, new_n27132_, new_n27133_, new_n27134_, new_n27135_,
    new_n27136_, new_n27137_, new_n27138_, new_n27139_, new_n27140_,
    new_n27141_, new_n27142_, new_n27143_, new_n27144_, new_n27145_,
    new_n27146_, new_n27147_, new_n27148_, new_n27149_, new_n27150_,
    new_n27151_, new_n27152_, new_n27153_, new_n27154_, new_n27155_,
    new_n27156_, new_n27157_, new_n27158_, new_n27159_, new_n27160_,
    new_n27161_, new_n27162_, new_n27163_, new_n27164_, new_n27165_,
    new_n27166_, new_n27167_, new_n27168_, new_n27169_, new_n27170_,
    new_n27171_, new_n27172_, new_n27173_, new_n27174_, new_n27175_,
    new_n27176_, new_n27177_, new_n27178_, new_n27179_, new_n27180_,
    new_n27181_, new_n27182_, new_n27183_, new_n27184_, new_n27185_,
    new_n27186_, new_n27187_, new_n27188_, new_n27189_, new_n27190_,
    new_n27191_, new_n27192_, new_n27193_, new_n27194_, new_n27195_,
    new_n27196_, new_n27197_, new_n27198_, new_n27199_, new_n27200_,
    new_n27201_, new_n27202_, new_n27203_, new_n27204_, new_n27205_,
    new_n27206_, new_n27207_, new_n27208_, new_n27209_, new_n27210_,
    new_n27211_, new_n27212_, new_n27213_, new_n27214_, new_n27215_,
    new_n27216_, new_n27217_, new_n27218_, new_n27219_, new_n27220_,
    new_n27221_, new_n27222_, new_n27223_, new_n27224_, new_n27225_,
    new_n27226_, new_n27227_, new_n27228_, new_n27229_, new_n27230_,
    new_n27231_, new_n27232_, new_n27233_, new_n27234_, new_n27235_,
    new_n27236_, new_n27237_, new_n27238_, new_n27239_, new_n27240_,
    new_n27241_, new_n27242_, new_n27243_, new_n27244_, new_n27245_,
    new_n27246_, new_n27247_, new_n27248_, new_n27249_, new_n27250_,
    new_n27251_, new_n27252_, new_n27253_, new_n27254_, new_n27255_,
    new_n27256_, new_n27257_, new_n27258_, new_n27259_, new_n27260_,
    new_n27261_, new_n27262_, new_n27263_, new_n27264_, new_n27265_,
    new_n27266_, new_n27267_, new_n27268_, new_n27269_, new_n27270_,
    new_n27271_, new_n27272_, new_n27273_, new_n27274_, new_n27275_,
    new_n27276_, new_n27277_, new_n27278_, new_n27279_, new_n27280_,
    new_n27281_, new_n27282_, new_n27283_, new_n27284_, new_n27285_,
    new_n27286_, new_n27287_, new_n27288_, new_n27289_, new_n27290_,
    new_n27291_, new_n27292_, new_n27293_, new_n27294_, new_n27295_,
    new_n27296_, new_n27297_, new_n27298_, new_n27299_, new_n27300_,
    new_n27301_, new_n27302_, new_n27303_, new_n27304_, new_n27305_,
    new_n27306_, new_n27307_, new_n27308_, new_n27309_, new_n27310_,
    new_n27311_, new_n27312_, new_n27313_, new_n27314_, new_n27315_,
    new_n27316_, new_n27317_, new_n27318_, new_n27319_, new_n27320_,
    new_n27321_, new_n27322_, new_n27323_, new_n27324_, new_n27325_,
    new_n27326_, new_n27327_, new_n27328_, new_n27329_, new_n27330_,
    new_n27331_, new_n27332_, new_n27333_, new_n27334_, new_n27335_,
    new_n27336_, new_n27337_, new_n27338_, new_n27339_, new_n27340_,
    new_n27341_, new_n27342_, new_n27343_, new_n27344_, new_n27345_,
    new_n27346_, new_n27347_, new_n27348_, new_n27349_, new_n27350_,
    new_n27351_, new_n27352_, new_n27353_, new_n27354_, new_n27355_,
    new_n27356_, new_n27357_, new_n27358_, new_n27359_, new_n27360_,
    new_n27361_, new_n27362_, new_n27363_, new_n27364_, new_n27365_,
    new_n27366_, new_n27367_, new_n27368_, new_n27369_, new_n27370_,
    new_n27371_, new_n27372_, new_n27373_, new_n27374_, new_n27375_,
    new_n27376_, new_n27377_, new_n27378_, new_n27379_, new_n27380_,
    new_n27381_, new_n27382_, new_n27383_, new_n27384_, new_n27385_,
    new_n27386_, new_n27387_, new_n27388_, new_n27389_, new_n27390_,
    new_n27391_, new_n27392_, new_n27393_, new_n27394_, new_n27395_,
    new_n27396_, new_n27397_, new_n27398_, new_n27399_, new_n27400_,
    new_n27401_, new_n27402_, new_n27403_, new_n27404_, new_n27405_,
    new_n27406_, new_n27407_, new_n27408_, new_n27409_, new_n27410_,
    new_n27411_, new_n27412_, new_n27413_, new_n27414_, new_n27415_,
    new_n27416_, new_n27417_, new_n27418_, new_n27419_, new_n27420_,
    new_n27421_, new_n27422_, new_n27423_, new_n27424_, new_n27425_,
    new_n27426_, new_n27427_, new_n27428_, new_n27429_, new_n27430_,
    new_n27431_, new_n27432_, new_n27433_, new_n27434_, new_n27435_,
    new_n27436_, new_n27437_, new_n27438_, new_n27439_, new_n27440_,
    new_n27441_, new_n27442_, new_n27443_, new_n27444_, new_n27445_,
    new_n27446_, new_n27447_, new_n27448_, new_n27449_, new_n27450_,
    new_n27451_, new_n27452_, new_n27453_, new_n27454_, new_n27455_,
    new_n27456_, new_n27457_, new_n27458_, new_n27459_, new_n27460_,
    new_n27461_, new_n27462_, new_n27463_, new_n27464_, new_n27465_,
    new_n27466_, new_n27467_, new_n27468_, new_n27469_, new_n27470_,
    new_n27471_, new_n27472_, new_n27473_, new_n27474_, new_n27475_,
    new_n27476_, new_n27477_, new_n27478_, new_n27479_, new_n27480_,
    new_n27481_, new_n27482_, new_n27483_, new_n27484_, new_n27485_,
    new_n27486_, new_n27487_, new_n27488_, new_n27489_, new_n27490_,
    new_n27491_, new_n27492_, new_n27493_, new_n27494_, new_n27495_,
    new_n27496_, new_n27497_, new_n27498_, new_n27499_, new_n27500_,
    new_n27501_, new_n27502_, new_n27503_, new_n27504_, new_n27505_,
    new_n27506_, new_n27507_, new_n27508_, new_n27509_, new_n27510_,
    new_n27511_, new_n27512_, new_n27513_, new_n27514_, new_n27515_,
    new_n27516_, new_n27517_, new_n27518_, new_n27519_, new_n27520_,
    new_n27521_, new_n27522_, new_n27523_, new_n27524_, new_n27525_,
    new_n27526_, new_n27527_, new_n27528_, new_n27529_, new_n27530_,
    new_n27531_, new_n27532_, new_n27533_, new_n27534_, new_n27535_,
    new_n27536_, new_n27537_, new_n27538_, new_n27539_, new_n27540_,
    new_n27541_, new_n27542_, new_n27543_, new_n27544_, new_n27545_,
    new_n27546_, new_n27547_, new_n27548_, new_n27549_, new_n27550_,
    new_n27551_, new_n27552_, new_n27553_, new_n27554_, new_n27555_,
    new_n27556_, new_n27557_, new_n27558_, new_n27559_, new_n27560_,
    new_n27561_, new_n27562_, new_n27563_, new_n27564_, new_n27565_,
    new_n27566_, new_n27567_, new_n27568_, new_n27569_, new_n27570_,
    new_n27571_, new_n27572_, new_n27573_, new_n27574_, new_n27575_,
    new_n27576_, new_n27577_, new_n27578_, new_n27579_, new_n27580_,
    new_n27581_, new_n27582_, new_n27583_, new_n27584_, new_n27585_,
    new_n27586_, new_n27587_, new_n27588_, new_n27589_, new_n27590_,
    new_n27591_, new_n27592_, new_n27593_, new_n27594_, new_n27595_,
    new_n27596_, new_n27597_, new_n27598_, new_n27599_, new_n27600_,
    new_n27601_, new_n27602_, new_n27603_, new_n27604_, new_n27605_,
    new_n27606_, new_n27607_, new_n27608_, new_n27609_, new_n27610_,
    new_n27611_, new_n27612_, new_n27613_, new_n27614_, new_n27615_,
    new_n27616_, new_n27617_, new_n27618_, new_n27619_, new_n27620_,
    new_n27621_, new_n27622_, new_n27623_, new_n27624_, new_n27625_,
    new_n27626_, new_n27627_, new_n27628_, new_n27629_, new_n27630_,
    new_n27631_, new_n27632_, new_n27633_, new_n27634_, new_n27635_,
    new_n27636_, new_n27637_, new_n27638_, new_n27639_, new_n27640_,
    new_n27641_, new_n27642_, new_n27643_, new_n27644_, new_n27645_,
    new_n27646_, new_n27647_, new_n27648_, new_n27649_, new_n27650_,
    new_n27651_, new_n27652_, new_n27653_, new_n27654_, new_n27655_,
    new_n27656_, new_n27657_, new_n27658_, new_n27659_, new_n27660_,
    new_n27661_, new_n27662_, new_n27663_, new_n27664_, new_n27665_,
    new_n27666_, new_n27667_, new_n27668_, new_n27669_, new_n27670_,
    new_n27671_, new_n27672_, new_n27673_, new_n27674_, new_n27675_,
    new_n27676_, new_n27677_, new_n27678_, new_n27679_, new_n27680_,
    new_n27681_, new_n27682_, new_n27683_, new_n27684_, new_n27685_,
    new_n27686_, new_n27687_, new_n27688_, new_n27689_, new_n27690_,
    new_n27691_, new_n27692_, new_n27693_, new_n27694_, new_n27695_,
    new_n27696_, new_n27697_, new_n27698_, new_n27699_, new_n27700_,
    new_n27701_, new_n27702_, new_n27703_, new_n27704_, new_n27705_,
    new_n27706_, new_n27707_, new_n27708_, new_n27709_, new_n27710_,
    new_n27711_, new_n27712_, new_n27713_, new_n27714_, new_n27715_,
    new_n27716_, new_n27717_, new_n27718_, new_n27719_, new_n27720_,
    new_n27721_, new_n27722_, new_n27723_, new_n27724_, new_n27725_,
    new_n27726_, new_n27727_, new_n27728_, new_n27729_, new_n27730_,
    new_n27731_, new_n27732_, new_n27733_, new_n27734_, new_n27735_,
    new_n27736_, new_n27737_, new_n27738_, new_n27739_, new_n27740_,
    new_n27741_, new_n27742_, new_n27743_, new_n27744_, new_n27745_,
    new_n27746_, new_n27747_, new_n27748_, new_n27749_, new_n27750_,
    new_n27751_, new_n27752_, new_n27753_, new_n27754_, new_n27755_,
    new_n27756_, new_n27757_, new_n27758_, new_n27759_, new_n27760_,
    new_n27761_, new_n27762_, new_n27763_, new_n27764_, new_n27765_,
    new_n27766_, new_n27767_, new_n27768_, new_n27769_, new_n27770_,
    new_n27771_, new_n27772_, new_n27773_, new_n27774_, new_n27775_,
    new_n27776_, new_n27777_, new_n27778_, new_n27779_, new_n27780_,
    new_n27781_, new_n27782_, new_n27783_, new_n27784_, new_n27785_,
    new_n27786_, new_n27787_, new_n27788_, new_n27789_, new_n27790_,
    new_n27791_, new_n27792_, new_n27793_, new_n27794_, new_n27795_,
    new_n27796_, new_n27797_, new_n27798_, new_n27799_, new_n27800_,
    new_n27801_, new_n27802_, new_n27803_, new_n27804_, new_n27805_,
    new_n27806_, new_n27807_, new_n27808_, new_n27809_, new_n27810_,
    new_n27811_, new_n27812_, new_n27813_, new_n27814_, new_n27815_,
    new_n27816_, new_n27817_, new_n27818_, new_n27819_, new_n27820_,
    new_n27821_, new_n27822_, new_n27823_, new_n27824_, new_n27825_,
    new_n27826_, new_n27827_, new_n27828_, new_n27829_, new_n27830_,
    new_n27831_, new_n27832_, new_n27833_, new_n27834_, new_n27835_,
    new_n27836_, new_n27837_, new_n27838_, new_n27839_, new_n27840_,
    new_n27841_, new_n27842_, new_n27843_, new_n27844_, new_n27845_,
    new_n27846_, new_n27847_, new_n27848_, new_n27849_, new_n27850_,
    new_n27851_, new_n27852_, new_n27853_, new_n27854_, new_n27855_,
    new_n27856_, new_n27857_, new_n27858_, new_n27859_, new_n27860_,
    new_n27861_, new_n27862_, new_n27863_, new_n27864_, new_n27865_,
    new_n27866_, new_n27867_, new_n27868_, new_n27869_, new_n27870_,
    new_n27871_, new_n27872_, new_n27873_, new_n27874_, new_n27875_,
    new_n27876_, new_n27877_, new_n27878_, new_n27879_, new_n27880_,
    new_n27881_, new_n27882_, new_n27883_, new_n27884_, new_n27885_,
    new_n27886_, new_n27887_, new_n27888_, new_n27889_, new_n27890_,
    new_n27891_, new_n27892_, new_n27893_, new_n27894_, new_n27895_,
    new_n27896_, new_n27897_, new_n27898_, new_n27899_, new_n27900_,
    new_n27901_, new_n27902_, new_n27903_, new_n27904_, new_n27905_,
    new_n27906_, new_n27907_, new_n27908_, new_n27909_, new_n27910_,
    new_n27911_, new_n27912_, new_n27913_, new_n27914_, new_n27915_,
    new_n27916_, new_n27917_, new_n27918_, new_n27919_, new_n27920_,
    new_n27921_, new_n27922_, new_n27923_, new_n27924_, new_n27925_,
    new_n27926_, new_n27927_, new_n27928_, new_n27929_, new_n27930_,
    new_n27931_, new_n27932_, new_n27933_, new_n27934_, new_n27935_,
    new_n27936_, new_n27937_, new_n27938_, new_n27939_, new_n27940_,
    new_n27941_, new_n27942_, new_n27943_, new_n27944_, new_n27945_,
    new_n27946_, new_n27947_, new_n27948_, new_n27949_, new_n27950_,
    new_n27951_, new_n27952_, new_n27953_, new_n27954_, new_n27955_,
    new_n27956_, new_n27957_, new_n27958_, new_n27959_, new_n27960_,
    new_n27961_, new_n27962_, new_n27963_, new_n27964_, new_n27965_,
    new_n27966_, new_n27967_, new_n27968_, new_n27969_, new_n27970_,
    new_n27971_, new_n27972_, new_n27973_, new_n27974_, new_n27975_,
    new_n27976_, new_n27977_, new_n27978_, new_n27979_, new_n27980_,
    new_n27981_, new_n27982_, new_n27983_, new_n27984_, new_n27985_,
    new_n27986_, new_n27987_, new_n27988_, new_n27989_, new_n27990_,
    new_n27991_, new_n27992_, new_n27993_, new_n27994_, new_n27995_,
    new_n27996_, new_n27997_, new_n27998_, new_n27999_, new_n28000_,
    new_n28001_, new_n28002_, new_n28003_, new_n28004_, new_n28005_,
    new_n28006_, new_n28007_, new_n28008_, new_n28009_, new_n28010_,
    new_n28011_, new_n28012_, new_n28013_, new_n28014_, new_n28015_,
    new_n28016_, new_n28017_, new_n28018_, new_n28019_, new_n28020_,
    new_n28021_, new_n28022_, new_n28023_, new_n28024_, new_n28025_,
    new_n28026_, new_n28027_, new_n28028_, new_n28029_, new_n28030_,
    new_n28031_, new_n28032_, new_n28033_, new_n28034_, new_n28035_,
    new_n28036_, new_n28037_, new_n28038_, new_n28039_, new_n28040_,
    new_n28041_, new_n28042_, new_n28043_, new_n28044_, new_n28045_,
    new_n28046_, new_n28047_, new_n28048_, new_n28049_, new_n28050_,
    new_n28051_, new_n28052_, new_n28053_, new_n28054_, new_n28055_,
    new_n28056_, new_n28057_, new_n28058_, new_n28059_, new_n28060_,
    new_n28061_, new_n28062_, new_n28063_, new_n28064_, new_n28065_,
    new_n28066_, new_n28067_, new_n28068_, new_n28069_, new_n28070_,
    new_n28071_, new_n28072_, new_n28073_, new_n28074_, new_n28075_,
    new_n28076_, new_n28077_, new_n28078_, new_n28079_, new_n28080_,
    new_n28081_, new_n28082_, new_n28083_, new_n28084_, new_n28085_,
    new_n28086_, new_n28087_, new_n28088_, new_n28089_, new_n28090_,
    new_n28091_, new_n28092_, new_n28093_, new_n28094_, new_n28095_,
    new_n28096_, new_n28097_, new_n28098_, new_n28099_, new_n28100_,
    new_n28101_, new_n28102_, new_n28103_, new_n28104_, new_n28105_,
    new_n28106_, new_n28107_, new_n28108_, new_n28109_, new_n28110_,
    new_n28111_, new_n28112_, new_n28113_, new_n28114_, new_n28115_,
    new_n28116_, new_n28117_, new_n28118_, new_n28119_, new_n28120_,
    new_n28121_, new_n28122_, new_n28123_, new_n28124_, new_n28125_,
    new_n28126_, new_n28127_, new_n28128_, new_n28129_, new_n28130_,
    new_n28131_, new_n28132_, new_n28133_, new_n28134_, new_n28135_,
    new_n28136_, new_n28137_, new_n28138_, new_n28139_, new_n28140_,
    new_n28141_, new_n28142_, new_n28143_, new_n28144_, new_n28145_,
    new_n28146_, new_n28147_, new_n28148_, new_n28149_, new_n28150_,
    new_n28151_, new_n28152_, new_n28153_, new_n28154_, new_n28155_,
    new_n28156_, new_n28157_, new_n28158_, new_n28159_, new_n28160_,
    new_n28161_, new_n28162_, new_n28163_, new_n28164_, new_n28165_,
    new_n28166_, new_n28167_, new_n28168_, new_n28169_, new_n28170_,
    new_n28171_, new_n28172_, new_n28173_, new_n28174_, new_n28175_,
    new_n28176_, new_n28177_, new_n28178_, new_n28179_, new_n28180_,
    new_n28181_, new_n28182_, new_n28183_, new_n28184_, new_n28185_,
    new_n28186_, new_n28187_, new_n28188_, new_n28189_, new_n28190_,
    new_n28191_, new_n28192_, new_n28193_, new_n28194_, new_n28195_,
    new_n28196_, new_n28197_, new_n28198_, new_n28199_, new_n28200_,
    new_n28201_, new_n28202_, new_n28203_, new_n28204_, new_n28205_,
    new_n28206_, new_n28207_, new_n28208_, new_n28209_, new_n28210_,
    new_n28211_, new_n28212_, new_n28213_, new_n28214_, new_n28215_,
    new_n28216_, new_n28217_, new_n28218_, new_n28219_, new_n28220_,
    new_n28221_, new_n28222_, new_n28223_, new_n28224_, new_n28225_,
    new_n28226_, new_n28227_, new_n28228_, new_n28229_, new_n28230_,
    new_n28231_, new_n28232_, new_n28233_, new_n28234_, new_n28235_,
    new_n28236_, new_n28237_, new_n28238_, new_n28239_, new_n28240_,
    new_n28241_, new_n28242_, new_n28243_, new_n28244_, new_n28245_,
    new_n28246_, new_n28247_, new_n28248_, new_n28249_, new_n28250_,
    new_n28251_, new_n28252_, new_n28253_, new_n28254_, new_n28255_,
    new_n28256_, new_n28257_, new_n28258_, new_n28259_, new_n28260_,
    new_n28261_, new_n28262_, new_n28263_, new_n28264_, new_n28265_,
    new_n28266_, new_n28267_, new_n28268_, new_n28269_, new_n28270_,
    new_n28271_, new_n28272_, new_n28273_, new_n28274_, new_n28275_,
    new_n28276_, new_n28277_, new_n28278_, new_n28279_, new_n28280_,
    new_n28281_, new_n28282_, new_n28283_, new_n28284_, new_n28285_,
    new_n28286_, new_n28287_, new_n28288_, new_n28289_, new_n28290_,
    new_n28291_, new_n28292_, new_n28293_, new_n28294_, new_n28295_,
    new_n28296_, new_n28297_, new_n28298_, new_n28299_, new_n28300_,
    new_n28301_, new_n28302_, new_n28303_, new_n28304_, new_n28305_,
    new_n28306_, new_n28307_, new_n28308_, new_n28309_, new_n28310_,
    new_n28311_, new_n28312_, new_n28313_, new_n28314_, new_n28315_,
    new_n28316_, new_n28317_, new_n28318_, new_n28319_, new_n28320_,
    new_n28321_, new_n28322_, new_n28323_, new_n28324_, new_n28325_,
    new_n28326_, new_n28327_, new_n28328_, new_n28329_, new_n28330_,
    new_n28331_, new_n28332_, new_n28333_, new_n28334_, new_n28335_,
    new_n28336_, new_n28337_, new_n28338_, new_n28339_, new_n28340_,
    new_n28341_, new_n28342_, new_n28343_, new_n28344_, new_n28345_,
    new_n28346_, new_n28347_, new_n28348_, new_n28349_, new_n28350_,
    new_n28351_, new_n28352_, new_n28353_, new_n28354_, new_n28355_,
    new_n28356_, new_n28357_, new_n28358_, new_n28359_, new_n28360_,
    new_n28361_, new_n28362_, new_n28363_, new_n28364_, new_n28365_,
    new_n28366_, new_n28367_, new_n28368_, new_n28369_, new_n28370_,
    new_n28371_, new_n28372_, new_n28373_, new_n28374_, new_n28375_,
    new_n28376_, new_n28377_, new_n28378_, new_n28379_, new_n28380_,
    new_n28381_, new_n28382_, new_n28383_, new_n28384_, new_n28385_,
    new_n28386_, new_n28387_, new_n28388_, new_n28389_, new_n28390_,
    new_n28391_, new_n28392_, new_n28393_, new_n28394_, new_n28395_,
    new_n28396_, new_n28397_, new_n28398_, new_n28399_, new_n28400_,
    new_n28401_, new_n28402_, new_n28403_, new_n28404_, new_n28405_,
    new_n28406_, new_n28407_, new_n28408_, new_n28409_, new_n28410_,
    new_n28411_, new_n28412_, new_n28413_, new_n28414_, new_n28415_,
    new_n28416_, new_n28417_, new_n28418_, new_n28419_, new_n28420_,
    new_n28421_, new_n28422_, new_n28423_, new_n28424_, new_n28425_,
    new_n28426_, new_n28427_, new_n28428_, new_n28429_, new_n28430_,
    new_n28431_, new_n28432_, new_n28433_, new_n28434_, new_n28435_,
    new_n28436_, new_n28437_, new_n28438_, new_n28439_, new_n28440_,
    new_n28441_, new_n28442_, new_n28443_, new_n28444_, new_n28445_,
    new_n28446_, new_n28447_, new_n28448_, new_n28449_, new_n28450_,
    new_n28451_, new_n28452_, new_n28453_, new_n28454_, new_n28455_,
    new_n28456_, new_n28457_, new_n28458_, new_n28459_, new_n28460_,
    new_n28461_, new_n28462_, new_n28463_, new_n28464_, new_n28465_,
    new_n28466_, new_n28467_, new_n28468_, new_n28469_, new_n28470_,
    new_n28471_, new_n28472_, new_n28473_, new_n28474_, new_n28475_,
    new_n28476_, new_n28477_, new_n28478_, new_n28479_, new_n28480_,
    new_n28481_, new_n28482_, new_n28483_, new_n28484_, new_n28485_,
    new_n28486_, new_n28487_, new_n28488_, new_n28489_, new_n28490_,
    new_n28491_, new_n28492_, new_n28493_, new_n28494_, new_n28495_,
    new_n28496_, new_n28497_, new_n28498_, new_n28499_, new_n28500_,
    new_n28501_, new_n28502_, new_n28503_, new_n28504_, new_n28505_,
    new_n28506_, new_n28507_, new_n28508_, new_n28509_, new_n28510_,
    new_n28511_, new_n28512_, new_n28513_, new_n28514_, new_n28515_,
    new_n28516_, new_n28517_, new_n28518_, new_n28519_, new_n28520_,
    new_n28521_, new_n28522_, new_n28523_, new_n28524_, new_n28525_,
    new_n28526_, new_n28527_, new_n28528_, new_n28529_, new_n28530_,
    new_n28531_, new_n28532_, new_n28533_, new_n28534_, new_n28535_,
    new_n28536_, new_n28537_, new_n28538_, new_n28539_, new_n28540_,
    new_n28541_, new_n28542_, new_n28543_, new_n28544_, new_n28545_,
    new_n28546_, new_n28547_, new_n28548_, new_n28549_, new_n28550_,
    new_n28551_, new_n28552_, new_n28553_, new_n28554_, new_n28555_,
    new_n28556_, new_n28557_, new_n28558_, new_n28559_, new_n28560_,
    new_n28561_, new_n28562_, new_n28563_, new_n28564_, new_n28565_,
    new_n28566_, new_n28567_, new_n28568_, new_n28569_, new_n28570_,
    new_n28571_, new_n28572_, new_n28573_, new_n28574_, new_n28575_,
    new_n28576_, new_n28577_, new_n28578_, new_n28579_, new_n28580_,
    new_n28581_, new_n28582_, new_n28583_, new_n28584_, new_n28585_,
    new_n28586_, new_n28587_, new_n28588_, new_n28589_, new_n28590_,
    new_n28591_, new_n28592_, new_n28593_, new_n28594_, new_n28595_,
    new_n28596_, new_n28597_, new_n28598_, new_n28599_, new_n28600_,
    new_n28601_, new_n28602_, new_n28603_, new_n28604_, new_n28605_,
    new_n28606_, new_n28607_, new_n28608_, new_n28609_, new_n28610_,
    new_n28611_, new_n28612_, new_n28613_, new_n28614_, new_n28615_,
    new_n28616_, new_n28617_, new_n28618_, new_n28619_, new_n28620_,
    new_n28621_, new_n28622_, new_n28623_, new_n28624_, new_n28625_,
    new_n28626_, new_n28627_, new_n28628_, new_n28629_, new_n28630_,
    new_n28631_, new_n28632_, new_n28633_, new_n28634_, new_n28635_,
    new_n28636_, new_n28637_, new_n28638_, new_n28639_, new_n28640_,
    new_n28641_, new_n28642_, new_n28643_, new_n28644_, new_n28645_,
    new_n28646_, new_n28647_, new_n28648_, new_n28649_, new_n28650_,
    new_n28651_, new_n28652_, new_n28653_, new_n28654_, new_n28655_,
    new_n28656_, new_n28657_, new_n28658_, new_n28659_, new_n28660_,
    new_n28661_, new_n28662_, new_n28663_, new_n28664_, new_n28665_,
    new_n28666_, new_n28667_, new_n28668_, new_n28669_, new_n28670_,
    new_n28671_, new_n28672_, new_n28673_, new_n28674_, new_n28675_,
    new_n28676_, new_n28677_, new_n28678_, new_n28679_, new_n28680_,
    new_n28681_, new_n28682_, new_n28683_, new_n28684_, new_n28685_,
    new_n28686_, new_n28687_, new_n28688_, new_n28689_, new_n28690_,
    new_n28691_, new_n28692_, new_n28693_, new_n28694_, new_n28695_,
    new_n28696_, new_n28697_, new_n28698_, new_n28699_, new_n28700_,
    new_n28701_, new_n28702_, new_n28703_, new_n28704_, new_n28705_,
    new_n28706_, new_n28707_, new_n28708_, new_n28709_, new_n28710_,
    new_n28711_, new_n28712_, new_n28713_, new_n28714_, new_n28715_,
    new_n28716_, new_n28717_, new_n28718_, new_n28719_, new_n28720_,
    new_n28721_, new_n28722_, new_n28723_, new_n28724_, new_n28725_,
    new_n28726_, new_n28727_, new_n28728_, new_n28729_, new_n28730_,
    new_n28731_, new_n28732_, new_n28733_, new_n28734_, new_n28735_,
    new_n28736_, new_n28737_, new_n28738_, new_n28739_, new_n28740_,
    new_n28741_, new_n28742_, new_n28743_, new_n28744_, new_n28745_,
    new_n28746_, new_n28747_, new_n28748_, new_n28749_, new_n28750_,
    new_n28751_, new_n28752_, new_n28753_, new_n28754_, new_n28755_,
    new_n28756_, new_n28757_, new_n28758_, new_n28759_, new_n28760_,
    new_n28761_, new_n28762_, new_n28763_, new_n28764_, new_n28765_,
    new_n28766_, new_n28767_, new_n28768_, new_n28769_, new_n28770_,
    new_n28771_, new_n28772_, new_n28773_, new_n28774_, new_n28775_,
    new_n28776_, new_n28777_, new_n28778_, new_n28779_, new_n28780_,
    new_n28781_, new_n28782_, new_n28783_, new_n28784_, new_n28785_,
    new_n28786_, new_n28787_, new_n28788_, new_n28789_, new_n28790_,
    new_n28791_, new_n28792_, new_n28793_, new_n28794_, new_n28795_,
    new_n28796_, new_n28797_, new_n28798_, new_n28799_, new_n28800_,
    new_n28801_, new_n28802_, new_n28803_, new_n28804_, new_n28805_,
    new_n28806_, new_n28807_, new_n28808_, new_n28809_, new_n28810_,
    new_n28811_, new_n28812_, new_n28813_, new_n28814_, new_n28815_,
    new_n28816_, new_n28817_, new_n28818_, new_n28819_, new_n28820_,
    new_n28821_, new_n28822_, new_n28823_, new_n28824_, new_n28825_,
    new_n28826_, new_n28827_, new_n28828_, new_n28829_, new_n28830_,
    new_n28831_, new_n28832_, new_n28833_, new_n28834_, new_n28835_,
    new_n28836_, new_n28837_, new_n28838_, new_n28839_, new_n28840_,
    new_n28841_, new_n28842_, new_n28843_, new_n28844_, new_n28845_,
    new_n28846_, new_n28847_, new_n28848_, new_n28849_, new_n28850_,
    new_n28851_, new_n28852_, new_n28853_, new_n28854_, new_n28855_,
    new_n28856_, new_n28857_, new_n28858_, new_n28859_, new_n28860_,
    new_n28861_, new_n28862_, new_n28863_, new_n28864_, new_n28865_,
    new_n28866_, new_n28867_, new_n28868_, new_n28869_, new_n28870_,
    new_n28871_, new_n28872_, new_n28873_, new_n28874_, new_n28875_,
    new_n28876_, new_n28877_, new_n28878_, new_n28879_, new_n28880_,
    new_n28881_, new_n28882_, new_n28883_, new_n28884_, new_n28885_,
    new_n28886_, new_n28887_, new_n28888_, new_n28889_, new_n28890_,
    new_n28891_, new_n28892_, new_n28893_, new_n28894_, new_n28895_,
    new_n28896_, new_n28897_, new_n28898_, new_n28899_, new_n28900_,
    new_n28901_, new_n28902_, new_n28903_, new_n28904_, new_n28905_,
    new_n28906_, new_n28907_, new_n28908_, new_n28909_, new_n28910_,
    new_n28911_, new_n28912_, new_n28913_, new_n28914_, new_n28915_,
    new_n28916_, new_n28917_, new_n28918_, new_n28919_, new_n28920_,
    new_n28921_, new_n28922_, new_n28923_, new_n28924_, new_n28925_,
    new_n28926_, new_n28927_, new_n28928_, new_n28929_, new_n28930_,
    new_n28931_, new_n28932_, new_n28933_, new_n28934_, new_n28935_,
    new_n28936_, new_n28937_, new_n28938_, new_n28939_, new_n28940_,
    new_n28941_, new_n28942_, new_n28943_, new_n28944_, new_n28945_,
    new_n28946_, new_n28947_, new_n28948_, new_n28949_, new_n28950_,
    new_n28951_, new_n28952_, new_n28953_, new_n28954_, new_n28955_,
    new_n28956_, new_n28957_, new_n28958_, new_n28959_, new_n28960_,
    new_n28961_, new_n28962_, new_n28963_, new_n28964_, new_n28965_,
    new_n28966_, new_n28967_, new_n28968_, new_n28969_, new_n28970_,
    new_n28971_, new_n28972_, new_n28973_, new_n28974_, new_n28975_,
    new_n28976_, new_n28977_, new_n28978_, new_n28979_, new_n28980_,
    new_n28981_, new_n28982_, new_n28983_, new_n28984_, new_n28985_,
    new_n28986_, new_n28987_, new_n28988_, new_n28989_, new_n28990_,
    new_n28991_, new_n28992_, new_n28993_, new_n28994_, new_n28995_,
    new_n28996_, new_n28997_, new_n28998_, new_n28999_, new_n29000_,
    new_n29001_, new_n29002_, new_n29003_, new_n29004_, new_n29005_,
    new_n29006_, new_n29007_, new_n29008_, new_n29009_, new_n29010_,
    new_n29011_, new_n29012_, new_n29013_, new_n29014_, new_n29015_,
    new_n29016_, new_n29017_, new_n29018_, new_n29019_, new_n29020_,
    new_n29021_, new_n29022_, new_n29023_, new_n29024_, new_n29025_,
    new_n29026_, new_n29027_, new_n29028_, new_n29029_, new_n29030_,
    new_n29031_, new_n29032_, new_n29033_, new_n29034_, new_n29035_,
    new_n29036_, new_n29037_, new_n29038_, new_n29039_, new_n29040_,
    new_n29041_, new_n29042_, new_n29043_, new_n29044_, new_n29045_,
    new_n29046_, new_n29047_, new_n29048_, new_n29049_, new_n29050_,
    new_n29051_, new_n29052_, new_n29053_, new_n29054_, new_n29055_,
    new_n29056_, new_n29057_, new_n29058_, new_n29059_, new_n29060_,
    new_n29061_, new_n29062_, new_n29063_, new_n29064_, new_n29065_,
    new_n29066_, new_n29067_, new_n29068_, new_n29069_, new_n29070_,
    new_n29071_, new_n29072_, new_n29073_, new_n29074_, new_n29075_,
    new_n29076_, new_n29077_, new_n29078_, new_n29079_, new_n29080_,
    new_n29081_, new_n29082_, new_n29083_, new_n29084_, new_n29085_,
    new_n29086_, new_n29087_, new_n29088_, new_n29089_, new_n29090_,
    new_n29091_, new_n29092_, new_n29093_, new_n29094_, new_n29095_,
    new_n29096_, new_n29097_, new_n29098_, new_n29099_, new_n29100_,
    new_n29101_, new_n29102_, new_n29103_, new_n29104_, new_n29105_,
    new_n29106_, new_n29107_, new_n29108_, new_n29109_, new_n29110_,
    new_n29111_, new_n29112_, new_n29113_, new_n29114_, new_n29115_,
    new_n29116_, new_n29117_, new_n29118_, new_n29119_, new_n29120_,
    new_n29121_, new_n29122_, new_n29123_, new_n29124_, new_n29125_,
    new_n29126_, new_n29127_, new_n29128_, new_n29129_, new_n29130_,
    new_n29131_, new_n29132_, new_n29133_, new_n29134_, new_n29135_,
    new_n29136_, new_n29137_, new_n29138_, new_n29139_, new_n29140_,
    new_n29141_, new_n29142_, new_n29143_, new_n29144_, new_n29145_,
    new_n29146_, new_n29147_, new_n29148_, new_n29149_, new_n29150_,
    new_n29151_, new_n29152_, new_n29153_, new_n29154_, new_n29155_,
    new_n29156_, new_n29157_, new_n29158_, new_n29159_, new_n29160_,
    new_n29161_, new_n29162_, new_n29163_, new_n29164_, new_n29165_,
    new_n29166_, new_n29167_, new_n29168_, new_n29169_, new_n29170_,
    new_n29171_, new_n29172_, new_n29173_, new_n29174_, new_n29175_,
    new_n29176_, new_n29177_, new_n29178_, new_n29179_, new_n29180_,
    new_n29181_, new_n29182_, new_n29183_, new_n29184_, new_n29185_,
    new_n29186_, new_n29187_, new_n29188_, new_n29189_, new_n29190_,
    new_n29191_, new_n29192_, new_n29193_, new_n29194_, new_n29195_,
    new_n29196_, new_n29197_, new_n29198_, new_n29199_, new_n29200_,
    new_n29201_, new_n29202_, new_n29203_, new_n29204_, new_n29205_,
    new_n29206_, new_n29207_, new_n29208_, new_n29209_, new_n29210_,
    new_n29211_, new_n29212_, new_n29213_, new_n29214_, new_n29215_,
    new_n29216_, new_n29217_, new_n29218_, new_n29219_, new_n29220_,
    new_n29221_, new_n29222_, new_n29223_, new_n29224_, new_n29225_,
    new_n29226_, new_n29227_, new_n29228_, new_n29229_, new_n29230_,
    new_n29231_, new_n29232_, new_n29233_, new_n29234_, new_n29235_,
    new_n29236_, new_n29237_, new_n29238_, new_n29239_, new_n29240_,
    new_n29241_, new_n29242_, new_n29243_, new_n29244_, new_n29245_,
    new_n29246_, new_n29247_, new_n29248_, new_n29249_, new_n29250_,
    new_n29251_, new_n29252_, new_n29253_, new_n29254_, new_n29255_,
    new_n29256_, new_n29257_, new_n29258_, new_n29259_, new_n29260_,
    new_n29261_, new_n29262_, new_n29263_, new_n29264_, new_n29265_,
    new_n29266_, new_n29267_, new_n29268_, new_n29269_, new_n29270_,
    new_n29271_, new_n29272_, new_n29273_, new_n29274_, new_n29275_,
    new_n29276_, new_n29277_, new_n29278_, new_n29279_, new_n29280_,
    new_n29281_, new_n29282_, new_n29283_, new_n29284_, new_n29285_,
    new_n29286_, new_n29287_, new_n29288_, new_n29289_, new_n29290_,
    new_n29291_, new_n29292_, new_n29293_, new_n29294_, new_n29295_,
    new_n29296_, new_n29297_, new_n29298_, new_n29299_, new_n29300_,
    new_n29301_, new_n29302_, new_n29303_, new_n29304_, new_n29305_,
    new_n29306_, new_n29307_, new_n29308_, new_n29309_, new_n29310_,
    new_n29311_, new_n29312_, new_n29313_, new_n29314_, new_n29315_,
    new_n29316_, new_n29317_, new_n29318_, new_n29319_, new_n29320_,
    new_n29321_, new_n29322_, new_n29323_, new_n29324_, new_n29325_,
    new_n29326_, new_n29327_, new_n29328_, new_n29329_, new_n29330_,
    new_n29331_, new_n29332_, new_n29333_, new_n29334_, new_n29335_,
    new_n29336_, new_n29337_, new_n29338_, new_n29339_, new_n29340_,
    new_n29341_, new_n29342_, new_n29343_, new_n29344_, new_n29345_,
    new_n29346_, new_n29347_, new_n29348_, new_n29349_, new_n29350_,
    new_n29351_, new_n29352_, new_n29353_, new_n29354_, new_n29355_,
    new_n29356_, new_n29357_, new_n29358_, new_n29359_, new_n29360_,
    new_n29361_, new_n29362_, new_n29363_, new_n29364_, new_n29365_,
    new_n29366_, new_n29367_, new_n29368_, new_n29369_, new_n29370_,
    new_n29371_, new_n29372_, new_n29373_, new_n29374_, new_n29375_,
    new_n29376_, new_n29377_, new_n29378_, new_n29379_, new_n29380_,
    new_n29381_, new_n29382_, new_n29383_, new_n29384_, new_n29385_,
    new_n29386_, new_n29387_, new_n29388_, new_n29389_, new_n29390_,
    new_n29391_, new_n29392_, new_n29393_, new_n29394_, new_n29395_,
    new_n29396_, new_n29397_, new_n29398_, new_n29399_, new_n29400_,
    new_n29401_, new_n29402_, new_n29403_, new_n29404_, new_n29405_,
    new_n29406_, new_n29407_, new_n29408_, new_n29409_, new_n29410_,
    new_n29411_, new_n29412_, new_n29413_, new_n29414_, new_n29415_,
    new_n29416_, new_n29417_, new_n29418_, new_n29419_, new_n29420_,
    new_n29421_, new_n29422_, new_n29423_, new_n29424_, new_n29425_,
    new_n29426_, new_n29427_, new_n29428_, new_n29429_, new_n29430_,
    new_n29431_, new_n29432_, new_n29433_, new_n29434_, new_n29435_,
    new_n29436_, new_n29437_, new_n29438_, new_n29439_, new_n29440_,
    new_n29441_, new_n29442_, new_n29443_, new_n29444_, new_n29445_,
    new_n29446_, new_n29447_, new_n29448_, new_n29449_, new_n29450_,
    new_n29451_, new_n29452_, new_n29453_, new_n29454_, new_n29455_,
    new_n29456_, new_n29457_, new_n29458_, new_n29459_, new_n29460_,
    new_n29461_, new_n29462_, new_n29463_, new_n29464_, new_n29465_,
    new_n29466_, new_n29467_, new_n29468_, new_n29469_, new_n29470_,
    new_n29471_, new_n29472_, new_n29473_, new_n29474_, new_n29475_,
    new_n29476_, new_n29477_, new_n29478_, new_n29479_, new_n29480_,
    new_n29481_, new_n29482_, new_n29483_, new_n29484_, new_n29485_,
    new_n29486_, new_n29487_, new_n29488_, new_n29489_, new_n29490_,
    new_n29491_, new_n29492_, new_n29493_, new_n29494_, new_n29495_,
    new_n29496_, new_n29497_, new_n29498_, new_n29499_, new_n29500_,
    new_n29501_, new_n29502_, new_n29503_, new_n29504_, new_n29505_,
    new_n29506_, new_n29507_, new_n29508_, new_n29509_, new_n29510_,
    new_n29511_, new_n29512_, new_n29513_, new_n29514_, new_n29515_,
    new_n29516_, new_n29517_, new_n29518_, new_n29519_, new_n29520_,
    new_n29521_, new_n29522_, new_n29523_, new_n29524_, new_n29525_,
    new_n29526_, new_n29527_, new_n29528_, new_n29529_, new_n29530_,
    new_n29531_, new_n29532_, new_n29533_, new_n29534_, new_n29535_,
    new_n29536_, new_n29537_, new_n29538_, new_n29539_, new_n29540_,
    new_n29541_, new_n29542_, new_n29543_, new_n29544_, new_n29545_,
    new_n29546_, new_n29547_, new_n29548_, new_n29549_, new_n29550_,
    new_n29551_, new_n29552_, new_n29553_, new_n29554_, new_n29555_,
    new_n29556_, new_n29557_, new_n29558_, new_n29559_, new_n29560_,
    new_n29561_, new_n29562_, new_n29563_, new_n29564_, new_n29565_,
    new_n29566_, new_n29567_, new_n29568_, new_n29569_, new_n29570_,
    new_n29571_, new_n29572_, new_n29573_, new_n29574_, new_n29575_,
    new_n29576_, new_n29577_, new_n29578_, new_n29579_, new_n29580_,
    new_n29581_, new_n29582_, new_n29583_, new_n29584_, new_n29585_,
    new_n29586_, new_n29587_, new_n29588_, new_n29589_, new_n29590_,
    new_n29591_, new_n29592_, new_n29593_, new_n29594_, new_n29595_,
    new_n29596_, new_n29597_, new_n29598_, new_n29599_, new_n29600_,
    new_n29601_, new_n29602_, new_n29603_, new_n29604_, new_n29605_,
    new_n29606_, new_n29607_, new_n29608_, new_n29609_, new_n29610_,
    new_n29611_, new_n29612_, new_n29613_, new_n29614_, new_n29615_,
    new_n29616_, new_n29617_, new_n29618_, new_n29619_, new_n29620_,
    new_n29621_, new_n29622_, new_n29623_, new_n29624_, new_n29625_,
    new_n29626_, new_n29627_, new_n29628_, new_n29629_, new_n29630_,
    new_n29631_, new_n29632_, new_n29633_, new_n29634_, new_n29635_,
    new_n29636_, new_n29637_, new_n29638_, new_n29639_, new_n29640_,
    new_n29641_, new_n29642_, new_n29643_, new_n29644_, new_n29645_,
    new_n29646_, new_n29647_, new_n29648_, new_n29649_, new_n29650_,
    new_n29651_, new_n29652_, new_n29653_, new_n29654_, new_n29655_,
    new_n29656_, new_n29657_, new_n29658_, new_n29659_, new_n29660_,
    new_n29661_, new_n29662_, new_n29663_, new_n29664_, new_n29665_,
    new_n29666_, new_n29667_, new_n29668_, new_n29669_, new_n29670_,
    new_n29671_, new_n29672_, new_n29673_, new_n29674_, new_n29675_,
    new_n29676_, new_n29677_, new_n29678_, new_n29679_, new_n29680_,
    new_n29681_, new_n29682_, new_n29683_, new_n29684_, new_n29685_,
    new_n29686_, new_n29687_, new_n29688_, new_n29689_, new_n29690_,
    new_n29691_, new_n29692_, new_n29693_, new_n29694_, new_n29695_,
    new_n29696_, new_n29697_, new_n29698_, new_n29699_, new_n29700_,
    new_n29701_, new_n29702_, new_n29703_, new_n29704_, new_n29705_,
    new_n29706_, new_n29707_, new_n29708_, new_n29709_, new_n29710_,
    new_n29711_, new_n29712_, new_n29713_, new_n29714_, new_n29715_,
    new_n29716_, new_n29717_, new_n29718_, new_n29719_, new_n29720_,
    new_n29721_, new_n29722_, new_n29723_, new_n29724_, new_n29725_,
    new_n29726_, new_n29727_, new_n29728_, new_n29729_, new_n29730_,
    new_n29731_, new_n29732_, new_n29733_, new_n29734_, new_n29735_,
    new_n29736_, new_n29737_, new_n29738_, new_n29739_, new_n29740_,
    new_n29741_, new_n29742_, new_n29743_, new_n29744_, new_n29745_,
    new_n29746_, new_n29747_, new_n29748_, new_n29749_, new_n29750_,
    new_n29751_, new_n29752_, new_n29753_, new_n29754_, new_n29755_,
    new_n29756_, new_n29757_, new_n29758_, new_n29759_, new_n29760_,
    new_n29761_, new_n29762_, new_n29763_, new_n29764_, new_n29765_,
    new_n29766_, new_n29767_, new_n29768_, new_n29769_, new_n29770_,
    new_n29771_, new_n29772_, new_n29773_, new_n29774_, new_n29775_,
    new_n29776_, new_n29777_, new_n29778_, new_n29779_, new_n29780_,
    new_n29781_, new_n29782_, new_n29783_, new_n29784_, new_n29785_,
    new_n29786_, new_n29787_, new_n29788_, new_n29789_, new_n29790_,
    new_n29791_, new_n29792_, new_n29793_, new_n29794_, new_n29795_,
    new_n29796_, new_n29797_, new_n29798_, new_n29799_, new_n29800_,
    new_n29801_, new_n29802_, new_n29803_, new_n29804_, new_n29805_,
    new_n29806_, new_n29807_, new_n29808_, new_n29809_, new_n29810_,
    new_n29811_, new_n29812_, new_n29813_, new_n29814_, new_n29815_,
    new_n29816_, new_n29817_, new_n29818_, new_n29819_, new_n29820_,
    new_n29821_, new_n29822_, new_n29823_, new_n29824_, new_n29825_,
    new_n29826_, new_n29827_, new_n29828_, new_n29829_, new_n29830_,
    new_n29831_, new_n29832_, new_n29833_, new_n29834_, new_n29835_,
    new_n29836_, new_n29837_, new_n29838_, new_n29839_, new_n29840_,
    new_n29841_, new_n29842_, new_n29843_, new_n29844_, new_n29845_,
    new_n29846_, new_n29847_, new_n29848_, new_n29849_, new_n29850_,
    new_n29851_, new_n29852_, new_n29853_, new_n29854_, new_n29855_,
    new_n29856_, new_n29857_, new_n29858_, new_n29859_, new_n29860_,
    new_n29861_, new_n29862_, new_n29863_, new_n29864_, new_n29865_,
    new_n29866_, new_n29867_, new_n29868_, new_n29869_, new_n29870_,
    new_n29871_, new_n29872_, new_n29873_, new_n29874_, new_n29875_,
    new_n29876_, new_n29877_, new_n29878_, new_n29879_, new_n29880_,
    new_n29881_, new_n29882_, new_n29883_, new_n29884_, new_n29885_,
    new_n29886_, new_n29887_, new_n29888_, new_n29889_, new_n29890_,
    new_n29891_, new_n29892_, new_n29893_, new_n29894_, new_n29895_,
    new_n29896_, new_n29897_, new_n29898_, new_n29899_, new_n29900_,
    new_n29901_, new_n29902_, new_n29903_, new_n29904_, new_n29905_,
    new_n29906_, new_n29907_, new_n29908_, new_n29909_, new_n29910_,
    new_n29911_, new_n29912_, new_n29913_, new_n29914_, new_n29915_,
    new_n29916_, new_n29917_, new_n29918_, new_n29919_, new_n29920_,
    new_n29921_, new_n29922_, new_n29923_, new_n29924_, new_n29925_,
    new_n29926_, new_n29927_, new_n29928_, new_n29929_, new_n29930_,
    new_n29931_, new_n29932_, new_n29933_, new_n29934_, new_n29935_,
    new_n29936_, new_n29937_, new_n29938_, new_n29939_, new_n29940_,
    new_n29941_, new_n29942_, new_n29943_, new_n29944_, new_n29945_,
    new_n29946_, new_n29947_, new_n29948_, new_n29949_, new_n29950_,
    new_n29951_, new_n29952_, new_n29953_, new_n29954_, new_n29955_,
    new_n29956_, new_n29957_, new_n29958_, new_n29959_, new_n29960_,
    new_n29961_, new_n29962_, new_n29963_, new_n29964_, new_n29965_,
    new_n29966_, new_n29967_, new_n29968_, new_n29969_, new_n29970_,
    new_n29971_, new_n29972_, new_n29973_, new_n29974_, new_n29975_,
    new_n29976_, new_n29977_, new_n29978_, new_n29979_, new_n29980_,
    new_n29981_, new_n29982_, new_n29983_, new_n29984_, new_n29985_,
    new_n29986_, new_n29987_, new_n29988_, new_n29989_, new_n29990_,
    new_n29991_, new_n29992_, new_n29993_, new_n29994_, new_n29995_,
    new_n29996_, new_n29997_, new_n29998_, new_n29999_, new_n30000_,
    new_n30001_, new_n30002_, new_n30003_, new_n30004_, new_n30005_,
    new_n30006_, new_n30007_, new_n30008_, new_n30009_, new_n30010_,
    new_n30011_, new_n30012_, new_n30013_, new_n30014_, new_n30015_,
    new_n30016_, new_n30017_, new_n30018_, new_n30019_, new_n30020_,
    new_n30021_, new_n30022_, new_n30023_, new_n30024_, new_n30025_,
    new_n30026_, new_n30027_, new_n30028_, new_n30029_, new_n30030_,
    new_n30031_, new_n30032_, new_n30033_, new_n30034_, new_n30035_,
    new_n30036_, new_n30037_, new_n30038_, new_n30039_, new_n30040_,
    new_n30041_, new_n30042_, new_n30043_, new_n30044_, new_n30045_,
    new_n30046_, new_n30047_, new_n30048_, new_n30049_, new_n30050_,
    new_n30051_, new_n30052_, new_n30053_, new_n30054_, new_n30055_,
    new_n30056_, new_n30057_, new_n30058_, new_n30059_, new_n30060_,
    new_n30061_, new_n30062_, new_n30063_, new_n30064_, new_n30065_,
    new_n30066_, new_n30067_, new_n30068_, new_n30069_, new_n30070_,
    new_n30071_, new_n30072_, new_n30073_, new_n30074_, new_n30075_,
    new_n30076_, new_n30077_, new_n30078_, new_n30079_, new_n30080_,
    new_n30081_, new_n30082_, new_n30083_, new_n30084_, new_n30085_,
    new_n30086_, new_n30087_, new_n30088_, new_n30089_, new_n30090_,
    new_n30091_, new_n30092_, new_n30093_, new_n30094_, new_n30095_,
    new_n30096_, new_n30097_, new_n30098_, new_n30099_, new_n30100_,
    new_n30101_, new_n30102_, new_n30103_, new_n30104_, new_n30105_,
    new_n30106_, new_n30107_, new_n30108_, new_n30109_, new_n30110_,
    new_n30111_, new_n30112_, new_n30113_, new_n30114_, new_n30115_,
    new_n30116_, new_n30117_, new_n30118_, new_n30119_, new_n30120_,
    new_n30121_, new_n30122_, new_n30123_, new_n30124_, new_n30125_,
    new_n30126_, new_n30127_, new_n30128_, new_n30129_, new_n30130_,
    new_n30131_, new_n30132_, new_n30133_, new_n30134_, new_n30135_,
    new_n30136_, new_n30137_, new_n30138_, new_n30139_, new_n30140_,
    new_n30141_, new_n30142_, new_n30143_, new_n30144_, new_n30145_,
    new_n30146_, new_n30147_, new_n30148_, new_n30149_, new_n30150_,
    new_n30151_, new_n30152_, new_n30153_, new_n30154_, new_n30155_,
    new_n30156_, new_n30157_, new_n30158_, new_n30159_, new_n30160_,
    new_n30161_, new_n30162_, new_n30163_, new_n30164_, new_n30165_,
    new_n30166_, new_n30167_, new_n30168_, new_n30169_, new_n30170_,
    new_n30171_, new_n30172_, new_n30173_, new_n30174_, new_n30175_,
    new_n30176_, new_n30177_, new_n30178_, new_n30179_, new_n30180_,
    new_n30181_, new_n30182_, new_n30183_, new_n30184_, new_n30185_,
    new_n30186_, new_n30187_, new_n30188_, new_n30189_, new_n30190_,
    new_n30191_, new_n30192_, new_n30193_, new_n30194_, new_n30195_,
    new_n30196_, new_n30197_, new_n30198_, new_n30199_, new_n30200_,
    new_n30201_, new_n30202_, new_n30203_, new_n30204_, new_n30205_,
    new_n30206_, new_n30207_, new_n30208_, new_n30209_, new_n30210_,
    new_n30211_, new_n30212_, new_n30213_, new_n30214_, new_n30215_,
    new_n30216_, new_n30217_, new_n30218_, new_n30219_, new_n30220_,
    new_n30221_, new_n30222_, new_n30223_, new_n30224_, new_n30225_,
    new_n30226_, new_n30227_, new_n30228_, new_n30229_, new_n30230_,
    new_n30231_, new_n30232_, new_n30233_, new_n30234_, new_n30235_,
    new_n30236_, new_n30237_, new_n30238_, new_n30239_, new_n30240_,
    new_n30241_, new_n30242_, new_n30243_, new_n30244_, new_n30245_,
    new_n30246_, new_n30247_, new_n30248_, new_n30249_, new_n30250_,
    new_n30251_, new_n30252_, new_n30253_, new_n30254_, new_n30255_,
    new_n30256_, new_n30257_, new_n30258_, new_n30259_, new_n30260_,
    new_n30261_, new_n30262_, new_n30263_, new_n30264_, new_n30265_,
    new_n30266_, new_n30267_, new_n30268_, new_n30269_, new_n30270_,
    new_n30271_, new_n30272_, new_n30273_, new_n30274_, new_n30275_,
    new_n30276_, new_n30277_, new_n30278_, new_n30279_, new_n30280_,
    new_n30281_, new_n30282_, new_n30283_, new_n30284_, new_n30285_,
    new_n30286_, new_n30287_, new_n30288_, new_n30289_, new_n30290_,
    new_n30291_, new_n30292_, new_n30293_, new_n30294_, new_n30295_,
    new_n30296_, new_n30297_, new_n30298_, new_n30299_, new_n30300_,
    new_n30301_, new_n30302_, new_n30303_, new_n30304_, new_n30305_,
    new_n30306_, new_n30307_, new_n30308_, new_n30309_, new_n30310_,
    new_n30311_, new_n30312_, new_n30313_, new_n30314_, new_n30315_,
    new_n30316_, new_n30317_, new_n30318_, new_n30319_, new_n30320_,
    new_n30321_, new_n30322_, new_n30323_, new_n30324_, new_n30325_,
    new_n30326_, new_n30327_, new_n30328_, new_n30329_, new_n30330_,
    new_n30331_, new_n30332_, new_n30333_, new_n30334_, new_n30335_,
    new_n30336_, new_n30337_, new_n30338_, new_n30339_, new_n30340_,
    new_n30341_, new_n30342_, new_n30343_, new_n30344_, new_n30345_,
    new_n30346_, new_n30347_, new_n30348_, new_n30349_, new_n30350_,
    new_n30351_, new_n30352_, new_n30353_, new_n30354_, new_n30355_,
    new_n30356_, new_n30357_, new_n30358_, new_n30359_, new_n30360_,
    new_n30361_, new_n30362_, new_n30363_, new_n30364_, new_n30365_,
    new_n30366_, new_n30367_, new_n30368_, new_n30369_, new_n30370_,
    new_n30371_, new_n30372_, new_n30373_, new_n30374_, new_n30375_,
    new_n30376_, new_n30377_, new_n30378_, new_n30379_, new_n30380_,
    new_n30381_, new_n30382_, new_n30383_, new_n30384_, new_n30385_,
    new_n30386_, new_n30387_, new_n30388_, new_n30389_, new_n30390_,
    new_n30391_, new_n30392_, new_n30393_, new_n30394_, new_n30395_,
    new_n30396_, new_n30397_, new_n30398_, new_n30399_, new_n30400_,
    new_n30401_, new_n30402_, new_n30403_, new_n30404_, new_n30405_,
    new_n30406_, new_n30407_, new_n30408_, new_n30409_, new_n30410_,
    new_n30411_, new_n30412_, new_n30413_, new_n30414_, new_n30415_,
    new_n30416_, new_n30417_, new_n30418_, new_n30419_, new_n30420_,
    new_n30421_, new_n30422_, new_n30423_, new_n30424_, new_n30425_,
    new_n30426_, new_n30427_, new_n30428_, new_n30429_, new_n30430_,
    new_n30431_, new_n30432_, new_n30433_, new_n30434_, new_n30435_,
    new_n30436_, new_n30437_, new_n30438_, new_n30439_, new_n30440_,
    new_n30441_, new_n30442_, new_n30443_, new_n30444_, new_n30445_,
    new_n30446_, new_n30447_, new_n30448_, new_n30449_, new_n30450_,
    new_n30451_, new_n30452_, new_n30453_, new_n30454_, new_n30455_,
    new_n30456_, new_n30457_, new_n30458_, new_n30459_, new_n30460_,
    new_n30461_, new_n30462_, new_n30463_, new_n30464_, new_n30465_,
    new_n30466_, new_n30467_, new_n30468_, new_n30469_, new_n30470_,
    new_n30471_, new_n30472_, new_n30473_, new_n30474_, new_n30475_,
    new_n30476_, new_n30477_, new_n30478_, new_n30479_, new_n30480_,
    new_n30481_, new_n30482_, new_n30483_, new_n30484_, new_n30485_,
    new_n30486_, new_n30487_, new_n30488_, new_n30489_, new_n30490_,
    new_n30491_, new_n30492_, new_n30493_, new_n30494_, new_n30495_,
    new_n30496_, new_n30497_, new_n30498_, new_n30499_, new_n30500_,
    new_n30501_, new_n30502_, new_n30503_, new_n30504_, new_n30505_,
    new_n30506_, new_n30507_, new_n30508_, new_n30509_, new_n30510_,
    new_n30511_, new_n30512_, new_n30513_, new_n30514_, new_n30515_,
    new_n30516_, new_n30517_, new_n30518_, new_n30519_, new_n30520_,
    new_n30521_, new_n30522_, new_n30523_, new_n30524_, new_n30525_,
    new_n30526_, new_n30527_, new_n30528_, new_n30529_, new_n30530_,
    new_n30531_, new_n30532_, new_n30533_, new_n30534_, new_n30535_,
    new_n30536_, new_n30537_, new_n30538_, new_n30539_, new_n30540_,
    new_n30541_, new_n30542_, new_n30543_, new_n30544_, new_n30545_,
    new_n30546_, new_n30547_, new_n30548_, new_n30549_, new_n30550_,
    new_n30551_, new_n30552_, new_n30553_, new_n30554_, new_n30555_,
    new_n30556_, new_n30557_, new_n30558_, new_n30559_, new_n30560_,
    new_n30561_, new_n30562_, new_n30563_, new_n30564_, new_n30565_,
    new_n30566_, new_n30567_, new_n30568_, new_n30569_, new_n30570_,
    new_n30571_, new_n30572_, new_n30573_, new_n30574_, new_n30575_,
    new_n30576_, new_n30577_, new_n30578_, new_n30579_, new_n30580_,
    new_n30581_, new_n30582_, new_n30583_, new_n30584_, new_n30585_,
    new_n30586_, new_n30587_, new_n30588_, new_n30589_, new_n30590_,
    new_n30591_, new_n30592_, new_n30593_, new_n30594_, new_n30595_,
    new_n30596_, new_n30597_, new_n30598_, new_n30599_, new_n30600_,
    new_n30601_, new_n30602_, new_n30603_, new_n30604_, new_n30605_,
    new_n30606_, new_n30607_, new_n30608_, new_n30609_, new_n30610_,
    new_n30611_, new_n30612_, new_n30613_, new_n30614_, new_n30615_,
    new_n30616_, new_n30617_, new_n30618_, new_n30619_, new_n30620_,
    new_n30621_, new_n30622_, new_n30623_, new_n30624_, new_n30625_,
    new_n30626_, new_n30627_, new_n30628_, new_n30629_, new_n30630_,
    new_n30631_, new_n30632_, new_n30633_, new_n30634_, new_n30635_,
    new_n30636_, new_n30637_, new_n30638_, new_n30639_, new_n30640_,
    new_n30641_, new_n30642_, new_n30643_, new_n30644_, new_n30645_,
    new_n30646_, new_n30647_, new_n30648_, new_n30649_, new_n30650_,
    new_n30651_, new_n30652_, new_n30653_, new_n30654_, new_n30655_,
    new_n30656_, new_n30657_, new_n30658_, new_n30659_, new_n30660_,
    new_n30661_, new_n30662_, new_n30663_, new_n30664_, new_n30665_,
    new_n30666_, new_n30667_, new_n30668_, new_n30669_, new_n30670_,
    new_n30671_, new_n30672_, new_n30673_, new_n30674_, new_n30675_,
    new_n30676_, new_n30677_, new_n30678_, new_n30679_, new_n30680_,
    new_n30681_, new_n30682_, new_n30683_, new_n30684_, new_n30685_,
    new_n30686_, new_n30687_, new_n30688_, new_n30689_, new_n30690_,
    new_n30691_, new_n30692_, new_n30693_, new_n30694_, new_n30695_,
    new_n30696_, new_n30697_, new_n30698_, new_n30699_, new_n30700_,
    new_n30701_, new_n30702_, new_n30703_, new_n30704_, new_n30705_,
    new_n30706_, new_n30707_, new_n30708_, new_n30709_, new_n30710_,
    new_n30711_, new_n30712_, new_n30713_, new_n30714_, new_n30715_,
    new_n30716_, new_n30717_, new_n30718_, new_n30719_, new_n30720_,
    new_n30721_, new_n30722_, new_n30723_, new_n30724_, new_n30725_,
    new_n30726_, new_n30727_, new_n30728_, new_n30729_, new_n30730_,
    new_n30731_, new_n30732_, new_n30733_, new_n30734_, new_n30735_,
    new_n30736_, new_n30737_, new_n30738_, new_n30739_, new_n30740_,
    new_n30741_, new_n30742_, new_n30743_, new_n30744_, new_n30745_,
    new_n30746_, new_n30747_, new_n30748_, new_n30749_, new_n30750_,
    new_n30751_, new_n30752_, new_n30753_, new_n30754_, new_n30755_,
    new_n30756_, new_n30757_, new_n30758_, new_n30759_, new_n30760_,
    new_n30761_, new_n30762_, new_n30763_, new_n30764_, new_n30765_,
    new_n30766_, new_n30767_, new_n30768_, new_n30769_, new_n30770_,
    new_n30771_, new_n30772_, new_n30773_, new_n30774_, new_n30775_,
    new_n30776_, new_n30777_, new_n30778_, new_n30779_, new_n30780_,
    new_n30781_, new_n30782_, new_n30783_, new_n30784_, new_n30785_,
    new_n30786_, new_n30787_, new_n30788_, new_n30789_, new_n30790_,
    new_n30791_, new_n30792_, new_n30793_, new_n30794_, new_n30795_,
    new_n30796_, new_n30797_, new_n30798_, new_n30799_, new_n30800_,
    new_n30801_, new_n30802_, new_n30803_, new_n30804_, new_n30805_,
    new_n30806_, new_n30807_, new_n30808_, new_n30809_, new_n30810_,
    new_n30811_, new_n30812_, new_n30813_, new_n30814_, new_n30815_,
    new_n30816_, new_n30817_, new_n30818_, new_n30819_, new_n30820_,
    new_n30821_, new_n30822_, new_n30823_, new_n30824_, new_n30825_,
    new_n30826_, new_n30827_, new_n30828_, new_n30829_, new_n30830_,
    new_n30831_, new_n30832_, new_n30833_, new_n30834_, new_n30835_,
    new_n30836_, new_n30837_, new_n30838_, new_n30839_, new_n30840_,
    new_n30841_, new_n30842_, new_n30843_, new_n30844_, new_n30845_,
    new_n30846_, new_n30847_, new_n30848_, new_n30849_, new_n30850_,
    new_n30851_, new_n30852_, new_n30853_, new_n30854_, new_n30855_,
    new_n30856_, new_n30857_, new_n30858_, new_n30859_, new_n30860_,
    new_n30861_, new_n30862_, new_n30863_, new_n30864_, new_n30865_,
    new_n30866_, new_n30867_, new_n30868_, new_n30869_, new_n30870_,
    new_n30871_, new_n30872_, new_n30873_, new_n30874_, new_n30875_,
    new_n30876_, new_n30877_, new_n30878_, new_n30879_, new_n30880_,
    new_n30881_, new_n30882_, new_n30883_, new_n30884_, new_n30885_,
    new_n30886_, new_n30887_, new_n30888_, new_n30889_, new_n30890_,
    new_n30891_, new_n30892_, new_n30893_, new_n30894_, new_n30895_,
    new_n30896_, new_n30897_, new_n30898_, new_n30899_, new_n30900_,
    new_n30901_, new_n30902_, new_n30903_, new_n30904_, new_n30905_,
    new_n30906_, new_n30907_, new_n30908_, new_n30909_, new_n30910_,
    new_n30911_, new_n30912_, new_n30913_, new_n30914_, new_n30915_,
    new_n30916_, new_n30917_, new_n30918_, new_n30919_, new_n30920_,
    new_n30921_, new_n30922_, new_n30923_, new_n30924_, new_n30925_,
    new_n30926_, new_n30927_, new_n30928_, new_n30929_, new_n30930_,
    new_n30931_, new_n30932_, new_n30933_, new_n30934_, new_n30935_,
    new_n30936_, new_n30937_, new_n30938_, new_n30939_, new_n30940_,
    new_n30941_, new_n30942_, new_n30943_, new_n30944_, new_n30945_,
    new_n30946_, new_n30947_, new_n30948_, new_n30949_, new_n30950_,
    new_n30951_, new_n30952_, new_n30953_, new_n30954_, new_n30955_,
    new_n30956_, new_n30957_, new_n30958_, new_n30959_, new_n30960_,
    new_n30961_, new_n30962_, new_n30963_, new_n30964_, new_n30965_,
    new_n30966_, new_n30967_, new_n30968_, new_n30969_, new_n30970_,
    new_n30971_, new_n30972_, new_n30973_, new_n30974_, new_n30975_,
    new_n30976_, new_n30977_, new_n30978_, new_n30979_, new_n30980_,
    new_n30981_, new_n30982_, new_n30983_, new_n30984_, new_n30985_,
    new_n30986_, new_n30987_, new_n30988_, new_n30989_, new_n30990_,
    new_n30991_, new_n30992_, new_n30993_, new_n30994_, new_n30995_,
    new_n30996_, new_n30997_, new_n30998_, new_n30999_, new_n31000_,
    new_n31001_, new_n31002_, new_n31003_, new_n31004_, new_n31005_,
    new_n31006_, new_n31007_, new_n31008_, new_n31009_, new_n31010_,
    new_n31011_, new_n31012_, new_n31013_, new_n31014_, new_n31015_,
    new_n31016_, new_n31017_, new_n31018_, new_n31019_, new_n31020_,
    new_n31021_, new_n31022_, new_n31023_, new_n31024_, new_n31025_,
    new_n31026_, new_n31027_, new_n31028_, new_n31029_, new_n31030_,
    new_n31031_, new_n31032_, new_n31033_, new_n31034_, new_n31035_,
    new_n31036_, new_n31037_, new_n31038_, new_n31039_, new_n31040_,
    new_n31041_, new_n31042_, new_n31043_, new_n31044_, new_n31045_,
    new_n31046_, new_n31047_, new_n31048_, new_n31049_, new_n31050_,
    new_n31051_, new_n31052_, new_n31053_, new_n31054_, new_n31055_,
    new_n31056_, new_n31057_, new_n31058_, new_n31059_, new_n31060_,
    new_n31061_, new_n31062_, new_n31063_, new_n31064_, new_n31065_,
    new_n31066_, new_n31067_, new_n31068_, new_n31069_, new_n31070_,
    new_n31071_, new_n31072_, new_n31073_, new_n31074_, new_n31075_,
    new_n31076_, new_n31077_, new_n31078_, new_n31079_, new_n31080_,
    new_n31081_, new_n31082_, new_n31083_, new_n31084_, new_n31085_,
    new_n31086_, new_n31087_, new_n31088_, new_n31089_, new_n31090_,
    new_n31091_, new_n31092_, new_n31093_, new_n31094_, new_n31095_,
    new_n31096_, new_n31097_, new_n31098_, new_n31099_, new_n31100_,
    new_n31101_, new_n31102_, new_n31103_, new_n31104_, new_n31105_,
    new_n31106_, new_n31107_, new_n31108_, new_n31109_, new_n31110_,
    new_n31111_, new_n31112_, new_n31113_, new_n31114_, new_n31115_,
    new_n31116_, new_n31117_, new_n31118_, new_n31119_, new_n31120_,
    new_n31121_, new_n31122_, new_n31123_, new_n31124_, new_n31125_,
    new_n31126_, new_n31127_, new_n31128_, new_n31129_, new_n31130_,
    new_n31131_, new_n31132_, new_n31133_, new_n31134_, new_n31135_,
    new_n31136_, new_n31137_, new_n31138_, new_n31139_, new_n31140_,
    new_n31141_, new_n31142_, new_n31143_, new_n31144_, new_n31145_,
    new_n31146_, new_n31147_, new_n31148_, new_n31149_, new_n31150_,
    new_n31151_, new_n31152_, new_n31153_, new_n31154_, new_n31155_,
    new_n31156_, new_n31157_, new_n31158_, new_n31159_, new_n31160_,
    new_n31161_, new_n31162_, new_n31163_, new_n31164_, new_n31165_,
    new_n31166_, new_n31167_, new_n31168_, new_n31169_, new_n31170_,
    new_n31171_, new_n31172_, new_n31173_, new_n31174_, new_n31175_,
    new_n31176_, new_n31177_, new_n31178_, new_n31179_, new_n31180_,
    new_n31181_, new_n31182_, new_n31183_, new_n31184_, new_n31185_,
    new_n31186_, new_n31187_, new_n31188_, new_n31189_, new_n31190_,
    new_n31191_, new_n31192_, new_n31193_, new_n31194_, new_n31195_,
    new_n31196_, new_n31197_, new_n31198_, new_n31199_, new_n31200_,
    new_n31201_, new_n31202_, new_n31203_, new_n31204_, new_n31205_,
    new_n31206_, new_n31207_, new_n31208_, new_n31209_, new_n31210_,
    new_n31211_, new_n31212_, new_n31213_, new_n31214_, new_n31215_,
    new_n31216_, new_n31217_, new_n31218_, new_n31219_, new_n31220_,
    new_n31221_, new_n31222_, new_n31223_, new_n31224_, new_n31225_,
    new_n31226_, new_n31227_, new_n31228_, new_n31229_, new_n31230_,
    new_n31231_, new_n31232_, new_n31233_, new_n31234_, new_n31235_,
    new_n31236_, new_n31237_, new_n31238_, new_n31239_, new_n31240_,
    new_n31241_, new_n31242_, new_n31243_, new_n31244_, new_n31245_,
    new_n31246_, new_n31247_, new_n31248_, new_n31249_, new_n31250_,
    new_n31251_, new_n31252_, new_n31253_, new_n31254_, new_n31255_,
    new_n31256_, new_n31257_, new_n31258_, new_n31259_, new_n31260_,
    new_n31261_, new_n31262_, new_n31263_, new_n31264_, new_n31265_,
    new_n31266_, new_n31267_, new_n31268_, new_n31269_, new_n31270_,
    new_n31271_, new_n31272_, new_n31273_, new_n31274_, new_n31275_,
    new_n31276_, new_n31277_, new_n31278_, new_n31279_, new_n31280_,
    new_n31281_, new_n31282_, new_n31283_, new_n31284_, new_n31285_,
    new_n31286_, new_n31287_, new_n31288_, new_n31289_, new_n31290_,
    new_n31291_, new_n31292_, new_n31293_, new_n31294_, new_n31295_,
    new_n31296_, new_n31297_, new_n31298_, new_n31299_, new_n31300_,
    new_n31301_, new_n31302_, new_n31303_, new_n31304_, new_n31305_,
    new_n31306_, new_n31307_, new_n31308_, new_n31309_, new_n31310_,
    new_n31311_, new_n31312_, new_n31313_, new_n31314_, new_n31315_,
    new_n31316_, new_n31317_, new_n31318_, new_n31319_, new_n31320_,
    new_n31321_, new_n31322_, new_n31323_, new_n31324_, new_n31325_,
    new_n31326_, new_n31327_, new_n31328_, new_n31329_, new_n31330_,
    new_n31331_, new_n31332_, new_n31333_, new_n31334_, new_n31335_,
    new_n31336_, new_n31337_, new_n31338_, new_n31339_, new_n31340_,
    new_n31341_, new_n31342_, new_n31343_, new_n31344_, new_n31345_,
    new_n31346_, new_n31347_, new_n31348_, new_n31349_, new_n31350_,
    new_n31351_, new_n31352_, new_n31353_, new_n31354_, new_n31355_,
    new_n31356_, new_n31357_, new_n31358_, new_n31359_, new_n31360_,
    new_n31361_, new_n31362_, new_n31363_, new_n31364_, new_n31365_,
    new_n31366_, new_n31367_, new_n31368_, new_n31369_, new_n31370_,
    new_n31371_, new_n31372_, new_n31373_, new_n31374_, new_n31375_,
    new_n31376_, new_n31377_, new_n31378_, new_n31379_, new_n31380_,
    new_n31381_, new_n31382_, new_n31383_, new_n31384_, new_n31385_,
    new_n31386_, new_n31387_, new_n31388_, new_n31389_, new_n31390_,
    new_n31391_, new_n31392_, new_n31393_, new_n31394_, new_n31395_,
    new_n31396_, new_n31397_, new_n31398_, new_n31399_, new_n31400_,
    new_n31401_, new_n31402_, new_n31403_, new_n31404_, new_n31405_,
    new_n31406_, new_n31407_, new_n31408_, new_n31409_, new_n31410_,
    new_n31411_, new_n31412_, new_n31413_, new_n31414_, new_n31415_,
    new_n31416_, new_n31417_, new_n31418_, new_n31419_, new_n31420_,
    new_n31421_, new_n31422_, new_n31423_, new_n31424_, new_n31425_,
    new_n31426_, new_n31427_, new_n31428_, new_n31429_, new_n31430_,
    new_n31431_, new_n31432_, new_n31433_, new_n31434_, new_n31435_,
    new_n31436_, new_n31437_, new_n31438_, new_n31439_, new_n31440_,
    new_n31441_, new_n31442_, new_n31443_, new_n31444_, new_n31445_,
    new_n31446_, new_n31447_, new_n31448_, new_n31449_, new_n31450_,
    new_n31451_, new_n31452_, new_n31453_, new_n31454_, new_n31455_,
    new_n31456_, new_n31457_, new_n31458_, new_n31459_, new_n31460_,
    new_n31461_, new_n31462_, new_n31463_, new_n31464_, new_n31465_,
    new_n31466_, new_n31467_, new_n31468_, new_n31469_, new_n31470_,
    new_n31471_, new_n31472_, new_n31473_, new_n31474_, new_n31475_,
    new_n31476_, new_n31477_, new_n31478_, new_n31479_, new_n31480_,
    new_n31481_, new_n31482_, new_n31483_, new_n31484_, new_n31485_,
    new_n31486_, new_n31487_, new_n31488_, new_n31489_, new_n31490_,
    new_n31491_, new_n31492_, new_n31493_, new_n31494_, new_n31495_,
    new_n31496_, new_n31497_, new_n31498_, new_n31499_, new_n31500_,
    new_n31501_, new_n31502_, new_n31503_, new_n31504_, new_n31505_,
    new_n31506_, new_n31507_, new_n31508_, new_n31509_, new_n31510_,
    new_n31511_, new_n31512_, new_n31513_, new_n31514_, new_n31515_,
    new_n31516_, new_n31517_, new_n31518_, new_n31519_, new_n31520_,
    new_n31521_, new_n31522_, new_n31523_, new_n31524_, new_n31525_,
    new_n31526_, new_n31527_, new_n31528_, new_n31529_, new_n31530_,
    new_n31531_, new_n31532_, new_n31533_, new_n31534_, new_n31535_,
    new_n31536_, new_n31537_, new_n31538_, new_n31539_, new_n31540_,
    new_n31541_, new_n31542_, new_n31543_, new_n31544_, new_n31545_,
    new_n31546_, new_n31547_, new_n31548_, new_n31549_, new_n31550_,
    new_n31551_, new_n31552_, new_n31553_, new_n31554_, new_n31555_,
    new_n31556_, new_n31557_, new_n31558_, new_n31559_, new_n31560_,
    new_n31561_, new_n31562_, new_n31563_, new_n31564_, new_n31565_,
    new_n31566_, new_n31567_, new_n31568_, new_n31569_, new_n31570_,
    new_n31571_, new_n31572_, new_n31573_, new_n31574_, new_n31575_,
    new_n31576_, new_n31577_, new_n31578_, new_n31579_, new_n31580_,
    new_n31581_, new_n31582_, new_n31583_, new_n31584_, new_n31585_,
    new_n31586_, new_n31587_, new_n31588_, new_n31589_, new_n31590_,
    new_n31591_, new_n31592_, new_n31593_, new_n31594_, new_n31595_,
    new_n31596_, new_n31597_, new_n31598_, new_n31599_, new_n31600_,
    new_n31601_, new_n31602_, new_n31603_, new_n31604_, new_n31605_,
    new_n31606_, new_n31607_, new_n31608_, new_n31609_, new_n31610_,
    new_n31611_, new_n31612_, new_n31613_, new_n31614_, new_n31615_,
    new_n31616_, new_n31617_, new_n31618_, new_n31619_, new_n31620_,
    new_n31621_, new_n31622_, new_n31623_, new_n31624_, new_n31625_,
    new_n31626_, new_n31627_, new_n31628_, new_n31629_, new_n31630_,
    new_n31631_, new_n31632_, new_n31633_, new_n31634_, new_n31635_,
    new_n31636_, new_n31637_, new_n31638_, new_n31639_, new_n31640_,
    new_n31641_, new_n31642_, new_n31643_, new_n31644_, new_n31645_,
    new_n31646_, new_n31647_, new_n31648_, new_n31649_, new_n31650_,
    new_n31651_, new_n31652_, new_n31653_, new_n31654_, new_n31655_,
    new_n31656_, new_n31657_, new_n31658_, new_n31659_, new_n31660_,
    new_n31661_, new_n31662_, new_n31663_, new_n31664_, new_n31665_,
    new_n31666_, new_n31667_, new_n31668_, new_n31669_, new_n31670_,
    new_n31671_, new_n31672_, new_n31673_, new_n31674_, new_n31675_,
    new_n31676_, new_n31677_, new_n31678_, new_n31679_, new_n31680_,
    new_n31681_, new_n31682_, new_n31683_, new_n31684_, new_n31685_,
    new_n31686_, new_n31687_, new_n31688_, new_n31689_, new_n31690_,
    new_n31691_, new_n31692_, new_n31693_, new_n31694_, new_n31695_,
    new_n31696_, new_n31697_, new_n31698_, new_n31699_, new_n31700_,
    new_n31701_, new_n31702_, new_n31703_, new_n31704_, new_n31705_,
    new_n31706_, new_n31707_, new_n31708_, new_n31709_, new_n31710_,
    new_n31711_, new_n31712_, new_n31713_, new_n31714_, new_n31715_,
    new_n31716_, new_n31717_, new_n31718_, new_n31719_, new_n31720_,
    new_n31721_, new_n31722_, new_n31723_, new_n31724_, new_n31725_,
    new_n31726_, new_n31727_, new_n31728_, new_n31729_, new_n31730_,
    new_n31731_, new_n31732_, new_n31733_, new_n31734_, new_n31735_,
    new_n31736_, new_n31737_, new_n31738_, new_n31739_, new_n31740_,
    new_n31741_, new_n31742_, new_n31743_, new_n31744_, new_n31745_,
    new_n31746_, new_n31747_, new_n31748_, new_n31749_, new_n31750_,
    new_n31751_, new_n31752_, new_n31753_, new_n31754_, new_n31755_,
    new_n31756_, new_n31757_, new_n31758_, new_n31759_, new_n31760_,
    new_n31761_, new_n31762_, new_n31763_, new_n31764_, new_n31765_,
    new_n31766_, new_n31767_, new_n31768_, new_n31769_, new_n31770_,
    new_n31771_, new_n31772_, new_n31773_, new_n31774_, new_n31775_,
    new_n31776_, new_n31777_, new_n31778_, new_n31779_, new_n31780_,
    new_n31781_, new_n31782_, new_n31783_, new_n31784_, new_n31785_,
    new_n31786_, new_n31787_, new_n31788_, new_n31789_, new_n31790_,
    new_n31791_, new_n31792_, new_n31793_, new_n31794_, new_n31795_,
    new_n31796_, new_n31797_, new_n31798_, new_n31799_, new_n31800_,
    new_n31801_, new_n31802_, new_n31803_, new_n31804_, new_n31805_,
    new_n31806_, new_n31807_, new_n31808_, new_n31809_, new_n31810_,
    new_n31811_, new_n31812_, new_n31813_, new_n31814_, new_n31815_,
    new_n31816_, new_n31817_, new_n31818_, new_n31819_, new_n31820_,
    new_n31821_, new_n31822_, new_n31823_, new_n31824_, new_n31825_,
    new_n31826_, new_n31827_, new_n31828_, new_n31829_, new_n31830_,
    new_n31831_, new_n31832_, new_n31833_, new_n31834_, new_n31835_,
    new_n31836_, new_n31837_, new_n31838_, new_n31839_, new_n31840_,
    new_n31841_, new_n31842_, new_n31843_, new_n31844_, new_n31845_,
    new_n31846_, new_n31847_, new_n31848_, new_n31849_, new_n31850_,
    new_n31851_, new_n31852_, new_n31853_, new_n31854_, new_n31855_,
    new_n31856_, new_n31857_, new_n31858_, new_n31859_, new_n31860_,
    new_n31861_, new_n31862_, new_n31863_, new_n31864_, new_n31865_,
    new_n31866_, new_n31867_, new_n31868_, new_n31869_, new_n31870_,
    new_n31871_, new_n31872_, new_n31873_, new_n31874_, new_n31875_,
    new_n31876_, new_n31877_, new_n31878_, new_n31879_, new_n31880_,
    new_n31881_, new_n31882_, new_n31883_, new_n31884_, new_n31885_,
    new_n31886_, new_n31887_, new_n31888_, new_n31889_, new_n31890_,
    new_n31891_, new_n31892_, new_n31893_, new_n31894_, new_n31895_,
    new_n31896_, new_n31897_, new_n31898_, new_n31899_, new_n31900_,
    new_n31901_, new_n31902_, new_n31903_, new_n31904_, new_n31905_,
    new_n31906_, new_n31907_, new_n31908_, new_n31909_, new_n31910_,
    new_n31911_, new_n31912_, new_n31913_, new_n31914_, new_n31915_,
    new_n31916_, new_n31917_, new_n31918_, new_n31919_, new_n31920_,
    new_n31921_, new_n31922_, new_n31923_, new_n31924_, new_n31925_,
    new_n31926_, new_n31927_, new_n31928_, new_n31929_, new_n31930_,
    new_n31931_, new_n31932_, new_n31933_, new_n31934_, new_n31935_,
    new_n31936_, new_n31937_, new_n31938_, new_n31939_, new_n31940_,
    new_n31941_, new_n31942_, new_n31943_, new_n31944_, new_n31945_,
    new_n31946_, new_n31947_, new_n31948_, new_n31949_, new_n31950_,
    new_n31951_, new_n31952_, new_n31953_, new_n31954_, new_n31955_,
    new_n31956_, new_n31957_, new_n31958_, new_n31959_, new_n31960_,
    new_n31961_, new_n31962_, new_n31963_, new_n31964_, new_n31965_,
    new_n31966_, new_n31967_, new_n31968_, new_n31969_, new_n31970_,
    new_n31971_, new_n31972_, new_n31973_, new_n31974_, new_n31975_,
    new_n31976_, new_n31977_, new_n31978_, new_n31979_, new_n31980_,
    new_n31981_, new_n31982_, new_n31983_, new_n31984_, new_n31985_,
    new_n31986_, new_n31987_, new_n31988_, new_n31989_, new_n31990_,
    new_n31991_, new_n31992_, new_n31993_, new_n31994_, new_n31995_,
    new_n31996_, new_n31997_, new_n31998_, new_n31999_, new_n32000_,
    new_n32001_, new_n32002_, new_n32003_, new_n32004_, new_n32005_,
    new_n32006_, new_n32007_, new_n32008_, new_n32009_, new_n32010_,
    new_n32011_, new_n32012_, new_n32013_, new_n32014_, new_n32015_,
    new_n32016_, new_n32017_, new_n32018_, new_n32019_, new_n32020_,
    new_n32021_, new_n32022_, new_n32023_, new_n32024_, new_n32025_,
    new_n32026_, new_n32027_, new_n32028_, new_n32029_, new_n32030_,
    new_n32031_, new_n32032_, new_n32033_, new_n32034_, new_n32035_,
    new_n32036_, new_n32037_, new_n32038_, new_n32039_, new_n32040_,
    new_n32041_, new_n32042_, new_n32043_, new_n32044_, new_n32045_,
    new_n32046_, new_n32047_, new_n32048_, new_n32049_, new_n32050_,
    new_n32051_, new_n32052_, new_n32053_, new_n32054_, new_n32055_,
    new_n32056_, new_n32057_, new_n32058_, new_n32059_, new_n32060_,
    new_n32061_, new_n32062_, new_n32063_, new_n32064_, new_n32065_,
    new_n32066_, new_n32067_, new_n32068_, new_n32069_, new_n32070_,
    new_n32071_, new_n32072_, new_n32073_, new_n32074_, new_n32075_,
    new_n32076_, new_n32077_, new_n32078_, new_n32079_, new_n32080_,
    new_n32081_, new_n32082_, new_n32083_, new_n32084_, new_n32085_,
    new_n32086_, new_n32087_, new_n32088_, new_n32089_, new_n32090_,
    new_n32091_, new_n32092_, new_n32093_, new_n32094_, new_n32095_,
    new_n32096_, new_n32097_, new_n32098_, new_n32099_, new_n32100_,
    new_n32101_, new_n32102_, new_n32103_, new_n32104_, new_n32105_,
    new_n32106_, new_n32107_, new_n32108_, new_n32109_, new_n32110_,
    new_n32111_, new_n32112_, new_n32113_, new_n32114_, new_n32115_,
    new_n32116_, new_n32117_, new_n32118_, new_n32119_, new_n32120_,
    new_n32121_, new_n32122_, new_n32123_, new_n32124_, new_n32125_,
    new_n32126_, new_n32127_, new_n32128_, new_n32129_, new_n32130_,
    new_n32131_, new_n32132_, new_n32133_, new_n32134_, new_n32135_,
    new_n32136_, new_n32137_, new_n32138_, new_n32139_, new_n32140_,
    new_n32141_, new_n32142_, new_n32143_, new_n32144_, new_n32145_,
    new_n32146_, new_n32147_, new_n32148_, new_n32149_, new_n32150_,
    new_n32151_, new_n32152_, new_n32153_, new_n32154_, new_n32155_,
    new_n32156_, new_n32157_, new_n32158_, new_n32159_, new_n32160_,
    new_n32161_, new_n32162_, new_n32163_, new_n32164_, new_n32165_,
    new_n32166_, new_n32167_, new_n32168_, new_n32169_, new_n32170_,
    new_n32171_, new_n32172_, new_n32173_, new_n32174_, new_n32175_,
    new_n32176_, new_n32177_, new_n32178_, new_n32179_, new_n32180_,
    new_n32181_, new_n32182_, new_n32183_, new_n32184_, new_n32185_,
    new_n32186_, new_n32187_, new_n32188_, new_n32189_, new_n32190_,
    new_n32191_, new_n32192_, new_n32193_, new_n32194_, new_n32195_,
    new_n32196_, new_n32197_, new_n32198_, new_n32199_, new_n32200_,
    new_n32201_, new_n32202_, new_n32203_, new_n32204_, new_n32205_,
    new_n32206_, new_n32207_, new_n32208_, new_n32209_, new_n32210_,
    new_n32211_, new_n32212_, new_n32213_, new_n32214_, new_n32215_,
    new_n32216_, new_n32217_, new_n32218_, new_n32219_, new_n32220_,
    new_n32221_, new_n32222_, new_n32223_, new_n32224_, new_n32225_,
    new_n32226_, new_n32227_, new_n32228_, new_n32229_, new_n32230_,
    new_n32231_, new_n32232_, new_n32233_, new_n32234_, new_n32235_,
    new_n32236_, new_n32237_, new_n32238_, new_n32239_, new_n32240_,
    new_n32241_, new_n32242_, new_n32243_, new_n32244_, new_n32245_,
    new_n32246_, new_n32247_, new_n32248_, new_n32249_, new_n32250_,
    new_n32251_, new_n32252_, new_n32253_, new_n32254_, new_n32255_,
    new_n32256_, new_n32257_, new_n32258_, new_n32259_, new_n32260_,
    new_n32261_, new_n32262_, new_n32263_, new_n32264_, new_n32265_,
    new_n32266_, new_n32267_, new_n32268_, new_n32269_, new_n32270_,
    new_n32271_, new_n32272_, new_n32273_, new_n32274_, new_n32275_,
    new_n32276_, new_n32277_, new_n32278_, new_n32279_, new_n32280_,
    new_n32281_, new_n32282_, new_n32283_, new_n32284_, new_n32285_,
    new_n32286_, new_n32287_, new_n32288_, new_n32289_, new_n32290_,
    new_n32291_, new_n32292_, new_n32293_, new_n32294_, new_n32295_,
    new_n32296_, new_n32297_, new_n32298_, new_n32299_, new_n32300_,
    new_n32301_, new_n32302_, new_n32303_, new_n32304_, new_n32305_,
    new_n32306_, new_n32307_, new_n32308_, new_n32309_, new_n32310_,
    new_n32311_, new_n32312_, new_n32313_, new_n32314_, new_n32315_,
    new_n32316_, new_n32317_, new_n32318_, new_n32319_, new_n32320_,
    new_n32321_, new_n32322_, new_n32323_, new_n32324_, new_n32325_,
    new_n32326_, new_n32327_, new_n32328_, new_n32329_, new_n32330_,
    new_n32331_, new_n32332_, new_n32333_, new_n32334_, new_n32335_,
    new_n32336_, new_n32337_, new_n32338_, new_n32339_, new_n32340_,
    new_n32341_, new_n32342_, new_n32343_, new_n32344_, new_n32345_,
    new_n32346_, new_n32347_, new_n32348_, new_n32349_, new_n32350_,
    new_n32351_, new_n32352_, new_n32353_, new_n32354_, new_n32355_,
    new_n32356_, new_n32357_, new_n32358_, new_n32359_, new_n32360_,
    new_n32361_, new_n32362_, new_n32363_, new_n32364_, new_n32365_,
    new_n32366_, new_n32367_, new_n32368_, new_n32369_, new_n32370_,
    new_n32371_, new_n32372_, new_n32373_, new_n32374_, new_n32375_,
    new_n32376_, new_n32377_, new_n32378_, new_n32379_, new_n32380_,
    new_n32381_, new_n32382_, new_n32383_, new_n32384_, new_n32385_,
    new_n32386_, new_n32387_, new_n32388_, new_n32389_, new_n32390_,
    new_n32391_, new_n32392_, new_n32393_, new_n32394_, new_n32395_,
    new_n32396_, new_n32397_, new_n32398_, new_n32399_, new_n32400_,
    new_n32401_, new_n32402_, new_n32403_, new_n32404_, new_n32405_,
    new_n32406_, new_n32407_, new_n32408_, new_n32409_, new_n32410_,
    new_n32411_, new_n32412_, new_n32413_, new_n32414_, new_n32415_,
    new_n32416_, new_n32417_, new_n32418_, new_n32419_, new_n32420_,
    new_n32421_, new_n32422_, new_n32423_, new_n32424_, new_n32425_,
    new_n32426_, new_n32427_, new_n32428_, new_n32429_, new_n32430_,
    new_n32431_, new_n32432_, new_n32433_, new_n32434_, new_n32435_,
    new_n32436_, new_n32437_, new_n32438_, new_n32439_, new_n32440_,
    new_n32441_, new_n32442_, new_n32443_, new_n32444_, new_n32445_,
    new_n32446_, new_n32447_, new_n32448_, new_n32449_, new_n32450_,
    new_n32451_, new_n32452_, new_n32453_, new_n32454_, new_n32455_,
    new_n32456_, new_n32457_, new_n32458_, new_n32459_, new_n32460_,
    new_n32461_, new_n32462_, new_n32463_, new_n32464_, new_n32465_,
    new_n32466_, new_n32467_, new_n32468_, new_n32469_, new_n32470_,
    new_n32471_, new_n32472_, new_n32473_, new_n32474_, new_n32475_,
    new_n32476_, new_n32477_, new_n32478_, new_n32479_, new_n32480_,
    new_n32481_, new_n32482_, new_n32483_, new_n32484_, new_n32485_,
    new_n32486_, new_n32487_, new_n32488_, new_n32489_, new_n32490_,
    new_n32491_, new_n32492_, new_n32493_, new_n32494_, new_n32495_,
    new_n32496_, new_n32497_, new_n32498_, new_n32499_, new_n32500_,
    new_n32501_, new_n32502_, new_n32503_, new_n32504_, new_n32505_,
    new_n32506_, new_n32507_, new_n32508_, new_n32509_, new_n32510_,
    new_n32511_, new_n32512_, new_n32513_, new_n32514_, new_n32515_,
    new_n32516_, new_n32517_, new_n32518_, new_n32519_, new_n32520_,
    new_n32521_, new_n32522_, new_n32523_, new_n32524_, new_n32525_,
    new_n32526_, new_n32527_, new_n32528_, new_n32529_, new_n32530_,
    new_n32531_, new_n32532_, new_n32533_, new_n32534_, new_n32535_,
    new_n32536_, new_n32537_, new_n32538_, new_n32539_, new_n32540_,
    new_n32541_, new_n32542_, new_n32543_, new_n32544_, new_n32545_,
    new_n32546_, new_n32547_, new_n32548_, new_n32549_, new_n32550_,
    new_n32551_, new_n32552_, new_n32553_, new_n32554_, new_n32555_,
    new_n32556_, new_n32557_, new_n32558_, new_n32559_, new_n32560_,
    new_n32561_, new_n32562_, new_n32563_, new_n32564_, new_n32565_,
    new_n32566_, new_n32567_, new_n32568_, new_n32569_, new_n32570_,
    new_n32571_, new_n32572_, new_n32573_, new_n32574_, new_n32575_,
    new_n32576_, new_n32577_, new_n32578_, new_n32579_, new_n32580_,
    new_n32581_, new_n32582_, new_n32583_, new_n32584_, new_n32585_,
    new_n32586_, new_n32587_, new_n32588_, new_n32589_, new_n32590_,
    new_n32591_, new_n32592_, new_n32593_, new_n32594_, new_n32595_,
    new_n32596_, new_n32597_, new_n32598_, new_n32599_, new_n32600_,
    new_n32601_, new_n32602_, new_n32603_, new_n32604_, new_n32605_,
    new_n32606_, new_n32607_, new_n32608_, new_n32609_, new_n32610_,
    new_n32611_, new_n32612_, new_n32613_, new_n32614_, new_n32615_,
    new_n32616_, new_n32617_, new_n32618_, new_n32619_, new_n32620_,
    new_n32621_, new_n32622_, new_n32623_, new_n32624_, new_n32625_,
    new_n32626_, new_n32627_, new_n32628_, new_n32629_, new_n32630_,
    new_n32631_, new_n32632_, new_n32633_, new_n32634_, new_n32635_,
    new_n32636_, new_n32637_, new_n32638_, new_n32639_, new_n32640_,
    new_n32641_, new_n32642_, new_n32643_, new_n32644_, new_n32645_,
    new_n32646_, new_n32647_, new_n32648_, new_n32649_, new_n32650_,
    new_n32651_, new_n32652_, new_n32653_, new_n32654_, new_n32655_,
    new_n32656_, new_n32657_, new_n32658_, new_n32659_, new_n32660_,
    new_n32661_, new_n32662_, new_n32663_, new_n32664_, new_n32665_,
    new_n32666_, new_n32667_, new_n32668_, new_n32669_, new_n32670_,
    new_n32671_, new_n32672_, new_n32673_, new_n32674_, new_n32675_,
    new_n32676_, new_n32677_, new_n32678_, new_n32679_, new_n32680_,
    new_n32681_, new_n32682_, new_n32683_, new_n32684_, new_n32685_,
    new_n32686_, new_n32687_, new_n32688_, new_n32689_, new_n32690_,
    new_n32691_, new_n32692_, new_n32693_, new_n32694_, new_n32695_,
    new_n32696_, new_n32697_, new_n32698_, new_n32699_, new_n32700_,
    new_n32701_, new_n32702_, new_n32703_, new_n32704_, new_n32705_,
    new_n32706_, new_n32707_, new_n32708_, new_n32709_, new_n32710_,
    new_n32711_, new_n32712_, new_n32713_, new_n32714_, new_n32715_,
    new_n32716_, new_n32717_, new_n32718_, new_n32719_, new_n32720_,
    new_n32721_, new_n32722_, new_n32723_, new_n32724_, new_n32725_,
    new_n32726_, new_n32727_, new_n32728_, new_n32729_, new_n32730_,
    new_n32731_, new_n32732_, new_n32733_, new_n32734_, new_n32735_,
    new_n32736_, new_n32737_, new_n32738_, new_n32739_, new_n32740_,
    new_n32741_, new_n32742_, new_n32743_, new_n32744_, new_n32745_,
    new_n32746_, new_n32747_, new_n32748_, new_n32749_, new_n32750_,
    new_n32751_, new_n32752_, new_n32753_, new_n32754_, new_n32755_,
    new_n32756_, new_n32757_, new_n32758_, new_n32759_, new_n32760_,
    new_n32761_, new_n32762_, new_n32763_, new_n32764_, new_n32765_,
    new_n32766_, new_n32767_, new_n32768_, new_n32769_, new_n32770_,
    new_n32771_, new_n32772_, new_n32773_, new_n32774_, new_n32775_,
    new_n32776_, new_n32777_, new_n32778_, new_n32779_, new_n32780_,
    new_n32781_, new_n32782_, new_n32783_, new_n32784_, new_n32785_,
    new_n32786_, new_n32787_, new_n32788_, new_n32789_, new_n32790_,
    new_n32791_, new_n32792_, new_n32793_, new_n32794_, new_n32795_,
    new_n32796_, new_n32797_, new_n32798_, new_n32799_, new_n32800_,
    new_n32801_, new_n32802_, new_n32803_, new_n32804_, new_n32805_,
    new_n32806_, new_n32807_, new_n32808_, new_n32809_, new_n32810_,
    new_n32811_, new_n32812_, new_n32813_, new_n32814_, new_n32815_,
    new_n32816_, new_n32817_, new_n32818_, new_n32819_, new_n32820_,
    new_n32821_, new_n32822_, new_n32823_, new_n32824_, new_n32825_,
    new_n32826_, new_n32827_, new_n32828_, new_n32829_, new_n32830_,
    new_n32831_, new_n32832_, new_n32833_, new_n32834_, new_n32835_,
    new_n32836_, new_n32837_, new_n32838_, new_n32839_, new_n32840_,
    new_n32841_, new_n32842_, new_n32843_, new_n32844_, new_n32845_,
    new_n32846_, new_n32847_, new_n32848_, new_n32849_, new_n32850_,
    new_n32851_, new_n32852_, new_n32853_, new_n32854_, new_n32855_,
    new_n32856_, new_n32857_, new_n32858_, new_n32859_, new_n32860_,
    new_n32861_, new_n32862_, new_n32863_, new_n32864_, new_n32865_,
    new_n32866_, new_n32867_, new_n32868_, new_n32869_, new_n32870_,
    new_n32871_, new_n32872_, new_n32873_, new_n32874_, new_n32875_,
    new_n32876_, new_n32877_, new_n32878_, new_n32879_, new_n32880_,
    new_n32881_, new_n32882_, new_n32883_, new_n32884_, new_n32885_,
    new_n32886_, new_n32887_, new_n32888_, new_n32889_, new_n32890_,
    new_n32891_, new_n32892_, new_n32893_, new_n32894_, new_n32895_,
    new_n32896_, new_n32897_, new_n32898_, new_n32899_, new_n32900_,
    new_n32901_, new_n32902_, new_n32903_, new_n32904_, new_n32905_,
    new_n32906_, new_n32907_, new_n32908_, new_n32909_, new_n32910_,
    new_n32911_, new_n32912_, new_n32913_, new_n32914_, new_n32915_,
    new_n32916_, new_n32917_, new_n32918_, new_n32919_, new_n32920_,
    new_n32921_, new_n32922_, new_n32923_, new_n32924_, new_n32925_,
    new_n32926_, new_n32927_, new_n32928_, new_n32929_, new_n32930_,
    new_n32931_, new_n32932_, new_n32933_, new_n32934_, new_n32935_,
    new_n32936_, new_n32937_, new_n32938_, new_n32939_, new_n32940_,
    new_n32941_, new_n32942_, new_n32943_, new_n32944_, new_n32945_,
    new_n32946_, new_n32947_, new_n32948_, new_n32949_, new_n32950_,
    new_n32951_, new_n32952_, new_n32953_, new_n32954_, new_n32955_,
    new_n32956_, new_n32957_, new_n32958_, new_n32959_, new_n32960_,
    new_n32961_, new_n32962_, new_n32963_, new_n32964_, new_n32965_,
    new_n32966_, new_n32967_, new_n32968_, new_n32969_, new_n32970_,
    new_n32971_, new_n32972_, new_n32973_, new_n32974_, new_n32975_,
    new_n32976_, new_n32977_, new_n32978_, new_n32979_, new_n32980_,
    new_n32981_, new_n32982_, new_n32983_, new_n32984_, new_n32985_,
    new_n32986_, new_n32987_, new_n32988_, new_n32989_, new_n32990_,
    new_n32991_, new_n32992_, new_n32993_, new_n32994_, new_n32995_,
    new_n32996_, new_n32997_, new_n32998_, new_n32999_, new_n33000_,
    new_n33001_, new_n33002_, new_n33003_, new_n33004_, new_n33005_,
    new_n33006_, new_n33007_, new_n33008_, new_n33009_, new_n33010_,
    new_n33011_, new_n33012_, new_n33013_, new_n33014_, new_n33015_,
    new_n33016_, new_n33017_, new_n33018_, new_n33019_, new_n33020_,
    new_n33021_, new_n33022_, new_n33023_, new_n33024_, new_n33025_,
    new_n33026_, new_n33027_, new_n33028_, new_n33029_, new_n33030_,
    new_n33031_, new_n33032_, new_n33033_, new_n33034_, new_n33035_,
    new_n33036_, new_n33037_, new_n33038_, new_n33039_, new_n33040_,
    new_n33041_, new_n33042_, new_n33043_, new_n33044_, new_n33045_,
    new_n33046_, new_n33047_, new_n33048_, new_n33049_, new_n33050_,
    new_n33051_, new_n33052_, new_n33053_, new_n33054_, new_n33055_,
    new_n33056_, new_n33057_, new_n33058_, new_n33059_, new_n33060_,
    new_n33061_, new_n33062_, new_n33063_, new_n33064_, new_n33065_,
    new_n33066_, new_n33067_, new_n33068_, new_n33069_, new_n33070_,
    new_n33071_, new_n33072_, new_n33073_, new_n33074_, new_n33075_,
    new_n33076_, new_n33077_, new_n33078_, new_n33079_, new_n33080_,
    new_n33081_, new_n33082_, new_n33083_, new_n33084_, new_n33085_,
    new_n33086_, new_n33087_, new_n33088_, new_n33089_, new_n33090_,
    new_n33091_, new_n33092_, new_n33093_, new_n33094_, new_n33095_,
    new_n33096_, new_n33097_, new_n33098_, new_n33099_, new_n33100_,
    new_n33101_, new_n33102_, new_n33103_, new_n33104_, new_n33105_,
    new_n33106_, new_n33107_, new_n33108_, new_n33109_, new_n33110_,
    new_n33111_, new_n33112_, new_n33113_, new_n33114_, new_n33115_,
    new_n33116_, new_n33117_, new_n33118_, new_n33119_, new_n33120_,
    new_n33121_, new_n33122_, new_n33123_, new_n33124_, new_n33125_,
    new_n33126_, new_n33127_, new_n33128_, new_n33129_, new_n33130_,
    new_n33131_, new_n33132_, new_n33133_, new_n33134_, new_n33135_,
    new_n33136_, new_n33137_, new_n33138_, new_n33139_, new_n33140_,
    new_n33141_, new_n33142_, new_n33143_, new_n33144_, new_n33145_,
    new_n33146_, new_n33147_, new_n33148_, new_n33149_, new_n33150_,
    new_n33151_, new_n33152_, new_n33153_, new_n33154_, new_n33155_,
    new_n33156_, new_n33157_, new_n33158_, new_n33159_, new_n33160_,
    new_n33161_, new_n33162_, new_n33163_, new_n33164_, new_n33165_,
    new_n33166_, new_n33167_, new_n33168_, new_n33169_, new_n33170_,
    new_n33171_, new_n33172_, new_n33173_, new_n33174_, new_n33175_,
    new_n33176_, new_n33177_, new_n33178_, new_n33179_, new_n33180_,
    new_n33181_, new_n33182_, new_n33183_, new_n33184_, new_n33185_,
    new_n33186_, new_n33187_, new_n33188_, new_n33189_, new_n33190_,
    new_n33191_, new_n33192_, new_n33193_, new_n33194_, new_n33195_,
    new_n33196_, new_n33197_, new_n33198_, new_n33199_, new_n33200_,
    new_n33201_, new_n33202_, new_n33203_, new_n33204_, new_n33205_,
    new_n33206_, new_n33207_, new_n33208_, new_n33209_, new_n33210_,
    new_n33211_, new_n33212_, new_n33213_, new_n33214_, new_n33215_,
    new_n33216_, new_n33217_, new_n33218_, new_n33219_, new_n33220_,
    new_n33221_, new_n33222_, new_n33223_, new_n33224_, new_n33225_,
    new_n33226_, new_n33227_, new_n33228_, new_n33229_, new_n33230_,
    new_n33231_, new_n33232_, new_n33233_, new_n33234_, new_n33235_,
    new_n33236_, new_n33237_, new_n33238_, new_n33239_, new_n33240_,
    new_n33241_, new_n33242_, new_n33243_, new_n33244_, new_n33245_,
    new_n33246_, new_n33247_, new_n33248_, new_n33249_, new_n33250_,
    new_n33251_, new_n33252_, new_n33253_, new_n33254_, new_n33255_,
    new_n33256_, new_n33257_, new_n33258_, new_n33259_, new_n33260_,
    new_n33261_, new_n33262_, new_n33263_, new_n33264_, new_n33265_,
    new_n33266_, new_n33267_, new_n33268_, new_n33269_, new_n33270_,
    new_n33271_, new_n33272_, new_n33273_, new_n33274_, new_n33275_,
    new_n33276_, new_n33277_, new_n33278_, new_n33279_, new_n33280_,
    new_n33281_, new_n33282_, new_n33283_, new_n33284_, new_n33285_,
    new_n33286_, new_n33287_, new_n33288_, new_n33289_, new_n33290_,
    new_n33291_, new_n33292_, new_n33293_, new_n33294_, new_n33295_,
    new_n33296_, new_n33297_, new_n33298_, new_n33299_, new_n33300_,
    new_n33301_, new_n33302_, new_n33303_, new_n33304_, new_n33305_,
    new_n33306_, new_n33307_, new_n33308_, new_n33309_, new_n33310_,
    new_n33311_, new_n33312_, new_n33313_, new_n33314_, new_n33315_,
    new_n33316_, new_n33317_, new_n33318_, new_n33319_, new_n33320_,
    new_n33321_, new_n33322_, new_n33323_, new_n33324_, new_n33325_,
    new_n33326_, new_n33327_, new_n33328_, new_n33329_, new_n33330_,
    new_n33331_, new_n33332_, new_n33333_, new_n33334_, new_n33335_,
    new_n33336_, new_n33337_, new_n33338_, new_n33339_, new_n33340_,
    new_n33341_, new_n33342_, new_n33343_, new_n33344_, new_n33345_,
    new_n33346_, new_n33347_, new_n33348_, new_n33349_, new_n33350_,
    new_n33351_, new_n33352_, new_n33353_, new_n33354_, new_n33355_,
    new_n33356_, new_n33357_, new_n33358_, new_n33359_, new_n33360_,
    new_n33361_, new_n33362_, new_n33363_, new_n33364_, new_n33365_,
    new_n33366_, new_n33367_, new_n33368_, new_n33369_, new_n33370_,
    new_n33371_, new_n33372_, new_n33373_, new_n33374_, new_n33375_,
    new_n33376_, new_n33377_, new_n33378_, new_n33379_, new_n33380_,
    new_n33381_, new_n33382_, new_n33383_, new_n33384_, new_n33385_,
    new_n33386_, new_n33387_, new_n33388_, new_n33389_, new_n33390_,
    new_n33391_, new_n33392_, new_n33393_, new_n33394_, new_n33395_,
    new_n33396_, new_n33397_, new_n33398_, new_n33399_, new_n33400_,
    new_n33401_, new_n33402_, new_n33403_, new_n33404_, new_n33405_,
    new_n33406_, new_n33407_, new_n33408_, new_n33409_, new_n33410_,
    new_n33411_, new_n33412_, new_n33413_, new_n33414_, new_n33415_,
    new_n33416_, new_n33417_, new_n33418_, new_n33419_, new_n33420_,
    new_n33421_, new_n33422_, new_n33423_, new_n33424_, new_n33425_,
    new_n33426_, new_n33427_, new_n33428_, new_n33429_, new_n33430_,
    new_n33431_, new_n33432_, new_n33433_, new_n33434_, new_n33435_,
    new_n33436_, new_n33437_, new_n33438_, new_n33439_, new_n33440_,
    new_n33441_, new_n33442_, new_n33443_, new_n33444_, new_n33445_,
    new_n33446_, new_n33447_, new_n33448_, new_n33449_, new_n33450_,
    new_n33451_, new_n33452_, new_n33453_, new_n33454_, new_n33455_,
    new_n33456_, new_n33457_, new_n33458_, new_n33459_, new_n33460_,
    new_n33461_, new_n33462_, new_n33463_, new_n33464_, new_n33465_,
    new_n33466_, new_n33467_, new_n33468_, new_n33469_, new_n33470_,
    new_n33471_, new_n33472_, new_n33473_, new_n33474_, new_n33475_,
    new_n33476_, new_n33477_, new_n33478_, new_n33479_, new_n33480_,
    new_n33481_, new_n33482_, new_n33483_, new_n33484_, new_n33485_,
    new_n33486_, new_n33487_, new_n33488_, new_n33489_, new_n33490_,
    new_n33491_, new_n33492_, new_n33493_, new_n33494_, new_n33495_,
    new_n33496_, new_n33497_, new_n33498_, new_n33499_, new_n33500_,
    new_n33501_, new_n33502_, new_n33503_, new_n33504_, new_n33505_,
    new_n33506_, new_n33507_, new_n33508_, new_n33509_, new_n33510_,
    new_n33511_, new_n33512_, new_n33513_, new_n33514_, new_n33515_,
    new_n33516_, new_n33517_, new_n33518_, new_n33519_, new_n33520_,
    new_n33521_, new_n33522_, new_n33523_, new_n33524_, new_n33525_,
    new_n33526_, new_n33527_, new_n33528_, new_n33529_, new_n33530_,
    new_n33531_, new_n33532_, new_n33533_, new_n33534_, new_n33535_,
    new_n33536_, new_n33537_, new_n33538_, new_n33539_, new_n33540_,
    new_n33541_, new_n33542_, new_n33543_, new_n33544_, new_n33545_,
    new_n33546_, new_n33547_, new_n33548_, new_n33549_, new_n33550_,
    new_n33551_, new_n33552_, new_n33553_, new_n33554_, new_n33555_,
    new_n33556_, new_n33557_, new_n33558_, new_n33559_, new_n33560_,
    new_n33561_, new_n33562_, new_n33563_, new_n33564_, new_n33565_,
    new_n33566_, new_n33567_, new_n33568_, new_n33569_, new_n33570_,
    new_n33571_, new_n33572_, new_n33573_, new_n33574_, new_n33575_,
    new_n33576_, new_n33577_, new_n33578_, new_n33579_, new_n33580_,
    new_n33581_, new_n33582_, new_n33583_, new_n33584_, new_n33585_,
    new_n33586_, new_n33587_, new_n33588_, new_n33589_, new_n33590_,
    new_n33591_, new_n33592_, new_n33593_, new_n33594_, new_n33595_,
    new_n33596_, new_n33597_, new_n33598_, new_n33599_, new_n33600_,
    new_n33601_, new_n33602_, new_n33603_, new_n33604_, new_n33605_,
    new_n33606_, new_n33607_, new_n33608_, new_n33609_, new_n33610_,
    new_n33611_, new_n33612_, new_n33613_, new_n33614_, new_n33615_,
    new_n33616_, new_n33617_, new_n33618_, new_n33619_, new_n33620_,
    new_n33621_, new_n33622_, new_n33623_, new_n33624_, new_n33625_,
    new_n33626_, new_n33627_, new_n33628_, new_n33629_, new_n33630_,
    new_n33631_, new_n33632_, new_n33633_, new_n33634_, new_n33635_,
    new_n33636_, new_n33637_, new_n33638_, new_n33639_, new_n33640_,
    new_n33641_, new_n33642_, new_n33643_, new_n33644_, new_n33645_,
    new_n33646_, new_n33647_, new_n33648_, new_n33649_, new_n33650_,
    new_n33651_, new_n33652_, new_n33653_, new_n33654_, new_n33655_,
    new_n33656_, new_n33657_, new_n33658_, new_n33659_, new_n33660_,
    new_n33661_, new_n33662_, new_n33663_, new_n33664_, new_n33665_,
    new_n33666_, new_n33667_, new_n33668_, new_n33669_, new_n33670_,
    new_n33671_, new_n33672_, new_n33673_, new_n33674_, new_n33675_,
    new_n33676_, new_n33677_, new_n33678_, new_n33679_, new_n33680_,
    new_n33681_, new_n33682_, new_n33683_, new_n33684_, new_n33685_,
    new_n33686_, new_n33687_, new_n33688_, new_n33689_, new_n33690_,
    new_n33691_, new_n33692_, new_n33693_, new_n33694_, new_n33695_,
    new_n33696_, new_n33697_, new_n33698_, new_n33699_, new_n33700_,
    new_n33701_, new_n33702_, new_n33703_, new_n33704_, new_n33705_,
    new_n33706_, new_n33707_, new_n33708_, new_n33709_, new_n33710_,
    new_n33711_, new_n33712_, new_n33713_, new_n33714_, new_n33715_,
    new_n33716_, new_n33717_, new_n33718_, new_n33719_, new_n33720_,
    new_n33721_, new_n33722_, new_n33723_, new_n33724_, new_n33725_,
    new_n33726_, new_n33727_, new_n33728_, new_n33729_, new_n33730_,
    new_n33731_, new_n33732_, new_n33733_, new_n33734_, new_n33735_,
    new_n33736_, new_n33737_, new_n33738_, new_n33739_, new_n33740_,
    new_n33741_, new_n33742_, new_n33743_, new_n33744_, new_n33745_,
    new_n33746_, new_n33747_, new_n33748_, new_n33749_, new_n33750_,
    new_n33751_, new_n33752_, new_n33753_, new_n33754_, new_n33755_,
    new_n33756_, new_n33757_, new_n33758_, new_n33759_, new_n33760_,
    new_n33761_, new_n33762_, new_n33763_, new_n33764_, new_n33765_,
    new_n33766_, new_n33767_, new_n33768_, new_n33769_, new_n33770_,
    new_n33771_, new_n33772_, new_n33773_, new_n33774_, new_n33775_,
    new_n33776_, new_n33777_, new_n33778_, new_n33779_, new_n33780_,
    new_n33781_, new_n33782_, new_n33783_, new_n33784_, new_n33785_,
    new_n33786_, new_n33787_, new_n33788_, new_n33789_, new_n33790_,
    new_n33791_, new_n33792_, new_n33793_, new_n33794_, new_n33795_,
    new_n33796_, new_n33797_, new_n33798_, new_n33799_, new_n33800_,
    new_n33801_, new_n33802_, new_n33803_, new_n33804_, new_n33805_,
    new_n33806_, new_n33807_, new_n33808_, new_n33809_, new_n33810_,
    new_n33811_, new_n33812_, new_n33813_, new_n33814_, new_n33815_,
    new_n33816_, new_n33817_, new_n33818_, new_n33819_, new_n33820_,
    new_n33821_, new_n33822_, new_n33823_, new_n33824_, new_n33825_,
    new_n33826_, new_n33827_, new_n33828_, new_n33829_, new_n33830_,
    new_n33831_, new_n33832_, new_n33833_, new_n33834_, new_n33835_,
    new_n33836_, new_n33837_, new_n33838_, new_n33839_, new_n33840_,
    new_n33841_, new_n33842_, new_n33843_, new_n33844_, new_n33845_,
    new_n33846_, new_n33847_, new_n33848_, new_n33849_, new_n33850_,
    new_n33851_, new_n33852_, new_n33853_, new_n33854_, new_n33855_,
    new_n33856_, new_n33857_, new_n33858_, new_n33859_, new_n33860_,
    new_n33861_, new_n33862_, new_n33863_, new_n33864_, new_n33865_,
    new_n33866_, new_n33867_, new_n33868_, new_n33869_, new_n33870_,
    new_n33871_, new_n33872_, new_n33873_, new_n33874_, new_n33875_,
    new_n33876_, new_n33877_, new_n33878_, new_n33879_, new_n33880_,
    new_n33881_, new_n33882_, new_n33883_, new_n33884_, new_n33885_,
    new_n33886_, new_n33887_, new_n33888_, new_n33889_, new_n33890_,
    new_n33891_, new_n33892_, new_n33893_, new_n33894_, new_n33895_,
    new_n33896_, new_n33897_, new_n33898_, new_n33899_, new_n33900_,
    new_n33901_, new_n33902_, new_n33903_, new_n33904_, new_n33905_,
    new_n33906_, new_n33907_, new_n33908_, new_n33909_, new_n33910_,
    new_n33911_, new_n33912_, new_n33913_, new_n33914_, new_n33915_,
    new_n33916_, new_n33917_, new_n33918_, new_n33919_, new_n33920_,
    new_n33921_, new_n33922_, new_n33923_, new_n33924_, new_n33925_,
    new_n33926_, new_n33927_, new_n33928_, new_n33929_, new_n33930_,
    new_n33931_, new_n33932_, new_n33933_, new_n33934_, new_n33935_,
    new_n33936_, new_n33937_, new_n33938_, new_n33939_, new_n33940_,
    new_n33941_, new_n33942_, new_n33943_, new_n33944_, new_n33945_,
    new_n33946_, new_n33947_, new_n33948_, new_n33949_, new_n33950_,
    new_n33951_, new_n33952_, new_n33953_, new_n33954_, new_n33955_,
    new_n33956_, new_n33957_, new_n33958_, new_n33959_, new_n33960_,
    new_n33961_, new_n33962_, new_n33963_, new_n33964_, new_n33965_,
    new_n33966_, new_n33967_, new_n33968_, new_n33969_, new_n33970_,
    new_n33971_, new_n33972_, new_n33973_, new_n33974_, new_n33975_,
    new_n33976_, new_n33977_, new_n33978_, new_n33979_, new_n33980_,
    new_n33981_, new_n33982_, new_n33983_, new_n33984_, new_n33985_,
    new_n33986_, new_n33987_, new_n33988_, new_n33989_, new_n33990_,
    new_n33991_, new_n33992_, new_n33993_, new_n33994_, new_n33995_,
    new_n33996_, new_n33997_, new_n33998_, new_n33999_, new_n34000_,
    new_n34001_, new_n34002_, new_n34003_, new_n34004_, new_n34005_,
    new_n34006_, new_n34007_, new_n34008_, new_n34009_, new_n34010_,
    new_n34011_, new_n34012_, new_n34013_, new_n34014_, new_n34015_,
    new_n34016_, new_n34017_, new_n34018_, new_n34019_, new_n34020_,
    new_n34021_, new_n34022_, new_n34023_, new_n34024_, new_n34025_,
    new_n34026_, new_n34027_, new_n34028_, new_n34029_, new_n34030_,
    new_n34031_, new_n34032_, new_n34033_, new_n34034_, new_n34035_,
    new_n34036_, new_n34037_, new_n34038_, new_n34039_, new_n34040_,
    new_n34041_, new_n34042_, new_n34043_, new_n34044_, new_n34045_,
    new_n34046_, new_n34047_, new_n34048_, new_n34049_, new_n34050_,
    new_n34051_, new_n34052_, new_n34053_, new_n34054_, new_n34055_,
    new_n34056_, new_n34057_, new_n34058_, new_n34059_, new_n34060_,
    new_n34061_, new_n34062_, new_n34063_, new_n34064_, new_n34065_,
    new_n34066_, new_n34067_, new_n34068_, new_n34069_, new_n34070_,
    new_n34071_, new_n34072_, new_n34073_, new_n34074_, new_n34075_,
    new_n34076_, new_n34077_, new_n34078_, new_n34079_, new_n34080_,
    new_n34081_, new_n34082_, new_n34083_, new_n34084_, new_n34085_,
    new_n34086_, new_n34087_, new_n34088_, new_n34089_, new_n34090_,
    new_n34091_, new_n34092_, new_n34093_, new_n34094_, new_n34095_,
    new_n34096_, new_n34097_, new_n34098_, new_n34099_, new_n34100_,
    new_n34101_, new_n34102_, new_n34103_, new_n34104_, new_n34105_,
    new_n34106_, new_n34107_, new_n34108_, new_n34109_, new_n34110_,
    new_n34111_, new_n34112_, new_n34113_, new_n34114_, new_n34115_,
    new_n34116_, new_n34117_, new_n34118_, new_n34119_, new_n34120_,
    new_n34121_, new_n34122_, new_n34123_, new_n34124_, new_n34125_,
    new_n34126_, new_n34127_, new_n34128_, new_n34129_, new_n34130_,
    new_n34131_, new_n34132_, new_n34133_, new_n34134_, new_n34135_,
    new_n34136_, new_n34137_, new_n34138_, new_n34139_, new_n34140_,
    new_n34141_, new_n34142_, new_n34143_, new_n34144_, new_n34145_,
    new_n34146_, new_n34147_, new_n34148_, new_n34149_, new_n34150_,
    new_n34151_, new_n34152_, new_n34153_, new_n34154_, new_n34155_,
    new_n34156_, new_n34157_, new_n34158_, new_n34159_, new_n34160_,
    new_n34161_, new_n34162_, new_n34163_, new_n34164_, new_n34165_,
    new_n34166_, new_n34167_, new_n34168_, new_n34169_, new_n34170_,
    new_n34171_, new_n34172_, new_n34173_, new_n34174_, new_n34175_,
    new_n34176_, new_n34177_, new_n34178_, new_n34179_, new_n34180_,
    new_n34181_, new_n34182_, new_n34183_, new_n34184_, new_n34185_,
    new_n34186_, new_n34187_, new_n34188_, new_n34189_, new_n34190_,
    new_n34191_, new_n34192_, new_n34193_, new_n34194_, new_n34195_,
    new_n34196_, new_n34197_, new_n34198_, new_n34199_, new_n34200_,
    new_n34201_, new_n34202_, new_n34203_, new_n34204_, new_n34205_,
    new_n34206_, new_n34207_, new_n34208_, new_n34209_, new_n34210_,
    new_n34211_, new_n34212_, new_n34213_, new_n34214_, new_n34215_,
    new_n34216_, new_n34217_, new_n34218_, new_n34219_, new_n34220_,
    new_n34221_, new_n34222_, new_n34223_, new_n34224_, new_n34225_,
    new_n34226_, new_n34227_, new_n34228_, new_n34229_, new_n34230_,
    new_n34231_, new_n34232_, new_n34233_, new_n34234_, new_n34235_,
    new_n34236_, new_n34237_, new_n34238_, new_n34239_, new_n34240_,
    new_n34241_, new_n34242_, new_n34243_, new_n34244_, new_n34245_,
    new_n34246_, new_n34247_, new_n34248_, new_n34249_, new_n34250_,
    new_n34251_, new_n34252_, new_n34253_, new_n34254_, new_n34255_,
    new_n34256_, new_n34257_, new_n34258_, new_n34259_, new_n34260_,
    new_n34261_, new_n34262_, new_n34263_, new_n34264_, new_n34265_,
    new_n34266_, new_n34267_, new_n34268_, new_n34269_, new_n34270_,
    new_n34271_, new_n34272_, new_n34273_, new_n34274_, new_n34275_,
    new_n34276_, new_n34277_, new_n34278_, new_n34279_, new_n34280_,
    new_n34281_, new_n34282_, new_n34283_, new_n34284_, new_n34285_,
    new_n34286_, new_n34287_, new_n34288_, new_n34289_, new_n34290_,
    new_n34291_, new_n34292_, new_n34293_, new_n34294_, new_n34295_,
    new_n34296_, new_n34297_, new_n34298_, new_n34299_, new_n34300_,
    new_n34301_, new_n34302_, new_n34303_, new_n34304_, new_n34305_,
    new_n34306_, new_n34307_, new_n34308_, new_n34309_, new_n34310_,
    new_n34311_, new_n34312_, new_n34313_, new_n34314_, new_n34315_,
    new_n34316_, new_n34317_, new_n34318_, new_n34319_, new_n34320_,
    new_n34321_, new_n34322_, new_n34323_, new_n34324_, new_n34325_,
    new_n34326_, new_n34327_, new_n34328_, new_n34329_, new_n34330_,
    new_n34331_, new_n34332_, new_n34333_, new_n34334_, new_n34335_,
    new_n34336_, new_n34337_, new_n34338_, new_n34339_, new_n34340_,
    new_n34341_, new_n34342_, new_n34343_, new_n34344_, new_n34345_,
    new_n34346_, new_n34347_, new_n34348_, new_n34349_, new_n34350_,
    new_n34351_, new_n34352_, new_n34353_, new_n34354_, new_n34355_,
    new_n34356_, new_n34357_, new_n34358_, new_n34359_, new_n34360_,
    new_n34361_, new_n34362_, new_n34363_, new_n34364_, new_n34365_,
    new_n34366_, new_n34367_, new_n34368_, new_n34369_, new_n34370_,
    new_n34371_, new_n34372_, new_n34373_, new_n34374_, new_n34375_,
    new_n34376_, new_n34377_, new_n34378_, new_n34379_, new_n34380_,
    new_n34381_, new_n34382_, new_n34383_, new_n34384_, new_n34385_,
    new_n34386_, new_n34387_, new_n34388_, new_n34389_, new_n34390_,
    new_n34391_, new_n34392_, new_n34393_, new_n34394_, new_n34395_,
    new_n34396_, new_n34397_, new_n34398_, new_n34399_, new_n34400_,
    new_n34401_, new_n34402_, new_n34403_, new_n34404_, new_n34405_,
    new_n34406_, new_n34407_, new_n34408_, new_n34409_, new_n34410_,
    new_n34411_, new_n34412_, new_n34413_, new_n34414_, new_n34415_,
    new_n34416_, new_n34417_, new_n34418_, new_n34419_, new_n34420_,
    new_n34421_, new_n34422_, new_n34423_, new_n34424_, new_n34425_,
    new_n34426_, new_n34427_, new_n34428_, new_n34429_, new_n34430_,
    new_n34431_, new_n34432_, new_n34433_, new_n34434_, new_n34435_,
    new_n34436_, new_n34437_, new_n34438_, new_n34439_, new_n34440_,
    new_n34441_, new_n34442_, new_n34443_, new_n34444_, new_n34445_,
    new_n34446_, new_n34447_, new_n34448_, new_n34449_, new_n34450_,
    new_n34451_, new_n34452_, new_n34453_, new_n34454_, new_n34455_,
    new_n34456_, new_n34457_, new_n34458_, new_n34459_, new_n34460_,
    new_n34461_, new_n34462_, new_n34463_, new_n34464_, new_n34465_,
    new_n34466_, new_n34467_, new_n34468_, new_n34469_, new_n34470_,
    new_n34471_, new_n34472_, new_n34473_, new_n34474_, new_n34475_,
    new_n34476_, new_n34477_, new_n34478_, new_n34479_, new_n34480_,
    new_n34481_, new_n34482_, new_n34483_, new_n34484_, new_n34485_,
    new_n34486_, new_n34487_, new_n34488_, new_n34489_, new_n34490_,
    new_n34491_, new_n34492_, new_n34493_, new_n34494_, new_n34495_,
    new_n34496_, new_n34497_, new_n34498_, new_n34499_, new_n34500_,
    new_n34501_, new_n34502_, new_n34503_, new_n34504_, new_n34505_,
    new_n34506_, new_n34507_, new_n34508_, new_n34509_, new_n34510_,
    new_n34511_, new_n34512_, new_n34513_, new_n34514_, new_n34515_,
    new_n34516_, new_n34517_, new_n34518_, new_n34519_, new_n34520_,
    new_n34521_, new_n34522_, new_n34523_, new_n34524_, new_n34525_,
    new_n34526_, new_n34527_, new_n34528_, new_n34529_, new_n34530_,
    new_n34531_, new_n34532_, new_n34533_, new_n34534_, new_n34535_,
    new_n34536_, new_n34537_, new_n34538_, new_n34539_, new_n34540_,
    new_n34541_, new_n34542_, new_n34543_, new_n34544_, new_n34545_,
    new_n34546_, new_n34547_, new_n34548_, new_n34549_, new_n34550_,
    new_n34551_, new_n34552_, new_n34553_, new_n34554_, new_n34555_,
    new_n34556_, new_n34557_, new_n34558_, new_n34559_, new_n34560_,
    new_n34561_, new_n34562_, new_n34563_, new_n34564_, new_n34565_,
    new_n34566_, new_n34567_, new_n34568_, new_n34569_, new_n34570_,
    new_n34571_, new_n34572_, new_n34573_, new_n34574_, new_n34575_,
    new_n34576_, new_n34577_, new_n34578_, new_n34579_, new_n34580_,
    new_n34581_, new_n34582_, new_n34583_, new_n34584_, new_n34585_,
    new_n34586_, new_n34587_, new_n34588_, new_n34589_, new_n34590_,
    new_n34591_, new_n34592_, new_n34593_, new_n34594_, new_n34595_,
    new_n34596_, new_n34597_, new_n34598_, new_n34599_, new_n34600_,
    new_n34601_, new_n34602_, new_n34603_, new_n34604_, new_n34605_,
    new_n34606_, new_n34607_, new_n34608_, new_n34609_, new_n34610_,
    new_n34611_, new_n34612_, new_n34613_, new_n34614_, new_n34615_,
    new_n34616_, new_n34617_, new_n34618_, new_n34619_, new_n34620_,
    new_n34621_, new_n34622_, new_n34623_, new_n34624_, new_n34625_,
    new_n34626_, new_n34627_, new_n34628_, new_n34629_, new_n34630_,
    new_n34631_, new_n34632_, new_n34633_, new_n34634_, new_n34635_,
    new_n34636_, new_n34637_, new_n34638_, new_n34639_, new_n34640_,
    new_n34641_, new_n34642_, new_n34643_, new_n34644_, new_n34645_,
    new_n34646_, new_n34647_, new_n34648_, new_n34649_, new_n34650_,
    new_n34651_, new_n34652_, new_n34653_, new_n34654_, new_n34655_,
    new_n34656_, new_n34657_, new_n34658_, new_n34659_, new_n34660_,
    new_n34661_, new_n34662_, new_n34663_, new_n34664_, new_n34665_,
    new_n34666_, new_n34667_, new_n34668_, new_n34669_, new_n34670_,
    new_n34671_, new_n34672_, new_n34673_, new_n34674_, new_n34675_,
    new_n34676_, new_n34677_, new_n34678_, new_n34679_, new_n34680_,
    new_n34681_, new_n34682_, new_n34683_, new_n34684_, new_n34685_,
    new_n34686_, new_n34687_, new_n34688_, new_n34689_, new_n34690_,
    new_n34691_, new_n34692_, new_n34693_, new_n34694_, new_n34695_,
    new_n34696_, new_n34697_, new_n34698_, new_n34699_, new_n34700_,
    new_n34701_, new_n34702_, new_n34703_, new_n34704_, new_n34705_,
    new_n34706_, new_n34707_, new_n34708_, new_n34709_, new_n34710_,
    new_n34711_, new_n34712_, new_n34713_, new_n34714_, new_n34715_,
    new_n34716_, new_n34717_, new_n34718_, new_n34719_, new_n34720_,
    new_n34721_, new_n34722_, new_n34723_, new_n34724_, new_n34725_,
    new_n34726_, new_n34727_, new_n34728_, new_n34729_, new_n34730_,
    new_n34731_, new_n34732_, new_n34733_, new_n34734_, new_n34735_,
    new_n34736_, new_n34737_, new_n34738_, new_n34739_, new_n34740_,
    new_n34741_, new_n34742_, new_n34743_, new_n34744_, new_n34745_,
    new_n34746_, new_n34747_, new_n34748_, new_n34749_, new_n34750_,
    new_n34751_, new_n34752_, new_n34753_, new_n34754_, new_n34755_,
    new_n34756_, new_n34757_, new_n34758_, new_n34759_, new_n34760_,
    new_n34761_, new_n34762_, new_n34763_, new_n34764_, new_n34765_,
    new_n34766_, new_n34767_, new_n34768_, new_n34769_, new_n34770_,
    new_n34771_, new_n34772_, new_n34773_, new_n34774_, new_n34775_,
    new_n34776_, new_n34777_, new_n34778_, new_n34779_, new_n34780_,
    new_n34781_, new_n34782_, new_n34783_, new_n34784_, new_n34785_,
    new_n34786_, new_n34787_, new_n34788_, new_n34789_, new_n34790_,
    new_n34791_, new_n34792_, new_n34793_, new_n34794_, new_n34795_,
    new_n34796_, new_n34797_, new_n34798_, new_n34799_, new_n34800_,
    new_n34801_, new_n34802_, new_n34803_, new_n34804_, new_n34805_,
    new_n34806_, new_n34807_, new_n34808_, new_n34809_, new_n34810_,
    new_n34811_, new_n34812_, new_n34813_, new_n34814_, new_n34815_,
    new_n34816_, new_n34817_, new_n34818_, new_n34819_, new_n34820_,
    new_n34821_, new_n34822_, new_n34823_, new_n34824_, new_n34825_,
    new_n34826_, new_n34827_, new_n34828_, new_n34829_, new_n34830_,
    new_n34831_, new_n34832_, new_n34833_, new_n34834_, new_n34835_,
    new_n34836_, new_n34837_, new_n34838_, new_n34839_, new_n34840_,
    new_n34841_, new_n34842_, new_n34843_, new_n34844_, new_n34845_,
    new_n34846_, new_n34847_, new_n34848_, new_n34849_, new_n34850_,
    new_n34851_, new_n34852_, new_n34853_, new_n34854_, new_n34855_,
    new_n34856_, new_n34857_, new_n34858_, new_n34859_, new_n34860_,
    new_n34861_, new_n34862_, new_n34863_, new_n34864_, new_n34865_,
    new_n34866_, new_n34867_, new_n34868_, new_n34869_, new_n34870_,
    new_n34871_, new_n34872_, new_n34873_, new_n34874_, new_n34875_,
    new_n34876_, new_n34877_, new_n34878_, new_n34879_, new_n34880_,
    new_n34881_, new_n34882_, new_n34883_, new_n34884_, new_n34885_,
    new_n34886_, new_n34887_, new_n34888_, new_n34889_, new_n34890_,
    new_n34891_, new_n34892_, new_n34893_, new_n34894_, new_n34895_,
    new_n34896_, new_n34897_, new_n34898_, new_n34899_, new_n34900_,
    new_n34901_, new_n34902_, new_n34903_, new_n34904_, new_n34905_,
    new_n34906_, new_n34907_, new_n34908_, new_n34909_, new_n34910_,
    new_n34911_, new_n34912_, new_n34913_, new_n34914_, new_n34915_,
    new_n34916_, new_n34917_, new_n34918_, new_n34919_, new_n34920_,
    new_n34921_, new_n34922_, new_n34923_, new_n34924_, new_n34925_,
    new_n34926_, new_n34927_, new_n34928_, new_n34929_, new_n34930_,
    new_n34931_, new_n34932_, new_n34933_, new_n34934_, new_n34935_,
    new_n34936_, new_n34937_, new_n34938_, new_n34939_, new_n34940_,
    new_n34941_, new_n34942_, new_n34943_, new_n34944_, new_n34945_,
    new_n34946_, new_n34947_, new_n34948_, new_n34949_, new_n34950_,
    new_n34951_, new_n34952_, new_n34953_, new_n34954_, new_n34955_,
    new_n34956_, new_n34957_, new_n34958_, new_n34959_, new_n34960_,
    new_n34961_, new_n34962_, new_n34963_, new_n34964_, new_n34965_,
    new_n34966_, new_n34967_, new_n34968_, new_n34969_, new_n34970_,
    new_n34971_, new_n34972_, new_n34973_, new_n34974_, new_n34975_,
    new_n34976_, new_n34977_, new_n34978_, new_n34979_, new_n34980_,
    new_n34981_, new_n34982_, new_n34983_, new_n34984_, new_n34985_,
    new_n34986_, new_n34987_, new_n34988_, new_n34989_, new_n34990_,
    new_n34991_, new_n34992_, new_n34993_, new_n34994_, new_n34995_,
    new_n34996_, new_n34997_, new_n34998_, new_n34999_, new_n35000_,
    new_n35001_, new_n35002_, new_n35003_, new_n35004_, new_n35005_,
    new_n35006_, new_n35007_, new_n35008_, new_n35009_, new_n35010_,
    new_n35011_, new_n35012_, new_n35013_, new_n35014_, new_n35015_,
    new_n35016_, new_n35017_, new_n35018_, new_n35019_, new_n35020_,
    new_n35021_, new_n35022_, new_n35023_, new_n35024_, new_n35025_,
    new_n35026_, new_n35027_, new_n35028_, new_n35029_, new_n35030_,
    new_n35031_, new_n35032_, new_n35033_, new_n35034_, new_n35035_,
    new_n35036_, new_n35037_, new_n35038_, new_n35039_, new_n35040_,
    new_n35041_, new_n35042_, new_n35043_, new_n35044_, new_n35045_,
    new_n35046_, new_n35047_, new_n35048_, new_n35049_, new_n35050_,
    new_n35051_, new_n35052_, new_n35053_, new_n35054_, new_n35055_,
    new_n35056_, new_n35057_, new_n35058_, new_n35059_, new_n35060_,
    new_n35061_, new_n35062_, new_n35063_, new_n35064_, new_n35065_,
    new_n35066_, new_n35067_, new_n35068_, new_n35069_, new_n35070_,
    new_n35071_, new_n35072_, new_n35073_, new_n35074_, new_n35075_,
    new_n35076_, new_n35077_, new_n35078_, new_n35079_, new_n35080_,
    new_n35081_, new_n35082_, new_n35083_, new_n35084_, new_n35085_,
    new_n35086_, new_n35087_, new_n35088_, new_n35089_, new_n35090_,
    new_n35091_, new_n35092_, new_n35093_, new_n35094_, new_n35095_,
    new_n35096_, new_n35097_, new_n35098_, new_n35099_, new_n35100_,
    new_n35101_, new_n35102_, new_n35103_, new_n35104_, new_n35105_,
    new_n35106_, new_n35107_, new_n35108_, new_n35109_, new_n35110_,
    new_n35111_, new_n35112_, new_n35113_, new_n35114_, new_n35115_,
    new_n35116_, new_n35117_, new_n35118_, new_n35119_, new_n35120_,
    new_n35121_, new_n35122_, new_n35123_, new_n35124_, new_n35125_,
    new_n35126_, new_n35127_, new_n35128_, new_n35129_, new_n35130_,
    new_n35131_, new_n35132_, new_n35133_, new_n35134_, new_n35135_,
    new_n35136_, new_n35137_, new_n35138_, new_n35139_, new_n35140_,
    new_n35141_, new_n35142_, new_n35143_, new_n35144_, new_n35145_,
    new_n35146_, new_n35147_, new_n35148_, new_n35149_, new_n35150_,
    new_n35151_, new_n35152_, new_n35153_, new_n35154_, new_n35155_,
    new_n35156_, new_n35157_, new_n35158_, new_n35159_, new_n35160_,
    new_n35161_, new_n35162_, new_n35163_, new_n35164_, new_n35165_,
    new_n35166_, new_n35167_, new_n35168_, new_n35169_, new_n35170_,
    new_n35171_, new_n35172_, new_n35173_, new_n35174_, new_n35175_,
    new_n35176_, new_n35177_, new_n35178_, new_n35179_, new_n35180_,
    new_n35181_, new_n35182_, new_n35183_, new_n35184_, new_n35185_,
    new_n35186_, new_n35187_, new_n35188_, new_n35189_, new_n35190_,
    new_n35191_, new_n35192_, new_n35193_, new_n35194_, new_n35195_,
    new_n35196_, new_n35197_, new_n35198_, new_n35199_, new_n35200_,
    new_n35201_, new_n35202_, new_n35203_, new_n35204_, new_n35205_,
    new_n35206_, new_n35207_, new_n35208_, new_n35209_, new_n35210_,
    new_n35211_, new_n35212_, new_n35213_, new_n35214_, new_n35215_,
    new_n35216_, new_n35217_, new_n35218_, new_n35219_, new_n35220_,
    new_n35221_, new_n35222_, new_n35223_, new_n35224_, new_n35225_,
    new_n35226_, new_n35227_, new_n35228_, new_n35229_, new_n35230_,
    new_n35231_, new_n35232_, new_n35233_, new_n35234_, new_n35235_,
    new_n35236_, new_n35237_, new_n35238_, new_n35239_, new_n35240_,
    new_n35241_, new_n35242_, new_n35243_, new_n35244_, new_n35245_,
    new_n35246_, new_n35247_, new_n35248_, new_n35249_, new_n35250_,
    new_n35251_, new_n35252_, new_n35253_, new_n35254_, new_n35255_,
    new_n35256_, new_n35257_, new_n35258_, new_n35259_, new_n35260_,
    new_n35261_, new_n35262_, new_n35263_, new_n35264_, new_n35265_,
    new_n35266_, new_n35267_, new_n35268_, new_n35269_, new_n35270_,
    new_n35271_, new_n35272_, new_n35273_, new_n35274_, new_n35275_,
    new_n35276_, new_n35277_, new_n35278_, new_n35279_, new_n35280_,
    new_n35281_, new_n35282_, new_n35283_, new_n35284_, new_n35285_,
    new_n35286_, new_n35287_, new_n35288_, new_n35289_, new_n35290_,
    new_n35291_, new_n35292_, new_n35293_, new_n35294_, new_n35295_,
    new_n35296_, new_n35297_, new_n35298_, new_n35299_, new_n35300_,
    new_n35301_, new_n35302_, new_n35303_, new_n35304_, new_n35305_,
    new_n35306_, new_n35307_, new_n35308_, new_n35309_, new_n35310_,
    new_n35311_, new_n35312_, new_n35313_, new_n35314_, new_n35315_,
    new_n35316_, new_n35317_, new_n35318_, new_n35319_, new_n35320_,
    new_n35321_, new_n35322_, new_n35323_, new_n35324_, new_n35325_,
    new_n35326_, new_n35327_, new_n35328_, new_n35329_, new_n35330_,
    new_n35331_, new_n35332_, new_n35333_, new_n35334_, new_n35335_,
    new_n35336_, new_n35337_, new_n35338_, new_n35339_, new_n35340_,
    new_n35341_, new_n35342_, new_n35343_, new_n35344_, new_n35345_,
    new_n35346_, new_n35347_, new_n35348_, new_n35349_, new_n35350_,
    new_n35351_, new_n35352_, new_n35353_, new_n35354_, new_n35355_,
    new_n35356_, new_n35357_, new_n35358_, new_n35359_, new_n35360_,
    new_n35361_, new_n35362_, new_n35363_, new_n35364_, new_n35365_,
    new_n35366_, new_n35367_, new_n35368_, new_n35369_, new_n35370_,
    new_n35371_, new_n35372_, new_n35373_, new_n35374_, new_n35375_,
    new_n35376_, new_n35377_, new_n35378_, new_n35379_, new_n35380_,
    new_n35381_, new_n35382_, new_n35383_, new_n35384_, new_n35385_,
    new_n35386_, new_n35387_, new_n35388_, new_n35389_, new_n35390_,
    new_n35391_, new_n35392_, new_n35393_, new_n35394_, new_n35395_,
    new_n35396_, new_n35397_, new_n35398_, new_n35399_, new_n35400_,
    new_n35401_, new_n35402_, new_n35403_, new_n35404_, new_n35405_,
    new_n35406_, new_n35407_, new_n35408_, new_n35409_, new_n35410_,
    new_n35411_, new_n35412_, new_n35413_, new_n35414_, new_n35415_,
    new_n35416_, new_n35417_, new_n35418_, new_n35419_, new_n35420_,
    new_n35421_, new_n35422_, new_n35423_, new_n35424_, new_n35425_,
    new_n35426_, new_n35427_, new_n35428_, new_n35429_, new_n35430_,
    new_n35431_, new_n35432_, new_n35433_, new_n35434_, new_n35435_,
    new_n35436_, new_n35437_, new_n35438_, new_n35439_, new_n35440_,
    new_n35441_, new_n35442_, new_n35443_, new_n35444_, new_n35445_,
    new_n35446_, new_n35447_, new_n35448_, new_n35449_, new_n35450_,
    new_n35451_, new_n35452_, new_n35453_, new_n35454_, new_n35455_,
    new_n35456_, new_n35457_, new_n35458_, new_n35459_, new_n35460_,
    new_n35461_, new_n35462_, new_n35463_, new_n35464_, new_n35465_,
    new_n35466_, new_n35467_, new_n35468_, new_n35469_, new_n35470_,
    new_n35471_, new_n35472_, new_n35473_, new_n35474_, new_n35475_,
    new_n35476_, new_n35477_, new_n35478_, new_n35479_, new_n35480_,
    new_n35481_, new_n35482_, new_n35483_, new_n35484_, new_n35485_,
    new_n35486_, new_n35487_, new_n35488_, new_n35489_, new_n35490_,
    new_n35491_, new_n35492_, new_n35493_, new_n35494_, new_n35495_,
    new_n35496_, new_n35497_, new_n35498_, new_n35499_, new_n35500_,
    new_n35501_, new_n35502_, new_n35503_, new_n35504_, new_n35505_,
    new_n35506_, new_n35507_, new_n35508_, new_n35509_, new_n35510_,
    new_n35511_, new_n35512_, new_n35513_, new_n35514_, new_n35515_,
    new_n35516_, new_n35517_, new_n35518_, new_n35519_, new_n35520_,
    new_n35521_, new_n35522_, new_n35523_, new_n35524_, new_n35525_,
    new_n35526_, new_n35527_, new_n35528_, new_n35529_, new_n35530_,
    new_n35531_, new_n35532_, new_n35533_, new_n35534_, new_n35535_,
    new_n35536_, new_n35537_, new_n35538_, new_n35539_, new_n35540_,
    new_n35541_, new_n35542_, new_n35543_, new_n35544_, new_n35545_,
    new_n35546_, new_n35547_, new_n35548_, new_n35549_, new_n35550_,
    new_n35551_, new_n35552_, new_n35553_, new_n35554_, new_n35555_,
    new_n35556_, new_n35557_, new_n35558_, new_n35559_, new_n35560_,
    new_n35561_, new_n35562_, new_n35563_, new_n35564_, new_n35565_,
    new_n35566_, new_n35567_, new_n35568_, new_n35569_, new_n35570_,
    new_n35571_, new_n35572_, new_n35573_, new_n35574_, new_n35575_,
    new_n35576_, new_n35577_, new_n35578_, new_n35579_, new_n35580_,
    new_n35581_, new_n35582_, new_n35583_, new_n35584_, new_n35585_,
    new_n35586_, new_n35587_, new_n35588_, new_n35589_, new_n35590_,
    new_n35591_, new_n35592_, new_n35593_, new_n35594_, new_n35595_,
    new_n35596_, new_n35597_, new_n35598_, new_n35599_, new_n35600_,
    new_n35601_, new_n35602_, new_n35603_, new_n35604_, new_n35605_,
    new_n35606_, new_n35607_, new_n35608_, new_n35609_, new_n35610_,
    new_n35611_, new_n35612_, new_n35613_, new_n35614_, new_n35615_,
    new_n35616_, new_n35617_, new_n35618_, new_n35619_, new_n35620_,
    new_n35621_, new_n35622_, new_n35623_, new_n35624_, new_n35625_,
    new_n35626_, new_n35627_, new_n35628_, new_n35629_, new_n35630_,
    new_n35631_, new_n35632_, new_n35633_, new_n35634_, new_n35635_,
    new_n35636_, new_n35637_, new_n35638_, new_n35639_, new_n35640_,
    new_n35641_, new_n35642_, new_n35643_, new_n35644_, new_n35645_,
    new_n35646_, new_n35647_, new_n35648_, new_n35649_, new_n35650_,
    new_n35651_, new_n35652_, new_n35653_, new_n35654_, new_n35655_,
    new_n35656_, new_n35657_, new_n35658_, new_n35659_, new_n35660_,
    new_n35661_, new_n35662_, new_n35663_, new_n35664_, new_n35665_,
    new_n35666_, new_n35667_, new_n35668_, new_n35669_, new_n35670_,
    new_n35671_, new_n35672_, new_n35673_, new_n35674_, new_n35675_,
    new_n35676_, new_n35677_, new_n35678_, new_n35679_, new_n35680_,
    new_n35681_, new_n35682_, new_n35683_, new_n35684_, new_n35685_,
    new_n35686_, new_n35687_, new_n35688_, new_n35689_, new_n35690_,
    new_n35691_, new_n35692_, new_n35693_, new_n35694_, new_n35695_,
    new_n35696_, new_n35697_, new_n35698_, new_n35699_, new_n35700_,
    new_n35701_, new_n35702_, new_n35703_, new_n35704_, new_n35705_,
    new_n35706_, new_n35707_, new_n35708_, new_n35709_, new_n35710_,
    new_n35711_, new_n35712_, new_n35713_, new_n35714_, new_n35715_,
    new_n35716_, new_n35717_, new_n35718_, new_n35719_, new_n35720_,
    new_n35721_, new_n35722_, new_n35723_, new_n35724_, new_n35725_,
    new_n35726_, new_n35727_, new_n35728_, new_n35729_, new_n35730_,
    new_n35731_, new_n35732_, new_n35733_, new_n35734_, new_n35735_,
    new_n35736_, new_n35737_, new_n35738_, new_n35739_, new_n35740_,
    new_n35741_, new_n35742_, new_n35743_, new_n35744_, new_n35745_,
    new_n35746_, new_n35747_, new_n35748_, new_n35749_, new_n35750_,
    new_n35751_, new_n35752_, new_n35753_, new_n35754_, new_n35755_,
    new_n35756_, new_n35757_, new_n35758_, new_n35759_, new_n35760_,
    new_n35761_, new_n35762_, new_n35763_, new_n35764_, new_n35765_,
    new_n35766_, new_n35767_, new_n35768_, new_n35769_, new_n35770_,
    new_n35771_, new_n35772_, new_n35773_, new_n35774_, new_n35775_,
    new_n35776_, new_n35777_, new_n35778_, new_n35779_, new_n35780_,
    new_n35781_, new_n35782_, new_n35783_, new_n35784_, new_n35785_,
    new_n35786_, new_n35787_, new_n35788_, new_n35789_, new_n35790_,
    new_n35791_, new_n35792_, new_n35793_, new_n35794_, new_n35795_,
    new_n35796_, new_n35797_, new_n35798_, new_n35799_, new_n35800_,
    new_n35801_, new_n35802_, new_n35803_, new_n35804_, new_n35805_,
    new_n35806_, new_n35807_, new_n35808_, new_n35809_, new_n35810_,
    new_n35811_, new_n35812_, new_n35813_, new_n35814_, new_n35815_,
    new_n35816_, new_n35817_, new_n35818_, new_n35819_, new_n35820_,
    new_n35821_, new_n35822_, new_n35823_, new_n35824_, new_n35825_,
    new_n35826_, new_n35827_, new_n35828_, new_n35829_, new_n35830_,
    new_n35831_, new_n35832_, new_n35833_, new_n35834_, new_n35835_,
    new_n35836_, new_n35837_, new_n35838_, new_n35839_, new_n35840_,
    new_n35841_, new_n35842_, new_n35843_, new_n35844_, new_n35845_,
    new_n35846_, new_n35847_, new_n35848_, new_n35849_, new_n35850_,
    new_n35851_, new_n35852_, new_n35853_, new_n35854_, new_n35855_,
    new_n35856_, new_n35857_, new_n35858_, new_n35859_, new_n35860_,
    new_n35861_, new_n35862_, new_n35863_, new_n35864_, new_n35865_,
    new_n35866_, new_n35867_, new_n35868_, new_n35869_, new_n35870_,
    new_n35871_, new_n35872_, new_n35873_, new_n35874_, new_n35875_,
    new_n35876_, new_n35877_, new_n35878_, new_n35879_, new_n35880_,
    new_n35881_, new_n35882_, new_n35883_, new_n35884_, new_n35885_,
    new_n35886_, new_n35887_, new_n35888_, new_n35889_, new_n35890_,
    new_n35891_, new_n35892_, new_n35893_, new_n35894_, new_n35895_,
    new_n35896_, new_n35897_, new_n35898_, new_n35899_, new_n35900_,
    new_n35901_, new_n35902_, new_n35903_, new_n35904_, new_n35905_,
    new_n35906_, new_n35907_, new_n35908_, new_n35909_, new_n35910_,
    new_n35911_, new_n35912_, new_n35913_, new_n35914_, new_n35915_,
    new_n35916_, new_n35917_, new_n35918_, new_n35919_, new_n35920_,
    new_n35921_, new_n35922_, new_n35923_, new_n35924_, new_n35925_,
    new_n35926_, new_n35927_, new_n35928_, new_n35929_, new_n35930_,
    new_n35931_, new_n35932_, new_n35933_, new_n35934_, new_n35935_,
    new_n35936_, new_n35937_, new_n35938_, new_n35939_, new_n35940_,
    new_n35941_, new_n35942_, new_n35943_, new_n35944_, new_n35945_,
    new_n35946_, new_n35947_, new_n35948_, new_n35949_, new_n35950_,
    new_n35951_, new_n35952_, new_n35953_, new_n35954_, new_n35955_,
    new_n35956_, new_n35957_, new_n35958_, new_n35959_, new_n35960_,
    new_n35961_, new_n35962_, new_n35963_, new_n35964_, new_n35965_,
    new_n35966_, new_n35967_, new_n35968_, new_n35969_, new_n35970_,
    new_n35971_, new_n35972_, new_n35973_, new_n35974_, new_n35975_,
    new_n35976_, new_n35977_, new_n35978_, new_n35979_, new_n35980_,
    new_n35981_, new_n35982_, new_n35983_, new_n35984_, new_n35985_,
    new_n35986_, new_n35987_, new_n35988_, new_n35989_, new_n35990_,
    new_n35991_, new_n35992_, new_n35993_, new_n35994_, new_n35995_,
    new_n35996_, new_n35997_, new_n35998_, new_n35999_, new_n36000_,
    new_n36001_, new_n36002_, new_n36003_, new_n36004_, new_n36005_,
    new_n36006_, new_n36007_, new_n36008_, new_n36009_, new_n36010_,
    new_n36011_, new_n36012_, new_n36013_, new_n36014_, new_n36015_,
    new_n36016_, new_n36017_, new_n36018_, new_n36019_, new_n36020_,
    new_n36021_, new_n36022_, new_n36023_, new_n36024_, new_n36025_,
    new_n36026_, new_n36027_, new_n36028_, new_n36029_, new_n36030_,
    new_n36031_, new_n36032_, new_n36033_, new_n36034_, new_n36035_,
    new_n36036_, new_n36037_, new_n36038_, new_n36039_, new_n36040_,
    new_n36041_, new_n36042_, new_n36043_, new_n36044_, new_n36045_,
    new_n36046_, new_n36047_, new_n36048_, new_n36049_, new_n36050_,
    new_n36051_, new_n36052_, new_n36053_, new_n36054_, new_n36055_,
    new_n36056_, new_n36057_, new_n36058_, new_n36059_, new_n36060_,
    new_n36061_, new_n36062_, new_n36063_, new_n36064_, new_n36065_,
    new_n36066_, new_n36067_, new_n36068_, new_n36069_, new_n36070_,
    new_n36071_, new_n36072_, new_n36073_, new_n36074_, new_n36075_,
    new_n36076_, new_n36077_, new_n36078_, new_n36079_, new_n36080_,
    new_n36081_, new_n36082_, new_n36083_, new_n36084_, new_n36085_,
    new_n36086_, new_n36087_, new_n36088_, new_n36089_, new_n36090_,
    new_n36091_, new_n36092_, new_n36093_, new_n36094_, new_n36095_,
    new_n36096_, new_n36097_, new_n36098_, new_n36099_, new_n36100_,
    new_n36101_, new_n36102_, new_n36103_, new_n36104_, new_n36105_,
    new_n36106_, new_n36107_, new_n36108_, new_n36109_, new_n36110_,
    new_n36111_, new_n36112_, new_n36113_, new_n36114_, new_n36115_,
    new_n36116_, new_n36117_, new_n36118_, new_n36119_, new_n36120_,
    new_n36121_, new_n36122_, new_n36123_, new_n36124_, new_n36125_,
    new_n36126_, new_n36127_, new_n36128_, new_n36129_, new_n36130_,
    new_n36131_, new_n36132_, new_n36133_, new_n36134_, new_n36135_,
    new_n36136_, new_n36137_, new_n36138_, new_n36139_, new_n36140_,
    new_n36141_, new_n36142_, new_n36143_, new_n36144_, new_n36145_,
    new_n36146_, new_n36147_, new_n36148_, new_n36149_, new_n36150_,
    new_n36151_, new_n36152_, new_n36153_, new_n36154_, new_n36155_,
    new_n36156_, new_n36157_, new_n36158_, new_n36159_, new_n36160_,
    new_n36161_, new_n36162_, new_n36163_, new_n36164_, new_n36165_,
    new_n36166_, new_n36167_, new_n36168_, new_n36169_, new_n36170_,
    new_n36171_, new_n36172_, new_n36173_, new_n36174_, new_n36175_,
    new_n36176_, new_n36177_, new_n36178_, new_n36179_, new_n36180_,
    new_n36181_, new_n36182_, new_n36183_, new_n36184_, new_n36185_,
    new_n36186_, new_n36187_, new_n36188_, new_n36189_, new_n36190_,
    new_n36191_, new_n36192_, new_n36193_, new_n36194_, new_n36195_,
    new_n36196_, new_n36197_, new_n36198_, new_n36199_, new_n36200_,
    new_n36201_, new_n36202_, new_n36203_, new_n36204_, new_n36205_,
    new_n36206_, new_n36207_, new_n36208_, new_n36209_, new_n36210_,
    new_n36211_, new_n36212_, new_n36213_, new_n36214_, new_n36215_,
    new_n36216_, new_n36217_, new_n36218_, new_n36219_, new_n36220_,
    new_n36221_, new_n36222_, new_n36223_, new_n36224_, new_n36225_,
    new_n36226_, new_n36227_, new_n36228_, new_n36229_, new_n36230_,
    new_n36231_, new_n36232_, new_n36233_, new_n36234_, new_n36235_,
    new_n36236_, new_n36237_, new_n36238_, new_n36239_, new_n36240_,
    new_n36241_, new_n36242_, new_n36243_, new_n36244_, new_n36245_,
    new_n36246_, new_n36247_, new_n36248_, new_n36249_, new_n36250_,
    new_n36251_, new_n36252_, new_n36253_, new_n36254_, new_n36255_,
    new_n36256_, new_n36257_, new_n36258_, new_n36259_, new_n36260_,
    new_n36261_, new_n36262_, new_n36263_, new_n36264_, new_n36265_,
    new_n36266_, new_n36267_, new_n36268_, new_n36269_, new_n36270_,
    new_n36271_, new_n36272_, new_n36273_, new_n36274_, new_n36275_,
    new_n36276_, new_n36277_, new_n36278_, new_n36279_, new_n36280_,
    new_n36281_, new_n36282_, new_n36283_, new_n36284_, new_n36285_,
    new_n36286_, new_n36287_, new_n36288_, new_n36289_, new_n36290_,
    new_n36291_, new_n36292_, new_n36293_, new_n36294_, new_n36295_,
    new_n36296_, new_n36297_, new_n36298_, new_n36299_, new_n36300_,
    new_n36301_, new_n36302_, new_n36303_, new_n36304_, new_n36305_,
    new_n36306_, new_n36307_, new_n36308_, new_n36309_, new_n36310_,
    new_n36311_, new_n36312_, new_n36313_, new_n36314_, new_n36315_,
    new_n36316_, new_n36317_, new_n36318_, new_n36319_, new_n36320_,
    new_n36321_, new_n36322_, new_n36323_, new_n36324_, new_n36325_,
    new_n36326_, new_n36327_, new_n36328_, new_n36329_, new_n36330_,
    new_n36331_, new_n36332_, new_n36333_, new_n36334_, new_n36335_,
    new_n36336_, new_n36337_, new_n36338_, new_n36339_, new_n36340_,
    new_n36341_, new_n36342_, new_n36343_, new_n36344_, new_n36345_,
    new_n36346_, new_n36347_, new_n36348_, new_n36349_, new_n36350_,
    new_n36351_, new_n36352_, new_n36353_, new_n36354_, new_n36355_,
    new_n36356_, new_n36357_, new_n36358_, new_n36359_, new_n36360_,
    new_n36361_, new_n36362_, new_n36363_, new_n36364_, new_n36365_,
    new_n36366_, new_n36367_, new_n36368_, new_n36369_, new_n36370_,
    new_n36371_, new_n36372_, new_n36373_, new_n36374_, new_n36375_,
    new_n36376_, new_n36377_, new_n36378_, new_n36379_, new_n36380_,
    new_n36381_, new_n36382_, new_n36383_, new_n36384_, new_n36385_,
    new_n36386_, new_n36387_, new_n36388_, new_n36389_, new_n36390_,
    new_n36391_, new_n36392_, new_n36393_, new_n36394_, new_n36395_,
    new_n36396_, new_n36397_, new_n36398_, new_n36399_, new_n36400_,
    new_n36401_, new_n36402_, new_n36403_, new_n36404_, new_n36405_,
    new_n36406_, new_n36407_, new_n36408_, new_n36409_, new_n36410_,
    new_n36411_, new_n36412_, new_n36413_, new_n36414_, new_n36415_,
    new_n36416_, new_n36417_, new_n36418_, new_n36419_, new_n36420_,
    new_n36421_, new_n36422_, new_n36423_, new_n36424_, new_n36425_,
    new_n36426_, new_n36427_, new_n36428_, new_n36429_, new_n36430_,
    new_n36431_, new_n36432_, new_n36433_, new_n36434_, new_n36435_,
    new_n36436_, new_n36437_, new_n36438_, new_n36439_, new_n36440_,
    new_n36441_, new_n36442_, new_n36443_, new_n36444_, new_n36445_,
    new_n36446_, new_n36447_, new_n36448_, new_n36449_, new_n36450_,
    new_n36451_, new_n36452_, new_n36453_, new_n36454_, new_n36455_,
    new_n36456_, new_n36457_, new_n36458_, new_n36459_, new_n36460_,
    new_n36461_, new_n36462_, new_n36463_, new_n36464_, new_n36465_,
    new_n36466_, new_n36467_, new_n36468_, new_n36469_, new_n36470_,
    new_n36471_, new_n36472_, new_n36473_, new_n36474_, new_n36475_,
    new_n36476_, new_n36477_, new_n36478_, new_n36479_, new_n36480_,
    new_n36481_, new_n36482_, new_n36483_, new_n36484_, new_n36485_,
    new_n36486_, new_n36487_, new_n36488_, new_n36489_, new_n36490_,
    new_n36491_, new_n36492_, new_n36493_, new_n36494_, new_n36495_,
    new_n36496_, new_n36497_, new_n36498_, new_n36499_, new_n36500_,
    new_n36501_, new_n36502_, new_n36503_, new_n36504_, new_n36505_,
    new_n36506_, new_n36507_, new_n36508_, new_n36509_, new_n36510_,
    new_n36511_, new_n36512_, new_n36513_, new_n36514_, new_n36515_,
    new_n36516_, new_n36517_, new_n36518_, new_n36519_, new_n36520_,
    new_n36521_, new_n36522_, new_n36523_, new_n36524_, new_n36525_,
    new_n36526_, new_n36527_, new_n36528_, new_n36529_, new_n36530_,
    new_n36531_, new_n36532_, new_n36533_, new_n36534_, new_n36535_,
    new_n36536_, new_n36537_, new_n36538_, new_n36539_, new_n36540_,
    new_n36541_, new_n36542_, new_n36543_, new_n36544_, new_n36545_,
    new_n36546_, new_n36547_, new_n36548_, new_n36549_, new_n36550_,
    new_n36551_, new_n36552_, new_n36553_, new_n36554_, new_n36555_,
    new_n36556_, new_n36557_, new_n36558_, new_n36559_, new_n36560_,
    new_n36561_, new_n36562_, new_n36563_, new_n36564_, new_n36565_,
    new_n36566_, new_n36567_, new_n36568_, new_n36569_, new_n36570_,
    new_n36571_, new_n36572_, new_n36573_, new_n36574_, new_n36575_,
    new_n36576_, new_n36577_, new_n36578_, new_n36579_, new_n36580_,
    new_n36581_, new_n36582_, new_n36583_, new_n36584_, new_n36585_,
    new_n36586_, new_n36587_, new_n36588_, new_n36589_, new_n36590_,
    new_n36591_, new_n36592_, new_n36593_, new_n36594_, new_n36595_,
    new_n36596_, new_n36597_, new_n36598_, new_n36599_, new_n36600_,
    new_n36601_, new_n36602_, new_n36603_, new_n36604_, new_n36605_,
    new_n36606_, new_n36607_, new_n36608_, new_n36609_, new_n36610_,
    new_n36611_, new_n36612_, new_n36613_, new_n36614_, new_n36615_,
    new_n36616_, new_n36617_, new_n36618_, new_n36619_, new_n36620_,
    new_n36621_, new_n36622_, new_n36623_, new_n36624_, new_n36625_,
    new_n36626_, new_n36627_, new_n36628_, new_n36629_, new_n36630_,
    new_n36631_, new_n36632_, new_n36633_, new_n36634_, new_n36635_,
    new_n36636_, new_n36637_, new_n36638_, new_n36639_, new_n36640_,
    new_n36641_, new_n36642_, new_n36643_, new_n36644_, new_n36645_,
    new_n36646_, new_n36647_, new_n36648_, new_n36649_, new_n36650_,
    new_n36651_, new_n36652_, new_n36653_, new_n36654_, new_n36655_,
    new_n36656_, new_n36657_, new_n36658_, new_n36659_, new_n36660_,
    new_n36661_, new_n36662_, new_n36663_, new_n36664_, new_n36665_,
    new_n36666_, new_n36667_, new_n36668_, new_n36669_, new_n36670_,
    new_n36671_, new_n36672_, new_n36673_, new_n36674_, new_n36675_,
    new_n36676_, new_n36677_, new_n36678_, new_n36679_, new_n36680_,
    new_n36681_, new_n36682_, new_n36683_, new_n36684_, new_n36685_,
    new_n36686_, new_n36687_, new_n36688_, new_n36689_, new_n36690_,
    new_n36691_, new_n36692_, new_n36693_, new_n36694_, new_n36695_,
    new_n36696_, new_n36697_, new_n36698_, new_n36699_, new_n36700_,
    new_n36701_, new_n36702_, new_n36703_, new_n36704_, new_n36705_,
    new_n36706_, new_n36707_, new_n36708_, new_n36709_, new_n36710_,
    new_n36711_, new_n36712_, new_n36713_, new_n36714_, new_n36715_,
    new_n36716_, new_n36717_, new_n36718_, new_n36719_, new_n36720_,
    new_n36721_, new_n36722_, new_n36723_, new_n36724_, new_n36725_,
    new_n36726_, new_n36727_, new_n36728_, new_n36729_, new_n36730_,
    new_n36731_, new_n36732_, new_n36733_, new_n36734_, new_n36735_,
    new_n36736_, new_n36737_, new_n36738_, new_n36739_, new_n36740_,
    new_n36741_, new_n36742_, new_n36743_, new_n36744_, new_n36745_,
    new_n36746_, new_n36747_, new_n36748_, new_n36749_, new_n36750_,
    new_n36751_, new_n36752_, new_n36753_, new_n36754_, new_n36755_,
    new_n36756_, new_n36757_, new_n36758_, new_n36759_, new_n36760_,
    new_n36761_, new_n36762_, new_n36763_, new_n36764_, new_n36765_,
    new_n36766_, new_n36767_, new_n36768_, new_n36769_, new_n36770_,
    new_n36771_, new_n36772_, new_n36773_, new_n36774_, new_n36775_,
    new_n36776_, new_n36777_, new_n36778_, new_n36779_, new_n36780_,
    new_n36781_, new_n36782_, new_n36783_, new_n36784_, new_n36785_,
    new_n36786_, new_n36787_, new_n36788_, new_n36789_, new_n36790_,
    new_n36791_, new_n36792_, new_n36793_, new_n36794_, new_n36795_,
    new_n36796_, new_n36797_, new_n36798_, new_n36799_, new_n36800_,
    new_n36801_, new_n36802_, new_n36803_, new_n36804_, new_n36805_,
    new_n36806_, new_n36807_, new_n36808_, new_n36809_, new_n36810_,
    new_n36811_, new_n36812_, new_n36813_, new_n36814_, new_n36815_,
    new_n36816_, new_n36817_, new_n36818_, new_n36819_, new_n36820_,
    new_n36821_, new_n36822_, new_n36823_, new_n36824_, new_n36825_,
    new_n36826_, new_n36827_, new_n36828_, new_n36829_, new_n36830_,
    new_n36831_, new_n36832_, new_n36833_, new_n36834_, new_n36835_,
    new_n36836_, new_n36837_, new_n36838_, new_n36839_, new_n36840_,
    new_n36841_, new_n36842_, new_n36843_, new_n36844_, new_n36845_,
    new_n36846_, new_n36847_, new_n36848_, new_n36849_, new_n36850_,
    new_n36851_, new_n36852_, new_n36853_, new_n36854_, new_n36855_,
    new_n36856_, new_n36857_, new_n36858_, new_n36859_, new_n36860_,
    new_n36861_, new_n36862_, new_n36863_, new_n36864_, new_n36865_,
    new_n36866_, new_n36867_, new_n36868_, new_n36869_, new_n36870_,
    new_n36871_, new_n36872_, new_n36873_, new_n36874_, new_n36875_,
    new_n36876_, new_n36877_, new_n36878_, new_n36879_, new_n36880_,
    new_n36881_, new_n36882_, new_n36883_, new_n36884_, new_n36885_,
    new_n36886_, new_n36887_, new_n36888_, new_n36889_, new_n36890_,
    new_n36891_, new_n36892_, new_n36893_, new_n36894_, new_n36895_,
    new_n36896_, new_n36897_, new_n36898_, new_n36899_, new_n36900_,
    new_n36901_, new_n36902_, new_n36903_, new_n36904_, new_n36905_,
    new_n36906_, new_n36907_, new_n36908_, new_n36909_, new_n36910_,
    new_n36911_, new_n36912_, new_n36913_, new_n36914_, new_n36915_,
    new_n36916_, new_n36917_, new_n36918_, new_n36919_, new_n36920_,
    new_n36921_, new_n36922_, new_n36923_, new_n36924_, new_n36925_,
    new_n36926_, new_n36927_, new_n36928_, new_n36929_, new_n36930_,
    new_n36931_, new_n36932_, new_n36933_, new_n36934_, new_n36935_,
    new_n36936_, new_n36937_, new_n36938_, new_n36939_, new_n36940_,
    new_n36941_, new_n36942_, new_n36943_, new_n36944_, new_n36945_,
    new_n36946_, new_n36947_, new_n36948_, new_n36949_, new_n36950_,
    new_n36951_, new_n36952_, new_n36953_, new_n36954_, new_n36955_,
    new_n36956_, new_n36957_, new_n36958_, new_n36959_, new_n36960_,
    new_n36961_, new_n36962_, new_n36963_, new_n36964_, new_n36965_,
    new_n36966_, new_n36967_, new_n36968_, new_n36969_, new_n36970_,
    new_n36971_, new_n36972_, new_n36973_, new_n36974_, new_n36975_,
    new_n36976_, new_n36977_, new_n36978_, new_n36979_, new_n36980_,
    new_n36981_, new_n36982_, new_n36983_, new_n36984_, new_n36985_,
    new_n36986_, new_n36987_, new_n36988_, new_n36989_, new_n36990_,
    new_n36991_, new_n36992_, new_n36993_, new_n36994_, new_n36995_,
    new_n36996_, new_n36997_, new_n36998_, new_n36999_, new_n37000_,
    new_n37001_, new_n37002_, new_n37003_, new_n37004_, new_n37005_,
    new_n37006_, new_n37007_, new_n37008_, new_n37009_, new_n37010_,
    new_n37011_, new_n37012_, new_n37013_, new_n37014_, new_n37015_,
    new_n37016_, new_n37017_, new_n37018_, new_n37019_, new_n37020_,
    new_n37021_, new_n37022_, new_n37023_, new_n37024_, new_n37025_,
    new_n37026_, new_n37027_, new_n37028_, new_n37029_, new_n37030_,
    new_n37031_, new_n37032_, new_n37033_, new_n37034_, new_n37035_,
    new_n37036_, new_n37037_, new_n37038_, new_n37039_, new_n37040_,
    new_n37041_, new_n37042_, new_n37043_, new_n37044_, new_n37045_,
    new_n37046_, new_n37047_, new_n37048_, new_n37049_, new_n37050_,
    new_n37051_, new_n37052_, new_n37053_, new_n37054_, new_n37055_,
    new_n37056_, new_n37057_, new_n37058_, new_n37059_, new_n37060_,
    new_n37061_, new_n37062_, new_n37063_, new_n37064_, new_n37065_,
    new_n37066_, new_n37067_, new_n37068_, new_n37069_, new_n37070_,
    new_n37071_, new_n37072_, new_n37073_, new_n37074_, new_n37075_,
    new_n37076_, new_n37077_, new_n37078_, new_n37079_, new_n37080_,
    new_n37081_, new_n37082_, new_n37083_, new_n37084_, new_n37085_,
    new_n37086_, new_n37087_, new_n37088_, new_n37089_, new_n37090_,
    new_n37091_, new_n37092_, new_n37093_, new_n37094_, new_n37095_,
    new_n37096_, new_n37097_, new_n37098_, new_n37099_, new_n37100_,
    new_n37101_, new_n37102_, new_n37103_, new_n37104_, new_n37105_,
    new_n37106_, new_n37107_, new_n37108_, new_n37109_, new_n37110_,
    new_n37111_, new_n37112_, new_n37113_, new_n37114_, new_n37115_,
    new_n37116_, new_n37117_, new_n37118_, new_n37119_, new_n37120_,
    new_n37121_, new_n37122_, new_n37123_, new_n37124_, new_n37125_,
    new_n37126_, new_n37127_, new_n37128_, new_n37129_, new_n37130_,
    new_n37131_, new_n37132_, new_n37133_, new_n37134_, new_n37135_,
    new_n37136_, new_n37137_, new_n37138_, new_n37139_, new_n37140_,
    new_n37141_, new_n37142_, new_n37143_, new_n37144_, new_n37145_,
    new_n37146_, new_n37147_, new_n37148_, new_n37149_, new_n37150_,
    new_n37151_, new_n37152_, new_n37153_, new_n37154_, new_n37155_,
    new_n37156_, new_n37157_, new_n37158_, new_n37159_, new_n37160_,
    new_n37161_, new_n37162_, new_n37163_, new_n37164_, new_n37165_,
    new_n37166_, new_n37167_, new_n37168_, new_n37169_, new_n37170_,
    new_n37171_, new_n37172_, new_n37173_, new_n37174_, new_n37175_,
    new_n37176_, new_n37177_, new_n37178_, new_n37179_, new_n37180_,
    new_n37181_, new_n37182_, new_n37183_, new_n37184_, new_n37185_,
    new_n37186_, new_n37187_, new_n37188_, new_n37189_, new_n37190_,
    new_n37191_, new_n37192_, new_n37193_, new_n37194_, new_n37195_,
    new_n37196_, new_n37197_, new_n37198_, new_n37199_, new_n37200_,
    new_n37201_, new_n37202_, new_n37203_, new_n37204_, new_n37205_,
    new_n37206_, new_n37207_, new_n37208_, new_n37209_, new_n37210_,
    new_n37211_, new_n37212_, new_n37213_, new_n37214_, new_n37215_,
    new_n37216_, new_n37217_, new_n37218_, new_n37219_, new_n37220_,
    new_n37221_, new_n37222_, new_n37223_, new_n37224_, new_n37225_,
    new_n37226_, new_n37227_, new_n37228_, new_n37229_, new_n37230_,
    new_n37231_, new_n37232_, new_n37233_, new_n37234_, new_n37235_,
    new_n37236_, new_n37237_, new_n37238_, new_n37239_, new_n37240_,
    new_n37241_, new_n37242_, new_n37243_, new_n37244_, new_n37245_,
    new_n37246_, new_n37247_, new_n37248_, new_n37249_, new_n37250_,
    new_n37251_, new_n37252_, new_n37253_, new_n37254_, new_n37255_,
    new_n37256_, new_n37257_, new_n37258_, new_n37259_, new_n37260_,
    new_n37261_, new_n37262_, new_n37263_, new_n37264_, new_n37265_,
    new_n37266_, new_n37267_, new_n37268_, new_n37269_, new_n37270_,
    new_n37271_, new_n37272_, new_n37273_, new_n37274_, new_n37275_,
    new_n37276_, new_n37277_, new_n37278_, new_n37279_, new_n37280_,
    new_n37281_, new_n37282_, new_n37283_, new_n37284_, new_n37285_,
    new_n37286_, new_n37287_, new_n37288_, new_n37289_, new_n37290_,
    new_n37291_, new_n37292_, new_n37293_, new_n37294_, new_n37295_,
    new_n37296_, new_n37297_, new_n37298_, new_n37299_, new_n37300_,
    new_n37301_, new_n37302_, new_n37303_, new_n37304_, new_n37305_,
    new_n37306_, new_n37307_, new_n37308_, new_n37309_, new_n37310_,
    new_n37311_, new_n37312_, new_n37313_, new_n37314_, new_n37315_,
    new_n37316_, new_n37317_, new_n37318_, new_n37319_, new_n37320_,
    new_n37321_, new_n37322_, new_n37323_, new_n37324_, new_n37325_,
    new_n37326_, new_n37327_, new_n37328_, new_n37329_, new_n37330_,
    new_n37331_, new_n37332_, new_n37333_, new_n37334_, new_n37335_,
    new_n37336_, new_n37337_, new_n37338_, new_n37339_, new_n37340_,
    new_n37341_, new_n37342_, new_n37343_, new_n37344_, new_n37345_,
    new_n37346_, new_n37347_, new_n37348_, new_n37349_, new_n37350_,
    new_n37351_, new_n37352_, new_n37353_, new_n37354_, new_n37355_,
    new_n37356_, new_n37357_, new_n37358_, new_n37359_, new_n37360_,
    new_n37361_, new_n37362_, new_n37363_, new_n37364_, new_n37365_,
    new_n37366_, new_n37367_, new_n37368_, new_n37369_, new_n37370_,
    new_n37371_, new_n37372_, new_n37373_, new_n37374_, new_n37375_,
    new_n37376_, new_n37377_, new_n37378_, new_n37379_, new_n37380_,
    new_n37381_, new_n37382_, new_n37383_, new_n37384_, new_n37385_,
    new_n37386_, new_n37387_, new_n37388_, new_n37389_, new_n37390_,
    new_n37391_, new_n37392_, new_n37393_, new_n37394_, new_n37395_,
    new_n37396_, new_n37397_, new_n37398_, new_n37399_, new_n37400_,
    new_n37401_, new_n37402_, new_n37403_, new_n37404_, new_n37405_,
    new_n37406_, new_n37407_, new_n37408_, new_n37409_, new_n37410_,
    new_n37411_, new_n37412_, new_n37413_, new_n37414_, new_n37415_,
    new_n37416_, new_n37417_, new_n37418_, new_n37419_, new_n37420_,
    new_n37421_, new_n37422_, new_n37423_, new_n37424_, new_n37425_,
    new_n37426_, new_n37427_, new_n37428_, new_n37429_, new_n37430_,
    new_n37431_, new_n37432_, new_n37433_, new_n37434_, new_n37435_,
    new_n37436_, new_n37437_, new_n37438_, new_n37439_, new_n37440_,
    new_n37441_, new_n37442_, new_n37443_, new_n37444_, new_n37445_,
    new_n37446_, new_n37447_, new_n37448_, new_n37449_, new_n37450_,
    new_n37451_, new_n37452_, new_n37453_, new_n37454_, new_n37455_,
    new_n37456_, new_n37457_, new_n37458_, new_n37459_, new_n37460_,
    new_n37461_, new_n37462_, new_n37463_, new_n37464_, new_n37465_,
    new_n37466_, new_n37467_, new_n37468_, new_n37469_, new_n37470_,
    new_n37471_, new_n37472_, new_n37473_, new_n37474_, new_n37475_,
    new_n37476_, new_n37477_, new_n37478_, new_n37479_, new_n37480_,
    new_n37481_, new_n37482_, new_n37483_, new_n37484_, new_n37485_,
    new_n37486_, new_n37487_, new_n37488_, new_n37489_, new_n37490_,
    new_n37491_, new_n37492_, new_n37493_, new_n37494_, new_n37495_,
    new_n37496_, new_n37497_, new_n37498_, new_n37499_, new_n37500_,
    new_n37501_, new_n37502_, new_n37503_, new_n37504_, new_n37505_,
    new_n37506_, new_n37507_, new_n37508_, new_n37509_, new_n37510_,
    new_n37511_, new_n37512_, new_n37513_, new_n37514_, new_n37515_,
    new_n37516_, new_n37517_, new_n37518_, new_n37519_, new_n37520_,
    new_n37521_, new_n37522_, new_n37523_, new_n37524_, new_n37525_,
    new_n37526_, new_n37527_, new_n37528_, new_n37529_, new_n37530_,
    new_n37531_, new_n37532_, new_n37533_, new_n37534_, new_n37535_,
    new_n37536_, new_n37537_, new_n37538_, new_n37539_, new_n37540_,
    new_n37541_, new_n37542_, new_n37543_, new_n37544_, new_n37545_,
    new_n37546_, new_n37547_, new_n37548_, new_n37549_, new_n37550_,
    new_n37551_, new_n37552_, new_n37553_, new_n37554_, new_n37555_,
    new_n37556_, new_n37557_, new_n37558_, new_n37559_, new_n37560_,
    new_n37561_, new_n37562_, new_n37563_, new_n37564_, new_n37565_,
    new_n37566_, new_n37567_, new_n37568_, new_n37569_, new_n37570_,
    new_n37571_, new_n37572_, new_n37573_, new_n37574_, new_n37575_,
    new_n37576_, new_n37577_, new_n37578_, new_n37579_, new_n37580_,
    new_n37581_, new_n37582_, new_n37583_, new_n37584_, new_n37585_,
    new_n37586_, new_n37587_, new_n37588_, new_n37589_, new_n37590_,
    new_n37591_, new_n37592_, new_n37593_, new_n37594_, new_n37595_,
    new_n37596_, new_n37597_, new_n37598_, new_n37599_, new_n37600_,
    new_n37601_, new_n37602_, new_n37603_, new_n37604_, new_n37605_,
    new_n37606_, new_n37607_, new_n37608_, new_n37609_, new_n37610_,
    new_n37611_, new_n37612_, new_n37613_, new_n37614_, new_n37615_,
    new_n37616_, new_n37617_, new_n37618_, new_n37619_, new_n37620_,
    new_n37621_, new_n37622_, new_n37623_, new_n37624_, new_n37625_,
    new_n37626_, new_n37627_, new_n37628_, new_n37629_, new_n37630_,
    new_n37631_, new_n37632_, new_n37633_, new_n37634_, new_n37635_,
    new_n37636_, new_n37637_, new_n37638_, new_n37639_, new_n37640_,
    new_n37641_, new_n37642_, new_n37643_, new_n37644_, new_n37645_,
    new_n37646_, new_n37647_, new_n37648_, new_n37649_, new_n37650_,
    new_n37651_, new_n37652_, new_n37653_, new_n37654_, new_n37655_,
    new_n37656_, new_n37657_, new_n37658_, new_n37659_, new_n37660_,
    new_n37661_, new_n37662_, new_n37663_, new_n37664_, new_n37665_,
    new_n37666_, new_n37667_, new_n37668_, new_n37669_, new_n37670_,
    new_n37671_, new_n37672_, new_n37673_, new_n37674_, new_n37675_,
    new_n37676_, new_n37677_, new_n37678_, new_n37679_, new_n37680_,
    new_n37681_, new_n37682_, new_n37683_, new_n37684_, new_n37685_,
    new_n37686_, new_n37687_, new_n37688_, new_n37689_, new_n37690_,
    new_n37691_, new_n37692_, new_n37693_, new_n37694_, new_n37695_,
    new_n37696_, new_n37697_, new_n37698_, new_n37699_, new_n37700_,
    new_n37701_, new_n37702_, new_n37703_, new_n37704_, new_n37705_,
    new_n37706_, new_n37707_, new_n37708_, new_n37709_, new_n37710_,
    new_n37711_, new_n37712_, new_n37713_, new_n37714_, new_n37715_,
    new_n37716_, new_n37717_, new_n37718_, new_n37719_, new_n37720_,
    new_n37721_, new_n37722_, new_n37723_, new_n37724_, new_n37725_,
    new_n37726_, new_n37727_, new_n37728_, new_n37729_, new_n37730_,
    new_n37731_, new_n37732_, new_n37733_, new_n37734_, new_n37735_,
    new_n37736_, new_n37737_, new_n37738_, new_n37739_, new_n37740_,
    new_n37741_, new_n37742_, new_n37743_, new_n37744_, new_n37745_,
    new_n37746_, new_n37747_, new_n37748_, new_n37749_, new_n37750_,
    new_n37751_, new_n37752_, new_n37753_, new_n37754_, new_n37755_,
    new_n37756_, new_n37757_, new_n37758_, new_n37759_, new_n37760_,
    new_n37761_, new_n37762_, new_n37763_, new_n37764_, new_n37765_,
    new_n37766_, new_n37767_, new_n37768_, new_n37769_, new_n37770_,
    new_n37771_, new_n37772_, new_n37773_, new_n37774_, new_n37775_,
    new_n37776_, new_n37777_, new_n37778_, new_n37779_, new_n37780_,
    new_n37781_, new_n37782_, new_n37783_, new_n37784_, new_n37785_,
    new_n37786_, new_n37787_, new_n37788_, new_n37789_, new_n37790_,
    new_n37791_, new_n37792_, new_n37793_, new_n37794_, new_n37795_,
    new_n37796_, new_n37797_, new_n37798_, new_n37799_, new_n37800_,
    new_n37801_, new_n37802_, new_n37803_, new_n37804_, new_n37805_,
    new_n37806_, new_n37807_, new_n37808_, new_n37809_, new_n37810_,
    new_n37811_, new_n37812_, new_n37813_, new_n37814_, new_n37815_,
    new_n37816_, new_n37817_, new_n37818_, new_n37819_, new_n37820_,
    new_n37821_, new_n37822_, new_n37823_, new_n37824_, new_n37825_,
    new_n37826_, new_n37827_, new_n37828_, new_n37829_, new_n37830_,
    new_n37831_, new_n37832_, new_n37833_, new_n37834_, new_n37835_,
    new_n37836_, new_n37837_, new_n37838_, new_n37839_, new_n37840_,
    new_n37841_, new_n37842_, new_n37843_, new_n37844_, new_n37845_,
    new_n37846_, new_n37847_, new_n37848_, new_n37849_, new_n37850_,
    new_n37851_, new_n37852_, new_n37853_, new_n37854_, new_n37855_,
    new_n37856_, new_n37857_, new_n37858_, new_n37859_, new_n37860_,
    new_n37861_, new_n37862_, new_n37863_, new_n37864_, new_n37865_,
    new_n37866_, new_n37867_, new_n37868_, new_n37869_, new_n37870_,
    new_n37871_, new_n37872_, new_n37873_, new_n37874_, new_n37875_,
    new_n37876_, new_n37877_, new_n37878_, new_n37879_, new_n37880_,
    new_n37881_, new_n37882_, new_n37883_, new_n37884_, new_n37885_,
    new_n37886_, new_n37887_, new_n37888_, new_n37889_, new_n37890_,
    new_n37891_, new_n37892_, new_n37893_, new_n37894_, new_n37895_,
    new_n37896_, new_n37897_, new_n37898_, new_n37899_, new_n37900_,
    new_n37901_, new_n37902_, new_n37903_, new_n37904_, new_n37905_,
    new_n37906_, new_n37907_, new_n37908_, new_n37909_, new_n37910_,
    new_n37911_, new_n37912_, new_n37913_, new_n37914_, new_n37915_,
    new_n37916_, new_n37917_, new_n37918_, new_n37919_, new_n37920_,
    new_n37921_, new_n37922_, new_n37923_, new_n37924_, new_n37925_,
    new_n37926_, new_n37927_, new_n37928_, new_n37929_, new_n37930_,
    new_n37931_, new_n37932_, new_n37933_, new_n37934_, new_n37935_,
    new_n37936_, new_n37937_, new_n37938_, new_n37939_, new_n37940_,
    new_n37941_, new_n37942_, new_n37943_, new_n37944_, new_n37945_,
    new_n37946_, new_n37947_, new_n37948_, new_n37949_, new_n37950_,
    new_n37951_, new_n37952_, new_n37953_, new_n37954_, new_n37955_,
    new_n37956_, new_n37957_, new_n37958_, new_n37959_, new_n37960_,
    new_n37961_, new_n37962_, new_n37963_, new_n37964_, new_n37965_,
    new_n37966_, new_n37967_, new_n37968_, new_n37969_, new_n37970_,
    new_n37971_, new_n37972_, new_n37973_, new_n37974_, new_n37975_,
    new_n37976_, new_n37977_, new_n37978_, new_n37979_, new_n37980_,
    new_n37981_, new_n37982_, new_n37983_, new_n37984_, new_n37985_,
    new_n37986_, new_n37987_, new_n37988_, new_n37989_, new_n37990_,
    new_n37991_, new_n37992_, new_n37993_, new_n37994_, new_n37995_,
    new_n37996_, new_n37997_, new_n37998_, new_n37999_, new_n38000_,
    new_n38001_, new_n38002_, new_n38003_, new_n38004_, new_n38005_,
    new_n38006_, new_n38007_, new_n38008_, new_n38009_, new_n38010_,
    new_n38011_, new_n38012_, new_n38013_, new_n38014_, new_n38015_,
    new_n38016_, new_n38017_, new_n38018_, new_n38019_, new_n38020_,
    new_n38021_, new_n38022_, new_n38023_, new_n38024_, new_n38025_,
    new_n38026_, new_n38027_, new_n38028_, new_n38029_, new_n38030_,
    new_n38031_, new_n38032_, new_n38033_, new_n38034_, new_n38035_,
    new_n38036_, new_n38037_, new_n38038_, new_n38039_, new_n38040_,
    new_n38041_, new_n38042_, new_n38043_, new_n38044_, new_n38045_,
    new_n38046_, new_n38047_, new_n38048_, new_n38049_, new_n38050_,
    new_n38051_, new_n38052_, new_n38053_, new_n38054_, new_n38055_,
    new_n38056_, new_n38057_, new_n38058_, new_n38059_, new_n38060_,
    new_n38061_, new_n38062_, new_n38063_, new_n38064_, new_n38065_,
    new_n38066_, new_n38067_, new_n38068_, new_n38069_, new_n38070_,
    new_n38071_, new_n38072_, new_n38073_, new_n38074_, new_n38075_,
    new_n38076_, new_n38077_, new_n38078_, new_n38079_, new_n38080_,
    new_n38081_, new_n38082_, new_n38083_, new_n38084_, new_n38085_,
    new_n38086_, new_n38087_, new_n38088_, new_n38089_, new_n38090_,
    new_n38091_, new_n38092_, new_n38093_, new_n38094_, new_n38095_,
    new_n38096_, new_n38097_, new_n38098_, new_n38099_, new_n38100_,
    new_n38101_, new_n38102_, new_n38103_, new_n38104_, new_n38105_,
    new_n38106_, new_n38107_, new_n38108_, new_n38109_, new_n38110_,
    new_n38111_, new_n38112_, new_n38113_, new_n38114_, new_n38115_,
    new_n38116_, new_n38117_, new_n38118_, new_n38119_, new_n38120_,
    new_n38121_, new_n38122_, new_n38123_, new_n38124_, new_n38125_,
    new_n38126_, new_n38127_, new_n38128_, new_n38129_, new_n38130_,
    new_n38131_, new_n38132_, new_n38133_, new_n38134_, new_n38135_,
    new_n38136_, new_n38137_, new_n38138_, new_n38139_, new_n38140_,
    new_n38141_, new_n38142_, new_n38143_, new_n38144_, new_n38145_,
    new_n38146_, new_n38147_, new_n38148_, new_n38149_, new_n38150_,
    new_n38151_, new_n38152_, new_n38153_, new_n38154_, new_n38155_,
    new_n38156_, new_n38157_, new_n38158_, new_n38159_, new_n38160_,
    new_n38161_, new_n38162_, new_n38163_, new_n38164_, new_n38165_,
    new_n38166_, new_n38167_, new_n38168_, new_n38169_, new_n38170_,
    new_n38171_, new_n38172_, new_n38173_, new_n38174_, new_n38175_,
    new_n38176_, new_n38177_, new_n38178_, new_n38179_, new_n38180_,
    new_n38181_, new_n38182_, new_n38183_, new_n38184_, new_n38185_,
    new_n38186_, new_n38187_, new_n38188_, new_n38189_, new_n38190_,
    new_n38191_, new_n38192_, new_n38193_, new_n38194_, new_n38195_,
    new_n38196_, new_n38197_, new_n38198_, new_n38199_, new_n38200_,
    new_n38201_, new_n38202_, new_n38203_, new_n38204_, new_n38205_,
    new_n38206_, new_n38207_, new_n38208_, new_n38209_, new_n38210_,
    new_n38211_, new_n38212_, new_n38213_, new_n38214_, new_n38215_,
    new_n38216_, new_n38217_, new_n38218_, new_n38219_, new_n38220_,
    new_n38221_, new_n38222_, new_n38223_, new_n38224_, new_n38225_,
    new_n38226_, new_n38227_, new_n38228_, new_n38229_, new_n38230_,
    new_n38231_, new_n38232_, new_n38233_, new_n38234_, new_n38235_,
    new_n38236_, new_n38237_, new_n38238_, new_n38239_, new_n38240_,
    new_n38241_, new_n38242_, new_n38243_, new_n38244_, new_n38245_,
    new_n38246_, new_n38247_, new_n38248_, new_n38249_, new_n38250_,
    new_n38251_, new_n38252_, new_n38253_, new_n38254_, new_n38255_,
    new_n38256_, new_n38257_, new_n38258_, new_n38259_, new_n38260_,
    new_n38261_, new_n38262_, new_n38263_, new_n38264_, new_n38265_,
    new_n38266_, new_n38267_, new_n38268_, new_n38269_, new_n38270_,
    new_n38271_, new_n38272_, new_n38273_, new_n38274_, new_n38275_,
    new_n38276_, new_n38277_, new_n38278_, new_n38279_, new_n38280_,
    new_n38281_, new_n38282_, new_n38283_, new_n38284_, new_n38285_,
    new_n38286_, new_n38287_, new_n38288_, new_n38289_, new_n38290_,
    new_n38291_, new_n38292_, new_n38293_, new_n38294_, new_n38295_,
    new_n38296_, new_n38297_, new_n38298_, new_n38299_, new_n38300_,
    new_n38301_, new_n38302_, new_n38303_, new_n38304_, new_n38305_,
    new_n38306_, new_n38307_, new_n38308_, new_n38309_, new_n38310_,
    new_n38311_, new_n38312_, new_n38313_, new_n38314_, new_n38315_,
    new_n38316_, new_n38317_, new_n38318_, new_n38319_, new_n38320_,
    new_n38321_, new_n38322_, new_n38323_, new_n38324_, new_n38325_,
    new_n38326_, new_n38327_, new_n38328_, new_n38329_, new_n38330_,
    new_n38331_, new_n38332_, new_n38333_, new_n38334_, new_n38335_,
    new_n38336_, new_n38337_, new_n38338_, new_n38339_, new_n38340_,
    new_n38341_, new_n38342_, new_n38343_, new_n38344_, new_n38345_,
    new_n38346_, new_n38347_, new_n38348_, new_n38349_, new_n38350_,
    new_n38351_, new_n38352_, new_n38353_, new_n38354_, new_n38355_,
    new_n38356_, new_n38357_, new_n38358_, new_n38359_, new_n38360_,
    new_n38361_, new_n38362_, new_n38363_, new_n38364_, new_n38365_,
    new_n38366_, new_n38367_, new_n38368_, new_n38369_, new_n38370_,
    new_n38371_, new_n38372_, new_n38373_, new_n38374_, new_n38375_,
    new_n38376_, new_n38377_, new_n38378_, new_n38379_, new_n38380_,
    new_n38381_, new_n38382_, new_n38383_, new_n38384_, new_n38385_,
    new_n38386_, new_n38387_, new_n38388_, new_n38389_, new_n38390_,
    new_n38391_, new_n38392_, new_n38393_, new_n38394_, new_n38395_,
    new_n38396_, new_n38397_, new_n38398_, new_n38399_, new_n38400_,
    new_n38401_, new_n38402_, new_n38403_, new_n38404_, new_n38405_,
    new_n38406_, new_n38407_, new_n38408_, new_n38409_, new_n38410_,
    new_n38411_, new_n38412_, new_n38413_, new_n38414_, new_n38415_,
    new_n38416_, new_n38417_, new_n38418_, new_n38419_, new_n38420_,
    new_n38421_, new_n38422_, new_n38423_, new_n38424_, new_n38425_,
    new_n38426_, new_n38427_, new_n38428_, new_n38429_, new_n38430_,
    new_n38431_, new_n38432_, new_n38433_, new_n38434_, new_n38435_,
    new_n38436_, new_n38437_, new_n38438_, new_n38439_, new_n38440_,
    new_n38441_, new_n38442_, new_n38443_, new_n38444_, new_n38445_,
    new_n38446_, new_n38447_, new_n38448_, new_n38449_, new_n38450_,
    new_n38451_, new_n38452_, new_n38453_, new_n38454_, new_n38455_,
    new_n38456_, new_n38457_, new_n38458_, new_n38459_, new_n38460_,
    new_n38461_, new_n38462_, new_n38463_, new_n38464_, new_n38465_,
    new_n38466_, new_n38467_, new_n38468_, new_n38469_, new_n38470_,
    new_n38471_, new_n38472_, new_n38473_, new_n38474_, new_n38475_,
    new_n38476_, new_n38477_, new_n38478_, new_n38479_, new_n38480_,
    new_n38481_, new_n38482_, new_n38483_, new_n38484_, new_n38485_,
    new_n38486_, new_n38487_, new_n38488_, new_n38489_, new_n38490_,
    new_n38491_, new_n38492_, new_n38493_, new_n38494_, new_n38495_,
    new_n38496_, new_n38497_, new_n38498_, new_n38499_, new_n38500_,
    new_n38501_, new_n38502_, new_n38503_, new_n38504_, new_n38505_,
    new_n38506_, new_n38507_, new_n38508_, new_n38509_, new_n38510_,
    new_n38511_, new_n38512_, new_n38513_, new_n38514_, new_n38515_,
    new_n38516_, new_n38517_, new_n38518_, new_n38519_, new_n38520_,
    new_n38521_, new_n38522_, new_n38523_, new_n38524_, new_n38525_,
    new_n38526_, new_n38527_, new_n38528_, new_n38529_, new_n38530_,
    new_n38531_, new_n38532_, new_n38533_, new_n38534_, new_n38535_,
    new_n38536_, new_n38537_, new_n38538_, new_n38539_, new_n38540_,
    new_n38541_, new_n38542_, new_n38543_, new_n38544_, new_n38545_,
    new_n38546_, new_n38547_, new_n38548_, new_n38549_, new_n38550_,
    new_n38551_, new_n38552_, new_n38553_, new_n38554_, new_n38555_,
    new_n38556_, new_n38557_, new_n38558_, new_n38559_, new_n38560_,
    new_n38561_, new_n38562_, new_n38563_, new_n38564_, new_n38565_,
    new_n38566_, new_n38567_, new_n38568_, new_n38569_, new_n38570_,
    new_n38571_, new_n38572_, new_n38573_, new_n38574_, new_n38575_,
    new_n38576_, new_n38577_, new_n38578_, new_n38579_, new_n38580_,
    new_n38581_, new_n38582_, new_n38583_, new_n38584_, new_n38585_,
    new_n38586_, new_n38587_, new_n38588_, new_n38589_, new_n38590_,
    new_n38591_, new_n38592_, new_n38593_, new_n38594_, new_n38595_,
    new_n38596_, new_n38597_, new_n38598_, new_n38599_, new_n38600_,
    new_n38601_, new_n38602_, new_n38603_, new_n38604_, new_n38605_,
    new_n38606_, new_n38607_, new_n38608_, new_n38609_, new_n38610_,
    new_n38611_, new_n38612_, new_n38613_, new_n38614_, new_n38615_,
    new_n38616_, new_n38617_, new_n38618_, new_n38619_, new_n38620_,
    new_n38621_, new_n38622_, new_n38623_, new_n38624_, new_n38625_,
    new_n38626_, new_n38627_, new_n38628_, new_n38629_, new_n38630_,
    new_n38631_, new_n38632_, new_n38633_, new_n38634_, new_n38635_,
    new_n38636_, new_n38637_, new_n38638_, new_n38639_, new_n38640_,
    new_n38641_, new_n38642_, new_n38643_, new_n38644_, new_n38645_,
    new_n38646_, new_n38647_, new_n38648_, new_n38649_, new_n38650_,
    new_n38651_, new_n38652_, new_n38653_, new_n38654_, new_n38655_,
    new_n38656_, new_n38657_, new_n38658_, new_n38659_, new_n38660_,
    new_n38661_, new_n38662_, new_n38663_, new_n38664_, new_n38665_,
    new_n38666_, new_n38667_, new_n38668_, new_n38669_, new_n38670_,
    new_n38671_, new_n38672_, new_n38673_, new_n38674_, new_n38675_,
    new_n38676_, new_n38677_, new_n38678_, new_n38679_, new_n38680_,
    new_n38681_, new_n38682_, new_n38683_, new_n38684_, new_n38685_,
    new_n38686_, new_n38687_, new_n38688_, new_n38689_, new_n38690_,
    new_n38691_, new_n38692_, new_n38693_, new_n38694_, new_n38695_,
    new_n38696_, new_n38697_, new_n38698_, new_n38699_, new_n38700_,
    new_n38701_, new_n38702_, new_n38703_, new_n38704_, new_n38705_,
    new_n38706_, new_n38707_, new_n38708_, new_n38709_, new_n38710_,
    new_n38711_, new_n38712_, new_n38713_, new_n38714_, new_n38715_,
    new_n38716_, new_n38717_, new_n38718_, new_n38719_, new_n38720_,
    new_n38721_, new_n38722_, new_n38723_, new_n38724_, new_n38725_,
    new_n38726_, new_n38727_, new_n38728_, new_n38729_, new_n38730_,
    new_n38731_, new_n38732_, new_n38733_, new_n38734_, new_n38735_,
    new_n38736_, new_n38737_, new_n38738_, new_n38739_, new_n38740_,
    new_n38741_, new_n38742_, new_n38743_, new_n38744_, new_n38745_,
    new_n38746_, new_n38747_, new_n38748_, new_n38749_, new_n38750_,
    new_n38751_, new_n38752_, new_n38753_, new_n38754_, new_n38755_,
    new_n38756_, new_n38757_, new_n38758_, new_n38759_, new_n38760_,
    new_n38761_, new_n38762_, new_n38763_, new_n38764_, new_n38765_,
    new_n38766_, new_n38767_, new_n38768_, new_n38769_, new_n38770_,
    new_n38771_, new_n38772_, new_n38773_, new_n38774_, new_n38775_,
    new_n38776_, new_n38777_, new_n38778_, new_n38779_, new_n38780_,
    new_n38781_, new_n38782_, new_n38783_, new_n38784_, new_n38785_,
    new_n38786_, new_n38787_, new_n38788_, new_n38789_, new_n38790_,
    new_n38791_, new_n38792_, new_n38793_, new_n38794_, new_n38795_,
    new_n38796_, new_n38797_, new_n38798_, new_n38799_, new_n38800_,
    new_n38801_, new_n38802_, new_n38803_, new_n38804_, new_n38805_,
    new_n38806_, new_n38807_, new_n38808_, new_n38809_, new_n38810_,
    new_n38811_, new_n38812_, new_n38813_, new_n38814_, new_n38815_,
    new_n38816_, new_n38817_, new_n38818_, new_n38819_, new_n38820_,
    new_n38821_, new_n38822_, new_n38823_, new_n38824_, new_n38825_,
    new_n38826_, new_n38827_, new_n38828_, new_n38829_, new_n38830_,
    new_n38831_, new_n38832_, new_n38833_, new_n38834_, new_n38835_,
    new_n38836_, new_n38837_, new_n38838_, new_n38839_, new_n38840_,
    new_n38841_, new_n38842_, new_n38843_, new_n38844_, new_n38845_,
    new_n38846_, new_n38847_, new_n38848_, new_n38849_, new_n38850_,
    new_n38851_, new_n38852_, new_n38853_, new_n38854_, new_n38855_,
    new_n38856_, new_n38857_, new_n38858_, new_n38859_, new_n38860_,
    new_n38861_, new_n38862_, new_n38863_, new_n38864_, new_n38865_,
    new_n38866_, new_n38867_, new_n38868_, new_n38869_, new_n38870_,
    new_n38871_, new_n38872_, new_n38873_, new_n38874_, new_n38875_,
    new_n38876_, new_n38877_, new_n38878_, new_n38879_, new_n38880_,
    new_n38881_, new_n38882_, new_n38883_, new_n38884_, new_n38885_,
    new_n38886_, new_n38887_, new_n38888_, new_n38889_, new_n38890_,
    new_n38891_, new_n38892_, new_n38893_, new_n38894_, new_n38895_,
    new_n38896_, new_n38897_, new_n38898_, new_n38899_, new_n38900_,
    new_n38901_, new_n38902_, new_n38903_, new_n38904_, new_n38905_,
    new_n38906_, new_n38907_, new_n38908_, new_n38909_, new_n38910_,
    new_n38911_, new_n38912_, new_n38913_, new_n38914_, new_n38915_,
    new_n38916_, new_n38917_, new_n38918_, new_n38919_, new_n38920_,
    new_n38921_, new_n38922_, new_n38923_, new_n38924_, new_n38925_,
    new_n38926_, new_n38927_, new_n38928_, new_n38929_, new_n38930_,
    new_n38931_, new_n38932_, new_n38933_, new_n38934_, new_n38935_,
    new_n38936_, new_n38937_, new_n38938_, new_n38939_, new_n38940_,
    new_n38941_, new_n38942_, new_n38943_, new_n38944_, new_n38945_,
    new_n38946_, new_n38947_, new_n38948_, new_n38949_, new_n38950_,
    new_n38951_, new_n38952_, new_n38953_, new_n38954_, new_n38955_,
    new_n38956_, new_n38957_, new_n38958_, new_n38959_, new_n38960_,
    new_n38961_, new_n38962_, new_n38963_, new_n38964_, new_n38965_,
    new_n38966_, new_n38967_, new_n38968_, new_n38969_, new_n38970_,
    new_n38971_, new_n38972_, new_n38973_, new_n38974_, new_n38975_,
    new_n38976_, new_n38977_, new_n38978_, new_n38979_, new_n38980_,
    new_n38981_, new_n38982_, new_n38983_, new_n38984_, new_n38985_,
    new_n38986_, new_n38987_, new_n38988_, new_n38989_, new_n38990_,
    new_n38991_, new_n38992_, new_n38993_, new_n38994_, new_n38995_,
    new_n38996_, new_n38997_, new_n38998_, new_n38999_, new_n39000_,
    new_n39001_, new_n39002_, new_n39003_, new_n39004_, new_n39005_,
    new_n39006_, new_n39007_, new_n39008_, new_n39009_, new_n39010_,
    new_n39011_, new_n39012_, new_n39013_, new_n39014_, new_n39015_,
    new_n39016_, new_n39017_, new_n39018_, new_n39019_, new_n39020_,
    new_n39021_, new_n39022_, new_n39023_, new_n39024_, new_n39025_,
    new_n39026_, new_n39027_, new_n39028_, new_n39029_, new_n39030_,
    new_n39031_, new_n39032_, new_n39033_, new_n39034_, new_n39035_,
    new_n39036_, new_n39037_, new_n39038_, new_n39039_, new_n39040_,
    new_n39041_, new_n39042_, new_n39043_, new_n39044_, new_n39045_,
    new_n39046_, new_n39047_, new_n39048_, new_n39049_, new_n39050_,
    new_n39051_, new_n39052_, new_n39053_, new_n39054_, new_n39055_,
    new_n39056_, new_n39057_, new_n39058_, new_n39059_, new_n39060_,
    new_n39061_, new_n39062_, new_n39063_, new_n39064_, new_n39065_,
    new_n39066_, new_n39067_, new_n39068_, new_n39069_, new_n39070_,
    new_n39071_, new_n39072_, new_n39073_, new_n39074_, new_n39075_,
    new_n39076_, new_n39077_, new_n39078_, new_n39079_, new_n39080_,
    new_n39081_, new_n39082_, new_n39083_, new_n39084_, new_n39085_,
    new_n39086_, new_n39087_, new_n39088_, new_n39089_, new_n39090_,
    new_n39091_, new_n39092_, new_n39093_, new_n39094_, new_n39095_,
    new_n39096_, new_n39097_, new_n39098_, new_n39099_, new_n39100_,
    new_n39101_, new_n39102_, new_n39103_, new_n39104_, new_n39105_,
    new_n39106_, new_n39107_, new_n39108_, new_n39109_, new_n39110_,
    new_n39111_, new_n39112_, new_n39113_, new_n39114_, new_n39115_,
    new_n39116_, new_n39117_, new_n39118_, new_n39119_, new_n39120_,
    new_n39121_, new_n39122_, new_n39123_, new_n39124_, new_n39125_,
    new_n39126_, new_n39127_, new_n39128_, new_n39129_, new_n39130_,
    new_n39131_, new_n39132_, new_n39133_, new_n39134_, new_n39135_,
    new_n39136_, new_n39137_, new_n39138_, new_n39139_, new_n39140_,
    new_n39141_, new_n39142_, new_n39143_, new_n39144_, new_n39145_,
    new_n39146_, new_n39147_, new_n39148_, new_n39149_, new_n39150_,
    new_n39151_, new_n39152_, new_n39153_, new_n39154_, new_n39155_,
    new_n39156_, new_n39157_, new_n39158_, new_n39159_, new_n39160_,
    new_n39161_, new_n39162_, new_n39163_, new_n39164_, new_n39165_,
    new_n39166_, new_n39167_, new_n39168_, new_n39169_, new_n39170_,
    new_n39171_, new_n39172_, new_n39173_, new_n39174_, new_n39175_,
    new_n39176_, new_n39177_, new_n39178_, new_n39179_, new_n39180_,
    new_n39181_, new_n39182_, new_n39183_, new_n39184_, new_n39185_,
    new_n39186_, new_n39187_, new_n39188_, new_n39189_, new_n39190_,
    new_n39191_, new_n39192_, new_n39193_, new_n39194_, new_n39195_,
    new_n39196_, new_n39197_, new_n39198_, new_n39199_, new_n39200_,
    new_n39201_, new_n39202_, new_n39203_, new_n39204_, new_n39205_,
    new_n39206_, new_n39207_, new_n39208_, new_n39209_, new_n39210_,
    new_n39211_, new_n39212_, new_n39213_, new_n39214_, new_n39215_,
    new_n39216_, new_n39217_, new_n39218_, new_n39219_, new_n39220_,
    new_n39221_, new_n39222_, new_n39223_, new_n39224_, new_n39225_,
    new_n39226_, new_n39227_, new_n39228_, new_n39229_, new_n39230_,
    new_n39231_, new_n39232_, new_n39233_, new_n39234_, new_n39235_,
    new_n39236_, new_n39237_, new_n39238_, new_n39239_, new_n39240_,
    new_n39241_, new_n39242_, new_n39243_, new_n39244_, new_n39245_,
    new_n39246_, new_n39247_, new_n39248_, new_n39249_, new_n39250_,
    new_n39251_, new_n39252_, new_n39253_, new_n39254_, new_n39255_,
    new_n39256_, new_n39257_, new_n39258_, new_n39259_, new_n39260_,
    new_n39261_, new_n39262_, new_n39263_, new_n39264_, new_n39265_,
    new_n39266_, new_n39267_, new_n39268_, new_n39269_, new_n39270_,
    new_n39271_, new_n39272_, new_n39273_, new_n39274_, new_n39275_,
    new_n39276_, new_n39277_, new_n39278_, new_n39279_, new_n39280_,
    new_n39281_, new_n39282_, new_n39283_, new_n39284_, new_n39285_,
    new_n39286_, new_n39287_, new_n39288_, new_n39289_, new_n39290_,
    new_n39291_, new_n39292_, new_n39293_, new_n39294_, new_n39295_,
    new_n39296_, new_n39297_, new_n39298_, new_n39299_, new_n39300_,
    new_n39301_, new_n39302_, new_n39303_, new_n39304_, new_n39305_,
    new_n39306_, new_n39307_, new_n39308_, new_n39309_, new_n39310_,
    new_n39311_, new_n39312_, new_n39313_, new_n39314_, new_n39315_,
    new_n39316_, new_n39317_, new_n39318_, new_n39319_, new_n39320_,
    new_n39321_, new_n39322_, new_n39323_, new_n39324_, new_n39325_,
    new_n39326_, new_n39327_, new_n39328_, new_n39329_, new_n39330_,
    new_n39331_, new_n39332_, new_n39333_, new_n39334_, new_n39335_,
    new_n39336_, new_n39337_, new_n39338_, new_n39339_, new_n39340_,
    new_n39341_, new_n39342_, new_n39343_, new_n39344_, new_n39345_,
    new_n39346_, new_n39347_, new_n39348_, new_n39349_, new_n39350_,
    new_n39351_, new_n39352_, new_n39353_, new_n39354_, new_n39355_,
    new_n39356_, new_n39357_, new_n39358_, new_n39359_, new_n39360_,
    new_n39361_, new_n39362_, new_n39363_, new_n39364_, new_n39365_,
    new_n39366_, new_n39367_, new_n39368_, new_n39369_, new_n39370_,
    new_n39371_, new_n39372_, new_n39373_, new_n39374_, new_n39375_,
    new_n39376_, new_n39377_, new_n39378_, new_n39379_, new_n39380_,
    new_n39381_, new_n39382_, new_n39383_, new_n39384_, new_n39385_,
    new_n39386_, new_n39387_, new_n39388_, new_n39389_, new_n39390_,
    new_n39391_, new_n39392_, new_n39393_, new_n39394_, new_n39395_,
    new_n39396_, new_n39397_, new_n39398_, new_n39399_, new_n39400_,
    new_n39401_, new_n39402_, new_n39403_, new_n39404_, new_n39405_,
    new_n39406_, new_n39407_, new_n39408_, new_n39409_, new_n39410_,
    new_n39411_, new_n39412_, new_n39413_, new_n39414_, new_n39415_,
    new_n39416_, new_n39417_, new_n39418_, new_n39419_, new_n39420_,
    new_n39421_, new_n39422_, new_n39423_, new_n39424_, new_n39425_,
    new_n39426_, new_n39427_, new_n39428_, new_n39429_, new_n39430_,
    new_n39431_, new_n39432_, new_n39433_, new_n39434_, new_n39435_,
    new_n39436_, new_n39437_, new_n39438_, new_n39439_, new_n39440_,
    new_n39441_, new_n39442_, new_n39443_, new_n39444_, new_n39445_,
    new_n39446_, new_n39447_, new_n39448_, new_n39449_, new_n39450_,
    new_n39451_, new_n39452_, new_n39453_, new_n39454_, new_n39455_,
    new_n39456_, new_n39457_, new_n39458_, new_n39459_, new_n39460_,
    new_n39461_, new_n39462_, new_n39463_, new_n39464_, new_n39465_,
    new_n39466_, new_n39467_, new_n39468_, new_n39469_, new_n39470_,
    new_n39471_, new_n39472_, new_n39473_, new_n39474_, new_n39475_,
    new_n39476_, new_n39477_, new_n39478_, new_n39479_, new_n39480_,
    new_n39481_, new_n39482_, new_n39483_, new_n39484_, new_n39485_,
    new_n39486_, new_n39487_, new_n39488_, new_n39489_, new_n39490_,
    new_n39491_, new_n39492_, new_n39493_, new_n39494_, new_n39495_,
    new_n39496_, new_n39497_, new_n39498_, new_n39499_, new_n39500_,
    new_n39501_, new_n39502_, new_n39503_, new_n39504_, new_n39505_,
    new_n39506_, new_n39507_, new_n39508_, new_n39509_, new_n39510_,
    new_n39511_, new_n39512_, new_n39513_, new_n39514_, new_n39515_,
    new_n39516_, new_n39517_, new_n39518_, new_n39519_, new_n39520_,
    new_n39521_, new_n39522_, new_n39523_, new_n39524_, new_n39525_,
    new_n39526_, new_n39527_, new_n39528_, new_n39529_, new_n39530_,
    new_n39531_, new_n39532_, new_n39533_, new_n39534_, new_n39535_,
    new_n39536_, new_n39537_, new_n39538_, new_n39539_, new_n39540_,
    new_n39541_, new_n39542_, new_n39543_, new_n39544_, new_n39545_,
    new_n39546_, new_n39547_, new_n39548_, new_n39549_, new_n39550_,
    new_n39551_, new_n39552_, new_n39553_, new_n39554_, new_n39555_,
    new_n39556_, new_n39557_, new_n39558_, new_n39559_, new_n39560_,
    new_n39561_, new_n39562_, new_n39563_, new_n39564_, new_n39565_,
    new_n39566_, new_n39567_, new_n39568_, new_n39569_, new_n39570_,
    new_n39571_, new_n39572_, new_n39573_, new_n39574_, new_n39575_,
    new_n39576_, new_n39577_, new_n39578_, new_n39579_, new_n39580_,
    new_n39581_, new_n39582_, new_n39583_, new_n39584_, new_n39585_,
    new_n39586_, new_n39587_, new_n39588_, new_n39589_, new_n39590_,
    new_n39591_, new_n39592_, new_n39593_, new_n39594_, new_n39595_,
    new_n39596_, new_n39597_, new_n39598_, new_n39599_, new_n39600_,
    new_n39601_, new_n39602_, new_n39603_, new_n39604_, new_n39605_,
    new_n39606_, new_n39607_, new_n39608_, new_n39609_, new_n39610_,
    new_n39611_, new_n39612_, new_n39613_, new_n39614_, new_n39615_,
    new_n39616_, new_n39617_, new_n39618_, new_n39619_, new_n39620_,
    new_n39621_, new_n39622_, new_n39623_, new_n39624_, new_n39625_,
    new_n39626_, new_n39627_, new_n39628_, new_n39629_, new_n39630_,
    new_n39631_, new_n39632_, new_n39633_, new_n39634_, new_n39635_,
    new_n39636_, new_n39637_, new_n39638_, new_n39639_, new_n39640_,
    new_n39641_, new_n39642_, new_n39643_, new_n39644_, new_n39645_,
    new_n39646_, new_n39647_, new_n39648_, new_n39649_, new_n39650_,
    new_n39651_, new_n39652_, new_n39653_, new_n39654_, new_n39655_,
    new_n39656_, new_n39657_, new_n39658_, new_n39659_, new_n39660_,
    new_n39661_, new_n39662_, new_n39663_, new_n39664_, new_n39665_,
    new_n39666_, new_n39667_, new_n39668_, new_n39669_, new_n39670_,
    new_n39671_, new_n39672_, new_n39673_, new_n39674_, new_n39675_,
    new_n39676_, new_n39677_, new_n39678_, new_n39679_, new_n39680_,
    new_n39681_, new_n39682_, new_n39683_, new_n39684_, new_n39685_,
    new_n39686_, new_n39687_, new_n39688_, new_n39689_, new_n39690_,
    new_n39691_, new_n39692_, new_n39693_, new_n39694_, new_n39695_,
    new_n39696_, new_n39697_, new_n39698_, new_n39699_, new_n39700_,
    new_n39701_, new_n39702_, new_n39703_, new_n39704_, new_n39705_,
    new_n39706_, new_n39707_, new_n39708_, new_n39709_, new_n39710_,
    new_n39711_, new_n39712_, new_n39713_, new_n39714_, new_n39715_,
    new_n39716_, new_n39717_, new_n39718_, new_n39719_, new_n39720_,
    new_n39721_, new_n39722_, new_n39723_, new_n39724_, new_n39725_,
    new_n39726_, new_n39727_, new_n39728_, new_n39729_, new_n39730_,
    new_n39731_, new_n39732_, new_n39733_, new_n39734_, new_n39735_,
    new_n39736_, new_n39737_, new_n39738_, new_n39739_, new_n39740_,
    new_n39741_, new_n39742_, new_n39743_, new_n39744_, new_n39745_,
    new_n39746_, new_n39747_, new_n39748_, new_n39749_, new_n39750_,
    new_n39751_, new_n39752_, new_n39753_, new_n39754_, new_n39755_,
    new_n39756_, new_n39757_, new_n39758_, new_n39759_, new_n39760_,
    new_n39761_, new_n39762_, new_n39763_, new_n39764_, new_n39765_,
    new_n39766_, new_n39767_, new_n39768_, new_n39769_, new_n39770_,
    new_n39771_, new_n39772_, new_n39773_, new_n39774_, new_n39775_,
    new_n39776_, new_n39777_, new_n39778_, new_n39779_, new_n39780_,
    new_n39781_, new_n39782_, new_n39783_, new_n39784_, new_n39785_,
    new_n39786_, new_n39787_, new_n39788_, new_n39789_, new_n39790_,
    new_n39791_, new_n39792_, new_n39793_, new_n39794_, new_n39795_,
    new_n39796_, new_n39797_, new_n39798_, new_n39799_, new_n39800_,
    new_n39801_, new_n39802_, new_n39803_, new_n39804_, new_n39805_,
    new_n39806_, new_n39807_, new_n39808_, new_n39809_, new_n39810_,
    new_n39811_, new_n39812_, new_n39813_, new_n39814_, new_n39815_,
    new_n39816_, new_n39817_, new_n39818_, new_n39819_, new_n39820_,
    new_n39821_, new_n39822_, new_n39823_, new_n39824_, new_n39825_,
    new_n39826_, new_n39827_, new_n39828_, new_n39829_, new_n39830_,
    new_n39831_, new_n39832_, new_n39833_, new_n39834_, new_n39835_,
    new_n39836_, new_n39837_, new_n39838_, new_n39839_, new_n39840_,
    new_n39841_, new_n39842_, new_n39843_, new_n39844_, new_n39845_,
    new_n39846_, new_n39847_, new_n39848_, new_n39849_, new_n39850_,
    new_n39851_, new_n39852_, new_n39853_, new_n39854_, new_n39855_,
    new_n39856_, new_n39857_, new_n39858_, new_n39859_, new_n39860_,
    new_n39861_, new_n39862_, new_n39863_, new_n39864_, new_n39865_,
    new_n39866_, new_n39867_, new_n39868_, new_n39869_, new_n39870_,
    new_n39871_, new_n39872_, new_n39873_, new_n39874_, new_n39875_,
    new_n39876_, new_n39877_, new_n39878_, new_n39879_, new_n39880_,
    new_n39881_, new_n39882_, new_n39883_, new_n39884_, new_n39885_,
    new_n39886_, new_n39887_, new_n39888_, new_n39889_, new_n39890_,
    new_n39891_, new_n39892_, new_n39893_, new_n39894_, new_n39895_,
    new_n39896_, new_n39897_, new_n39898_, new_n39899_, new_n39900_,
    new_n39901_, new_n39902_, new_n39903_, new_n39904_, new_n39905_,
    new_n39906_, new_n39907_, new_n39908_, new_n39909_, new_n39910_,
    new_n39911_, new_n39912_, new_n39913_, new_n39914_, new_n39915_,
    new_n39916_, new_n39917_, new_n39918_, new_n39919_, new_n39920_,
    new_n39921_, new_n39922_, new_n39923_, new_n39924_, new_n39925_,
    new_n39926_, new_n39927_, new_n39928_, new_n39929_, new_n39930_,
    new_n39931_, new_n39932_, new_n39933_, new_n39934_, new_n39935_,
    new_n39936_, new_n39937_, new_n39938_, new_n39939_, new_n39940_,
    new_n39941_, new_n39942_, new_n39943_, new_n39944_, new_n39945_,
    new_n39946_, new_n39947_, new_n39948_, new_n39949_, new_n39950_,
    new_n39951_, new_n39952_, new_n39953_, new_n39954_, new_n39955_,
    new_n39956_, new_n39957_, new_n39958_, new_n39959_, new_n39960_,
    new_n39961_, new_n39962_, new_n39963_, new_n39964_, new_n39965_,
    new_n39966_, new_n39967_, new_n39968_, new_n39969_, new_n39970_,
    new_n39971_, new_n39972_, new_n39973_, new_n39974_, new_n39975_,
    new_n39976_, new_n39977_, new_n39978_, new_n39979_, new_n39980_,
    new_n39981_, new_n39982_, new_n39983_, new_n39984_, new_n39985_,
    new_n39986_, new_n39987_, new_n39988_, new_n39989_, new_n39990_,
    new_n39991_, new_n39992_, new_n39993_, new_n39994_, new_n39995_,
    new_n39996_, new_n39997_, new_n39998_, new_n39999_, new_n40000_,
    new_n40001_, new_n40002_, new_n40003_, new_n40004_, new_n40005_,
    new_n40006_, new_n40007_, new_n40008_, new_n40009_, new_n40010_,
    new_n40011_, new_n40012_, new_n40013_, new_n40014_, new_n40015_,
    new_n40016_, new_n40017_, new_n40018_, new_n40019_, new_n40020_,
    new_n40021_, new_n40022_, new_n40023_, new_n40024_, new_n40025_,
    new_n40026_, new_n40027_, new_n40028_, new_n40029_, new_n40030_,
    new_n40031_, new_n40032_, new_n40033_, new_n40034_, new_n40035_,
    new_n40036_, new_n40037_, new_n40038_, new_n40039_, new_n40040_,
    new_n40041_, new_n40042_, new_n40043_, new_n40044_, new_n40045_,
    new_n40046_, new_n40047_, new_n40048_, new_n40049_, new_n40050_,
    new_n40051_, new_n40052_, new_n40053_, new_n40054_, new_n40055_,
    new_n40056_, new_n40057_, new_n40058_, new_n40059_, new_n40060_,
    new_n40061_, new_n40062_, new_n40063_, new_n40064_, new_n40065_,
    new_n40066_, new_n40067_, new_n40068_, new_n40069_, new_n40070_,
    new_n40071_, new_n40072_, new_n40073_, new_n40074_, new_n40075_,
    new_n40076_, new_n40077_, new_n40078_, new_n40079_, new_n40080_,
    new_n40081_, new_n40082_, new_n40083_, new_n40084_, new_n40085_,
    new_n40086_, new_n40087_, new_n40088_, new_n40089_, new_n40090_,
    new_n40091_, new_n40092_, new_n40093_, new_n40094_, new_n40095_,
    new_n40096_, new_n40097_, new_n40098_, new_n40099_, new_n40100_,
    new_n40101_, new_n40102_, new_n40103_, new_n40104_, new_n40105_,
    new_n40106_, new_n40107_, new_n40108_, new_n40109_, new_n40110_,
    new_n40111_, new_n40112_, new_n40113_, new_n40114_, new_n40115_,
    new_n40116_, new_n40117_, new_n40118_, new_n40119_, new_n40120_,
    new_n40121_, new_n40122_, new_n40123_, new_n40124_, new_n40125_,
    new_n40126_, new_n40127_, new_n40128_, new_n40129_, new_n40130_,
    new_n40131_, new_n40132_, new_n40133_, new_n40134_, new_n40135_,
    new_n40136_, new_n40137_, new_n40138_, new_n40139_, new_n40140_,
    new_n40141_, new_n40142_, new_n40143_, new_n40144_, new_n40145_,
    new_n40146_, new_n40147_, new_n40148_, new_n40149_, new_n40150_,
    new_n40151_, new_n40152_, new_n40153_, new_n40154_, new_n40155_,
    new_n40156_, new_n40157_, new_n40158_, new_n40159_, new_n40160_,
    new_n40161_, new_n40162_, new_n40163_, new_n40164_, new_n40165_,
    new_n40166_, new_n40167_, new_n40168_, new_n40169_, new_n40170_,
    new_n40171_, new_n40172_, new_n40173_, new_n40174_, new_n40175_,
    new_n40176_, new_n40177_, new_n40178_, new_n40179_, new_n40180_,
    new_n40181_, new_n40182_, new_n40183_, new_n40184_, new_n40185_,
    new_n40186_, new_n40187_, new_n40188_, new_n40189_, new_n40190_,
    new_n40191_, new_n40192_, new_n40193_, new_n40194_, new_n40195_,
    new_n40196_, new_n40197_, new_n40198_, new_n40199_, new_n40200_,
    new_n40201_, new_n40202_, new_n40203_, new_n40204_, new_n40205_,
    new_n40206_, new_n40207_, new_n40208_, new_n40209_, new_n40210_,
    new_n40211_, new_n40212_, new_n40213_, new_n40214_, new_n40215_,
    new_n40216_, new_n40217_, new_n40218_, new_n40219_, new_n40220_,
    new_n40221_, new_n40222_, new_n40223_, new_n40224_, new_n40225_,
    new_n40226_, new_n40227_, new_n40228_, new_n40229_, new_n40230_,
    new_n40231_, new_n40232_, new_n40233_, new_n40234_, new_n40235_,
    new_n40236_, new_n40237_, new_n40238_, new_n40239_, new_n40240_,
    new_n40241_, new_n40242_, new_n40243_, new_n40244_, new_n40245_,
    new_n40246_, new_n40247_, new_n40248_, new_n40249_, new_n40250_,
    new_n40251_, new_n40252_, new_n40253_, new_n40254_, new_n40255_,
    new_n40256_, new_n40257_, new_n40258_, new_n40259_, new_n40260_,
    new_n40261_, new_n40262_, new_n40263_, new_n40264_, new_n40265_,
    new_n40266_, new_n40267_, new_n40268_, new_n40269_, new_n40270_,
    new_n40271_, new_n40272_, new_n40273_, new_n40274_, new_n40275_,
    new_n40276_, new_n40277_, new_n40278_, new_n40279_, new_n40280_,
    new_n40281_, new_n40282_, new_n40283_, new_n40284_, new_n40285_,
    new_n40286_, new_n40287_, new_n40288_, new_n40289_, new_n40290_,
    new_n40291_, new_n40292_, new_n40293_, new_n40294_, new_n40295_,
    new_n40296_, new_n40297_, new_n40298_, new_n40299_, new_n40300_,
    new_n40301_, new_n40302_, new_n40303_, new_n40304_, new_n40305_,
    new_n40306_, new_n40307_, new_n40308_, new_n40309_, new_n40310_,
    new_n40311_, new_n40312_, new_n40313_, new_n40314_, new_n40315_,
    new_n40316_, new_n40317_, new_n40318_, new_n40319_, new_n40320_,
    new_n40321_, new_n40322_, new_n40323_, new_n40324_, new_n40325_,
    new_n40326_, new_n40327_, new_n40328_, new_n40329_, new_n40330_,
    new_n40331_, new_n40332_, new_n40333_, new_n40334_, new_n40335_,
    new_n40336_, new_n40337_, new_n40338_, new_n40339_, new_n40340_,
    new_n40341_, new_n40342_, new_n40343_, new_n40344_, new_n40345_,
    new_n40346_, new_n40347_, new_n40348_, new_n40349_, new_n40350_,
    new_n40351_, new_n40352_, new_n40353_, new_n40354_, new_n40355_,
    new_n40356_, new_n40357_, new_n40358_, new_n40359_, new_n40360_,
    new_n40361_, new_n40362_, new_n40363_, new_n40364_, new_n40365_,
    new_n40366_, new_n40367_, new_n40368_, new_n40369_, new_n40370_,
    new_n40371_, new_n40372_, new_n40373_, new_n40374_, new_n40375_,
    new_n40376_, new_n40377_, new_n40378_, new_n40379_, new_n40380_,
    new_n40381_, new_n40382_, new_n40383_, new_n40384_, new_n40385_,
    new_n40386_, new_n40387_, new_n40388_, new_n40389_, new_n40390_,
    new_n40391_, new_n40392_, new_n40393_, new_n40394_, new_n40395_,
    new_n40396_, new_n40397_, new_n40398_, new_n40399_, new_n40400_,
    new_n40401_, new_n40402_, new_n40403_, new_n40404_, new_n40405_,
    new_n40406_, new_n40407_, new_n40408_, new_n40409_, new_n40410_,
    new_n40411_, new_n40412_, new_n40413_, new_n40414_, new_n40415_,
    new_n40416_, new_n40417_, new_n40418_, new_n40419_, new_n40420_,
    new_n40421_, new_n40422_, new_n40423_, new_n40424_, new_n40425_,
    new_n40426_, new_n40427_, new_n40428_, new_n40429_, new_n40430_,
    new_n40431_, new_n40432_, new_n40433_, new_n40434_, new_n40435_,
    new_n40436_, new_n40437_, new_n40438_, new_n40439_, new_n40440_,
    new_n40441_, new_n40442_, new_n40443_, new_n40444_, new_n40445_,
    new_n40446_, new_n40447_, new_n40448_, new_n40449_, new_n40450_,
    new_n40451_, new_n40452_, new_n40453_, new_n40454_, new_n40455_,
    new_n40456_, new_n40457_, new_n40458_, new_n40459_, new_n40460_,
    new_n40461_, new_n40462_, new_n40463_, new_n40464_, new_n40465_,
    new_n40466_, new_n40467_, new_n40468_, new_n40469_, new_n40470_,
    new_n40471_, new_n40472_, new_n40473_, new_n40474_, new_n40475_,
    new_n40476_, new_n40477_, new_n40478_, new_n40479_, new_n40480_,
    new_n40481_, new_n40482_, new_n40483_, new_n40484_, new_n40485_,
    new_n40486_, new_n40487_, new_n40488_, new_n40489_, new_n40490_,
    new_n40491_, new_n40492_, new_n40493_, new_n40494_, new_n40495_,
    new_n40496_, new_n40497_, new_n40498_, new_n40499_, new_n40500_,
    new_n40501_, new_n40502_, new_n40503_, new_n40504_, new_n40505_,
    new_n40506_, new_n40507_, new_n40508_, new_n40509_, new_n40510_,
    new_n40511_, new_n40512_, new_n40513_, new_n40514_, new_n40515_,
    new_n40516_, new_n40517_, new_n40518_, new_n40519_, new_n40520_,
    new_n40521_, new_n40522_, new_n40523_, new_n40524_, new_n40525_,
    new_n40526_, new_n40527_, new_n40528_, new_n40529_, new_n40530_,
    new_n40531_, new_n40532_, new_n40533_, new_n40534_, new_n40535_,
    new_n40536_, new_n40537_, new_n40538_, new_n40539_, new_n40540_,
    new_n40541_, new_n40542_, new_n40543_, new_n40544_, new_n40545_,
    new_n40546_, new_n40547_, new_n40548_, new_n40549_, new_n40550_,
    new_n40551_, new_n40552_, new_n40553_, new_n40554_, new_n40555_,
    new_n40556_, new_n40557_, new_n40558_, new_n40559_, new_n40560_,
    new_n40561_, new_n40562_, new_n40563_, new_n40564_, new_n40565_,
    new_n40566_, new_n40567_, new_n40568_, new_n40569_, new_n40570_,
    new_n40571_, new_n40572_, new_n40573_, new_n40574_, new_n40575_,
    new_n40576_, new_n40577_, new_n40578_, new_n40579_, new_n40580_,
    new_n40581_, new_n40582_, new_n40583_, new_n40584_, new_n40585_,
    new_n40586_, new_n40587_, new_n40588_, new_n40589_, new_n40590_,
    new_n40591_, new_n40592_, new_n40593_, new_n40594_, new_n40595_,
    new_n40596_, new_n40597_, new_n40598_, new_n40599_, new_n40600_,
    new_n40601_, new_n40602_, new_n40603_, new_n40604_, new_n40605_,
    new_n40606_, new_n40607_, new_n40608_, new_n40609_, new_n40610_,
    new_n40611_, new_n40612_, new_n40613_, new_n40614_, new_n40615_,
    new_n40616_, new_n40617_, new_n40618_, new_n40619_, new_n40620_,
    new_n40621_, new_n40622_, new_n40623_, new_n40624_, new_n40625_,
    new_n40626_, new_n40627_, new_n40628_, new_n40629_, new_n40630_,
    new_n40631_, new_n40632_, new_n40633_, new_n40634_, new_n40635_,
    new_n40636_, new_n40637_, new_n40638_, new_n40639_, new_n40640_,
    new_n40641_, new_n40642_, new_n40643_, new_n40644_, new_n40645_,
    new_n40646_, new_n40647_, new_n40648_, new_n40649_, new_n40650_,
    new_n40651_, new_n40652_, new_n40653_, new_n40654_, new_n40655_,
    new_n40656_, new_n40657_, new_n40658_, new_n40659_, new_n40660_,
    new_n40661_, new_n40662_, new_n40663_, new_n40664_, new_n40665_,
    new_n40666_, new_n40667_, new_n40668_, new_n40669_, new_n40670_,
    new_n40671_, new_n40672_, new_n40673_, new_n40674_, new_n40675_,
    new_n40676_, new_n40677_, new_n40678_, new_n40679_, new_n40680_,
    new_n40681_, new_n40682_, new_n40683_, new_n40684_, new_n40685_,
    new_n40686_, new_n40687_, new_n40688_, new_n40689_, new_n40690_,
    new_n40691_, new_n40692_, new_n40693_, new_n40694_, new_n40695_,
    new_n40696_, new_n40697_, new_n40698_, new_n40699_, new_n40700_,
    new_n40701_, new_n40702_, new_n40703_, new_n40704_, new_n40705_,
    new_n40706_, new_n40707_, new_n40708_, new_n40709_, new_n40710_,
    new_n40711_, new_n40712_, new_n40713_, new_n40714_, new_n40715_,
    new_n40716_, new_n40717_, new_n40718_, new_n40719_, new_n40720_,
    new_n40721_, new_n40722_, new_n40723_, new_n40724_, new_n40725_,
    new_n40726_, new_n40727_, new_n40728_, new_n40729_, new_n40730_,
    new_n40731_, new_n40732_, new_n40733_, new_n40734_, new_n40735_,
    new_n40736_, new_n40737_, new_n40738_, new_n40739_, new_n40740_,
    new_n40741_, new_n40742_, new_n40743_, new_n40744_, new_n40745_,
    new_n40746_, new_n40747_, new_n40748_, new_n40749_, new_n40750_,
    new_n40751_, new_n40752_, new_n40753_, new_n40754_, new_n40755_,
    new_n40756_, new_n40757_, new_n40758_, new_n40759_, new_n40760_,
    new_n40761_, new_n40762_, new_n40763_, new_n40764_, new_n40765_,
    new_n40766_, new_n40767_, new_n40768_, new_n40769_, new_n40770_,
    new_n40771_, new_n40772_, new_n40773_, new_n40774_, new_n40775_,
    new_n40776_, new_n40777_, new_n40778_, new_n40779_, new_n40780_,
    new_n40781_, new_n40782_, new_n40783_, new_n40784_, new_n40785_,
    new_n40786_, new_n40787_, new_n40788_, new_n40789_, new_n40790_,
    new_n40791_, new_n40792_, new_n40793_, new_n40794_, new_n40795_,
    new_n40796_, new_n40797_, new_n40798_, new_n40799_, new_n40800_,
    new_n40801_, new_n40802_, new_n40803_, new_n40804_, new_n40805_,
    new_n40806_, new_n40807_, new_n40808_, new_n40809_, new_n40810_,
    new_n40811_, new_n40812_, new_n40813_, new_n40814_, new_n40815_,
    new_n40816_, new_n40817_, new_n40818_, new_n40819_, new_n40820_,
    new_n40821_, new_n40822_, new_n40823_, new_n40824_, new_n40825_,
    new_n40826_, new_n40827_, new_n40828_, new_n40829_, new_n40830_,
    new_n40831_, new_n40832_, new_n40833_, new_n40834_, new_n40835_,
    new_n40836_, new_n40837_, new_n40838_, new_n40839_, new_n40840_,
    new_n40841_, new_n40842_, new_n40843_, new_n40844_, new_n40845_,
    new_n40846_, new_n40847_, new_n40848_, new_n40849_, new_n40850_,
    new_n40851_, new_n40852_, new_n40853_, new_n40854_, new_n40855_,
    new_n40856_, new_n40857_, new_n40858_, new_n40859_, new_n40860_,
    new_n40861_, new_n40862_, new_n40863_, new_n40864_, new_n40865_,
    new_n40866_, new_n40867_, new_n40868_, new_n40869_, new_n40870_,
    new_n40871_, new_n40872_, new_n40873_, new_n40874_, new_n40875_,
    new_n40876_, new_n40877_, new_n40878_, new_n40879_, new_n40880_,
    new_n40881_, new_n40882_, new_n40883_, new_n40884_, new_n40885_,
    new_n40886_, new_n40887_, new_n40888_, new_n40889_, new_n40890_,
    new_n40891_, new_n40892_, new_n40893_, new_n40894_, new_n40895_,
    new_n40896_, new_n40897_, new_n40898_, new_n40899_, new_n40900_,
    new_n40901_, new_n40902_, new_n40903_, new_n40904_, new_n40905_,
    new_n40906_, new_n40907_, new_n40908_, new_n40909_, new_n40910_,
    new_n40911_, new_n40912_, new_n40913_, new_n40914_, new_n40915_,
    new_n40916_, new_n40917_, new_n40918_, new_n40919_, new_n40920_,
    new_n40921_, new_n40922_, new_n40923_, new_n40924_, new_n40925_,
    new_n40926_, new_n40927_, new_n40928_, new_n40929_, new_n40930_,
    new_n40931_, new_n40932_, new_n40933_, new_n40934_, new_n40935_,
    new_n40936_, new_n40937_, new_n40938_, new_n40939_, new_n40940_,
    new_n40941_, new_n40942_, new_n40943_, new_n40944_, new_n40945_,
    new_n40946_, new_n40947_, new_n40948_, new_n40949_, new_n40950_,
    new_n40951_, new_n40952_, new_n40953_, new_n40954_, new_n40955_,
    new_n40956_, new_n40957_, new_n40958_, new_n40959_, new_n40960_,
    new_n40961_, new_n40962_, new_n40963_, new_n40964_, new_n40965_,
    new_n40966_, new_n40967_, new_n40968_, new_n40969_, new_n40970_,
    new_n40971_, new_n40972_, new_n40973_, new_n40974_, new_n40975_,
    new_n40976_, new_n40977_, new_n40978_, new_n40979_, new_n40980_,
    new_n40981_, new_n40982_, new_n40983_, new_n40984_, new_n40985_,
    new_n40986_, new_n40987_, new_n40988_, new_n40989_, new_n40990_,
    new_n40991_, new_n40992_, new_n40993_, new_n40994_, new_n40995_,
    new_n40996_, new_n40997_, new_n40998_, new_n40999_, new_n41000_,
    new_n41001_, new_n41002_, new_n41003_, new_n41004_, new_n41005_,
    new_n41006_, new_n41007_, new_n41008_, new_n41009_, new_n41010_,
    new_n41011_, new_n41012_, new_n41013_, new_n41014_, new_n41015_,
    new_n41016_, new_n41017_, new_n41018_, new_n41019_, new_n41020_,
    new_n41021_, new_n41022_, new_n41023_, new_n41024_, new_n41025_,
    new_n41026_, new_n41027_, new_n41028_, new_n41029_, new_n41030_,
    new_n41031_, new_n41032_, new_n41033_, new_n41034_, new_n41035_,
    new_n41036_, new_n41037_, new_n41038_, new_n41039_, new_n41040_,
    new_n41041_, new_n41042_, new_n41043_, new_n41044_, new_n41045_,
    new_n41046_, new_n41047_, new_n41048_, new_n41049_, new_n41050_,
    new_n41051_, new_n41052_, new_n41053_, new_n41054_, new_n41055_,
    new_n41056_, new_n41057_, new_n41058_, new_n41059_, new_n41060_,
    new_n41061_, new_n41062_, new_n41063_, new_n41064_, new_n41065_,
    new_n41066_, new_n41067_, new_n41068_, new_n41069_, new_n41070_,
    new_n41071_, new_n41072_, new_n41073_, new_n41074_, new_n41075_,
    new_n41076_, new_n41077_, new_n41078_, new_n41079_, new_n41080_,
    new_n41081_, new_n41082_, new_n41083_, new_n41084_, new_n41085_,
    new_n41086_, new_n41087_, new_n41088_, new_n41089_, new_n41090_,
    new_n41091_, new_n41092_, new_n41093_, new_n41094_, new_n41095_,
    new_n41096_, new_n41097_, new_n41098_, new_n41099_, new_n41100_,
    new_n41101_, new_n41102_, new_n41103_, new_n41104_, new_n41105_,
    new_n41106_, new_n41107_, new_n41108_, new_n41109_, new_n41110_,
    new_n41111_, new_n41112_, new_n41113_, new_n41114_, new_n41115_,
    new_n41116_, new_n41117_, new_n41118_, new_n41119_, new_n41120_,
    new_n41121_, new_n41122_, new_n41123_, new_n41124_, new_n41125_,
    new_n41126_, new_n41127_, new_n41128_, new_n41129_, new_n41130_,
    new_n41131_, new_n41132_, new_n41133_, new_n41134_, new_n41135_,
    new_n41136_, new_n41137_, new_n41138_, new_n41139_, new_n41140_,
    new_n41141_, new_n41142_, new_n41143_, new_n41144_, new_n41145_,
    new_n41146_, new_n41147_, new_n41148_, new_n41149_, new_n41150_,
    new_n41151_, new_n41152_, new_n41153_, new_n41154_, new_n41155_,
    new_n41156_, new_n41157_, new_n41158_, new_n41159_, new_n41160_,
    new_n41161_, new_n41162_, new_n41163_, new_n41164_, new_n41165_,
    new_n41166_, new_n41167_, new_n41168_, new_n41169_, new_n41170_,
    new_n41171_, new_n41172_, new_n41173_, new_n41174_, new_n41175_,
    new_n41176_, new_n41177_, new_n41178_, new_n41179_, new_n41180_,
    new_n41181_, new_n41182_, new_n41183_, new_n41184_, new_n41185_,
    new_n41186_, new_n41187_, new_n41188_, new_n41189_, new_n41190_,
    new_n41191_, new_n41192_, new_n41193_, new_n41194_, new_n41195_,
    new_n41196_, new_n41197_, new_n41198_, new_n41199_, new_n41200_,
    new_n41201_, new_n41202_, new_n41203_, new_n41204_, new_n41205_,
    new_n41206_, new_n41207_, new_n41208_, new_n41209_, new_n41210_,
    new_n41211_, new_n41212_, new_n41213_, new_n41214_, new_n41215_,
    new_n41216_, new_n41217_, new_n41218_, new_n41219_, new_n41220_,
    new_n41221_, new_n41222_, new_n41223_, new_n41224_, new_n41225_,
    new_n41226_, new_n41227_, new_n41228_, new_n41229_, new_n41230_,
    new_n41231_, new_n41232_, new_n41233_, new_n41234_, new_n41235_,
    new_n41236_, new_n41237_, new_n41238_, new_n41239_, new_n41240_,
    new_n41241_, new_n41242_, new_n41243_, new_n41244_, new_n41245_,
    new_n41246_, new_n41247_, new_n41248_, new_n41249_, new_n41250_,
    new_n41251_, new_n41252_, new_n41253_, new_n41254_, new_n41255_,
    new_n41256_, new_n41257_, new_n41258_, new_n41259_, new_n41260_,
    new_n41261_, new_n41262_, new_n41263_, new_n41264_, new_n41265_,
    new_n41266_, new_n41267_, new_n41268_, new_n41269_, new_n41270_,
    new_n41271_, new_n41272_, new_n41273_, new_n41274_, new_n41275_,
    new_n41276_, new_n41277_, new_n41278_, new_n41279_, new_n41280_,
    new_n41281_, new_n41282_, new_n41283_, new_n41284_, new_n41285_,
    new_n41286_, new_n41287_, new_n41288_, new_n41289_, new_n41290_,
    new_n41291_, new_n41292_, new_n41293_, new_n41294_, new_n41295_,
    new_n41296_, new_n41297_, new_n41298_, new_n41299_, new_n41300_,
    new_n41301_, new_n41302_, new_n41303_, new_n41304_, new_n41305_,
    new_n41306_, new_n41307_, new_n41308_, new_n41309_, new_n41310_,
    new_n41311_, new_n41312_, new_n41313_, new_n41314_, new_n41315_,
    new_n41316_, new_n41317_, new_n41318_, new_n41319_, new_n41320_,
    new_n41321_, new_n41322_, new_n41323_, new_n41324_, new_n41325_,
    new_n41326_, new_n41327_, new_n41328_, new_n41329_, new_n41330_,
    new_n41331_, new_n41332_, new_n41333_, new_n41334_, new_n41335_,
    new_n41336_, new_n41337_, new_n41338_, new_n41339_, new_n41340_,
    new_n41341_, new_n41342_, new_n41343_, new_n41344_, new_n41345_,
    new_n41346_, new_n41347_, new_n41348_, new_n41349_, new_n41350_,
    new_n41351_, new_n41352_, new_n41353_, new_n41354_, new_n41355_,
    new_n41356_, new_n41357_, new_n41358_, new_n41359_, new_n41360_,
    new_n41361_, new_n41362_, new_n41363_, new_n41364_, new_n41365_,
    new_n41366_, new_n41367_, new_n41368_, new_n41369_, new_n41370_,
    new_n41371_, new_n41372_, new_n41373_, new_n41374_, new_n41375_,
    new_n41376_, new_n41377_, new_n41378_, new_n41379_, new_n41380_,
    new_n41381_, new_n41382_, new_n41383_, new_n41384_, new_n41385_,
    new_n41386_, new_n41387_, new_n41388_, new_n41389_, new_n41390_,
    new_n41391_, new_n41392_, new_n41393_, new_n41394_, new_n41395_,
    new_n41396_, new_n41397_, new_n41398_, new_n41399_, new_n41400_,
    new_n41401_, new_n41402_, new_n41403_, new_n41404_, new_n41405_,
    new_n41406_, new_n41407_, new_n41408_, new_n41409_, new_n41410_,
    new_n41411_, new_n41412_, new_n41413_, new_n41414_, new_n41415_,
    new_n41416_, new_n41417_, new_n41418_, new_n41419_, new_n41420_,
    new_n41421_, new_n41422_, new_n41423_, new_n41424_, new_n41425_,
    new_n41426_, new_n41427_, new_n41428_, new_n41429_, new_n41430_,
    new_n41431_, new_n41432_, new_n41433_, new_n41434_, new_n41435_,
    new_n41436_, new_n41437_, new_n41438_, new_n41439_, new_n41440_,
    new_n41441_, new_n41442_, new_n41443_, new_n41444_, new_n41445_,
    new_n41446_, new_n41447_, new_n41448_, new_n41449_, new_n41450_,
    new_n41451_, new_n41452_, new_n41453_, new_n41454_, new_n41455_,
    new_n41456_, new_n41457_, new_n41458_, new_n41459_, new_n41460_,
    new_n41461_, new_n41462_, new_n41463_, new_n41464_, new_n41465_,
    new_n41466_, new_n41467_, new_n41468_, new_n41469_, new_n41470_,
    new_n41471_, new_n41472_, new_n41473_, new_n41474_, new_n41475_,
    new_n41476_, new_n41477_, new_n41478_, new_n41479_, new_n41480_,
    new_n41481_, new_n41482_, new_n41483_, new_n41484_, new_n41485_,
    new_n41486_, new_n41487_, new_n41488_, new_n41489_, new_n41490_,
    new_n41491_, new_n41492_, new_n41493_, new_n41494_, new_n41495_,
    new_n41496_, new_n41497_, new_n41498_, new_n41499_, new_n41500_,
    new_n41501_, new_n41502_, new_n41503_, new_n41504_, new_n41505_,
    new_n41506_, new_n41507_, new_n41508_, new_n41509_, new_n41510_,
    new_n41511_, new_n41512_, new_n41513_, new_n41514_, new_n41515_,
    new_n41516_, new_n41517_, new_n41518_, new_n41519_, new_n41520_,
    new_n41521_, new_n41522_, new_n41523_, new_n41524_, new_n41525_,
    new_n41526_, new_n41527_, new_n41528_, new_n41529_, new_n41530_,
    new_n41531_, new_n41532_, new_n41533_, new_n41534_, new_n41535_,
    new_n41536_, new_n41537_, new_n41538_, new_n41539_, new_n41540_,
    new_n41541_, new_n41542_, new_n41543_, new_n41544_, new_n41545_,
    new_n41546_, new_n41547_, new_n41548_, new_n41549_, new_n41550_,
    new_n41551_, new_n41552_, new_n41553_, new_n41554_, new_n41555_,
    new_n41556_, new_n41557_, new_n41558_, new_n41559_, new_n41560_,
    new_n41561_, new_n41562_, new_n41563_, new_n41564_, new_n41565_,
    new_n41566_, new_n41567_, new_n41568_, new_n41569_, new_n41570_,
    new_n41571_, new_n41572_, new_n41573_, new_n41574_, new_n41575_,
    new_n41576_, new_n41577_, new_n41578_, new_n41579_, new_n41580_,
    new_n41581_, new_n41582_, new_n41583_, new_n41584_, new_n41585_,
    new_n41586_, new_n41587_, new_n41588_, new_n41589_, new_n41590_,
    new_n41591_, new_n41592_, new_n41593_, new_n41594_, new_n41595_,
    new_n41596_, new_n41597_, new_n41598_, new_n41599_, new_n41600_,
    new_n41601_, new_n41602_, new_n41603_, new_n41604_, new_n41605_,
    new_n41606_, new_n41607_, new_n41608_, new_n41609_, new_n41610_,
    new_n41611_, new_n41612_, new_n41613_, new_n41614_, new_n41615_,
    new_n41616_, new_n41617_, new_n41618_, new_n41619_, new_n41620_,
    new_n41621_, new_n41622_, new_n41623_, new_n41624_, new_n41625_,
    new_n41626_, new_n41627_, new_n41628_, new_n41629_, new_n41630_,
    new_n41631_, new_n41632_, new_n41633_, new_n41634_, new_n41635_,
    new_n41636_, new_n41637_, new_n41638_, new_n41639_, new_n41640_,
    new_n41641_, new_n41642_, new_n41643_, new_n41644_, new_n41645_,
    new_n41646_, new_n41647_, new_n41648_, new_n41649_, new_n41650_,
    new_n41651_, new_n41652_, new_n41653_, new_n41654_, new_n41655_,
    new_n41656_, new_n41657_, new_n41658_, new_n41659_, new_n41660_,
    new_n41661_, new_n41662_, new_n41663_, new_n41664_, new_n41665_,
    new_n41666_, new_n41667_, new_n41668_, new_n41669_, new_n41670_,
    new_n41671_, new_n41672_, new_n41673_, new_n41674_, new_n41675_,
    new_n41676_, new_n41677_, new_n41678_, new_n41679_, new_n41680_,
    new_n41681_, new_n41682_, new_n41683_, new_n41684_, new_n41685_,
    new_n41686_, new_n41687_, new_n41688_, new_n41689_, new_n41690_,
    new_n41691_, new_n41692_, new_n41693_, new_n41694_, new_n41695_,
    new_n41696_, new_n41697_, new_n41698_, new_n41699_, new_n41700_,
    new_n41701_, new_n41702_, new_n41703_, new_n41704_, new_n41705_,
    new_n41706_, new_n41707_, new_n41708_, new_n41709_, new_n41710_,
    new_n41711_, new_n41712_, new_n41713_, new_n41714_, new_n41715_,
    new_n41716_, new_n41717_, new_n41718_, new_n41719_, new_n41720_,
    new_n41721_, new_n41722_, new_n41723_, new_n41724_, new_n41725_,
    new_n41726_, new_n41727_, new_n41728_, new_n41729_, new_n41730_,
    new_n41731_, new_n41732_, new_n41733_, new_n41734_, new_n41735_,
    new_n41736_, new_n41737_, new_n41738_, new_n41739_, new_n41740_,
    new_n41741_, new_n41742_, new_n41743_, new_n41744_, new_n41745_,
    new_n41746_, new_n41747_, new_n41748_, new_n41749_, new_n41750_,
    new_n41751_, new_n41752_, new_n41753_, new_n41754_, new_n41755_,
    new_n41756_, new_n41757_, new_n41758_, new_n41759_, new_n41760_,
    new_n41761_, new_n41762_, new_n41763_, new_n41764_, new_n41765_,
    new_n41766_, new_n41767_, new_n41768_, new_n41769_, new_n41770_,
    new_n41771_, new_n41772_, new_n41773_, new_n41774_, new_n41775_,
    new_n41776_, new_n41777_, new_n41778_, new_n41779_, new_n41780_,
    new_n41781_, new_n41782_, new_n41783_, new_n41784_, new_n41785_,
    new_n41786_, new_n41787_, new_n41788_, new_n41789_, new_n41790_,
    new_n41791_, new_n41792_, new_n41793_, new_n41794_, new_n41795_,
    new_n41796_, new_n41797_, new_n41798_, new_n41799_, new_n41800_,
    new_n41801_, new_n41802_, new_n41803_, new_n41804_, new_n41805_,
    new_n41806_, new_n41807_, new_n41808_, new_n41809_, new_n41810_,
    new_n41811_, new_n41812_, new_n41813_, new_n41814_, new_n41815_,
    new_n41816_, new_n41817_, new_n41818_, new_n41819_, new_n41820_,
    new_n41821_, new_n41822_, new_n41823_, new_n41824_, new_n41825_,
    new_n41826_, new_n41827_, new_n41828_, new_n41829_, new_n41830_,
    new_n41831_, new_n41832_, new_n41833_, new_n41834_, new_n41835_,
    new_n41836_, new_n41837_, new_n41838_, new_n41839_, new_n41840_,
    new_n41841_, new_n41842_, new_n41843_, new_n41844_, new_n41845_,
    new_n41846_, new_n41847_, new_n41848_, new_n41849_, new_n41850_,
    new_n41851_, new_n41852_, new_n41853_, new_n41854_, new_n41855_,
    new_n41856_, new_n41857_, new_n41858_, new_n41859_, new_n41860_,
    new_n41861_, new_n41862_, new_n41863_, new_n41864_, new_n41865_,
    new_n41866_, new_n41867_, new_n41868_, new_n41869_, new_n41870_,
    new_n41871_, new_n41872_, new_n41873_, new_n41874_, new_n41875_,
    new_n41876_, new_n41877_, new_n41878_, new_n41879_, new_n41880_,
    new_n41881_, new_n41882_, new_n41883_, new_n41884_, new_n41885_,
    new_n41886_, new_n41887_, new_n41888_, new_n41889_, new_n41890_,
    new_n41891_, new_n41892_, new_n41893_, new_n41894_, new_n41895_,
    new_n41896_, new_n41897_, new_n41898_, new_n41899_, new_n41900_,
    new_n41901_, new_n41902_, new_n41903_, new_n41904_, new_n41905_,
    new_n41906_, new_n41907_, new_n41908_, new_n41909_, new_n41910_,
    new_n41911_, new_n41912_, new_n41913_, new_n41914_, new_n41915_,
    new_n41916_, new_n41917_, new_n41918_, new_n41919_, new_n41920_,
    new_n41921_, new_n41922_, new_n41923_, new_n41924_, new_n41925_,
    new_n41926_, new_n41927_, new_n41928_, new_n41929_, new_n41930_,
    new_n41931_, new_n41932_, new_n41933_, new_n41934_, new_n41935_,
    new_n41936_, new_n41937_, new_n41938_, new_n41939_, new_n41940_,
    new_n41941_, new_n41942_, new_n41943_, new_n41944_, new_n41945_,
    new_n41946_, new_n41947_, new_n41948_, new_n41949_, new_n41950_,
    new_n41951_, new_n41952_, new_n41953_, new_n41954_, new_n41955_,
    new_n41956_, new_n41957_, new_n41958_, new_n41959_, new_n41960_,
    new_n41961_, new_n41962_, new_n41963_, new_n41964_, new_n41965_,
    new_n41966_, new_n41967_, new_n41968_, new_n41969_, new_n41970_,
    new_n41971_, new_n41972_, new_n41973_, new_n41974_, new_n41975_,
    new_n41976_, new_n41977_, new_n41978_, new_n41979_, new_n41980_,
    new_n41981_, new_n41982_, new_n41983_, new_n41984_, new_n41985_,
    new_n41986_, new_n41987_, new_n41988_, new_n41989_, new_n41990_,
    new_n41991_, new_n41992_, new_n41993_, new_n41994_, new_n41995_,
    new_n41996_, new_n41997_, new_n41998_, new_n41999_, new_n42000_,
    new_n42001_, new_n42002_, new_n42003_, new_n42004_, new_n42005_,
    new_n42006_, new_n42007_, new_n42008_, new_n42009_, new_n42010_,
    new_n42011_, new_n42012_, new_n42013_, new_n42014_, new_n42015_,
    new_n42016_, new_n42017_, new_n42018_, new_n42019_, new_n42020_,
    new_n42021_, new_n42022_, new_n42023_, new_n42024_, new_n42025_,
    new_n42026_, new_n42027_, new_n42028_, new_n42029_, new_n42030_,
    new_n42031_, new_n42032_, new_n42033_, new_n42034_, new_n42035_,
    new_n42036_, new_n42037_, new_n42038_, new_n42039_, new_n42040_,
    new_n42041_, new_n42042_, new_n42043_, new_n42044_, new_n42045_,
    new_n42046_, new_n42047_, new_n42048_, new_n42049_, new_n42050_,
    new_n42051_, new_n42052_, new_n42053_, new_n42054_, new_n42055_,
    new_n42056_, new_n42057_, new_n42058_, new_n42059_, new_n42060_,
    new_n42061_, new_n42062_, new_n42063_, new_n42064_, new_n42065_,
    new_n42066_, new_n42067_, new_n42068_, new_n42069_, new_n42070_,
    new_n42071_, new_n42072_, new_n42073_, new_n42074_, new_n42075_,
    new_n42076_, new_n42077_, new_n42078_, new_n42079_, new_n42080_,
    new_n42081_, new_n42082_, new_n42083_, new_n42084_, new_n42085_,
    new_n42086_, new_n42087_, new_n42088_, new_n42089_, new_n42090_,
    new_n42091_, new_n42092_, new_n42093_, new_n42094_, new_n42095_,
    new_n42096_, new_n42097_, new_n42098_, new_n42099_, new_n42100_,
    new_n42101_, new_n42102_, new_n42103_, new_n42104_, new_n42105_,
    new_n42106_, new_n42107_, new_n42108_, new_n42109_, new_n42110_,
    new_n42111_, new_n42112_, new_n42113_, new_n42114_, new_n42115_,
    new_n42116_, new_n42117_, new_n42118_, new_n42119_, new_n42120_,
    new_n42121_, new_n42122_, new_n42123_, new_n42124_, new_n42125_,
    new_n42126_, new_n42127_, new_n42128_, new_n42129_, new_n42130_,
    new_n42131_, new_n42132_, new_n42133_, new_n42134_, new_n42135_,
    new_n42136_, new_n42137_, new_n42138_, new_n42139_, new_n42140_,
    new_n42141_, new_n42142_, new_n42143_, new_n42144_, new_n42145_,
    new_n42146_, new_n42147_, new_n42148_, new_n42149_, new_n42150_,
    new_n42151_, new_n42152_, new_n42153_, new_n42154_, new_n42155_,
    new_n42156_, new_n42157_, new_n42158_, new_n42159_, new_n42160_,
    new_n42161_, new_n42162_, new_n42163_, new_n42164_, new_n42165_,
    new_n42166_, new_n42167_, new_n42168_, new_n42169_, new_n42170_,
    new_n42171_, new_n42172_, new_n42173_, new_n42174_, new_n42175_,
    new_n42176_, new_n42177_, new_n42178_, new_n42179_, new_n42180_,
    new_n42181_, new_n42182_, new_n42183_, new_n42184_, new_n42185_,
    new_n42186_, new_n42187_, new_n42188_, new_n42189_, new_n42190_,
    new_n42191_, new_n42192_, new_n42193_, new_n42194_, new_n42195_,
    new_n42196_, new_n42197_, new_n42198_, new_n42199_, new_n42200_,
    new_n42201_, new_n42202_, new_n42203_, new_n42204_, new_n42205_,
    new_n42206_, new_n42207_, new_n42208_, new_n42209_, new_n42210_,
    new_n42211_, new_n42212_, new_n42213_, new_n42214_, new_n42215_,
    new_n42216_, new_n42217_, new_n42218_, new_n42219_, new_n42220_,
    new_n42221_, new_n42222_, new_n42223_, new_n42224_, new_n42225_,
    new_n42226_, new_n42227_, new_n42228_, new_n42229_, new_n42230_,
    new_n42231_, new_n42232_, new_n42233_, new_n42234_, new_n42235_,
    new_n42236_, new_n42237_, new_n42238_, new_n42239_, new_n42240_,
    new_n42241_, new_n42242_, new_n42243_, new_n42244_, new_n42245_,
    new_n42246_, new_n42247_, new_n42248_, new_n42249_, new_n42250_,
    new_n42251_, new_n42252_, new_n42253_, new_n42254_, new_n42255_,
    new_n42256_, new_n42257_, new_n42258_, new_n42259_, new_n42260_,
    new_n42261_, new_n42262_, new_n42263_, new_n42264_, new_n42265_,
    new_n42266_, new_n42267_, new_n42268_, new_n42269_, new_n42270_,
    new_n42271_, new_n42272_, new_n42273_, new_n42274_, new_n42275_,
    new_n42276_, new_n42277_, new_n42278_, new_n42279_, new_n42280_,
    new_n42281_, new_n42282_, new_n42283_, new_n42284_, new_n42285_,
    new_n42286_, new_n42287_, new_n42288_, new_n42289_, new_n42290_,
    new_n42291_, new_n42292_, new_n42293_, new_n42294_, new_n42295_,
    new_n42296_, new_n42297_, new_n42298_, new_n42299_, new_n42300_,
    new_n42301_, new_n42302_, new_n42303_, new_n42304_, new_n42305_,
    new_n42306_, new_n42307_, new_n42308_, new_n42309_, new_n42310_,
    new_n42311_, new_n42312_, new_n42313_, new_n42314_, new_n42315_,
    new_n42316_, new_n42317_, new_n42318_, new_n42319_, new_n42320_,
    new_n42321_, new_n42322_, new_n42323_, new_n42324_, new_n42325_,
    new_n42326_, new_n42327_, new_n42328_, new_n42329_, new_n42330_,
    new_n42331_, new_n42332_, new_n42333_, new_n42334_, new_n42335_,
    new_n42336_, new_n42337_, new_n42338_, new_n42339_, new_n42340_,
    new_n42341_, new_n42342_, new_n42343_, new_n42344_, new_n42345_,
    new_n42346_, new_n42347_, new_n42348_, new_n42349_, new_n42350_,
    new_n42351_, new_n42352_, new_n42353_, new_n42354_, new_n42355_,
    new_n42356_, new_n42357_, new_n42358_, new_n42359_, new_n42360_,
    new_n42361_, new_n42362_, new_n42363_, new_n42364_, new_n42365_,
    new_n42366_, new_n42367_, new_n42368_, new_n42369_, new_n42370_,
    new_n42371_, new_n42372_, new_n42373_, new_n42374_, new_n42375_,
    new_n42376_, new_n42377_, new_n42378_, new_n42379_, new_n42380_,
    new_n42381_, new_n42382_, new_n42383_, new_n42384_, new_n42385_,
    new_n42386_, new_n42387_, new_n42388_, new_n42389_, new_n42390_,
    new_n42391_, new_n42392_, new_n42393_, new_n42394_, new_n42395_,
    new_n42396_, new_n42397_, new_n42398_, new_n42399_, new_n42400_,
    new_n42401_, new_n42402_, new_n42403_, new_n42404_, new_n42405_,
    new_n42406_, new_n42407_, new_n42408_, new_n42409_, new_n42410_,
    new_n42411_, new_n42412_, new_n42413_, new_n42414_, new_n42415_,
    new_n42416_, new_n42417_, new_n42418_, new_n42419_, new_n42420_,
    new_n42421_, new_n42422_, new_n42423_, new_n42424_, new_n42425_,
    new_n42426_, new_n42427_, new_n42428_, new_n42429_, new_n42430_,
    new_n42431_, new_n42432_, new_n42433_, new_n42434_, new_n42435_,
    new_n42436_, new_n42437_, new_n42438_, new_n42439_, new_n42440_,
    new_n42441_, new_n42442_, new_n42443_, new_n42444_, new_n42445_,
    new_n42446_, new_n42447_, new_n42448_, new_n42449_, new_n42450_,
    new_n42451_, new_n42452_, new_n42453_, new_n42454_, new_n42455_,
    new_n42456_, new_n42457_, new_n42458_, new_n42459_, new_n42460_,
    new_n42461_, new_n42462_, new_n42463_, new_n42464_, new_n42465_,
    new_n42466_, new_n42467_, new_n42468_, new_n42469_, new_n42470_,
    new_n42471_, new_n42472_, new_n42473_, new_n42474_, new_n42475_,
    new_n42476_, new_n42477_, new_n42478_, new_n42479_, new_n42480_,
    new_n42481_, new_n42482_, new_n42483_, new_n42484_, new_n42485_,
    new_n42486_, new_n42487_, new_n42488_, new_n42489_, new_n42490_,
    new_n42491_, new_n42492_, new_n42493_, new_n42494_, new_n42495_,
    new_n42496_, new_n42497_, new_n42498_, new_n42499_, new_n42500_,
    new_n42501_, new_n42502_, new_n42503_, new_n42504_, new_n42505_,
    new_n42506_, new_n42507_, new_n42508_, new_n42509_, new_n42510_,
    new_n42511_, new_n42512_, new_n42513_, new_n42514_, new_n42515_,
    new_n42516_, new_n42517_, new_n42518_, new_n42519_, new_n42520_,
    new_n42521_, new_n42522_, new_n42523_, new_n42524_, new_n42525_,
    new_n42526_, new_n42527_, new_n42528_, new_n42529_, new_n42530_,
    new_n42531_, new_n42532_, new_n42533_, new_n42534_, new_n42535_,
    new_n42536_, new_n42537_, new_n42538_, new_n42539_, new_n42540_,
    new_n42541_, new_n42542_, new_n42543_, new_n42544_, new_n42545_,
    new_n42546_, new_n42547_, new_n42548_, new_n42549_, new_n42550_,
    new_n42551_, new_n42552_, new_n42553_, new_n42554_, new_n42555_,
    new_n42556_, new_n42557_, new_n42558_, new_n42559_, new_n42560_,
    new_n42561_, new_n42562_, new_n42563_, new_n42564_, new_n42565_,
    new_n42566_, new_n42567_, new_n42568_, new_n42569_, new_n42570_,
    new_n42571_, new_n42572_, new_n42573_, new_n42574_, new_n42575_,
    new_n42576_, new_n42577_, new_n42578_, new_n42579_, new_n42580_,
    new_n42581_, new_n42582_, new_n42583_, new_n42584_, new_n42585_,
    new_n42586_, new_n42587_, new_n42588_, new_n42589_, new_n42590_,
    new_n42591_, new_n42592_, new_n42593_, new_n42594_, new_n42595_,
    new_n42596_, new_n42597_, new_n42598_, new_n42599_, new_n42600_,
    new_n42601_, new_n42602_, new_n42603_, new_n42604_, new_n42605_,
    new_n42606_, new_n42607_, new_n42608_, new_n42609_, new_n42610_,
    new_n42611_, new_n42612_, new_n42613_, new_n42614_, new_n42615_,
    new_n42616_, new_n42617_, new_n42618_, new_n42619_, new_n42620_,
    new_n42621_, new_n42622_, new_n42623_, new_n42624_, new_n42625_,
    new_n42626_, new_n42627_, new_n42628_, new_n42629_, new_n42630_,
    new_n42631_, new_n42632_, new_n42633_, new_n42634_, new_n42635_,
    new_n42636_, new_n42637_, new_n42638_, new_n42639_, new_n42640_,
    new_n42641_, new_n42642_, new_n42643_, new_n42644_, new_n42645_,
    new_n42646_, new_n42647_, new_n42648_, new_n42649_, new_n42650_,
    new_n42651_, new_n42652_, new_n42653_, new_n42654_, new_n42655_,
    new_n42656_, new_n42657_, new_n42658_, new_n42659_, new_n42660_,
    new_n42661_, new_n42662_, new_n42663_, new_n42664_, new_n42665_,
    new_n42666_, new_n42667_, new_n42668_, new_n42669_, new_n42670_,
    new_n42671_, new_n42672_, new_n42673_, new_n42674_, new_n42675_,
    new_n42676_, new_n42677_, new_n42678_, new_n42679_, new_n42680_,
    new_n42681_, new_n42682_, new_n42683_, new_n42684_, new_n42685_,
    new_n42686_, new_n42687_, new_n42688_, new_n42689_, new_n42690_,
    new_n42691_, new_n42692_, new_n42693_, new_n42694_, new_n42695_,
    new_n42696_, new_n42697_, new_n42698_, new_n42699_, new_n42700_,
    new_n42701_, new_n42702_, new_n42703_, new_n42704_, new_n42705_,
    new_n42706_, new_n42707_, new_n42708_, new_n42709_, new_n42710_,
    new_n42711_, new_n42712_, new_n42713_, new_n42714_, new_n42715_,
    new_n42716_, new_n42717_, new_n42718_, new_n42719_, new_n42720_,
    new_n42721_, new_n42722_, new_n42723_, new_n42724_, new_n42725_,
    new_n42726_, new_n42727_, new_n42728_, new_n42729_, new_n42730_,
    new_n42731_, new_n42732_, new_n42733_, new_n42734_, new_n42735_,
    new_n42736_, new_n42737_, new_n42738_, new_n42739_, new_n42740_,
    new_n42741_, new_n42742_, new_n42743_, new_n42744_, new_n42745_,
    new_n42746_, new_n42747_, new_n42748_, new_n42749_, new_n42750_,
    new_n42751_, new_n42752_, new_n42753_, new_n42754_, new_n42755_,
    new_n42756_, new_n42757_, new_n42758_, new_n42759_, new_n42760_,
    new_n42761_, new_n42762_, new_n42763_, new_n42764_, new_n42765_,
    new_n42766_, new_n42767_, new_n42768_, new_n42769_, new_n42770_,
    new_n42771_, new_n42772_, new_n42773_, new_n42774_, new_n42775_,
    new_n42776_, new_n42777_, new_n42778_, new_n42779_, new_n42780_,
    new_n42781_, new_n42782_, new_n42783_, new_n42784_, new_n42785_,
    new_n42786_, new_n42787_, new_n42788_, new_n42789_, new_n42790_,
    new_n42791_, new_n42792_, new_n42793_, new_n42794_, new_n42795_,
    new_n42796_, new_n42797_, new_n42798_, new_n42799_, new_n42800_,
    new_n42801_, new_n42802_, new_n42803_, new_n42804_, new_n42805_,
    new_n42806_, new_n42807_, new_n42808_, new_n42809_, new_n42810_,
    new_n42811_, new_n42812_, new_n42813_, new_n42814_, new_n42815_,
    new_n42816_, new_n42817_, new_n42818_, new_n42819_, new_n42820_,
    new_n42821_, new_n42822_, new_n42823_, new_n42824_, new_n42825_,
    new_n42826_, new_n42827_, new_n42828_, new_n42829_, new_n42830_,
    new_n42831_, new_n42832_, new_n42833_, new_n42834_, new_n42835_,
    new_n42836_, new_n42837_, new_n42838_, new_n42839_, new_n42840_,
    new_n42841_, new_n42842_, new_n42843_, new_n42844_, new_n42845_,
    new_n42846_, new_n42847_, new_n42848_, new_n42849_, new_n42850_,
    new_n42851_, new_n42852_, new_n42853_, new_n42854_, new_n42855_,
    new_n42856_, new_n42857_, new_n42858_, new_n42859_, new_n42860_,
    new_n42861_, new_n42862_, new_n42863_, new_n42864_, new_n42865_,
    new_n42866_, new_n42867_, new_n42868_, new_n42869_, new_n42870_,
    new_n42871_, new_n42872_, new_n42873_, new_n42874_, new_n42875_,
    new_n42876_, new_n42877_, new_n42878_, new_n42879_, new_n42880_,
    new_n42881_, new_n42882_, new_n42883_, new_n42884_, new_n42885_,
    new_n42886_, new_n42887_, new_n42888_, new_n42889_, new_n42890_,
    new_n42891_, new_n42892_, new_n42893_, new_n42894_, new_n42895_,
    new_n42896_, new_n42897_, new_n42898_, new_n42899_, new_n42900_,
    new_n42901_, new_n42902_, new_n42903_, new_n42904_, new_n42905_,
    new_n42906_, new_n42907_, new_n42908_, new_n42909_, new_n42910_,
    new_n42911_, new_n42912_, new_n42913_, new_n42914_, new_n42915_,
    new_n42916_, new_n42917_, new_n42918_, new_n42919_, new_n42920_,
    new_n42921_, new_n42922_, new_n42923_, new_n42924_, new_n42925_,
    new_n42926_, new_n42927_, new_n42928_, new_n42929_, new_n42930_,
    new_n42931_, new_n42932_, new_n42933_, new_n42934_, new_n42935_,
    new_n42936_, new_n42937_, new_n42938_, new_n42939_, new_n42940_,
    new_n42941_, new_n42942_, new_n42943_, new_n42944_, new_n42945_,
    new_n42946_, new_n42947_, new_n42948_, new_n42949_, new_n42950_,
    new_n42951_, new_n42952_, new_n42953_, new_n42954_, new_n42955_,
    new_n42956_, new_n42957_, new_n42958_, new_n42959_, new_n42960_,
    new_n42961_, new_n42962_, new_n42963_, new_n42964_, new_n42965_,
    new_n42966_, new_n42967_, new_n42968_, new_n42969_, new_n42970_,
    new_n42971_, new_n42972_, new_n42973_, new_n42974_, new_n42975_,
    new_n42976_, new_n42977_, new_n42978_, new_n42979_, new_n42980_,
    new_n42981_, new_n42982_, new_n42983_, new_n42984_, new_n42985_,
    new_n42986_, new_n42987_, new_n42988_, new_n42989_, new_n42990_,
    new_n42991_, new_n42992_, new_n42993_, new_n42994_, new_n42995_,
    new_n42996_, new_n42997_, new_n42998_, new_n42999_, new_n43000_,
    new_n43001_, new_n43002_, new_n43003_, new_n43004_, new_n43005_,
    new_n43006_, new_n43007_, new_n43008_, new_n43009_, new_n43010_,
    new_n43011_, new_n43012_, new_n43013_, new_n43014_, new_n43015_,
    new_n43016_, new_n43017_, new_n43018_, new_n43019_, new_n43020_,
    new_n43021_, new_n43022_, new_n43023_, new_n43024_, new_n43025_,
    new_n43026_, new_n43027_, new_n43028_, new_n43029_, new_n43030_,
    new_n43031_, new_n43032_, new_n43033_, new_n43034_, new_n43035_,
    new_n43036_, new_n43037_, new_n43038_, new_n43039_, new_n43040_,
    new_n43041_, new_n43042_, new_n43043_, new_n43044_, new_n43045_,
    new_n43046_, new_n43047_, new_n43048_, new_n43049_, new_n43050_,
    new_n43051_, new_n43052_, new_n43053_, new_n43054_, new_n43055_,
    new_n43056_, new_n43057_, new_n43058_, new_n43059_, new_n43060_,
    new_n43061_, new_n43062_, new_n43063_, new_n43064_, new_n43065_,
    new_n43066_, new_n43067_, new_n43068_, new_n43069_, new_n43070_,
    new_n43071_, new_n43072_, new_n43073_, new_n43074_, new_n43075_,
    new_n43076_, new_n43077_, new_n43078_, new_n43079_, new_n43080_,
    new_n43081_, new_n43082_, new_n43083_, new_n43084_, new_n43085_,
    new_n43086_, new_n43087_, new_n43088_, new_n43089_, new_n43090_,
    new_n43091_, new_n43092_, new_n43093_, new_n43094_, new_n43095_,
    new_n43096_, new_n43097_, new_n43098_, new_n43099_, new_n43100_,
    new_n43101_, new_n43102_, new_n43103_, new_n43104_, new_n43105_,
    new_n43106_, new_n43107_, new_n43108_, new_n43109_, new_n43110_,
    new_n43111_, new_n43112_, new_n43113_, new_n43114_, new_n43115_,
    new_n43116_, new_n43117_, new_n43118_, new_n43119_, new_n43120_,
    new_n43121_, new_n43122_, new_n43123_, new_n43124_, new_n43125_,
    new_n43126_, new_n43127_, new_n43128_, new_n43129_, new_n43130_,
    new_n43131_, new_n43132_, new_n43133_, new_n43134_, new_n43135_,
    new_n43136_, new_n43137_, new_n43138_, new_n43139_, new_n43140_,
    new_n43141_, new_n43142_, new_n43143_, new_n43144_, new_n43145_,
    new_n43146_, new_n43147_, new_n43148_, new_n43149_, new_n43150_,
    new_n43151_, new_n43152_, new_n43153_, new_n43154_, new_n43155_,
    new_n43156_, new_n43157_, new_n43158_, new_n43159_, new_n43160_,
    new_n43161_, new_n43162_, new_n43163_, new_n43164_, new_n43165_,
    new_n43166_, new_n43167_, new_n43168_, new_n43169_, new_n43170_,
    new_n43171_, new_n43172_, new_n43173_, new_n43174_, new_n43175_,
    new_n43176_, new_n43177_, new_n43178_, new_n43179_, new_n43180_,
    new_n43181_, new_n43182_, new_n43183_, new_n43184_, new_n43185_,
    new_n43186_, new_n43187_, new_n43188_, new_n43189_, new_n43190_,
    new_n43191_, new_n43192_, new_n43193_, new_n43194_, new_n43195_,
    new_n43196_, new_n43197_, new_n43198_, new_n43199_, new_n43200_,
    new_n43201_, new_n43202_, new_n43203_, new_n43204_, new_n43205_,
    new_n43206_, new_n43207_, new_n43208_, new_n43209_, new_n43210_,
    new_n43211_, new_n43212_, new_n43213_, new_n43214_, new_n43215_,
    new_n43216_, new_n43217_, new_n43218_, new_n43219_, new_n43220_,
    new_n43221_, new_n43222_, new_n43223_, new_n43224_, new_n43225_,
    new_n43226_, new_n43227_, new_n43228_, new_n43229_, new_n43230_,
    new_n43231_, new_n43232_, new_n43233_, new_n43234_, new_n43235_,
    new_n43236_, new_n43237_, new_n43238_, new_n43239_, new_n43240_,
    new_n43241_, new_n43242_, new_n43243_, new_n43244_, new_n43245_,
    new_n43246_, new_n43247_, new_n43248_, new_n43249_, new_n43250_,
    new_n43251_, new_n43252_, new_n43253_, new_n43254_, new_n43255_,
    new_n43256_, new_n43257_, new_n43258_, new_n43259_, new_n43260_,
    new_n43261_, new_n43262_, new_n43263_, new_n43264_, new_n43265_,
    new_n43266_, new_n43267_, new_n43268_, new_n43269_, new_n43270_,
    new_n43271_, new_n43272_, new_n43273_, new_n43274_, new_n43275_,
    new_n43276_, new_n43277_, new_n43278_, new_n43279_, new_n43280_,
    new_n43281_, new_n43282_, new_n43283_, new_n43284_, new_n43285_,
    new_n43286_, new_n43287_, new_n43288_, new_n43289_, new_n43290_,
    new_n43291_, new_n43292_, new_n43293_, new_n43294_, new_n43295_,
    new_n43296_, new_n43297_, new_n43298_, new_n43299_, new_n43300_,
    new_n43301_, new_n43302_, new_n43303_, new_n43304_, new_n43305_,
    new_n43306_, new_n43307_, new_n43308_, new_n43309_, new_n43310_,
    new_n43311_, new_n43312_, new_n43313_, new_n43314_, new_n43315_,
    new_n43316_, new_n43317_, new_n43318_, new_n43319_, new_n43320_,
    new_n43321_, new_n43322_, new_n43323_, new_n43324_, new_n43325_,
    new_n43326_, new_n43327_, new_n43328_, new_n43329_, new_n43330_,
    new_n43331_, new_n43332_, new_n43333_, new_n43334_, new_n43335_,
    new_n43336_, new_n43337_, new_n43338_, new_n43339_, new_n43340_,
    new_n43341_, new_n43342_, new_n43343_, new_n43344_, new_n43345_,
    new_n43346_, new_n43347_, new_n43348_, new_n43349_, new_n43350_,
    new_n43351_, new_n43352_, new_n43353_, new_n43354_, new_n43355_,
    new_n43356_, new_n43357_, new_n43358_, new_n43359_, new_n43360_,
    new_n43361_, new_n43362_, new_n43363_, new_n43364_, new_n43365_,
    new_n43366_, new_n43367_, new_n43368_, new_n43369_, new_n43370_,
    new_n43371_, new_n43372_, new_n43373_, new_n43374_, new_n43375_,
    new_n43376_, new_n43377_, new_n43378_, new_n43379_, new_n43380_,
    new_n43381_, new_n43382_, new_n43383_, new_n43384_, new_n43385_,
    new_n43386_, new_n43387_, new_n43388_, new_n43389_, new_n43390_,
    new_n43391_, new_n43392_, new_n43393_, new_n43394_, new_n43395_,
    new_n43396_, new_n43397_, new_n43398_, new_n43399_, new_n43400_,
    new_n43401_, new_n43402_, new_n43403_, new_n43404_, new_n43405_,
    new_n43406_, new_n43407_, new_n43408_, new_n43409_, new_n43410_,
    new_n43411_, new_n43412_, new_n43413_, new_n43414_, new_n43415_,
    new_n43416_, new_n43417_, new_n43418_, new_n43419_, new_n43420_,
    new_n43421_, new_n43422_, new_n43423_, new_n43424_, new_n43425_,
    new_n43426_, new_n43427_, new_n43428_, new_n43429_, new_n43430_,
    new_n43431_, new_n43432_, new_n43433_, new_n43434_, new_n43435_,
    new_n43436_, new_n43437_, new_n43438_, new_n43439_, new_n43440_,
    new_n43441_, new_n43442_, new_n43443_, new_n43444_, new_n43445_,
    new_n43446_, new_n43447_, new_n43448_, new_n43449_, new_n43450_,
    new_n43451_, new_n43452_, new_n43453_, new_n43454_, new_n43455_,
    new_n43456_, new_n43457_, new_n43458_, new_n43459_, new_n43460_,
    new_n43461_, new_n43462_, new_n43463_, new_n43464_, new_n43465_,
    new_n43466_, new_n43467_, new_n43468_, new_n43469_, new_n43470_,
    new_n43471_, new_n43472_, new_n43473_, new_n43474_, new_n43475_,
    new_n43476_, new_n43477_, new_n43478_, new_n43479_, new_n43480_,
    new_n43481_, new_n43482_, new_n43483_, new_n43484_, new_n43485_,
    new_n43486_, new_n43487_, new_n43488_, new_n43489_, new_n43490_,
    new_n43491_, new_n43492_, new_n43493_, new_n43494_, new_n43495_,
    new_n43496_, new_n43497_, new_n43498_, new_n43499_, new_n43500_,
    new_n43501_, new_n43502_, new_n43503_, new_n43504_, new_n43505_,
    new_n43506_, new_n43507_, new_n43508_, new_n43509_, new_n43510_,
    new_n43511_, new_n43512_, new_n43513_, new_n43514_, new_n43515_,
    new_n43516_, new_n43517_, new_n43518_, new_n43519_, new_n43520_,
    new_n43521_, new_n43522_, new_n43523_, new_n43524_, new_n43525_,
    new_n43526_, new_n43527_, new_n43528_, new_n43529_, new_n43530_,
    new_n43531_, new_n43532_, new_n43533_, new_n43534_, new_n43535_,
    new_n43536_, new_n43537_, new_n43538_, new_n43539_, new_n43540_,
    new_n43541_, new_n43542_, new_n43543_, new_n43544_, new_n43545_,
    new_n43546_, new_n43547_, new_n43548_, new_n43549_, new_n43550_,
    new_n43551_, new_n43552_, new_n43553_, new_n43554_, new_n43555_,
    new_n43556_, new_n43557_, new_n43558_, new_n43559_, new_n43560_,
    new_n43561_, new_n43562_, new_n43563_, new_n43564_, new_n43565_,
    new_n43566_, new_n43567_, new_n43568_, new_n43569_, new_n43570_,
    new_n43571_, new_n43572_, new_n43573_, new_n43574_, new_n43575_,
    new_n43576_, new_n43577_, new_n43578_, new_n43579_, new_n43580_,
    new_n43581_, new_n43582_, new_n43583_, new_n43584_, new_n43585_,
    new_n43586_, new_n43587_, new_n43588_, new_n43589_, new_n43590_,
    new_n43591_, new_n43592_, new_n43593_, new_n43594_, new_n43595_,
    new_n43596_, new_n43597_, new_n43598_, new_n43599_, new_n43600_,
    new_n43601_, new_n43602_, new_n43603_, new_n43604_, new_n43605_,
    new_n43606_, new_n43607_, new_n43608_, new_n43609_, new_n43610_,
    new_n43611_, new_n43612_, new_n43613_, new_n43614_, new_n43615_,
    new_n43616_, new_n43617_, new_n43618_, new_n43619_, new_n43620_,
    new_n43621_, new_n43622_, new_n43623_, new_n43624_, new_n43625_,
    new_n43626_, new_n43627_, new_n43628_, new_n43629_, new_n43630_,
    new_n43631_, new_n43632_, new_n43633_, new_n43634_, new_n43635_,
    new_n43636_, new_n43637_, new_n43638_, new_n43639_, new_n43640_,
    new_n43641_, new_n43642_, new_n43643_, new_n43644_, new_n43645_,
    new_n43646_, new_n43647_, new_n43648_, new_n43649_, new_n43650_,
    new_n43651_, new_n43652_, new_n43653_, new_n43654_, new_n43655_,
    new_n43656_, new_n43657_, new_n43658_, new_n43659_, new_n43660_,
    new_n43661_, new_n43662_, new_n43663_, new_n43664_, new_n43665_,
    new_n43666_, new_n43667_, new_n43668_, new_n43669_, new_n43670_,
    new_n43671_, new_n43672_, new_n43673_, new_n43674_, new_n43675_,
    new_n43676_, new_n43677_, new_n43678_, new_n43679_, new_n43680_,
    new_n43681_, new_n43682_, new_n43683_, new_n43684_, new_n43685_,
    new_n43686_, new_n43687_, new_n43688_, new_n43689_, new_n43690_,
    new_n43691_, new_n43692_, new_n43693_, new_n43694_, new_n43695_,
    new_n43696_, new_n43697_, new_n43698_, new_n43699_, new_n43700_,
    new_n43701_, new_n43702_, new_n43703_, new_n43704_, new_n43705_,
    new_n43706_, new_n43707_, new_n43708_, new_n43709_, new_n43710_,
    new_n43711_, new_n43712_, new_n43713_, new_n43714_, new_n43715_,
    new_n43716_, new_n43717_, new_n43718_, new_n43719_, new_n43720_,
    new_n43721_, new_n43722_, new_n43723_, new_n43724_, new_n43725_,
    new_n43726_, new_n43727_, new_n43728_, new_n43729_, new_n43730_,
    new_n43731_, new_n43732_, new_n43733_, new_n43734_, new_n43735_,
    new_n43736_, new_n43737_, new_n43738_, new_n43739_, new_n43740_,
    new_n43741_, new_n43742_, new_n43743_, new_n43744_, new_n43745_,
    new_n43746_, new_n43747_, new_n43748_, new_n43749_, new_n43750_,
    new_n43751_, new_n43752_, new_n43753_, new_n43754_, new_n43755_,
    new_n43756_, new_n43757_, new_n43758_, new_n43759_, new_n43760_,
    new_n43761_, new_n43762_, new_n43763_, new_n43764_, new_n43765_,
    new_n43766_, new_n43767_, new_n43768_, new_n43769_, new_n43770_,
    new_n43771_, new_n43772_, new_n43773_, new_n43774_, new_n43775_,
    new_n43776_, new_n43777_, new_n43778_, new_n43779_, new_n43780_,
    new_n43781_, new_n43782_, new_n43783_, new_n43784_, new_n43785_,
    new_n43786_, new_n43787_, new_n43788_, new_n43789_, new_n43790_,
    new_n43791_, new_n43792_, new_n43793_, new_n43794_, new_n43795_,
    new_n43796_, new_n43797_, new_n43798_, new_n43799_, new_n43800_,
    new_n43801_, new_n43802_, new_n43803_, new_n43804_, new_n43805_,
    new_n43806_, new_n43807_, new_n43808_, new_n43809_, new_n43810_,
    new_n43811_, new_n43812_, new_n43813_, new_n43814_, new_n43815_,
    new_n43816_, new_n43817_, new_n43818_, new_n43819_, new_n43820_,
    new_n43821_, new_n43822_, new_n43823_, new_n43824_, new_n43825_,
    new_n43826_, new_n43827_, new_n43828_, new_n43829_, new_n43830_,
    new_n43831_, new_n43832_, new_n43833_, new_n43834_, new_n43835_,
    new_n43836_, new_n43837_, new_n43838_, new_n43839_, new_n43840_,
    new_n43841_, new_n43842_, new_n43843_, new_n43844_, new_n43845_,
    new_n43846_, new_n43847_, new_n43848_, new_n43849_, new_n43850_,
    new_n43851_, new_n43852_, new_n43853_, new_n43854_, new_n43855_,
    new_n43856_, new_n43857_, new_n43858_, new_n43859_, new_n43860_,
    new_n43861_, new_n43862_, new_n43863_, new_n43864_, new_n43865_,
    new_n43866_, new_n43867_, new_n43868_, new_n43869_, new_n43870_,
    new_n43871_, new_n43872_, new_n43873_, new_n43874_, new_n43875_,
    new_n43876_, new_n43877_, new_n43878_, new_n43879_, new_n43880_,
    new_n43881_, new_n43882_, new_n43883_, new_n43884_, new_n43885_,
    new_n43886_, new_n43887_, new_n43888_, new_n43889_, new_n43890_,
    new_n43891_, new_n43892_, new_n43893_, new_n43894_, new_n43895_,
    new_n43896_, new_n43897_, new_n43898_, new_n43899_, new_n43900_,
    new_n43901_, new_n43902_, new_n43903_, new_n43904_, new_n43905_,
    new_n43906_, new_n43907_, new_n43908_, new_n43909_, new_n43910_,
    new_n43911_, new_n43912_, new_n43913_, new_n43914_, new_n43915_,
    new_n43916_, new_n43917_, new_n43918_, new_n43919_, new_n43920_,
    new_n43921_, new_n43922_, new_n43923_, new_n43924_, new_n43925_,
    new_n43926_, new_n43927_, new_n43928_, new_n43929_, new_n43930_,
    new_n43931_, new_n43932_, new_n43933_, new_n43934_, new_n43935_,
    new_n43936_, new_n43937_, new_n43938_, new_n43939_, new_n43940_,
    new_n43941_, new_n43942_, new_n43943_, new_n43944_, new_n43945_,
    new_n43946_, new_n43947_, new_n43948_, new_n43949_, new_n43950_,
    new_n43951_, new_n43952_, new_n43953_, new_n43954_, new_n43955_,
    new_n43956_, new_n43957_, new_n43958_, new_n43959_, new_n43960_,
    new_n43961_, new_n43962_, new_n43963_, new_n43964_, new_n43965_,
    new_n43966_, new_n43967_, new_n43968_, new_n43969_, new_n43970_,
    new_n43971_, new_n43972_, new_n43973_, new_n43974_, new_n43975_,
    new_n43976_, new_n43977_, new_n43978_, new_n43979_, new_n43980_,
    new_n43981_, new_n43982_, new_n43983_, new_n43984_, new_n43985_,
    new_n43986_, new_n43987_, new_n43988_, new_n43989_, new_n43990_,
    new_n43991_, new_n43992_, new_n43993_, new_n43994_, new_n43995_,
    new_n43996_, new_n43997_, new_n43998_, new_n43999_, new_n44000_,
    new_n44001_, new_n44002_, new_n44003_, new_n44004_, new_n44005_,
    new_n44006_, new_n44007_, new_n44008_, new_n44009_, new_n44010_,
    new_n44011_, new_n44012_, new_n44013_, new_n44014_, new_n44015_,
    new_n44016_, new_n44017_, new_n44018_, new_n44019_, new_n44020_,
    new_n44021_, new_n44022_, new_n44023_, new_n44024_, new_n44025_,
    new_n44026_, new_n44027_, new_n44028_, new_n44029_, new_n44030_,
    new_n44031_, new_n44032_, new_n44033_, new_n44034_, new_n44035_,
    new_n44036_, new_n44037_, new_n44038_, new_n44039_, new_n44040_,
    new_n44041_, new_n44042_, new_n44043_, new_n44044_, new_n44045_,
    new_n44046_, new_n44047_, new_n44048_, new_n44049_, new_n44050_,
    new_n44051_, new_n44052_, new_n44053_, new_n44054_, new_n44055_,
    new_n44056_, new_n44057_, new_n44058_, new_n44059_, new_n44060_,
    new_n44061_, new_n44062_, new_n44063_, new_n44064_, new_n44065_,
    new_n44066_, new_n44067_, new_n44068_, new_n44069_, new_n44070_,
    new_n44071_, new_n44072_, new_n44073_, new_n44074_, new_n44075_,
    new_n44076_, new_n44077_, new_n44078_, new_n44079_, new_n44080_,
    new_n44081_, new_n44082_, new_n44083_, new_n44084_, new_n44085_,
    new_n44086_, new_n44087_, new_n44088_, new_n44089_, new_n44090_,
    new_n44091_, new_n44092_, new_n44093_, new_n44094_, new_n44095_,
    new_n44096_, new_n44097_, new_n44098_, new_n44099_, new_n44100_,
    new_n44101_, new_n44102_, new_n44103_, new_n44104_, new_n44105_,
    new_n44106_, new_n44107_, new_n44108_, new_n44109_, new_n44110_,
    new_n44111_, new_n44112_, new_n44113_, new_n44114_, new_n44115_,
    new_n44116_, new_n44117_, new_n44118_, new_n44119_, new_n44120_,
    new_n44121_, new_n44122_, new_n44123_, new_n44124_, new_n44125_,
    new_n44126_, new_n44127_, new_n44128_, new_n44129_, new_n44130_,
    new_n44131_, new_n44132_, new_n44133_, new_n44134_, new_n44135_,
    new_n44136_, new_n44137_, new_n44138_, new_n44139_, new_n44140_,
    new_n44141_, new_n44142_, new_n44143_, new_n44144_, new_n44145_,
    new_n44146_, new_n44147_, new_n44148_, new_n44149_, new_n44150_,
    new_n44151_, new_n44152_, new_n44153_, new_n44154_, new_n44155_,
    new_n44156_, new_n44157_, new_n44158_, new_n44159_, new_n44160_,
    new_n44161_, new_n44162_, new_n44163_, new_n44164_, new_n44165_,
    new_n44166_, new_n44167_, new_n44168_, new_n44169_, new_n44170_,
    new_n44171_, new_n44172_, new_n44173_, new_n44174_, new_n44175_,
    new_n44176_, new_n44177_, new_n44178_, new_n44179_, new_n44180_,
    new_n44181_, new_n44182_, new_n44183_, new_n44184_, new_n44185_,
    new_n44186_, new_n44187_, new_n44188_, new_n44189_, new_n44190_,
    new_n44191_, new_n44192_, new_n44193_, new_n44194_, new_n44195_,
    new_n44196_, new_n44197_, new_n44198_, new_n44199_, new_n44200_,
    new_n44201_, new_n44202_, new_n44203_, new_n44204_, new_n44205_,
    new_n44206_, new_n44207_, new_n44208_, new_n44209_, new_n44210_,
    new_n44211_, new_n44212_, new_n44213_, new_n44214_, new_n44215_,
    new_n44216_, new_n44217_, new_n44218_, new_n44219_, new_n44220_,
    new_n44221_, new_n44222_, new_n44223_, new_n44224_, new_n44225_,
    new_n44226_, new_n44227_, new_n44228_, new_n44229_, new_n44230_,
    new_n44231_, new_n44232_, new_n44233_, new_n44234_, new_n44235_,
    new_n44236_, new_n44237_, new_n44238_, new_n44239_, new_n44240_,
    new_n44241_, new_n44242_, new_n44243_, new_n44244_, new_n44245_,
    new_n44246_, new_n44247_, new_n44248_, new_n44249_, new_n44250_,
    new_n44251_, new_n44252_, new_n44253_, new_n44254_, new_n44255_,
    new_n44256_, new_n44257_, new_n44258_, new_n44259_, new_n44260_,
    new_n44261_, new_n44262_, new_n44263_, new_n44264_, new_n44265_,
    new_n44266_, new_n44267_, new_n44268_, new_n44269_, new_n44270_,
    new_n44271_, new_n44272_, new_n44273_, new_n44274_, new_n44275_,
    new_n44276_, new_n44277_, new_n44278_, new_n44279_, new_n44280_,
    new_n44281_, new_n44282_, new_n44283_, new_n44284_, new_n44285_,
    new_n44286_, new_n44287_, new_n44288_, new_n44289_, new_n44290_,
    new_n44291_, new_n44292_, new_n44293_, new_n44294_, new_n44295_,
    new_n44296_, new_n44297_, new_n44298_, new_n44299_, new_n44300_,
    new_n44301_, new_n44302_, new_n44303_, new_n44304_, new_n44305_,
    new_n44306_, new_n44307_, new_n44308_, new_n44309_, new_n44310_,
    new_n44311_, new_n44312_, new_n44313_, new_n44314_, new_n44315_,
    new_n44316_, new_n44317_, new_n44318_, new_n44319_, new_n44320_,
    new_n44321_, new_n44322_, new_n44323_, new_n44324_, new_n44325_,
    new_n44326_, new_n44327_, new_n44328_, new_n44329_, new_n44330_,
    new_n44331_, new_n44332_, new_n44333_, new_n44334_, new_n44335_,
    new_n44336_, new_n44337_, new_n44338_, new_n44339_, new_n44340_,
    new_n44341_, new_n44342_, new_n44343_, new_n44344_, new_n44345_,
    new_n44346_, new_n44347_, new_n44348_, new_n44349_, new_n44350_,
    new_n44351_, new_n44352_, new_n44353_, new_n44354_, new_n44355_,
    new_n44356_, new_n44357_, new_n44358_, new_n44359_, new_n44360_,
    new_n44361_, new_n44362_, new_n44363_, new_n44364_, new_n44365_,
    new_n44366_, new_n44367_, new_n44368_, new_n44369_, new_n44370_,
    new_n44371_, new_n44372_, new_n44373_, new_n44374_, new_n44375_,
    new_n44376_, new_n44377_, new_n44378_, new_n44379_, new_n44380_,
    new_n44381_, new_n44382_, new_n44383_, new_n44384_, new_n44385_,
    new_n44386_, new_n44387_, new_n44388_, new_n44389_, new_n44390_,
    new_n44391_, new_n44392_, new_n44393_, new_n44394_, new_n44395_,
    new_n44396_, new_n44397_, new_n44398_, new_n44399_, new_n44400_,
    new_n44401_, new_n44402_, new_n44403_, new_n44404_, new_n44405_,
    new_n44406_, new_n44407_, new_n44408_, new_n44409_, new_n44410_,
    new_n44411_, new_n44412_, new_n44413_, new_n44414_, new_n44415_,
    new_n44416_, new_n44417_, new_n44418_, new_n44419_, new_n44420_,
    new_n44421_, new_n44422_, new_n44423_, new_n44424_, new_n44425_,
    new_n44426_, new_n44427_, new_n44428_, new_n44429_, new_n44430_,
    new_n44431_, new_n44432_, new_n44433_, new_n44434_, new_n44435_,
    new_n44436_, new_n44437_, new_n44438_, new_n44439_, new_n44440_,
    new_n44441_, new_n44442_, new_n44443_, new_n44444_, new_n44445_,
    new_n44446_, new_n44447_, new_n44448_, new_n44449_, new_n44450_,
    new_n44451_, new_n44452_, new_n44453_, new_n44454_, new_n44455_,
    new_n44456_, new_n44457_, new_n44458_, new_n44459_, new_n44460_,
    new_n44461_, new_n44462_, new_n44463_, new_n44464_, new_n44465_,
    new_n44466_, new_n44467_, new_n44468_, new_n44469_, new_n44470_,
    new_n44471_, new_n44472_, new_n44473_, new_n44474_, new_n44475_,
    new_n44476_, new_n44477_, new_n44478_, new_n44479_, new_n44480_,
    new_n44481_, new_n44482_, new_n44483_, new_n44484_, new_n44485_,
    new_n44486_, new_n44487_, new_n44488_, new_n44489_, new_n44490_,
    new_n44491_, new_n44492_, new_n44493_, new_n44494_, new_n44495_,
    new_n44496_, new_n44497_, new_n44498_, new_n44499_, new_n44500_,
    new_n44501_, new_n44502_, new_n44503_, new_n44504_, new_n44505_,
    new_n44506_, new_n44507_, new_n44508_, new_n44509_, new_n44510_,
    new_n44511_, new_n44512_, new_n44513_, new_n44514_, new_n44515_,
    new_n44516_, new_n44517_, new_n44518_, new_n44519_, new_n44520_,
    new_n44521_, new_n44522_, new_n44523_, new_n44524_, new_n44525_,
    new_n44526_, new_n44527_, new_n44528_, new_n44529_, new_n44530_,
    new_n44531_, new_n44532_, new_n44533_, new_n44534_, new_n44535_,
    new_n44536_, new_n44537_, new_n44538_, new_n44539_, new_n44540_,
    new_n44541_, new_n44542_, new_n44543_, new_n44544_, new_n44545_,
    new_n44546_, new_n44547_, new_n44548_, new_n44549_, new_n44550_,
    new_n44551_, new_n44552_, new_n44553_, new_n44554_, new_n44555_,
    new_n44556_, new_n44557_, new_n44558_, new_n44559_, new_n44560_,
    new_n44561_, new_n44562_, new_n44563_, new_n44564_, new_n44565_,
    new_n44566_, new_n44567_, new_n44568_, new_n44569_, new_n44570_,
    new_n44571_, new_n44572_, new_n44573_, new_n44574_, new_n44575_,
    new_n44576_, new_n44577_, new_n44578_, new_n44579_, new_n44580_,
    new_n44581_, new_n44582_, new_n44583_, new_n44584_, new_n44585_,
    new_n44586_, new_n44587_, new_n44588_, new_n44589_, new_n44590_,
    new_n44591_, new_n44592_, new_n44593_, new_n44594_, new_n44595_,
    new_n44596_, new_n44597_, new_n44598_, new_n44599_, new_n44600_,
    new_n44601_, new_n44602_, new_n44603_, new_n44604_, new_n44605_,
    new_n44606_, new_n44607_, new_n44608_, new_n44609_, new_n44610_,
    new_n44611_, new_n44612_, new_n44613_, new_n44614_, new_n44615_,
    new_n44616_, new_n44617_, new_n44618_, new_n44619_, new_n44620_,
    new_n44621_, new_n44622_, new_n44623_, new_n44624_, new_n44625_,
    new_n44626_, new_n44627_, new_n44628_, new_n44629_, new_n44630_,
    new_n44631_, new_n44632_, new_n44633_, new_n44634_, new_n44635_,
    new_n44636_, new_n44637_, new_n44638_, new_n44639_, new_n44640_,
    new_n44641_, new_n44642_, new_n44643_, new_n44644_, new_n44645_,
    new_n44646_, new_n44647_, new_n44648_, new_n44649_, new_n44650_,
    new_n44651_, new_n44652_, new_n44653_, new_n44654_, new_n44655_,
    new_n44656_, new_n44657_, new_n44658_, new_n44659_, new_n44660_,
    new_n44661_, new_n44662_, new_n44663_, new_n44664_, new_n44665_,
    new_n44666_, new_n44667_, new_n44668_, new_n44669_, new_n44670_,
    new_n44671_, new_n44672_, new_n44673_, new_n44674_, new_n44675_,
    new_n44676_, new_n44677_, new_n44678_, new_n44679_, new_n44680_,
    new_n44681_, new_n44682_, new_n44683_, new_n44684_, new_n44685_,
    new_n44686_, new_n44687_, new_n44688_, new_n44689_, new_n44690_,
    new_n44691_, new_n44692_, new_n44693_, new_n44694_, new_n44695_,
    new_n44696_, new_n44697_, new_n44698_, new_n44699_, new_n44700_,
    new_n44701_, new_n44702_, new_n44703_, new_n44704_, new_n44705_,
    new_n44706_, new_n44707_, new_n44708_, new_n44709_, new_n44710_,
    new_n44711_, new_n44712_, new_n44713_, new_n44714_, new_n44715_,
    new_n44716_, new_n44717_, new_n44718_, new_n44719_, new_n44720_,
    new_n44721_, new_n44722_, new_n44723_, new_n44724_, new_n44725_,
    new_n44726_, new_n44727_, new_n44728_, new_n44729_, new_n44730_,
    new_n44731_, new_n44732_, new_n44733_, new_n44734_, new_n44735_,
    new_n44736_, new_n44737_, new_n44738_, new_n44739_, new_n44740_,
    new_n44741_, new_n44742_, new_n44743_, new_n44744_, new_n44745_,
    new_n44746_, new_n44747_, new_n44748_, new_n44749_, new_n44750_,
    new_n44751_, new_n44752_, new_n44753_, new_n44754_, new_n44755_,
    new_n44756_, new_n44757_, new_n44758_, new_n44759_, new_n44760_,
    new_n44761_, new_n44762_, new_n44763_, new_n44764_, new_n44765_,
    new_n44766_, new_n44767_, new_n44768_, new_n44769_, new_n44770_,
    new_n44771_, new_n44772_, new_n44773_, new_n44774_, new_n44775_,
    new_n44776_, new_n44777_, new_n44778_, new_n44779_, new_n44780_,
    new_n44781_, new_n44782_, new_n44783_, new_n44784_, new_n44785_,
    new_n44786_, new_n44787_, new_n44788_, new_n44789_, new_n44790_,
    new_n44791_, new_n44792_, new_n44793_, new_n44794_, new_n44795_,
    new_n44796_, new_n44797_, new_n44798_, new_n44799_, new_n44800_,
    new_n44801_, new_n44802_, new_n44803_, new_n44804_, new_n44805_,
    new_n44806_, new_n44807_, new_n44808_, new_n44809_, new_n44810_,
    new_n44811_, new_n44812_, new_n44813_, new_n44814_, new_n44815_,
    new_n44816_, new_n44817_, new_n44818_, new_n44819_, new_n44820_,
    new_n44821_, new_n44822_, new_n44823_, new_n44824_, new_n44825_,
    new_n44826_, new_n44827_, new_n44828_, new_n44829_, new_n44830_,
    new_n44831_, new_n44832_, new_n44833_, new_n44834_, new_n44835_,
    new_n44836_, new_n44837_, new_n44838_, new_n44839_, new_n44840_,
    new_n44841_, new_n44842_, new_n44843_, new_n44844_, new_n44845_,
    new_n44846_, new_n44847_, new_n44848_, new_n44849_, new_n44850_,
    new_n44851_, new_n44852_, new_n44853_, new_n44854_, new_n44855_,
    new_n44856_, new_n44857_, new_n44858_, new_n44859_, new_n44860_,
    new_n44861_, new_n44862_, new_n44863_, new_n44864_, new_n44865_,
    new_n44866_, new_n44867_, new_n44868_, new_n44869_, new_n44870_,
    new_n44871_, new_n44872_, new_n44873_, new_n44874_, new_n44875_,
    new_n44876_, new_n44877_, new_n44878_, new_n44879_, new_n44880_,
    new_n44881_, new_n44882_, new_n44883_, new_n44884_, new_n44885_,
    new_n44886_, new_n44887_, new_n44888_, new_n44889_, new_n44890_,
    new_n44891_, new_n44892_, new_n44893_, new_n44894_, new_n44895_,
    new_n44896_, new_n44897_, new_n44898_, new_n44899_, new_n44900_,
    new_n44901_, new_n44902_, new_n44903_, new_n44904_, new_n44905_,
    new_n44906_, new_n44907_, new_n44908_, new_n44909_, new_n44910_,
    new_n44911_, new_n44912_, new_n44913_, new_n44914_, new_n44915_,
    new_n44916_, new_n44917_, new_n44918_, new_n44919_, new_n44920_,
    new_n44921_, new_n44922_, new_n44923_, new_n44924_, new_n44925_,
    new_n44926_, new_n44927_, new_n44928_, new_n44929_, new_n44930_,
    new_n44931_, new_n44932_, new_n44933_, new_n44934_, new_n44935_,
    new_n44936_, new_n44937_, new_n44938_, new_n44939_, new_n44940_,
    new_n44941_, new_n44942_, new_n44943_, new_n44944_, new_n44945_,
    new_n44946_, new_n44947_, new_n44948_, new_n44949_, new_n44950_,
    new_n44951_, new_n44952_, new_n44953_, new_n44954_, new_n44955_,
    new_n44956_, new_n44957_, new_n44958_, new_n44959_, new_n44960_,
    new_n44961_, new_n44962_, new_n44963_, new_n44964_, new_n44965_,
    new_n44966_, new_n44967_, new_n44968_, new_n44969_, new_n44970_,
    new_n44971_, new_n44972_, new_n44973_, new_n44974_, new_n44975_,
    new_n44976_, new_n44977_, new_n44978_, new_n44979_, new_n44980_,
    new_n44981_, new_n44982_, new_n44983_, new_n44984_, new_n44985_,
    new_n44986_, new_n44987_, new_n44988_, new_n44989_, new_n44990_,
    new_n44991_, new_n44992_, new_n44993_, new_n44994_, new_n44995_,
    new_n44996_, new_n44997_, new_n44998_, new_n44999_, new_n45000_,
    new_n45001_, new_n45002_, new_n45003_, new_n45004_, new_n45005_,
    new_n45006_, new_n45007_, new_n45008_, new_n45009_, new_n45010_,
    new_n45011_, new_n45012_, new_n45013_, new_n45014_, new_n45015_,
    new_n45016_, new_n45017_, new_n45018_, new_n45019_, new_n45020_,
    new_n45021_, new_n45022_, new_n45023_, new_n45024_, new_n45025_,
    new_n45026_, new_n45027_, new_n45028_, new_n45029_, new_n45030_,
    new_n45031_, new_n45032_, new_n45033_, new_n45034_, new_n45035_,
    new_n45036_, new_n45037_, new_n45038_, new_n45039_, new_n45040_,
    new_n45041_, new_n45042_, new_n45043_, new_n45044_, new_n45045_,
    new_n45046_, new_n45047_, new_n45048_, new_n45049_, new_n45050_,
    new_n45051_, new_n45052_, new_n45053_, new_n45054_, new_n45055_,
    new_n45056_, new_n45057_, new_n45058_, new_n45059_, new_n45060_,
    new_n45061_, new_n45062_, new_n45063_, new_n45064_, new_n45065_,
    new_n45066_, new_n45067_, new_n45068_, new_n45069_, new_n45070_,
    new_n45071_, new_n45072_, new_n45073_, new_n45074_, new_n45075_,
    new_n45076_, new_n45077_, new_n45078_, new_n45079_, new_n45080_,
    new_n45081_, new_n45082_, new_n45083_, new_n45084_, new_n45085_,
    new_n45086_, new_n45087_, new_n45088_, new_n45089_, new_n45090_,
    new_n45091_, new_n45092_, new_n45093_, new_n45094_, new_n45095_,
    new_n45096_, new_n45097_, new_n45098_, new_n45099_, new_n45100_,
    new_n45101_, new_n45102_, new_n45103_, new_n45104_, new_n45105_,
    new_n45106_, new_n45107_, new_n45108_, new_n45109_, new_n45110_,
    new_n45111_, new_n45112_, new_n45113_, new_n45114_, new_n45115_,
    new_n45116_, new_n45117_, new_n45118_, new_n45119_, new_n45120_,
    new_n45121_, new_n45122_, new_n45123_, new_n45124_, new_n45125_,
    new_n45126_, new_n45127_, new_n45128_, new_n45129_, new_n45130_,
    new_n45131_, new_n45132_, new_n45133_, new_n45134_, new_n45135_,
    new_n45136_, new_n45137_, new_n45138_, new_n45139_, new_n45140_,
    new_n45141_, new_n45142_, new_n45143_, new_n45144_, new_n45145_,
    new_n45146_, new_n45147_, new_n45148_, new_n45149_, new_n45150_,
    new_n45151_, new_n45152_, new_n45153_, new_n45154_, new_n45155_,
    new_n45156_, new_n45157_, new_n45158_, new_n45159_, new_n45160_,
    new_n45161_, new_n45162_, new_n45163_, new_n45164_, new_n45165_,
    new_n45166_, new_n45167_, new_n45168_, new_n45169_, new_n45170_,
    new_n45171_, new_n45172_, new_n45173_, new_n45174_, new_n45175_,
    new_n45176_, new_n45177_, new_n45178_, new_n45179_, new_n45180_,
    new_n45181_, new_n45182_, new_n45183_, new_n45184_, new_n45185_,
    new_n45186_, new_n45187_, new_n45188_, new_n45189_, new_n45190_,
    new_n45191_, new_n45192_, new_n45193_, new_n45194_, new_n45195_,
    new_n45196_, new_n45197_, new_n45198_, new_n45199_, new_n45200_,
    new_n45201_, new_n45202_, new_n45203_, new_n45204_, new_n45205_,
    new_n45206_, new_n45207_, new_n45208_, new_n45209_, new_n45210_,
    new_n45211_, new_n45212_, new_n45213_, new_n45214_, new_n45215_,
    new_n45216_, new_n45217_, new_n45218_, new_n45219_, new_n45220_,
    new_n45221_, new_n45222_, new_n45223_, new_n45224_, new_n45225_,
    new_n45226_, new_n45227_, new_n45228_, new_n45229_, new_n45230_,
    new_n45231_, new_n45232_, new_n45233_, new_n45234_, new_n45235_,
    new_n45236_, new_n45237_, new_n45238_, new_n45239_, new_n45240_,
    new_n45241_, new_n45242_, new_n45243_, new_n45244_, new_n45245_,
    new_n45246_, new_n45247_, new_n45248_, new_n45249_, new_n45250_,
    new_n45251_, new_n45252_, new_n45253_, new_n45254_, new_n45255_,
    new_n45256_, new_n45257_, new_n45258_, new_n45259_, new_n45260_,
    new_n45261_, new_n45262_, new_n45263_, new_n45264_, new_n45265_,
    new_n45266_, new_n45267_, new_n45268_, new_n45269_, new_n45270_,
    new_n45271_, new_n45272_, new_n45273_, new_n45274_, new_n45275_,
    new_n45276_, new_n45277_, new_n45278_, new_n45279_, new_n45280_,
    new_n45281_, new_n45282_, new_n45283_, new_n45284_, new_n45285_,
    new_n45286_, new_n45287_, new_n45288_, new_n45289_, new_n45290_,
    new_n45291_, new_n45292_, new_n45293_, new_n45294_, new_n45295_,
    new_n45296_, new_n45297_, new_n45298_, new_n45299_, new_n45300_,
    new_n45301_, new_n45302_, new_n45303_, new_n45304_, new_n45305_,
    new_n45306_, new_n45307_, new_n45308_, new_n45309_, new_n45310_,
    new_n45311_, new_n45312_, new_n45313_, new_n45314_, new_n45315_,
    new_n45316_, new_n45317_, new_n45318_, new_n45319_, new_n45320_,
    new_n45321_, new_n45322_, new_n45323_, new_n45324_, new_n45325_,
    new_n45326_, new_n45327_, new_n45328_, new_n45329_, new_n45330_,
    new_n45331_, new_n45332_, new_n45333_, new_n45334_, new_n45335_,
    new_n45336_, new_n45337_, new_n45338_, new_n45339_, new_n45340_,
    new_n45341_, new_n45342_, new_n45343_, new_n45344_, new_n45345_,
    new_n45346_, new_n45347_, new_n45348_, new_n45349_, new_n45350_,
    new_n45351_, new_n45352_, new_n45353_, new_n45354_, new_n45355_,
    new_n45356_, new_n45357_, new_n45358_, new_n45359_, new_n45360_,
    new_n45361_, new_n45362_, new_n45363_, new_n45364_, new_n45365_,
    new_n45366_, new_n45367_, new_n45368_, new_n45369_, new_n45370_,
    new_n45371_, new_n45372_, new_n45373_, new_n45374_, new_n45375_,
    new_n45376_, new_n45377_, new_n45378_, new_n45379_, new_n45380_,
    new_n45381_, new_n45382_, new_n45383_, new_n45384_, new_n45385_,
    new_n45386_, new_n45387_, new_n45388_, new_n45389_, new_n45390_,
    new_n45391_, new_n45392_, new_n45393_, new_n45394_, new_n45395_,
    new_n45396_, new_n45397_, new_n45398_, new_n45399_, new_n45400_,
    new_n45401_, new_n45402_, new_n45403_, new_n45404_, new_n45405_,
    new_n45406_, new_n45407_, new_n45408_, new_n45409_, new_n45410_,
    new_n45411_, new_n45412_, new_n45413_, new_n45414_, new_n45415_,
    new_n45416_, new_n45417_, new_n45418_, new_n45419_, new_n45420_,
    new_n45421_, new_n45422_, new_n45423_, new_n45424_, new_n45425_,
    new_n45426_, new_n45427_, new_n45428_, new_n45429_, new_n45430_,
    new_n45431_, new_n45432_, new_n45433_, new_n45434_, new_n45435_,
    new_n45436_, new_n45437_, new_n45438_, new_n45439_, new_n45440_,
    new_n45441_, new_n45442_, new_n45443_, new_n45444_, new_n45445_,
    new_n45446_, new_n45447_, new_n45448_, new_n45449_, new_n45450_,
    new_n45451_, new_n45452_, new_n45453_, new_n45454_, new_n45455_,
    new_n45456_, new_n45457_, new_n45458_, new_n45459_, new_n45460_,
    new_n45461_, new_n45462_, new_n45463_, new_n45464_, new_n45465_,
    new_n45466_, new_n45467_, new_n45468_, new_n45469_, new_n45470_,
    new_n45471_, new_n45472_, new_n45473_, new_n45474_, new_n45475_,
    new_n45476_, new_n45477_, new_n45478_, new_n45479_, new_n45480_,
    new_n45481_, new_n45482_, new_n45483_, new_n45484_, new_n45485_,
    new_n45486_, new_n45487_, new_n45488_, new_n45489_, new_n45490_,
    new_n45491_, new_n45492_, new_n45493_, new_n45494_, new_n45495_,
    new_n45496_, new_n45497_, new_n45498_, new_n45499_, new_n45500_,
    new_n45501_, new_n45502_, new_n45503_, new_n45504_, new_n45505_,
    new_n45506_, new_n45507_, new_n45508_, new_n45509_, new_n45510_,
    new_n45511_, new_n45512_, new_n45513_, new_n45514_, new_n45515_,
    new_n45516_, new_n45517_, new_n45518_, new_n45519_, new_n45520_,
    new_n45521_, new_n45522_, new_n45523_, new_n45524_, new_n45525_,
    new_n45526_, new_n45527_, new_n45528_, new_n45529_, new_n45530_,
    new_n45531_, new_n45532_, new_n45533_, new_n45534_, new_n45535_,
    new_n45536_, new_n45537_, new_n45538_, new_n45539_, new_n45540_,
    new_n45541_, new_n45542_, new_n45543_, new_n45544_, new_n45545_,
    new_n45546_, new_n45547_, new_n45548_, new_n45549_, new_n45550_,
    new_n45551_, new_n45552_, new_n45553_, new_n45554_, new_n45555_,
    new_n45556_, new_n45557_, new_n45558_, new_n45559_, new_n45560_,
    new_n45561_, new_n45562_, new_n45563_, new_n45564_, new_n45565_,
    new_n45566_, new_n45567_, new_n45568_, new_n45569_, new_n45570_,
    new_n45571_, new_n45572_, new_n45573_, new_n45574_, new_n45575_,
    new_n45576_, new_n45577_, new_n45578_, new_n45579_, new_n45580_,
    new_n45581_, new_n45582_, new_n45583_, new_n45584_, new_n45585_,
    new_n45586_, new_n45587_, new_n45588_, new_n45589_, new_n45590_,
    new_n45591_, new_n45592_, new_n45593_, new_n45594_, new_n45595_,
    new_n45596_, new_n45597_, new_n45598_, new_n45599_, new_n45600_,
    new_n45601_, new_n45602_, new_n45603_, new_n45604_, new_n45605_,
    new_n45606_, new_n45607_, new_n45608_, new_n45609_, new_n45610_,
    new_n45611_, new_n45612_, new_n45613_, new_n45614_, new_n45615_,
    new_n45616_, new_n45617_, new_n45618_, new_n45619_, new_n45620_,
    new_n45621_, new_n45622_, new_n45623_, new_n45624_, new_n45625_,
    new_n45626_, new_n45627_, new_n45628_, new_n45629_, new_n45630_,
    new_n45631_, new_n45632_, new_n45633_, new_n45634_, new_n45635_,
    new_n45636_, new_n45637_, new_n45638_, new_n45639_, new_n45640_,
    new_n45641_, new_n45642_, new_n45643_, new_n45644_, new_n45645_,
    new_n45646_, new_n45647_, new_n45648_, new_n45649_, new_n45650_,
    new_n45651_, new_n45652_, new_n45653_, new_n45654_, new_n45655_,
    new_n45656_, new_n45657_, new_n45658_, new_n45659_, new_n45660_,
    new_n45661_, new_n45662_, new_n45663_, new_n45664_, new_n45665_,
    new_n45666_, new_n45667_, new_n45668_, new_n45669_, new_n45670_,
    new_n45671_, new_n45672_, new_n45673_, new_n45674_, new_n45675_,
    new_n45676_, new_n45677_, new_n45678_, new_n45679_, new_n45680_,
    new_n45681_, new_n45682_, new_n45683_, new_n45684_, new_n45685_,
    new_n45686_, new_n45687_, new_n45688_, new_n45689_, new_n45690_,
    new_n45691_, new_n45692_, new_n45693_, new_n45694_, new_n45695_,
    new_n45696_, new_n45697_, new_n45698_, new_n45699_, new_n45700_,
    new_n45701_, new_n45702_, new_n45703_, new_n45704_, new_n45705_,
    new_n45706_, new_n45707_, new_n45708_, new_n45709_, new_n45710_,
    new_n45711_, new_n45712_, new_n45713_, new_n45714_, new_n45715_,
    new_n45716_, new_n45717_, new_n45718_, new_n45719_, new_n45720_,
    new_n45721_, new_n45722_, new_n45723_, new_n45724_, new_n45725_,
    new_n45726_, new_n45727_, new_n45728_, new_n45729_, new_n45730_,
    new_n45731_, new_n45732_, new_n45733_, new_n45734_, new_n45735_,
    new_n45736_, new_n45737_, new_n45738_, new_n45739_, new_n45740_,
    new_n45741_, new_n45742_, new_n45743_, new_n45744_, new_n45745_,
    new_n45746_, new_n45747_, new_n45748_, new_n45749_, new_n45750_,
    new_n45751_, new_n45752_, new_n45753_, new_n45754_, new_n45755_,
    new_n45756_, new_n45757_, new_n45758_, new_n45759_, new_n45760_,
    new_n45761_, new_n45762_, new_n45763_, new_n45764_, new_n45765_,
    new_n45766_, new_n45767_, new_n45768_, new_n45769_, new_n45770_,
    new_n45771_, new_n45772_, new_n45773_, new_n45774_, new_n45775_,
    new_n45776_, new_n45777_, new_n45778_, new_n45779_, new_n45780_,
    new_n45781_, new_n45782_, new_n45783_, new_n45784_, new_n45785_,
    new_n45786_, new_n45787_, new_n45788_, new_n45789_, new_n45790_,
    new_n45791_, new_n45792_, new_n45793_, new_n45794_, new_n45795_,
    new_n45796_, new_n45797_, new_n45798_, new_n45799_, new_n45800_,
    new_n45801_, new_n45802_, new_n45803_, new_n45804_, new_n45805_,
    new_n45806_, new_n45807_, new_n45808_, new_n45809_, new_n45810_,
    new_n45811_, new_n45812_, new_n45813_, new_n45814_, new_n45815_,
    new_n45816_, new_n45817_, new_n45818_, new_n45819_, new_n45820_,
    new_n45821_, new_n45822_, new_n45823_, new_n45824_, new_n45825_,
    new_n45826_, new_n45827_, new_n45828_, new_n45829_, new_n45830_,
    new_n45831_, new_n45832_, new_n45833_, new_n45834_, new_n45835_,
    new_n45836_, new_n45837_, new_n45838_, new_n45839_, new_n45840_,
    new_n45841_, new_n45842_, new_n45843_, new_n45844_, new_n45845_,
    new_n45846_, new_n45847_, new_n45848_, new_n45849_, new_n45850_,
    new_n45851_, new_n45852_, new_n45853_, new_n45854_, new_n45855_,
    new_n45856_, new_n45857_, new_n45858_, new_n45859_, new_n45860_,
    new_n45861_, new_n45862_, new_n45863_, new_n45864_, new_n45865_,
    new_n45866_, new_n45867_, new_n45868_, new_n45869_, new_n45870_,
    new_n45871_, new_n45872_, new_n45873_, new_n45874_, new_n45875_,
    new_n45876_, new_n45877_, new_n45878_, new_n45879_, new_n45880_,
    new_n45881_, new_n45882_, new_n45883_, new_n45884_, new_n45885_,
    new_n45886_, new_n45887_, new_n45888_, new_n45889_, new_n45890_,
    new_n45891_, new_n45892_, new_n45893_, new_n45894_, new_n45895_,
    new_n45896_, new_n45897_, new_n45898_, new_n45899_, new_n45900_,
    new_n45901_, new_n45902_, new_n45903_, new_n45904_, new_n45905_,
    new_n45906_, new_n45907_, new_n45908_, new_n45909_, new_n45910_,
    new_n45911_, new_n45912_, new_n45913_, new_n45914_, new_n45915_,
    new_n45916_, new_n45917_, new_n45918_, new_n45919_, new_n45920_,
    new_n45921_, new_n45922_, new_n45923_, new_n45924_, new_n45925_,
    new_n45926_, new_n45927_, new_n45928_, new_n45929_, new_n45930_,
    new_n45931_, new_n45932_, new_n45933_, new_n45934_, new_n45935_,
    new_n45936_, new_n45937_, new_n45938_, new_n45939_, new_n45940_,
    new_n45941_, new_n45942_, new_n45943_, new_n45944_, new_n45945_,
    new_n45946_, new_n45947_, new_n45948_, new_n45949_, new_n45950_,
    new_n45951_, new_n45952_, new_n45953_, new_n45954_, new_n45955_,
    new_n45956_, new_n45957_, new_n45958_, new_n45959_, new_n45960_,
    new_n45961_, new_n45962_, new_n45963_, new_n45964_, new_n45965_,
    new_n45966_, new_n45967_, new_n45968_, new_n45969_, new_n45970_,
    new_n45971_, new_n45972_, new_n45973_, new_n45974_, new_n45975_,
    new_n45976_, new_n45977_, new_n45978_, new_n45979_, new_n45980_,
    new_n45981_, new_n45982_, new_n45983_, new_n45984_, new_n45985_,
    new_n45986_, new_n45987_, new_n45988_, new_n45989_, new_n45990_,
    new_n45991_, new_n45992_, new_n45993_, new_n45994_, new_n45995_,
    new_n45996_, new_n45997_, new_n45998_, new_n45999_, new_n46000_,
    new_n46001_, new_n46002_, new_n46003_, new_n46004_, new_n46005_,
    new_n46006_, new_n46007_, new_n46008_, new_n46009_, new_n46010_,
    new_n46011_, new_n46012_, new_n46013_, new_n46014_, new_n46015_,
    new_n46016_, new_n46017_, new_n46018_, new_n46019_, new_n46020_,
    new_n46021_, new_n46022_, new_n46023_, new_n46024_, new_n46025_,
    new_n46026_, new_n46027_, new_n46028_, new_n46029_, new_n46030_,
    new_n46031_, new_n46032_, new_n46033_, new_n46034_, new_n46035_,
    new_n46036_, new_n46037_, new_n46038_, new_n46039_, new_n46040_,
    new_n46041_, new_n46042_, new_n46043_, new_n46044_, new_n46045_,
    new_n46046_, new_n46047_, new_n46048_, new_n46049_, new_n46050_,
    new_n46051_, new_n46052_, new_n46053_, new_n46054_, new_n46055_,
    new_n46056_, new_n46057_, new_n46058_, new_n46059_, new_n46060_,
    new_n46061_, new_n46062_, new_n46063_, new_n46064_, new_n46065_,
    new_n46066_, new_n46067_, new_n46068_, new_n46069_, new_n46070_,
    new_n46071_, new_n46072_, new_n46073_, new_n46074_, new_n46075_,
    new_n46076_, new_n46077_, new_n46078_, new_n46079_, new_n46080_,
    new_n46081_, new_n46082_, new_n46083_, new_n46084_, new_n46085_,
    new_n46086_, new_n46087_, new_n46088_, new_n46089_, new_n46090_,
    new_n46091_, new_n46092_, new_n46093_, new_n46094_, new_n46095_,
    new_n46096_, new_n46097_, new_n46098_, new_n46099_, new_n46100_,
    new_n46101_, new_n46102_, new_n46103_, new_n46104_, new_n46105_,
    new_n46106_, new_n46107_, new_n46108_, new_n46109_, new_n46110_,
    new_n46111_, new_n46112_, new_n46113_, new_n46114_, new_n46115_,
    new_n46116_, new_n46117_, new_n46118_, new_n46119_, new_n46120_,
    new_n46121_, new_n46122_, new_n46123_, new_n46124_, new_n46125_,
    new_n46126_, new_n46127_, new_n46128_, new_n46129_, new_n46130_,
    new_n46131_, new_n46132_, new_n46133_, new_n46134_, new_n46135_,
    new_n46136_, new_n46137_, new_n46138_, new_n46139_, new_n46140_,
    new_n46141_, new_n46142_, new_n46143_, new_n46144_, new_n46145_,
    new_n46146_, new_n46147_, new_n46148_, new_n46149_, new_n46150_,
    new_n46151_, new_n46152_, new_n46153_, new_n46154_, new_n46155_,
    new_n46156_, new_n46157_, new_n46158_, new_n46159_, new_n46160_,
    new_n46161_, new_n46162_, new_n46163_, new_n46164_, new_n46165_,
    new_n46166_, new_n46167_, new_n46168_, new_n46169_, new_n46170_,
    new_n46171_, new_n46172_, new_n46173_, new_n46174_, new_n46175_,
    new_n46176_, new_n46177_, new_n46178_, new_n46179_, new_n46180_,
    new_n46181_, new_n46182_, new_n46183_, new_n46184_, new_n46185_,
    new_n46186_, new_n46187_, new_n46188_, new_n46189_, new_n46190_,
    new_n46191_, new_n46192_, new_n46193_, new_n46194_, new_n46195_,
    new_n46196_, new_n46197_, new_n46198_, new_n46199_, new_n46200_,
    new_n46201_, new_n46202_, new_n46203_, new_n46204_, new_n46205_,
    new_n46206_, new_n46207_, new_n46208_, new_n46209_, new_n46210_,
    new_n46211_, new_n46212_, new_n46213_, new_n46214_, new_n46215_,
    new_n46216_, new_n46217_, new_n46218_, new_n46219_, new_n46220_,
    new_n46221_, new_n46222_, new_n46223_, new_n46224_, new_n46225_,
    new_n46226_, new_n46227_, new_n46228_, new_n46229_, new_n46230_,
    new_n46231_, new_n46232_, new_n46233_, new_n46234_, new_n46235_,
    new_n46236_, new_n46237_, new_n46238_, new_n46239_, new_n46240_,
    new_n46241_, new_n46242_, new_n46243_, new_n46244_, new_n46245_,
    new_n46246_, new_n46247_, new_n46248_, new_n46249_, new_n46250_,
    new_n46251_, new_n46252_, new_n46253_, new_n46254_, new_n46255_,
    new_n46256_, new_n46257_, new_n46258_, new_n46259_, new_n46260_,
    new_n46261_, new_n46262_, new_n46263_, new_n46264_, new_n46265_,
    new_n46266_, new_n46267_, new_n46268_, new_n46269_, new_n46270_,
    new_n46271_, new_n46272_, new_n46273_, new_n46274_, new_n46275_,
    new_n46276_, new_n46277_, new_n46278_, new_n46279_, new_n46280_,
    new_n46281_, new_n46282_, new_n46283_, new_n46284_, new_n46285_,
    new_n46286_, new_n46287_, new_n46288_, new_n46289_, new_n46290_,
    new_n46291_, new_n46292_, new_n46293_, new_n46294_, new_n46295_,
    new_n46296_, new_n46297_, new_n46298_, new_n46299_, new_n46300_,
    new_n46301_, new_n46302_, new_n46303_, new_n46304_, new_n46305_,
    new_n46306_, new_n46307_, new_n46308_, new_n46309_, new_n46310_,
    new_n46311_, new_n46312_, new_n46313_, new_n46314_, new_n46315_,
    new_n46316_, new_n46317_, new_n46318_, new_n46319_, new_n46320_,
    new_n46321_, new_n46322_, new_n46323_, new_n46324_, new_n46325_,
    new_n46326_, new_n46327_, new_n46328_, new_n46329_, new_n46330_,
    new_n46331_, new_n46332_, new_n46333_, new_n46334_, new_n46335_,
    new_n46336_, new_n46337_, new_n46338_, new_n46339_, new_n46340_,
    new_n46341_, new_n46342_, new_n46343_, new_n46344_, new_n46345_,
    new_n46346_, new_n46347_, new_n46348_, new_n46349_, new_n46350_,
    new_n46351_, new_n46352_, new_n46353_, new_n46354_, new_n46355_,
    new_n46356_, new_n46357_, new_n46358_, new_n46359_, new_n46360_,
    new_n46361_, new_n46362_, new_n46363_, new_n46364_, new_n46365_,
    new_n46366_, new_n46367_, new_n46368_, new_n46369_, new_n46370_,
    new_n46371_, new_n46372_, new_n46373_, new_n46374_, new_n46375_,
    new_n46376_, new_n46377_, new_n46378_, new_n46379_, new_n46380_,
    new_n46381_, new_n46382_, new_n46383_, new_n46384_, new_n46385_,
    new_n46386_, new_n46387_, new_n46388_, new_n46389_, new_n46390_,
    new_n46391_, new_n46392_, new_n46393_, new_n46394_, new_n46395_,
    new_n46396_, new_n46397_, new_n46398_, new_n46399_, new_n46400_,
    new_n46401_, new_n46402_, new_n46403_, new_n46404_, new_n46405_,
    new_n46406_, new_n46407_, new_n46408_, new_n46409_, new_n46410_,
    new_n46411_, new_n46412_, new_n46413_, new_n46414_, new_n46415_,
    new_n46416_, new_n46417_, new_n46418_, new_n46419_, new_n46420_,
    new_n46421_, new_n46422_, new_n46423_, new_n46424_, new_n46425_,
    new_n46426_, new_n46427_, new_n46428_, new_n46429_, new_n46430_,
    new_n46431_, new_n46432_, new_n46433_, new_n46434_, new_n46435_,
    new_n46436_, new_n46437_, new_n46438_, new_n46439_, new_n46440_,
    new_n46441_, new_n46442_, new_n46443_, new_n46444_, new_n46445_,
    new_n46446_, new_n46447_, new_n46448_, new_n46449_, new_n46450_,
    new_n46451_, new_n46452_, new_n46453_, new_n46454_, new_n46455_,
    new_n46456_, new_n46457_, new_n46458_, new_n46459_, new_n46460_,
    new_n46461_, new_n46462_, new_n46463_, new_n46464_, new_n46465_,
    new_n46466_, new_n46467_, new_n46468_, new_n46469_, new_n46470_,
    new_n46471_, new_n46472_, new_n46473_, new_n46474_, new_n46475_,
    new_n46476_, new_n46477_, new_n46478_, new_n46479_, new_n46480_,
    new_n46481_, new_n46482_, new_n46483_, new_n46484_, new_n46485_,
    new_n46486_, new_n46487_, new_n46488_, new_n46489_, new_n46490_,
    new_n46491_, new_n46492_, new_n46493_, new_n46494_, new_n46495_,
    new_n46496_, new_n46497_, new_n46498_, new_n46499_, new_n46500_,
    new_n46501_, new_n46502_, new_n46503_, new_n46504_, new_n46505_,
    new_n46506_, new_n46507_, new_n46508_, new_n46509_, new_n46510_,
    new_n46511_, new_n46512_, new_n46513_, new_n46514_, new_n46515_,
    new_n46516_, new_n46517_, new_n46518_, new_n46519_, new_n46520_,
    new_n46521_, new_n46522_, new_n46523_, new_n46524_, new_n46525_,
    new_n46526_, new_n46527_, new_n46528_, new_n46529_, new_n46530_,
    new_n46531_, new_n46532_, new_n46533_, new_n46534_, new_n46535_,
    new_n46536_, new_n46537_, new_n46538_, new_n46539_, new_n46540_,
    new_n46541_, new_n46542_, new_n46543_, new_n46544_, new_n46545_,
    new_n46546_, new_n46547_, new_n46548_, new_n46549_, new_n46550_,
    new_n46551_, new_n46552_, new_n46553_, new_n46554_, new_n46555_,
    new_n46556_, new_n46557_, new_n46558_, new_n46559_, new_n46560_,
    new_n46561_, new_n46562_, new_n46563_, new_n46564_, new_n46565_,
    new_n46566_, new_n46567_, new_n46568_, new_n46569_, new_n46570_,
    new_n46571_, new_n46572_, new_n46573_, new_n46574_, new_n46575_,
    new_n46576_, new_n46577_, new_n46578_, new_n46579_, new_n46580_,
    new_n46581_, new_n46582_, new_n46583_, new_n46584_, new_n46585_,
    new_n46586_, new_n46587_, new_n46588_, new_n46589_, new_n46590_,
    new_n46591_, new_n46592_, new_n46593_, new_n46594_, new_n46595_,
    new_n46596_, new_n46597_, new_n46598_, new_n46599_, new_n46600_,
    new_n46601_, new_n46602_, new_n46603_, new_n46604_, new_n46605_,
    new_n46606_, new_n46607_, new_n46608_, new_n46609_, new_n46610_,
    new_n46611_, new_n46612_, new_n46613_, new_n46614_, new_n46615_,
    new_n46616_, new_n46617_, new_n46618_, new_n46619_, new_n46620_,
    new_n46621_, new_n46622_, new_n46623_, new_n46624_, new_n46625_,
    new_n46626_, new_n46627_, new_n46628_, new_n46629_, new_n46630_,
    new_n46631_, new_n46632_, new_n46633_, new_n46634_, new_n46635_,
    new_n46636_, new_n46637_, new_n46638_, new_n46639_, new_n46640_,
    new_n46641_, new_n46642_, new_n46643_, new_n46644_, new_n46645_,
    new_n46646_, new_n46647_, new_n46648_, new_n46649_, new_n46650_,
    new_n46651_, new_n46652_, new_n46653_, new_n46654_, new_n46655_,
    new_n46656_, new_n46657_, new_n46658_, new_n46659_, new_n46660_,
    new_n46661_, new_n46662_, new_n46663_, new_n46664_, new_n46665_,
    new_n46666_, new_n46667_, new_n46668_, new_n46669_, new_n46670_,
    new_n46671_, new_n46672_, new_n46673_, new_n46674_, new_n46675_,
    new_n46676_, new_n46677_, new_n46678_, new_n46679_, new_n46680_,
    new_n46681_, new_n46682_, new_n46683_, new_n46684_, new_n46685_,
    new_n46686_, new_n46687_, new_n46688_, new_n46689_, new_n46690_,
    new_n46691_, new_n46692_, new_n46693_, new_n46694_, new_n46695_,
    new_n46696_, new_n46697_, new_n46698_, new_n46699_, new_n46700_,
    new_n46701_, new_n46702_, new_n46703_, new_n46704_, new_n46705_,
    new_n46706_, new_n46707_, new_n46708_, new_n46709_, new_n46710_,
    new_n46711_, new_n46712_, new_n46713_, new_n46714_, new_n46715_,
    new_n46716_, new_n46717_, new_n46718_, new_n46719_, new_n46720_,
    new_n46721_, new_n46722_, new_n46723_, new_n46724_, new_n46725_,
    new_n46726_, new_n46727_, new_n46728_, new_n46729_, new_n46730_,
    new_n46731_, new_n46732_, new_n46733_, new_n46734_, new_n46735_,
    new_n46736_, new_n46737_, new_n46738_, new_n46739_, new_n46740_,
    new_n46741_, new_n46742_, new_n46743_, new_n46744_, new_n46745_,
    new_n46746_, new_n46747_, new_n46748_, new_n46749_, new_n46750_,
    new_n46751_, new_n46752_, new_n46753_, new_n46754_, new_n46755_,
    new_n46756_, new_n46757_, new_n46758_, new_n46759_, new_n46760_,
    new_n46761_, new_n46762_, new_n46763_, new_n46764_, new_n46765_,
    new_n46766_, new_n46767_, new_n46768_, new_n46769_, new_n46770_,
    new_n46771_, new_n46772_, new_n46773_, new_n46774_, new_n46775_,
    new_n46776_, new_n46777_, new_n46778_, new_n46779_, new_n46780_,
    new_n46781_, new_n46782_, new_n46783_, new_n46784_, new_n46785_,
    new_n46786_, new_n46787_, new_n46788_, new_n46789_, new_n46790_,
    new_n46791_, new_n46792_, new_n46793_, new_n46794_, new_n46795_,
    new_n46796_, new_n46797_, new_n46798_, new_n46799_, new_n46800_,
    new_n46801_, new_n46802_, new_n46803_, new_n46804_, new_n46805_,
    new_n46806_, new_n46807_, new_n46808_, new_n46809_, new_n46810_,
    new_n46811_, new_n46812_, new_n46813_, new_n46814_, new_n46815_,
    new_n46816_, new_n46817_, new_n46818_, new_n46819_, new_n46820_,
    new_n46821_, new_n46822_, new_n46823_, new_n46824_, new_n46825_,
    new_n46826_, new_n46827_, new_n46828_, new_n46829_, new_n46830_,
    new_n46831_, new_n46832_, new_n46833_, new_n46834_, new_n46835_,
    new_n46836_, new_n46837_, new_n46838_, new_n46839_, new_n46840_,
    new_n46841_, new_n46842_, new_n46843_, new_n46844_, new_n46845_,
    new_n46846_, new_n46847_, new_n46848_, new_n46849_, new_n46850_,
    new_n46851_, new_n46852_, new_n46853_, new_n46854_, new_n46855_,
    new_n46856_, new_n46857_, new_n46858_, new_n46859_, new_n46860_,
    new_n46861_, new_n46862_, new_n46863_, new_n46864_, new_n46865_,
    new_n46866_, new_n46867_, new_n46868_, new_n46869_, new_n46870_,
    new_n46871_, new_n46872_, new_n46873_, new_n46874_, new_n46875_,
    new_n46876_, new_n46877_, new_n46878_, new_n46879_, new_n46880_,
    new_n46881_, new_n46882_, new_n46883_, new_n46884_, new_n46885_,
    new_n46886_, new_n46887_, new_n46888_, new_n46889_, new_n46890_,
    new_n46891_, new_n46892_, new_n46893_, new_n46894_, new_n46895_,
    new_n46896_, new_n46897_, new_n46898_, new_n46899_, new_n46900_,
    new_n46901_, new_n46902_, new_n46903_, new_n46904_, new_n46905_,
    new_n46906_, new_n46907_, new_n46908_, new_n46909_, new_n46910_,
    new_n46911_, new_n46912_, new_n46913_, new_n46914_, new_n46915_,
    new_n46916_, new_n46917_, new_n46918_, new_n46919_, new_n46920_,
    new_n46921_, new_n46922_, new_n46923_, new_n46924_, new_n46925_,
    new_n46926_, new_n46927_, new_n46928_, new_n46929_, new_n46930_,
    new_n46931_, new_n46932_, new_n46933_, new_n46934_, new_n46935_,
    new_n46936_, new_n46937_, new_n46938_, new_n46939_, new_n46940_,
    new_n46941_, new_n46942_, new_n46943_, new_n46944_, new_n46945_,
    new_n46946_, new_n46947_, new_n46948_, new_n46949_, new_n46950_,
    new_n46951_, new_n46952_, new_n46953_, new_n46954_, new_n46955_,
    new_n46956_, new_n46957_, new_n46958_, new_n46959_, new_n46960_,
    new_n46961_, new_n46962_, new_n46963_, new_n46964_, new_n46965_,
    new_n46966_, new_n46967_, new_n46968_, new_n46969_, new_n46970_,
    new_n46971_, new_n46972_, new_n46973_, new_n46974_, new_n46975_,
    new_n46976_, new_n46977_, new_n46978_, new_n46979_, new_n46980_,
    new_n46981_, new_n46982_, new_n46983_, new_n46984_, new_n46985_,
    new_n46986_, new_n46987_, new_n46988_, new_n46989_, new_n46990_,
    new_n46991_, new_n46992_, new_n46993_, new_n46994_, new_n46995_,
    new_n46996_, new_n46997_, new_n46998_, new_n46999_, new_n47000_,
    new_n47001_, new_n47002_, new_n47003_, new_n47004_, new_n47005_,
    new_n47006_, new_n47007_, new_n47008_, new_n47009_, new_n47010_,
    new_n47011_, new_n47012_, new_n47013_, new_n47014_, new_n47015_,
    new_n47016_, new_n47017_, new_n47018_, new_n47019_, new_n47020_,
    new_n47021_, new_n47022_, new_n47023_, new_n47024_, new_n47025_,
    new_n47026_, new_n47027_, new_n47028_, new_n47029_, new_n47030_,
    new_n47031_, new_n47032_, new_n47033_, new_n47034_, new_n47035_,
    new_n47036_, new_n47037_, new_n47038_, new_n47039_, new_n47040_,
    new_n47041_, new_n47042_, new_n47043_, new_n47044_, new_n47045_,
    new_n47046_, new_n47047_, new_n47048_, new_n47049_, new_n47050_,
    new_n47051_, new_n47052_, new_n47053_, new_n47054_, new_n47055_,
    new_n47056_, new_n47057_, new_n47058_, new_n47059_, new_n47060_,
    new_n47061_, new_n47062_, new_n47063_, new_n47064_, new_n47065_,
    new_n47066_, new_n47067_, new_n47068_, new_n47069_, new_n47070_,
    new_n47071_, new_n47072_, new_n47073_, new_n47074_, new_n47075_,
    new_n47076_, new_n47077_, new_n47078_, new_n47079_, new_n47080_,
    new_n47081_, new_n47082_, new_n47083_, new_n47084_, new_n47085_,
    new_n47086_, new_n47087_, new_n47088_, new_n47089_, new_n47090_,
    new_n47091_, new_n47092_, new_n47093_, new_n47094_, new_n47095_,
    new_n47096_, new_n47097_, new_n47098_, new_n47099_, new_n47100_,
    new_n47101_, new_n47102_, new_n47103_, new_n47104_, new_n47105_,
    new_n47106_, new_n47107_, new_n47108_, new_n47109_, new_n47110_,
    new_n47111_, new_n47112_, new_n47113_, new_n47114_, new_n47115_,
    new_n47116_, new_n47117_, new_n47118_, new_n47119_, new_n47120_,
    new_n47121_, new_n47122_, new_n47123_, new_n47124_, new_n47125_,
    new_n47126_, new_n47127_, new_n47128_, new_n47129_, new_n47130_,
    new_n47131_, new_n47132_, new_n47133_, new_n47134_, new_n47135_,
    new_n47136_, new_n47137_, new_n47138_, new_n47139_, new_n47140_,
    new_n47141_, new_n47142_, new_n47143_, new_n47144_, new_n47145_,
    new_n47146_, new_n47147_, new_n47148_, new_n47149_, new_n47150_,
    new_n47151_, new_n47152_, new_n47153_, new_n47154_, new_n47155_,
    new_n47156_, new_n47157_, new_n47158_, new_n47159_, new_n47160_,
    new_n47161_, new_n47162_, new_n47163_, new_n47164_, new_n47165_,
    new_n47166_, new_n47167_, new_n47168_, new_n47169_, new_n47170_,
    new_n47171_, new_n47172_, new_n47173_, new_n47174_, new_n47175_,
    new_n47176_, new_n47177_, new_n47178_, new_n47179_, new_n47180_,
    new_n47181_, new_n47182_, new_n47183_, new_n47184_, new_n47185_,
    new_n47186_, new_n47187_, new_n47188_, new_n47189_, new_n47190_,
    new_n47191_, new_n47192_, new_n47193_, new_n47194_, new_n47195_,
    new_n47196_, new_n47197_, new_n47198_, new_n47199_, new_n47200_,
    new_n47201_, new_n47202_, new_n47203_, new_n47204_, new_n47205_,
    new_n47206_, new_n47207_, new_n47208_, new_n47209_, new_n47210_,
    new_n47211_, new_n47212_, new_n47213_, new_n47214_, new_n47215_,
    new_n47216_, new_n47217_, new_n47218_, new_n47219_, new_n47220_,
    new_n47221_, new_n47222_, new_n47223_, new_n47224_, new_n47225_,
    new_n47226_, new_n47227_, new_n47228_, new_n47229_, new_n47230_,
    new_n47231_, new_n47232_, new_n47233_, new_n47234_, new_n47235_,
    new_n47236_, new_n47237_, new_n47238_, new_n47239_, new_n47240_,
    new_n47241_, new_n47242_, new_n47243_, new_n47244_, new_n47245_,
    new_n47246_, new_n47247_, new_n47248_, new_n47249_, new_n47250_,
    new_n47251_, new_n47252_, new_n47253_, new_n47254_, new_n47255_,
    new_n47256_, new_n47257_, new_n47258_, new_n47259_, new_n47260_,
    new_n47261_, new_n47262_, new_n47263_, new_n47264_, new_n47265_,
    new_n47266_, new_n47267_, new_n47268_, new_n47269_, new_n47270_,
    new_n47271_, new_n47272_, new_n47273_, new_n47274_, new_n47275_,
    new_n47276_, new_n47277_, new_n47278_, new_n47279_, new_n47280_,
    new_n47281_, new_n47282_, new_n47283_, new_n47284_, new_n47285_,
    new_n47286_, new_n47287_, new_n47288_, new_n47289_, new_n47290_,
    new_n47291_, new_n47292_, new_n47293_, new_n47294_, new_n47295_,
    new_n47296_, new_n47297_, new_n47298_, new_n47299_, new_n47300_,
    new_n47301_, new_n47302_, new_n47303_, new_n47304_, new_n47305_,
    new_n47306_, new_n47307_, new_n47308_, new_n47309_, new_n47310_,
    new_n47311_, new_n47312_, new_n47313_, new_n47314_, new_n47315_,
    new_n47316_, new_n47317_, new_n47318_, new_n47319_, new_n47320_,
    new_n47321_, new_n47322_, new_n47323_, new_n47324_, new_n47325_,
    new_n47326_, new_n47327_, new_n47328_, new_n47329_, new_n47330_,
    new_n47331_, new_n47332_, new_n47333_, new_n47334_, new_n47335_,
    new_n47336_, new_n47337_, new_n47338_, new_n47339_, new_n47340_,
    new_n47341_, new_n47342_, new_n47343_, new_n47344_, new_n47345_,
    new_n47346_, new_n47347_, new_n47348_, new_n47349_, new_n47350_,
    new_n47351_, new_n47352_, new_n47353_, new_n47354_, new_n47355_,
    new_n47356_, new_n47357_, new_n47358_, new_n47359_, new_n47360_,
    new_n47361_, new_n47362_, new_n47363_, new_n47364_, new_n47365_,
    new_n47366_, new_n47367_, new_n47368_, new_n47369_, new_n47370_,
    new_n47371_, new_n47372_, new_n47373_, new_n47374_, new_n47375_,
    new_n47376_, new_n47377_, new_n47378_, new_n47379_, new_n47380_,
    new_n47381_, new_n47382_, new_n47383_, new_n47384_, new_n47385_,
    new_n47386_, new_n47387_, new_n47388_, new_n47389_, new_n47390_,
    new_n47391_, new_n47392_, new_n47393_, new_n47394_, new_n47395_,
    new_n47396_, new_n47397_, new_n47398_, new_n47399_, new_n47400_,
    new_n47401_, new_n47402_, new_n47403_, new_n47404_, new_n47405_,
    new_n47406_, new_n47407_, new_n47408_, new_n47409_, new_n47410_,
    new_n47411_, new_n47412_, new_n47413_, new_n47414_, new_n47415_,
    new_n47416_, new_n47417_, new_n47418_, new_n47419_, new_n47420_,
    new_n47421_, new_n47422_, new_n47423_, new_n47424_, new_n47425_,
    new_n47426_, new_n47427_, new_n47428_, new_n47429_, new_n47430_,
    new_n47431_, new_n47432_, new_n47433_, new_n47434_, new_n47435_,
    new_n47436_, new_n47437_, new_n47438_, new_n47439_, new_n47440_,
    new_n47441_, new_n47442_, new_n47443_, new_n47444_, new_n47445_,
    new_n47446_, new_n47447_, new_n47448_, new_n47449_, new_n47450_,
    new_n47451_, new_n47452_, new_n47453_, new_n47454_, new_n47455_,
    new_n47456_, new_n47457_, new_n47458_, new_n47459_, new_n47460_,
    new_n47461_, new_n47462_, new_n47463_, new_n47464_, new_n47465_,
    new_n47466_, new_n47467_, new_n47468_, new_n47469_, new_n47470_,
    new_n47471_, new_n47472_, new_n47473_, new_n47474_, new_n47475_,
    new_n47476_, new_n47477_, new_n47478_, new_n47479_, new_n47480_,
    new_n47481_, new_n47482_, new_n47483_, new_n47484_, new_n47485_,
    new_n47486_, new_n47487_, new_n47488_, new_n47489_, new_n47490_,
    new_n47491_, new_n47492_, new_n47493_, new_n47494_, new_n47495_,
    new_n47496_, new_n47497_, new_n47498_, new_n47499_, new_n47500_,
    new_n47501_, new_n47502_, new_n47503_, new_n47504_, new_n47505_,
    new_n47506_, new_n47507_, new_n47508_, new_n47509_, new_n47510_,
    new_n47511_, new_n47512_, new_n47513_, new_n47514_, new_n47515_,
    new_n47516_, new_n47517_, new_n47518_, new_n47519_, new_n47520_,
    new_n47521_, new_n47522_, new_n47523_, new_n47524_, new_n47525_,
    new_n47526_, new_n47527_, new_n47528_, new_n47529_, new_n47530_,
    new_n47531_, new_n47532_, new_n47533_, new_n47534_, new_n47535_,
    new_n47536_, new_n47537_, new_n47538_, new_n47539_, new_n47540_,
    new_n47541_, new_n47542_, new_n47543_, new_n47544_, new_n47545_,
    new_n47546_, new_n47547_, new_n47548_, new_n47549_, new_n47550_,
    new_n47551_, new_n47552_, new_n47553_, new_n47554_, new_n47555_,
    new_n47556_, new_n47557_, new_n47558_, new_n47559_, new_n47560_,
    new_n47561_, new_n47562_, new_n47563_, new_n47564_, new_n47565_,
    new_n47566_, new_n47567_, new_n47568_, new_n47569_, new_n47570_,
    new_n47571_, new_n47572_, new_n47573_, new_n47574_, new_n47575_,
    new_n47576_, new_n47577_, new_n47578_, new_n47579_, new_n47580_,
    new_n47581_, new_n47582_, new_n47583_, new_n47584_, new_n47585_,
    new_n47586_, new_n47587_, new_n47588_, new_n47589_, new_n47590_,
    new_n47591_, new_n47592_, new_n47593_, new_n47594_, new_n47595_,
    new_n47596_, new_n47597_, new_n47598_, new_n47599_, new_n47600_,
    new_n47601_, new_n47602_, new_n47603_, new_n47604_, new_n47605_,
    new_n47606_, new_n47607_, new_n47608_, new_n47609_, new_n47610_,
    new_n47611_, new_n47612_, new_n47613_, new_n47614_, new_n47615_,
    new_n47616_, new_n47617_, new_n47618_, new_n47619_, new_n47620_,
    new_n47621_, new_n47622_, new_n47623_, new_n47624_, new_n47625_,
    new_n47626_, new_n47627_, new_n47628_, new_n47629_, new_n47630_,
    new_n47631_, new_n47632_, new_n47633_, new_n47634_, new_n47635_,
    new_n47636_, new_n47637_, new_n47638_, new_n47639_, new_n47640_,
    new_n47641_, new_n47642_, new_n47643_, new_n47644_, new_n47645_,
    new_n47646_, new_n47647_, new_n47648_, new_n47649_, new_n47650_,
    new_n47651_, new_n47652_, new_n47653_, new_n47654_, new_n47655_,
    new_n47656_, new_n47657_, new_n47658_, new_n47659_, new_n47660_,
    new_n47661_, new_n47662_, new_n47663_, new_n47664_, new_n47665_,
    new_n47666_, new_n47667_, new_n47668_, new_n47669_, new_n47670_,
    new_n47671_, new_n47672_, new_n47673_, new_n47674_, new_n47675_,
    new_n47676_, new_n47677_, new_n47678_, new_n47679_, new_n47680_,
    new_n47681_, new_n47682_, new_n47683_, new_n47684_, new_n47685_,
    new_n47686_, new_n47687_, new_n47688_, new_n47689_, new_n47690_,
    new_n47691_, new_n47692_, new_n47693_, new_n47694_, new_n47695_,
    new_n47696_, new_n47697_, new_n47698_, new_n47699_, new_n47700_,
    new_n47701_, new_n47702_, new_n47703_, new_n47704_, new_n47705_,
    new_n47706_, new_n47707_, new_n47708_, new_n47709_, new_n47710_,
    new_n47711_, new_n47712_, new_n47713_, new_n47714_, new_n47715_,
    new_n47716_, new_n47717_, new_n47718_, new_n47719_, new_n47720_,
    new_n47721_, new_n47722_, new_n47723_, new_n47724_, new_n47725_,
    new_n47726_, new_n47727_, new_n47728_, new_n47729_, new_n47730_,
    new_n47731_, new_n47732_, new_n47733_, new_n47734_, new_n47735_,
    new_n47736_, new_n47737_, new_n47738_, new_n47739_, new_n47740_,
    new_n47741_, new_n47742_, new_n47743_, new_n47744_, new_n47745_,
    new_n47746_, new_n47747_, new_n47748_, new_n47749_, new_n47750_,
    new_n47751_, new_n47752_, new_n47753_, new_n47754_, new_n47755_,
    new_n47756_, new_n47757_, new_n47758_, new_n47759_, new_n47760_,
    new_n47761_, new_n47762_, new_n47763_, new_n47764_, new_n47765_,
    new_n47766_, new_n47767_, new_n47768_, new_n47769_, new_n47770_,
    new_n47771_, new_n47772_, new_n47773_, new_n47774_, new_n47775_,
    new_n47776_, new_n47777_, new_n47778_, new_n47779_, new_n47780_,
    new_n47781_, new_n47782_, new_n47783_, new_n47784_, new_n47785_,
    new_n47786_, new_n47787_, new_n47788_, new_n47789_, new_n47790_,
    new_n47791_, new_n47792_, new_n47793_, new_n47794_, new_n47795_,
    new_n47796_, new_n47797_, new_n47798_, new_n47799_, new_n47800_,
    new_n47801_, new_n47802_, new_n47803_, new_n47804_, new_n47805_,
    new_n47806_, new_n47807_, new_n47808_, new_n47809_, new_n47810_,
    new_n47811_, new_n47812_, new_n47813_, new_n47814_, new_n47815_,
    new_n47816_, new_n47817_, new_n47818_, new_n47819_, new_n47820_,
    new_n47821_, new_n47822_, new_n47823_, new_n47824_, new_n47825_,
    new_n47826_, new_n47827_, new_n47828_, new_n47829_, new_n47830_,
    new_n47831_, new_n47832_, new_n47833_, new_n47834_, new_n47835_,
    new_n47836_, new_n47837_, new_n47838_, new_n47839_, new_n47840_,
    new_n47841_, new_n47842_, new_n47843_, new_n47844_, new_n47845_,
    new_n47846_, new_n47847_, new_n47848_, new_n47849_, new_n47850_,
    new_n47851_, new_n47852_, new_n47853_, new_n47854_, new_n47855_,
    new_n47856_, new_n47857_, new_n47858_, new_n47859_, new_n47860_,
    new_n47861_, new_n47862_, new_n47863_, new_n47864_, new_n47865_,
    new_n47866_, new_n47867_, new_n47868_, new_n47869_, new_n47870_,
    new_n47871_, new_n47872_, new_n47873_, new_n47874_, new_n47875_,
    new_n47876_, new_n47877_, new_n47878_, new_n47879_, new_n47880_,
    new_n47881_, new_n47882_, new_n47883_, new_n47884_, new_n47885_,
    new_n47886_, new_n47887_, new_n47888_, new_n47889_, new_n47890_,
    new_n47891_, new_n47892_, new_n47893_, new_n47894_, new_n47895_,
    new_n47896_, new_n47897_, new_n47898_, new_n47899_, new_n47900_,
    new_n47901_, new_n47902_, new_n47903_, new_n47904_, new_n47905_,
    new_n47906_, new_n47907_, new_n47908_, new_n47909_, new_n47910_,
    new_n47911_, new_n47912_, new_n47913_, new_n47914_, new_n47915_,
    new_n47916_, new_n47917_, new_n47918_, new_n47919_, new_n47920_,
    new_n47921_, new_n47922_, new_n47923_, new_n47924_, new_n47925_,
    new_n47926_, new_n47927_, new_n47928_, new_n47929_, new_n47930_,
    new_n47931_, new_n47932_, new_n47933_, new_n47934_, new_n47935_,
    new_n47936_, new_n47937_, new_n47938_, new_n47939_, new_n47940_,
    new_n47941_, new_n47942_, new_n47943_, new_n47944_, new_n47945_,
    new_n47946_, new_n47947_, new_n47948_, new_n47949_, new_n47950_,
    new_n47951_, new_n47952_, new_n47953_, new_n47954_, new_n47955_,
    new_n47956_, new_n47957_, new_n47958_, new_n47959_, new_n47960_,
    new_n47961_, new_n47962_, new_n47963_, new_n47964_, new_n47965_,
    new_n47966_, new_n47967_, new_n47968_, new_n47969_, new_n47970_,
    new_n47971_, new_n47972_, new_n47973_, new_n47974_, new_n47975_,
    new_n47976_, new_n47977_, new_n47978_, new_n47979_, new_n47980_,
    new_n47981_, new_n47982_, new_n47983_, new_n47984_, new_n47985_,
    new_n47986_, new_n47987_, new_n47988_, new_n47989_, new_n47990_,
    new_n47991_, new_n47992_, new_n47993_, new_n47994_, new_n47995_,
    new_n47996_, new_n47997_, new_n47998_, new_n47999_, new_n48000_,
    new_n48001_, new_n48002_, new_n48003_, new_n48004_, new_n48005_,
    new_n48006_, new_n48007_, new_n48008_, new_n48009_, new_n48010_,
    new_n48011_, new_n48012_, new_n48013_, new_n48014_, new_n48015_,
    new_n48016_, new_n48017_, new_n48018_, new_n48019_, new_n48020_,
    new_n48021_, new_n48022_, new_n48023_, new_n48024_, new_n48025_,
    new_n48026_, new_n48027_, new_n48028_, new_n48029_, new_n48030_,
    new_n48031_, new_n48032_, new_n48033_, new_n48034_, new_n48035_,
    new_n48036_, new_n48037_, new_n48038_, new_n48039_, new_n48040_,
    new_n48041_, new_n48042_, new_n48043_, new_n48044_, new_n48045_,
    new_n48046_, new_n48047_, new_n48048_, new_n48049_, new_n48050_,
    new_n48051_, new_n48052_, new_n48053_, new_n48054_, new_n48055_,
    new_n48056_, new_n48057_, new_n48058_, new_n48059_, new_n48060_,
    new_n48061_, new_n48062_, new_n48063_, new_n48064_, new_n48065_,
    new_n48066_, new_n48067_, new_n48068_, new_n48069_, new_n48070_,
    new_n48071_, new_n48072_, new_n48073_, new_n48074_, new_n48075_,
    new_n48076_, new_n48077_, new_n48078_, new_n48079_, new_n48080_,
    new_n48081_, new_n48082_, new_n48083_, new_n48084_, new_n48085_,
    new_n48086_, new_n48087_, new_n48088_, new_n48089_, new_n48090_,
    new_n48091_, new_n48092_, new_n48093_, new_n48094_, new_n48095_,
    new_n48096_, new_n48097_, new_n48098_, new_n48099_, new_n48100_,
    new_n48101_, new_n48102_, new_n48103_, new_n48104_, new_n48105_,
    new_n48106_, new_n48107_, new_n48108_, new_n48109_, new_n48110_,
    new_n48111_, new_n48112_, new_n48113_, new_n48114_, new_n48115_,
    new_n48116_, new_n48117_, new_n48118_, new_n48119_, new_n48120_,
    new_n48121_, new_n48122_, new_n48123_, new_n48124_, new_n48125_,
    new_n48126_, new_n48127_, new_n48128_, new_n48129_, new_n48130_,
    new_n48131_, new_n48132_, new_n48133_, new_n48134_, new_n48135_,
    new_n48136_, new_n48137_, new_n48138_, new_n48139_, new_n48140_,
    new_n48141_, new_n48142_, new_n48143_, new_n48144_, new_n48145_,
    new_n48146_, new_n48147_, new_n48148_, new_n48149_, new_n48150_,
    new_n48151_, new_n48152_, new_n48153_, new_n48154_, new_n48155_,
    new_n48156_, new_n48157_, new_n48158_, new_n48159_, new_n48160_,
    new_n48161_, new_n48162_, new_n48163_, new_n48164_, new_n48165_,
    new_n48166_, new_n48167_, new_n48168_, new_n48169_, new_n48170_,
    new_n48171_, new_n48172_, new_n48173_, new_n48174_, new_n48175_,
    new_n48176_, new_n48177_, new_n48178_, new_n48179_, new_n48180_,
    new_n48181_, new_n48182_, new_n48183_, new_n48184_, new_n48185_,
    new_n48186_, new_n48187_, new_n48188_, new_n48189_, new_n48190_,
    new_n48191_, new_n48192_, new_n48193_, new_n48194_, new_n48195_,
    new_n48196_, new_n48197_, new_n48198_, new_n48199_, new_n48200_,
    new_n48201_, new_n48202_, new_n48203_, new_n48204_, new_n48205_,
    new_n48206_, new_n48207_, new_n48208_, new_n48209_, new_n48210_,
    new_n48211_, new_n48212_, new_n48213_, new_n48214_, new_n48215_,
    new_n48216_, new_n48217_, new_n48218_, new_n48219_, new_n48220_,
    new_n48221_, new_n48222_, new_n48223_, new_n48224_, new_n48225_,
    new_n48226_, new_n48227_, new_n48228_, new_n48229_, new_n48230_,
    new_n48231_, new_n48232_, new_n48233_, new_n48234_, new_n48235_,
    new_n48236_, new_n48237_, new_n48238_, new_n48239_, new_n48240_,
    new_n48241_, new_n48242_, new_n48243_, new_n48244_, new_n48245_,
    new_n48246_, new_n48247_, new_n48248_, new_n48249_, new_n48250_,
    new_n48251_, new_n48252_, new_n48253_, new_n48254_, new_n48255_,
    new_n48256_, new_n48257_, new_n48258_, new_n48259_, new_n48260_,
    new_n48261_, new_n48262_, new_n48263_, new_n48264_, new_n48265_,
    new_n48266_, new_n48267_, new_n48268_, new_n48269_, new_n48270_,
    new_n48271_, new_n48272_, new_n48273_, new_n48274_, new_n48275_,
    new_n48276_, new_n48277_, new_n48278_, new_n48279_, new_n48280_,
    new_n48281_, new_n48282_, new_n48283_, new_n48284_, new_n48285_,
    new_n48286_, new_n48287_, new_n48288_, new_n48289_, new_n48290_,
    new_n48291_, new_n48292_, new_n48293_, new_n48294_, new_n48295_,
    new_n48296_, new_n48297_, new_n48298_, new_n48299_, new_n48300_,
    new_n48301_, new_n48302_, new_n48303_, new_n48304_, new_n48305_,
    new_n48306_, new_n48307_, new_n48308_, new_n48309_, new_n48310_,
    new_n48311_, new_n48312_, new_n48313_, new_n48314_, new_n48315_,
    new_n48316_, new_n48317_, new_n48318_, new_n48319_, new_n48320_,
    new_n48321_, new_n48322_, new_n48323_, new_n48324_, new_n48325_,
    new_n48326_, new_n48327_, new_n48328_, new_n48329_, new_n48330_,
    new_n48331_, new_n48332_, new_n48333_, new_n48334_, new_n48335_,
    new_n48336_, new_n48337_, new_n48338_, new_n48339_, new_n48340_,
    new_n48341_, new_n48342_, new_n48343_, new_n48344_, new_n48345_,
    new_n48346_, new_n48347_, new_n48348_, new_n48349_, new_n48350_,
    new_n48351_, new_n48352_, new_n48353_, new_n48354_, new_n48355_,
    new_n48356_, new_n48357_, new_n48358_, new_n48359_, new_n48360_,
    new_n48361_, new_n48362_, new_n48363_, new_n48364_, new_n48365_,
    new_n48366_, new_n48367_, new_n48368_, new_n48369_, new_n48370_,
    new_n48371_, new_n48372_, new_n48373_, new_n48374_, new_n48375_,
    new_n48376_, new_n48377_, new_n48378_, new_n48379_, new_n48380_,
    new_n48381_, new_n48382_, new_n48383_, new_n48384_, new_n48385_,
    new_n48386_, new_n48387_, new_n48388_, new_n48389_, new_n48390_,
    new_n48391_, new_n48392_, new_n48393_, new_n48394_, new_n48395_,
    new_n48396_, new_n48397_, new_n48398_, new_n48399_, new_n48400_,
    new_n48401_, new_n48402_, new_n48403_, new_n48404_, new_n48405_,
    new_n48406_, new_n48407_, new_n48408_, new_n48409_, new_n48410_,
    new_n48411_, new_n48412_, new_n48413_, new_n48414_, new_n48415_,
    new_n48416_, new_n48417_, new_n48418_, new_n48419_, new_n48420_,
    new_n48421_, new_n48422_, new_n48423_, new_n48424_, new_n48425_,
    new_n48426_, new_n48427_, new_n48428_, new_n48429_, new_n48430_,
    new_n48431_, new_n48432_, new_n48433_, new_n48434_, new_n48435_,
    new_n48436_, new_n48437_, new_n48438_, new_n48439_, new_n48440_,
    new_n48441_, new_n48442_, new_n48443_, new_n48444_, new_n48445_,
    new_n48446_, new_n48447_, new_n48448_, new_n48449_, new_n48450_,
    new_n48451_, new_n48452_, new_n48453_, new_n48454_, new_n48455_,
    new_n48456_, new_n48457_, new_n48458_, new_n48459_, new_n48460_,
    new_n48461_, new_n48462_, new_n48463_, new_n48464_, new_n48465_,
    new_n48466_, new_n48467_, new_n48468_, new_n48469_, new_n48470_,
    new_n48471_, new_n48472_, new_n48473_, new_n48474_, new_n48475_,
    new_n48476_, new_n48477_, new_n48478_, new_n48479_, new_n48480_,
    new_n48481_, new_n48482_, new_n48483_, new_n48484_, new_n48485_,
    new_n48486_, new_n48487_, new_n48488_, new_n48489_, new_n48490_,
    new_n48491_, new_n48492_, new_n48493_, new_n48494_, new_n48495_,
    new_n48496_, new_n48497_, new_n48498_, new_n48499_, new_n48500_,
    new_n48501_, new_n48502_, new_n48503_, new_n48504_, new_n48505_,
    new_n48506_, new_n48507_, new_n48508_, new_n48509_, new_n48510_,
    new_n48511_, new_n48512_, new_n48513_, new_n48514_, new_n48515_,
    new_n48516_, new_n48517_, new_n48518_, new_n48519_, new_n48520_,
    new_n48521_, new_n48522_, new_n48523_, new_n48524_, new_n48525_,
    new_n48526_, new_n48527_, new_n48528_, new_n48529_, new_n48530_,
    new_n48531_, new_n48532_, new_n48533_, new_n48534_, new_n48535_,
    new_n48536_, new_n48537_, new_n48538_, new_n48539_, new_n48540_,
    new_n48541_, new_n48542_, new_n48543_, new_n48544_, new_n48545_,
    new_n48546_, new_n48547_, new_n48548_, new_n48549_, new_n48550_,
    new_n48551_, new_n48552_, new_n48553_, new_n48554_, new_n48555_,
    new_n48556_, new_n48557_, new_n48558_, new_n48559_, new_n48560_,
    new_n48561_, new_n48562_, new_n48563_, new_n48564_, new_n48565_,
    new_n48566_, new_n48567_, new_n48568_, new_n48569_, new_n48570_,
    new_n48571_, new_n48572_, new_n48573_, new_n48574_, new_n48575_,
    new_n48576_, new_n48577_, new_n48578_, new_n48579_, new_n48580_,
    new_n48581_, new_n48582_, new_n48583_, new_n48584_, new_n48585_,
    new_n48586_, new_n48587_, new_n48588_, new_n48589_, new_n48590_,
    new_n48591_, new_n48592_, new_n48593_, new_n48594_, new_n48595_,
    new_n48596_, new_n48597_, new_n48598_, new_n48599_, new_n48600_,
    new_n48601_, new_n48602_, new_n48603_, new_n48604_, new_n48605_,
    new_n48606_, new_n48607_, new_n48608_, new_n48609_, new_n48610_,
    new_n48611_, new_n48612_, new_n48613_, new_n48614_, new_n48615_,
    new_n48616_, new_n48617_, new_n48618_, new_n48619_, new_n48620_,
    new_n48621_, new_n48622_, new_n48623_, new_n48624_, new_n48625_,
    new_n48626_, new_n48627_, new_n48628_, new_n48629_, new_n48630_,
    new_n48631_, new_n48632_, new_n48633_, new_n48634_, new_n48635_,
    new_n48636_, new_n48637_, new_n48638_, new_n48639_, new_n48640_,
    new_n48641_, new_n48642_, new_n48643_, new_n48644_, new_n48645_,
    new_n48646_, new_n48647_, new_n48648_, new_n48649_, new_n48650_,
    new_n48651_, new_n48652_, new_n48653_, new_n48654_, new_n48655_,
    new_n48656_, new_n48657_, new_n48658_, new_n48659_, new_n48660_,
    new_n48661_, new_n48662_, new_n48663_, new_n48664_, new_n48665_,
    new_n48666_, new_n48667_, new_n48668_, new_n48669_, new_n48670_,
    new_n48671_, new_n48672_, new_n48673_, new_n48674_, new_n48675_,
    new_n48676_, new_n48677_, new_n48678_, new_n48679_, new_n48680_,
    new_n48681_, new_n48682_, new_n48683_, new_n48684_, new_n48685_,
    new_n48686_, new_n48687_, new_n48688_, new_n48689_, new_n48690_,
    new_n48691_, new_n48692_, new_n48693_, new_n48694_, new_n48695_,
    new_n48696_, new_n48697_, new_n48698_, new_n48699_, new_n48700_,
    new_n48701_, new_n48702_, new_n48703_, new_n48704_, new_n48705_,
    new_n48706_, new_n48707_, new_n48708_, new_n48709_, new_n48710_,
    new_n48711_, new_n48712_, new_n48713_, new_n48714_, new_n48715_,
    new_n48716_, new_n48717_, new_n48718_, new_n48719_, new_n48720_,
    new_n48721_, new_n48722_, new_n48723_, new_n48724_, new_n48725_,
    new_n48726_, new_n48727_, new_n48728_, new_n48729_, new_n48730_,
    new_n48731_, new_n48732_, new_n48733_, new_n48734_, new_n48735_,
    new_n48736_, new_n48737_, new_n48738_, new_n48739_, new_n48740_,
    new_n48741_, new_n48742_, new_n48743_, new_n48744_, new_n48745_,
    new_n48746_, new_n48747_, new_n48748_, new_n48749_, new_n48750_,
    new_n48751_, new_n48752_, new_n48753_, new_n48754_, new_n48755_,
    new_n48756_, new_n48757_, new_n48758_, new_n48759_, new_n48760_,
    new_n48761_, new_n48762_, new_n48763_, new_n48764_, new_n48765_,
    new_n48766_, new_n48767_, new_n48768_, new_n48769_, new_n48770_,
    new_n48771_, new_n48772_, new_n48773_, new_n48774_, new_n48775_,
    new_n48776_, new_n48777_, new_n48778_, new_n48779_, new_n48780_,
    new_n48781_, new_n48782_, new_n48783_, new_n48784_, new_n48785_,
    new_n48786_, new_n48787_, new_n48788_, new_n48789_, new_n48790_,
    new_n48791_, new_n48792_, new_n48793_, new_n48794_, new_n48795_,
    new_n48796_, new_n48797_, new_n48798_, new_n48799_, new_n48800_,
    new_n48801_, new_n48802_, new_n48803_, new_n48804_, new_n48805_,
    new_n48806_, new_n48807_, new_n48808_, new_n48809_, new_n48810_,
    new_n48811_, new_n48812_, new_n48813_, new_n48814_, new_n48815_,
    new_n48816_, new_n48817_, new_n48818_, new_n48819_, new_n48820_,
    new_n48821_, new_n48822_, new_n48823_, new_n48824_, new_n48825_,
    new_n48826_, new_n48827_, new_n48828_, new_n48829_, new_n48830_,
    new_n48831_, new_n48832_, new_n48833_, new_n48834_, new_n48835_,
    new_n48836_, new_n48837_, new_n48838_, new_n48839_, new_n48840_,
    new_n48841_, new_n48842_, new_n48843_, new_n48844_, new_n48845_,
    new_n48846_, new_n48847_, new_n48848_, new_n48849_, new_n48850_,
    new_n48851_, new_n48852_, new_n48853_, new_n48854_, new_n48855_,
    new_n48856_, new_n48857_, new_n48858_, new_n48859_, new_n48860_,
    new_n48861_, new_n48862_, new_n48863_, new_n48864_, new_n48865_,
    new_n48866_, new_n48867_, new_n48868_, new_n48869_, new_n48870_,
    new_n48871_, new_n48872_, new_n48873_, new_n48874_, new_n48875_,
    new_n48876_, new_n48877_, new_n48878_, new_n48879_, new_n48880_,
    new_n48881_, new_n48882_, new_n48883_, new_n48884_, new_n48885_,
    new_n48886_, new_n48887_, new_n48888_, new_n48889_, new_n48890_,
    new_n48891_, new_n48892_, new_n48893_, new_n48894_, new_n48895_,
    new_n48896_, new_n48897_, new_n48898_, new_n48899_, new_n48900_,
    new_n48901_, new_n48902_, new_n48903_, new_n48904_, new_n48905_,
    new_n48906_, new_n48907_, new_n48908_, new_n48909_, new_n48910_,
    new_n48911_, new_n48912_, new_n48913_, new_n48914_, new_n48915_,
    new_n48916_, new_n48917_, new_n48918_, new_n48919_, new_n48920_,
    new_n48921_, new_n48922_, new_n48923_, new_n48924_, new_n48925_,
    new_n48926_, new_n48927_, new_n48928_, new_n48929_, new_n48930_,
    new_n48931_, new_n48932_, new_n48933_, new_n48934_, new_n48935_,
    new_n48936_, new_n48937_, new_n48938_, new_n48939_, new_n48940_,
    new_n48941_, new_n48942_, new_n48943_, new_n48944_, new_n48945_,
    new_n48946_, new_n48947_, new_n48948_, new_n48949_, new_n48950_,
    new_n48951_, new_n48952_, new_n48953_, new_n48954_, new_n48955_,
    new_n48956_, new_n48957_, new_n48958_, new_n48959_, new_n48960_,
    new_n48961_, new_n48962_, new_n48963_, new_n48964_, new_n48965_,
    new_n48966_, new_n48967_, new_n48968_, new_n48969_, new_n48970_,
    new_n48971_, new_n48972_, new_n48973_, new_n48974_, new_n48975_,
    new_n48976_, new_n48977_, new_n48978_, new_n48979_, new_n48980_,
    new_n48981_, new_n48982_, new_n48983_, new_n48984_, new_n48985_,
    new_n48986_, new_n48987_, new_n48988_, new_n48989_, new_n48990_,
    new_n48991_, new_n48992_, new_n48993_, new_n48994_, new_n48995_,
    new_n48996_, new_n48997_, new_n48998_, new_n48999_, new_n49000_,
    new_n49001_, new_n49002_, new_n49003_, new_n49004_, new_n49005_,
    new_n49006_, new_n49007_, new_n49008_, new_n49009_, new_n49010_,
    new_n49011_, new_n49012_, new_n49013_, new_n49014_, new_n49015_,
    new_n49016_, new_n49017_, new_n49018_, new_n49019_, new_n49020_,
    new_n49021_, new_n49022_, new_n49023_, new_n49024_, new_n49025_,
    new_n49026_, new_n49027_, new_n49028_, new_n49029_, new_n49030_,
    new_n49031_, new_n49032_, new_n49033_, new_n49034_, new_n49035_,
    new_n49036_, new_n49037_, new_n49038_, new_n49039_, new_n49040_,
    new_n49041_, new_n49042_, new_n49043_, new_n49044_, new_n49045_,
    new_n49046_, new_n49047_, new_n49048_, new_n49049_, new_n49050_,
    new_n49051_, new_n49052_, new_n49053_, new_n49054_, new_n49055_,
    new_n49056_, new_n49057_, new_n49058_, new_n49059_, new_n49060_,
    new_n49061_, new_n49062_, new_n49063_, new_n49064_, new_n49065_,
    new_n49066_, new_n49067_, new_n49068_, new_n49069_, new_n49070_,
    new_n49071_, new_n49072_, new_n49073_, new_n49074_, new_n49075_,
    new_n49076_, new_n49077_, new_n49078_, new_n49079_, new_n49080_,
    new_n49081_, new_n49082_, new_n49083_, new_n49084_, new_n49085_,
    new_n49086_, new_n49087_, new_n49088_, new_n49089_, new_n49090_,
    new_n49091_, new_n49092_, new_n49093_, new_n49094_, new_n49095_,
    new_n49096_, new_n49097_, new_n49098_, new_n49099_, new_n49100_,
    new_n49101_, new_n49102_, new_n49103_, new_n49104_, new_n49105_,
    new_n49106_, new_n49107_, new_n49108_, new_n49109_, new_n49110_,
    new_n49111_, new_n49112_, new_n49113_, new_n49114_, new_n49115_,
    new_n49116_, new_n49117_, new_n49118_, new_n49119_, new_n49120_,
    new_n49121_, new_n49122_, new_n49123_, new_n49124_, new_n49125_,
    new_n49126_, new_n49127_, new_n49128_, new_n49129_, new_n49130_,
    new_n49131_, new_n49132_, new_n49133_, new_n49134_, new_n49135_,
    new_n49136_, new_n49137_, new_n49138_, new_n49139_, new_n49140_,
    new_n49141_, new_n49142_, new_n49143_, new_n49144_, new_n49145_,
    new_n49146_, new_n49147_, new_n49148_, new_n49149_, new_n49150_,
    new_n49151_, new_n49152_, new_n49153_, new_n49154_, new_n49155_,
    new_n49156_, new_n49157_, new_n49158_, new_n49159_, new_n49160_,
    new_n49161_, new_n49162_, new_n49163_, new_n49164_, new_n49165_,
    new_n49166_, new_n49167_, new_n49168_, new_n49169_, new_n49170_,
    new_n49171_, new_n49172_, new_n49173_, new_n49174_, new_n49175_,
    new_n49176_, new_n49177_, new_n49178_, new_n49179_, new_n49180_,
    new_n49181_, new_n49182_, new_n49183_, new_n49184_, new_n49185_,
    new_n49186_, new_n49187_, new_n49188_, new_n49189_, new_n49190_,
    new_n49191_, new_n49192_, new_n49193_, new_n49194_, new_n49195_,
    new_n49196_, new_n49197_, new_n49198_, new_n49199_, new_n49200_,
    new_n49201_, new_n49202_, new_n49203_, new_n49204_, new_n49205_,
    new_n49206_, new_n49207_, new_n49208_, new_n49209_, new_n49210_,
    new_n49211_, new_n49212_, new_n49213_, new_n49214_, new_n49215_,
    new_n49216_, new_n49217_, new_n49218_, new_n49219_, new_n49220_,
    new_n49221_, new_n49222_, new_n49223_, new_n49224_, new_n49225_,
    new_n49226_, new_n49227_, new_n49228_, new_n49229_, new_n49230_,
    new_n49231_, new_n49232_, new_n49233_, new_n49234_, new_n49235_,
    new_n49236_, new_n49237_, new_n49238_, new_n49239_, new_n49240_,
    new_n49241_, new_n49242_, new_n49243_, new_n49244_, new_n49245_,
    new_n49246_, new_n49247_, new_n49248_, new_n49249_, new_n49250_,
    new_n49251_, new_n49252_, new_n49253_, new_n49254_, new_n49255_,
    new_n49256_, new_n49257_, new_n49258_, new_n49259_, new_n49260_,
    new_n49261_, new_n49262_, new_n49263_, new_n49264_, new_n49265_,
    new_n49266_, new_n49267_, new_n49268_, new_n49269_, new_n49270_,
    new_n49271_, new_n49272_, new_n49273_, new_n49274_, new_n49275_,
    new_n49276_, new_n49277_, new_n49278_, new_n49279_, new_n49280_,
    new_n49281_, new_n49282_, new_n49283_, new_n49284_, new_n49285_,
    new_n49286_, new_n49287_, new_n49288_, new_n49289_, new_n49290_,
    new_n49291_, new_n49292_, new_n49293_, new_n49294_, new_n49295_,
    new_n49296_, new_n49297_, new_n49298_, new_n49299_, new_n49300_,
    new_n49301_, new_n49302_, new_n49303_, new_n49304_, new_n49305_,
    new_n49306_, new_n49307_, new_n49308_, new_n49309_, new_n49310_,
    new_n49311_, new_n49312_, new_n49313_, new_n49314_, new_n49315_,
    new_n49316_, new_n49317_, new_n49318_, new_n49319_, new_n49320_,
    new_n49321_, new_n49322_, new_n49323_, new_n49324_, new_n49325_,
    new_n49326_, new_n49327_, new_n49328_, new_n49329_, new_n49330_,
    new_n49331_, new_n49332_, new_n49333_, new_n49334_, new_n49335_,
    new_n49336_, new_n49337_, new_n49338_, new_n49339_, new_n49340_,
    new_n49341_, new_n49342_, new_n49343_, new_n49344_, new_n49345_,
    new_n49346_, new_n49347_, new_n49348_, new_n49349_, new_n49350_,
    new_n49351_, new_n49352_, new_n49353_, new_n49354_, new_n49355_,
    new_n49356_, new_n49357_, new_n49358_, new_n49359_, new_n49360_,
    new_n49361_, new_n49362_, new_n49363_, new_n49364_, new_n49365_,
    new_n49366_, new_n49367_, new_n49368_, new_n49369_, new_n49370_,
    new_n49371_, new_n49372_, new_n49373_, new_n49374_, new_n49375_,
    new_n49376_, new_n49377_, new_n49378_, new_n49379_, new_n49380_,
    new_n49381_, new_n49382_, new_n49383_, new_n49384_, new_n49385_,
    new_n49386_, new_n49387_, new_n49388_, new_n49389_, new_n49390_,
    new_n49391_, new_n49392_, new_n49393_, new_n49394_, new_n49395_,
    new_n49396_, new_n49397_, new_n49398_, new_n49399_, new_n49400_,
    new_n49401_, new_n49402_, new_n49403_, new_n49404_, new_n49405_,
    new_n49406_, new_n49407_, new_n49408_, new_n49409_, new_n49410_,
    new_n49411_, new_n49412_, new_n49413_, new_n49414_, new_n49415_,
    new_n49416_, new_n49417_, new_n49418_, new_n49419_, new_n49420_,
    new_n49421_, new_n49422_, new_n49423_, new_n49424_, new_n49425_,
    new_n49426_, new_n49427_, new_n49428_, new_n49429_, new_n49430_,
    new_n49431_, new_n49432_, new_n49433_, new_n49434_, new_n49435_,
    new_n49436_, new_n49437_, new_n49438_, new_n49439_, new_n49440_,
    new_n49441_, new_n49442_, new_n49443_, new_n49444_, new_n49445_,
    new_n49446_, new_n49447_, new_n49448_, new_n49449_, new_n49450_,
    new_n49451_, new_n49452_, new_n49453_, new_n49454_, new_n49455_,
    new_n49456_, new_n49457_, new_n49458_, new_n49459_, new_n49460_,
    new_n49461_, new_n49462_, new_n49463_, new_n49464_, new_n49465_,
    new_n49466_, new_n49467_, new_n49468_, new_n49469_, new_n49470_,
    new_n49471_, new_n49472_, new_n49473_, new_n49474_, new_n49475_,
    new_n49476_, new_n49477_, new_n49478_, new_n49479_, new_n49480_,
    new_n49481_, new_n49482_, new_n49483_, new_n49484_, new_n49485_,
    new_n49486_, new_n49487_, new_n49488_, new_n49489_, new_n49490_,
    new_n49491_, new_n49492_, new_n49493_, new_n49494_, new_n49495_,
    new_n49496_, new_n49497_, new_n49498_, new_n49499_, new_n49500_,
    new_n49501_, new_n49502_, new_n49503_, new_n49504_, new_n49505_,
    new_n49506_, new_n49507_, new_n49508_, new_n49509_, new_n49510_,
    new_n49511_, new_n49512_, new_n49513_, new_n49514_, new_n49515_,
    new_n49516_, new_n49517_, new_n49518_, new_n49519_, new_n49520_,
    new_n49521_, new_n49522_, new_n49523_, new_n49524_, new_n49525_,
    new_n49526_, new_n49527_, new_n49528_, new_n49529_, new_n49530_,
    new_n49531_, new_n49532_, new_n49533_, new_n49534_, new_n49535_,
    new_n49536_, new_n49537_, new_n49538_, new_n49539_, new_n49540_,
    new_n49541_, new_n49542_, new_n49543_, new_n49544_, new_n49545_,
    new_n49546_, new_n49547_, new_n49548_, new_n49549_, new_n49550_,
    new_n49551_, new_n49552_, new_n49553_, new_n49554_, new_n49555_,
    new_n49556_, new_n49557_, new_n49558_, new_n49559_, new_n49560_,
    new_n49561_, new_n49562_, new_n49563_, new_n49564_, new_n49565_,
    new_n49566_, new_n49567_, new_n49568_, new_n49569_, new_n49570_,
    new_n49571_, new_n49572_, new_n49573_, new_n49574_, new_n49575_,
    new_n49576_, new_n49577_, new_n49578_, new_n49579_, new_n49580_,
    new_n49581_, new_n49582_, new_n49583_, new_n49584_, new_n49585_,
    new_n49586_, new_n49587_, new_n49588_, new_n49589_, new_n49590_,
    new_n49591_, new_n49592_, new_n49593_, new_n49594_, new_n49595_,
    new_n49596_, new_n49597_, new_n49598_, new_n49599_, new_n49600_,
    new_n49601_, new_n49602_, new_n49603_, new_n49604_, new_n49605_,
    new_n49606_, new_n49607_, new_n49608_, new_n49609_, new_n49610_,
    new_n49611_, new_n49612_, new_n49613_, new_n49614_, new_n49615_,
    new_n49616_, new_n49617_, new_n49618_, new_n49619_, new_n49620_,
    new_n49621_, new_n49622_, new_n49623_, new_n49624_, new_n49625_,
    new_n49626_, new_n49627_, new_n49628_, new_n49629_, new_n49630_,
    new_n49631_, new_n49632_, new_n49633_, new_n49634_, new_n49635_,
    new_n49636_, new_n49637_, new_n49638_, new_n49639_, new_n49640_,
    new_n49641_, new_n49642_, new_n49643_, new_n49644_, new_n49645_,
    new_n49646_, new_n49647_, new_n49648_, new_n49649_, new_n49650_,
    new_n49651_, new_n49652_, new_n49653_, new_n49654_, new_n49655_,
    new_n49656_, new_n49657_, new_n49658_, new_n49659_, new_n49660_,
    new_n49661_, new_n49662_, new_n49663_, new_n49664_, new_n49665_,
    new_n49666_, new_n49667_, new_n49668_, new_n49669_, new_n49670_,
    new_n49671_, new_n49672_, new_n49673_, new_n49674_, new_n49675_,
    new_n49676_, new_n49677_, new_n49678_, new_n49679_, new_n49680_,
    new_n49681_, new_n49682_, new_n49683_, new_n49684_, new_n49685_,
    new_n49686_, new_n49687_, new_n49688_, new_n49689_, new_n49690_,
    new_n49691_, new_n49692_, new_n49693_, new_n49694_, new_n49695_,
    new_n49696_, new_n49697_, new_n49698_, new_n49699_, new_n49700_,
    new_n49701_, new_n49702_, new_n49703_, new_n49704_, new_n49705_,
    new_n49706_, new_n49707_, new_n49708_, new_n49709_, new_n49710_,
    new_n49711_, new_n49712_, new_n49713_, new_n49714_, new_n49715_,
    new_n49716_, new_n49717_, new_n49718_, new_n49719_, new_n49720_,
    new_n49721_, new_n49722_, new_n49723_, new_n49724_, new_n49725_,
    new_n49726_, new_n49727_, new_n49728_, new_n49729_, new_n49730_,
    new_n49731_, new_n49732_, new_n49733_, new_n49734_, new_n49735_,
    new_n49736_, new_n49737_, new_n49738_, new_n49739_, new_n49740_,
    new_n49741_, new_n49742_, new_n49743_, new_n49744_, new_n49745_,
    new_n49746_, new_n49747_, new_n49748_, new_n49749_, new_n49750_,
    new_n49751_, new_n49752_, new_n49753_, new_n49754_, new_n49755_,
    new_n49756_, new_n49757_, new_n49758_, new_n49759_, new_n49760_,
    new_n49761_, new_n49762_, new_n49763_, new_n49764_, new_n49765_,
    new_n49766_, new_n49767_, new_n49768_, new_n49769_, new_n49770_,
    new_n49771_, new_n49772_, new_n49773_, new_n49774_, new_n49775_,
    new_n49776_, new_n49777_, new_n49778_, new_n49779_, new_n49780_,
    new_n49781_, new_n49782_, new_n49783_, new_n49784_, new_n49785_,
    new_n49786_, new_n49787_, new_n49788_, new_n49789_, new_n49790_,
    new_n49791_, new_n49792_, new_n49793_, new_n49794_, new_n49795_,
    new_n49796_, new_n49797_, new_n49798_, new_n49799_, new_n49800_,
    new_n49801_, new_n49802_, new_n49803_, new_n49804_, new_n49805_,
    new_n49806_, new_n49807_, new_n49808_, new_n49809_, new_n49810_,
    new_n49811_, new_n49812_, new_n49813_, new_n49814_, new_n49815_,
    new_n49816_, new_n49817_, new_n49818_, new_n49819_, new_n49820_,
    new_n49821_, new_n49822_, new_n49823_, new_n49824_, new_n49825_,
    new_n49826_, new_n49827_, new_n49828_, new_n49829_, new_n49830_,
    new_n49831_, new_n49832_, new_n49833_, new_n49834_, new_n49835_,
    new_n49836_, new_n49837_, new_n49838_, new_n49839_, new_n49840_,
    new_n49841_, new_n49842_, new_n49843_, new_n49844_, new_n49845_,
    new_n49846_, new_n49847_, new_n49848_, new_n49849_, new_n49850_,
    new_n49851_, new_n49852_, new_n49853_, new_n49854_, new_n49855_,
    new_n49856_, new_n49857_, new_n49858_, new_n49859_, new_n49860_,
    new_n49861_, new_n49862_, new_n49863_, new_n49864_, new_n49865_,
    new_n49866_, new_n49867_, new_n49868_, new_n49869_, new_n49870_,
    new_n49871_, new_n49872_, new_n49873_, new_n49874_, new_n49875_,
    new_n49876_, new_n49877_, new_n49878_, new_n49879_, new_n49880_,
    new_n49881_, new_n49882_, new_n49883_, new_n49884_, new_n49885_,
    new_n49886_, new_n49887_, new_n49888_, new_n49889_, new_n49890_,
    new_n49891_, new_n49892_, new_n49893_, new_n49894_, new_n49895_,
    new_n49896_, new_n49897_, new_n49898_, new_n49899_, new_n49900_,
    new_n49901_, new_n49902_, new_n49903_, new_n49904_, new_n49905_,
    new_n49906_, new_n49907_, new_n49908_, new_n49909_, new_n49910_,
    new_n49911_, new_n49912_, new_n49913_, new_n49914_, new_n49915_,
    new_n49916_, new_n49917_, new_n49918_, new_n49919_, new_n49920_,
    new_n49921_, new_n49922_, new_n49923_, new_n49924_, new_n49925_,
    new_n49926_, new_n49927_, new_n49928_, new_n49929_, new_n49930_,
    new_n49931_, new_n49932_, new_n49933_, new_n49934_, new_n49935_,
    new_n49936_, new_n49937_, new_n49938_, new_n49939_, new_n49940_,
    new_n49941_, new_n49942_, new_n49943_, new_n49944_, new_n49945_,
    new_n49946_, new_n49947_, new_n49948_, new_n49949_, new_n49950_,
    new_n49951_, new_n49952_, new_n49953_, new_n49954_, new_n49955_,
    new_n49956_, new_n49957_, new_n49958_, new_n49959_, new_n49960_,
    new_n49961_, new_n49962_, new_n49963_, new_n49964_, new_n49965_,
    new_n49966_, new_n49967_, new_n49968_, new_n49969_, new_n49970_,
    new_n49971_, new_n49972_, new_n49973_, new_n49974_, new_n49975_,
    new_n49976_, new_n49977_, new_n49978_, new_n49979_, new_n49980_,
    new_n49981_, new_n49982_, new_n49983_, new_n49984_, new_n49985_,
    new_n49986_, new_n49987_, new_n49988_, new_n49989_, new_n49990_,
    new_n49991_, new_n49992_, new_n49993_, new_n49994_, new_n49995_,
    new_n49996_, new_n49997_, new_n49998_, new_n49999_, new_n50000_,
    new_n50001_, new_n50002_, new_n50003_, new_n50004_, new_n50005_,
    new_n50006_, new_n50007_, new_n50008_, new_n50009_, new_n50010_,
    new_n50011_, new_n50012_, new_n50013_, new_n50014_, new_n50015_,
    new_n50016_, new_n50017_, new_n50018_, new_n50019_, new_n50020_,
    new_n50021_, new_n50022_, new_n50023_, new_n50024_, new_n50025_,
    new_n50026_, new_n50027_, new_n50028_, new_n50029_, new_n50030_,
    new_n50031_, new_n50032_, new_n50033_, new_n50034_, new_n50035_,
    new_n50036_, new_n50037_, new_n50038_, new_n50039_, new_n50040_,
    new_n50041_, new_n50042_, new_n50043_, new_n50044_, new_n50045_,
    new_n50046_, new_n50047_, new_n50048_, new_n50049_, new_n50050_,
    new_n50051_, new_n50052_, new_n50053_, new_n50054_, new_n50055_,
    new_n50056_, new_n50057_, new_n50058_, new_n50059_, new_n50060_,
    new_n50061_, new_n50062_, new_n50063_, new_n50064_, new_n50065_,
    new_n50066_, new_n50067_, new_n50068_, new_n50069_, new_n50070_,
    new_n50071_, new_n50072_, new_n50073_, new_n50074_, new_n50075_,
    new_n50076_, new_n50077_, new_n50078_, new_n50079_, new_n50080_,
    new_n50081_, new_n50082_, new_n50083_, new_n50084_, new_n50085_,
    new_n50086_, new_n50087_, new_n50088_, new_n50089_, new_n50090_,
    new_n50091_, new_n50092_, new_n50093_, new_n50094_, new_n50095_,
    new_n50096_, new_n50097_, new_n50098_, new_n50099_, new_n50100_,
    new_n50101_, new_n50102_, new_n50103_, new_n50104_, new_n50105_,
    new_n50106_, new_n50107_, new_n50108_, new_n50109_, new_n50110_,
    new_n50111_, new_n50112_, new_n50113_, new_n50114_, new_n50115_,
    new_n50116_, new_n50117_, new_n50118_, new_n50119_, new_n50120_,
    new_n50121_, new_n50122_, new_n50123_, new_n50124_, new_n50125_,
    new_n50126_, new_n50127_, new_n50128_, new_n50129_, new_n50130_,
    new_n50131_, new_n50132_, new_n50133_, new_n50134_, new_n50135_,
    new_n50136_, new_n50137_, new_n50138_, new_n50139_, new_n50140_,
    new_n50141_, new_n50142_, new_n50143_, new_n50144_, new_n50145_,
    new_n50146_, new_n50147_, new_n50148_, new_n50149_, new_n50150_,
    new_n50151_, new_n50152_, new_n50153_, new_n50154_, new_n50155_,
    new_n50156_, new_n50157_, new_n50158_, new_n50159_, new_n50160_,
    new_n50161_, new_n50162_, new_n50163_, new_n50164_, new_n50165_,
    new_n50166_, new_n50167_, new_n50168_, new_n50169_, new_n50170_,
    new_n50171_, new_n50172_, new_n50173_, new_n50174_, new_n50175_,
    new_n50176_, new_n50177_, new_n50178_, new_n50179_, new_n50180_,
    new_n50181_, new_n50182_, new_n50183_, new_n50184_, new_n50185_,
    new_n50186_, new_n50187_, new_n50188_, new_n50189_, new_n50190_,
    new_n50191_, new_n50192_, new_n50193_, new_n50194_, new_n50195_,
    new_n50196_, new_n50197_, new_n50198_, new_n50199_, new_n50200_,
    new_n50201_, new_n50202_, new_n50203_, new_n50204_, new_n50205_,
    new_n50206_, new_n50207_, new_n50208_, new_n50209_, new_n50210_,
    new_n50211_, new_n50212_, new_n50213_, new_n50214_, new_n50215_,
    new_n50216_, new_n50217_, new_n50218_, new_n50219_, new_n50220_,
    new_n50221_, new_n50222_, new_n50223_, new_n50224_, new_n50225_,
    new_n50226_, new_n50227_, new_n50228_, new_n50229_, new_n50230_,
    new_n50231_, new_n50232_, new_n50233_, new_n50234_, new_n50235_,
    new_n50236_, new_n50237_, new_n50238_, new_n50239_, new_n50240_,
    new_n50241_, new_n50242_, new_n50243_, new_n50244_, new_n50245_,
    new_n50246_, new_n50247_, new_n50248_, new_n50249_, new_n50250_,
    new_n50251_, new_n50252_, new_n50253_, new_n50254_, new_n50255_,
    new_n50256_, new_n50257_, new_n50258_, new_n50259_, new_n50260_,
    new_n50261_, new_n50262_, new_n50263_, new_n50264_, new_n50265_,
    new_n50266_, new_n50267_, new_n50268_, new_n50269_, new_n50270_,
    new_n50271_, new_n50272_, new_n50273_, new_n50274_, new_n50275_,
    new_n50276_, new_n50277_, new_n50278_, new_n50279_, new_n50280_,
    new_n50281_, new_n50282_, new_n50283_, new_n50284_, new_n50285_,
    new_n50286_, new_n50287_, new_n50288_, new_n50289_, new_n50290_,
    new_n50291_, new_n50292_, new_n50293_, new_n50294_, new_n50295_,
    new_n50296_, new_n50297_, new_n50298_, new_n50299_, new_n50300_,
    new_n50301_, new_n50302_, new_n50303_, new_n50304_, new_n50305_,
    new_n50306_, new_n50307_, new_n50308_, new_n50309_, new_n50310_,
    new_n50311_, new_n50312_, new_n50313_, new_n50314_, new_n50315_,
    new_n50316_, new_n50317_, new_n50318_, new_n50319_, new_n50320_,
    new_n50321_, new_n50322_, new_n50323_, new_n50324_, new_n50325_,
    new_n50326_, new_n50327_, new_n50328_, new_n50329_, new_n50330_,
    new_n50331_, new_n50332_, new_n50333_, new_n50334_, new_n50335_,
    new_n50336_, new_n50337_, new_n50338_, new_n50339_, new_n50340_,
    new_n50341_, new_n50342_, new_n50343_, new_n50344_, new_n50345_,
    new_n50346_, new_n50347_, new_n50348_, new_n50349_, new_n50350_,
    new_n50351_, new_n50352_, new_n50353_, new_n50354_, new_n50355_,
    new_n50356_, new_n50357_, new_n50358_, new_n50359_, new_n50360_,
    new_n50361_, new_n50362_, new_n50363_, new_n50364_, new_n50365_,
    new_n50366_, new_n50367_, new_n50368_, new_n50369_, new_n50370_,
    new_n50371_, new_n50372_, new_n50373_, new_n50374_, new_n50375_,
    new_n50376_, new_n50377_, new_n50378_, new_n50379_, new_n50380_,
    new_n50381_, new_n50382_, new_n50383_, new_n50384_, new_n50385_,
    new_n50386_, new_n50387_, new_n50388_, new_n50389_, new_n50390_,
    new_n50391_, new_n50392_, new_n50393_, new_n50394_, new_n50395_,
    new_n50396_, new_n50397_, new_n50398_, new_n50399_, new_n50400_,
    new_n50401_, new_n50402_, new_n50403_, new_n50404_, new_n50405_,
    new_n50406_, new_n50407_, new_n50408_, new_n50409_, new_n50410_,
    new_n50411_, new_n50412_, new_n50413_, new_n50414_, new_n50415_,
    new_n50416_, new_n50417_, new_n50418_, new_n50419_, new_n50420_,
    new_n50421_, new_n50422_, new_n50423_, new_n50424_, new_n50425_,
    new_n50426_, new_n50427_, new_n50428_, new_n50429_, new_n50430_,
    new_n50431_, new_n50432_, new_n50433_, new_n50434_, new_n50435_,
    new_n50436_, new_n50437_, new_n50438_, new_n50439_, new_n50440_,
    new_n50441_, new_n50442_, new_n50443_, new_n50444_, new_n50445_,
    new_n50446_, new_n50447_, new_n50448_, new_n50449_, new_n50450_,
    new_n50451_, new_n50452_, new_n50453_, new_n50454_, new_n50455_,
    new_n50456_, new_n50457_, new_n50458_, new_n50459_, new_n50460_,
    new_n50461_, new_n50462_, new_n50463_, new_n50464_, new_n50465_,
    new_n50466_, new_n50467_, new_n50468_, new_n50469_, new_n50470_,
    new_n50471_, new_n50472_, new_n50473_, new_n50474_, new_n50475_,
    new_n50476_, new_n50477_, new_n50478_, new_n50479_, new_n50480_,
    new_n50481_, new_n50482_, new_n50483_, new_n50484_, new_n50485_,
    new_n50486_, new_n50487_, new_n50488_, new_n50489_, new_n50490_,
    new_n50491_, new_n50492_, new_n50493_, new_n50494_, new_n50495_,
    new_n50496_, new_n50497_, new_n50498_, new_n50499_, new_n50500_,
    new_n50501_, new_n50502_, new_n50503_, new_n50504_, new_n50505_,
    new_n50506_, new_n50507_, new_n50508_, new_n50509_, new_n50510_,
    new_n50511_, new_n50512_, new_n50513_, new_n50514_, new_n50515_,
    new_n50516_, new_n50517_, new_n50518_, new_n50519_, new_n50520_,
    new_n50521_, new_n50522_, new_n50523_, new_n50524_, new_n50525_,
    new_n50526_, new_n50527_, new_n50528_, new_n50529_, new_n50530_,
    new_n50531_, new_n50532_, new_n50533_, new_n50534_, new_n50535_,
    new_n50536_, new_n50537_, new_n50538_, new_n50539_, new_n50540_,
    new_n50541_, new_n50542_, new_n50543_, new_n50544_, new_n50545_,
    new_n50546_, new_n50547_, new_n50548_, new_n50549_, new_n50550_,
    new_n50551_, new_n50552_, new_n50553_, new_n50554_, new_n50555_,
    new_n50556_, new_n50557_, new_n50558_, new_n50559_, new_n50560_,
    new_n50561_, new_n50562_, new_n50563_, new_n50564_, new_n50565_,
    new_n50566_, new_n50567_, new_n50568_, new_n50569_, new_n50570_,
    new_n50571_, new_n50572_, new_n50573_, new_n50574_, new_n50575_,
    new_n50576_, new_n50577_, new_n50578_, new_n50579_, new_n50580_,
    new_n50581_, new_n50582_, new_n50583_, new_n50584_, new_n50585_,
    new_n50586_, new_n50587_, new_n50588_, new_n50589_, new_n50590_,
    new_n50591_, new_n50592_, new_n50593_, new_n50594_, new_n50595_,
    new_n50596_, new_n50597_, new_n50598_, new_n50599_, new_n50600_,
    new_n50601_, new_n50602_, new_n50603_, new_n50604_, new_n50605_,
    new_n50606_, new_n50607_, new_n50608_, new_n50609_, new_n50610_,
    new_n50611_, new_n50612_, new_n50613_, new_n50614_, new_n50615_,
    new_n50616_, new_n50617_, new_n50618_, new_n50619_, new_n50620_,
    new_n50621_, new_n50622_, new_n50623_, new_n50624_, new_n50625_,
    new_n50626_, new_n50627_, new_n50628_, new_n50629_, new_n50630_,
    new_n50631_, new_n50632_, new_n50633_, new_n50634_, new_n50635_,
    new_n50636_, new_n50637_, new_n50638_, new_n50639_, new_n50640_,
    new_n50641_, new_n50642_, new_n50643_, new_n50644_, new_n50645_,
    new_n50646_, new_n50647_, new_n50648_, new_n50649_, new_n50650_,
    new_n50651_, new_n50652_, new_n50653_, new_n50654_, new_n50655_,
    new_n50656_, new_n50657_, new_n50658_, new_n50659_, new_n50660_,
    new_n50661_, new_n50662_, new_n50663_, new_n50664_, new_n50665_,
    new_n50666_, new_n50667_, new_n50668_, new_n50669_, new_n50670_,
    new_n50671_, new_n50672_, new_n50673_, new_n50674_, new_n50675_,
    new_n50676_, new_n50677_, new_n50678_, new_n50679_, new_n50680_,
    new_n50681_, new_n50682_, new_n50683_, new_n50684_, new_n50685_,
    new_n50686_, new_n50687_, new_n50688_, new_n50689_, new_n50690_,
    new_n50691_, new_n50692_, new_n50693_, new_n50694_, new_n50695_,
    new_n50696_, new_n50697_, new_n50698_, new_n50699_, new_n50700_,
    new_n50701_, new_n50702_, new_n50703_, new_n50704_, new_n50705_,
    new_n50706_, new_n50707_, new_n50708_, new_n50709_, new_n50710_,
    new_n50711_, new_n50712_, new_n50713_, new_n50714_, new_n50715_,
    new_n50716_, new_n50717_, new_n50718_, new_n50719_, new_n50720_,
    new_n50721_, new_n50722_, new_n50723_, new_n50724_, new_n50725_,
    new_n50726_, new_n50727_, new_n50728_, new_n50729_, new_n50730_,
    new_n50731_, new_n50732_, new_n50733_, new_n50734_, new_n50735_,
    new_n50736_, new_n50737_, new_n50738_, new_n50739_, new_n50740_,
    new_n50741_, new_n50742_, new_n50743_, new_n50744_, new_n50745_,
    new_n50746_, new_n50747_, new_n50748_, new_n50749_, new_n50750_,
    new_n50751_, new_n50752_, new_n50753_, new_n50754_, new_n50755_,
    new_n50756_, new_n50757_, new_n50758_, new_n50759_, new_n50760_,
    new_n50761_, new_n50762_, new_n50763_, new_n50764_, new_n50765_,
    new_n50766_, new_n50767_, new_n50768_, new_n50769_, new_n50770_,
    new_n50771_, new_n50772_, new_n50773_, new_n50774_, new_n50775_,
    new_n50776_, new_n50777_, new_n50778_, new_n50779_, new_n50780_,
    new_n50781_, new_n50782_, new_n50783_, new_n50784_, new_n50785_,
    new_n50786_, new_n50787_, new_n50788_, new_n50789_, new_n50790_,
    new_n50791_, new_n50792_, new_n50793_, new_n50794_, new_n50795_,
    new_n50796_, new_n50797_, new_n50798_, new_n50799_, new_n50800_,
    new_n50801_, new_n50802_, new_n50803_, new_n50804_, new_n50805_,
    new_n50806_, new_n50807_, new_n50808_, new_n50809_, new_n50810_,
    new_n50811_, new_n50812_, new_n50813_, new_n50814_, new_n50815_,
    new_n50816_, new_n50817_, new_n50818_, new_n50819_, new_n50820_,
    new_n50821_, new_n50822_, new_n50823_, new_n50824_, new_n50825_,
    new_n50826_, new_n50827_, new_n50828_, new_n50829_, new_n50830_,
    new_n50831_, new_n50832_, new_n50833_, new_n50834_, new_n50835_,
    new_n50836_, new_n50837_, new_n50838_, new_n50839_, new_n50840_,
    new_n50841_, new_n50842_, new_n50843_, new_n50844_, new_n50845_,
    new_n50846_, new_n50847_, new_n50848_, new_n50849_, new_n50850_,
    new_n50851_, new_n50852_, new_n50853_, new_n50854_, new_n50855_,
    new_n50856_, new_n50857_, new_n50858_, new_n50859_, new_n50860_,
    new_n50861_, new_n50862_, new_n50863_, new_n50864_, new_n50865_,
    new_n50866_, new_n50867_, new_n50868_, new_n50869_, new_n50870_,
    new_n50871_, new_n50872_, new_n50873_, new_n50874_, new_n50875_,
    new_n50876_, new_n50877_, new_n50878_, new_n50879_, new_n50880_,
    new_n50881_, new_n50882_, new_n50883_, new_n50884_, new_n50885_,
    new_n50886_, new_n50887_, new_n50888_, new_n50889_, new_n50890_,
    new_n50891_, new_n50892_, new_n50893_, new_n50894_, new_n50895_,
    new_n50896_, new_n50897_, new_n50898_, new_n50899_, new_n50900_,
    new_n50901_, new_n50902_, new_n50903_, new_n50904_, new_n50905_,
    new_n50906_, new_n50907_, new_n50908_, new_n50909_, new_n50910_,
    new_n50911_, new_n50912_, new_n50913_, new_n50914_, new_n50915_,
    new_n50916_, new_n50917_, new_n50918_, new_n50919_, new_n50920_,
    new_n50921_, new_n50922_, new_n50923_, new_n50924_, new_n50925_,
    new_n50926_, new_n50927_, new_n50928_, new_n50929_, new_n50930_,
    new_n50931_, new_n50932_, new_n50933_, new_n50934_, new_n50935_,
    new_n50936_, new_n50937_, new_n50938_, new_n50939_, new_n50940_,
    new_n50941_, new_n50942_, new_n50943_, new_n50944_, new_n50945_,
    new_n50946_, new_n50947_, new_n50948_, new_n50949_, new_n50950_,
    new_n50951_, new_n50952_, new_n50953_, new_n50954_, new_n50955_,
    new_n50956_, new_n50957_, new_n50958_, new_n50959_, new_n50960_,
    new_n50961_, new_n50962_, new_n50963_, new_n50964_, new_n50965_,
    new_n50966_, new_n50967_, new_n50968_, new_n50969_, new_n50970_,
    new_n50971_, new_n50972_, new_n50973_, new_n50974_, new_n50975_,
    new_n50976_, new_n50977_, new_n50978_, new_n50979_, new_n50980_,
    new_n50981_, new_n50982_, new_n50983_, new_n50984_, new_n50985_,
    new_n50986_, new_n50987_, new_n50988_, new_n50989_, new_n50990_,
    new_n50991_, new_n50992_, new_n50993_, new_n50994_, new_n50995_,
    new_n50996_, new_n50997_, new_n50998_, new_n50999_, new_n51000_,
    new_n51001_, new_n51002_, new_n51003_, new_n51004_, new_n51005_,
    new_n51006_, new_n51007_, new_n51008_, new_n51009_, new_n51010_,
    new_n51011_, new_n51012_, new_n51013_, new_n51014_, new_n51015_,
    new_n51016_, new_n51017_, new_n51018_, new_n51019_, new_n51020_,
    new_n51021_, new_n51022_, new_n51023_, new_n51024_, new_n51025_,
    new_n51026_, new_n51027_, new_n51028_, new_n51029_, new_n51030_,
    new_n51031_, new_n51032_, new_n51033_, new_n51034_, new_n51035_,
    new_n51036_, new_n51037_, new_n51038_, new_n51039_, new_n51040_,
    new_n51041_, new_n51042_, new_n51043_, new_n51044_, new_n51045_,
    new_n51046_, new_n51047_, new_n51048_, new_n51049_, new_n51050_,
    new_n51051_, new_n51052_, new_n51053_, new_n51054_, new_n51055_,
    new_n51056_, new_n51057_, new_n51058_, new_n51059_, new_n51060_,
    new_n51061_, new_n51062_, new_n51063_, new_n51064_, new_n51065_,
    new_n51066_, new_n51067_, new_n51068_, new_n51069_, new_n51070_,
    new_n51071_, new_n51072_, new_n51073_, new_n51074_, new_n51075_,
    new_n51076_, new_n51077_, new_n51078_, new_n51079_, new_n51080_,
    new_n51081_, new_n51082_, new_n51083_, new_n51084_, new_n51085_,
    new_n51086_, new_n51087_, new_n51088_, new_n51089_, new_n51090_,
    new_n51091_, new_n51092_, new_n51093_, new_n51094_, new_n51095_,
    new_n51096_, new_n51097_, new_n51098_, new_n51099_, new_n51100_,
    new_n51101_, new_n51102_, new_n51103_, new_n51104_, new_n51105_,
    new_n51106_, new_n51107_, new_n51108_, new_n51109_, new_n51110_,
    new_n51111_, new_n51112_, new_n51113_, new_n51114_, new_n51115_,
    new_n51116_, new_n51117_, new_n51118_, new_n51119_, new_n51120_,
    new_n51121_, new_n51122_, new_n51123_, new_n51124_, new_n51125_,
    new_n51126_, new_n51127_, new_n51128_, new_n51129_, new_n51130_,
    new_n51131_, new_n51132_, new_n51133_, new_n51134_, new_n51135_,
    new_n51136_, new_n51137_, new_n51138_, new_n51139_, new_n51140_,
    new_n51141_, new_n51142_, new_n51143_, new_n51144_, new_n51145_,
    new_n51146_, new_n51147_, new_n51148_, new_n51149_, new_n51150_,
    new_n51151_, new_n51152_, new_n51153_, new_n51154_, new_n51155_,
    new_n51156_, new_n51157_, new_n51158_, new_n51159_, new_n51160_,
    new_n51161_, new_n51162_, new_n51163_, new_n51164_, new_n51165_,
    new_n51166_, new_n51167_, new_n51168_, new_n51169_, new_n51170_,
    new_n51171_, new_n51172_, new_n51173_, new_n51174_, new_n51175_,
    new_n51176_, new_n51177_, new_n51178_, new_n51179_, new_n51180_,
    new_n51181_, new_n51182_, new_n51183_, new_n51184_, new_n51185_,
    new_n51186_, new_n51187_, new_n51188_, new_n51189_, new_n51190_,
    new_n51191_, new_n51192_, new_n51193_, new_n51194_, new_n51195_,
    new_n51196_, new_n51197_, new_n51198_, new_n51199_, new_n51200_,
    new_n51201_, new_n51202_, new_n51203_, new_n51204_, new_n51205_,
    new_n51206_, new_n51207_, new_n51208_, new_n51209_, new_n51210_,
    new_n51211_, new_n51212_, new_n51213_, new_n51214_, new_n51215_,
    new_n51216_, new_n51217_, new_n51218_, new_n51219_, new_n51220_,
    new_n51221_, new_n51222_, new_n51223_, new_n51224_, new_n51225_,
    new_n51226_, new_n51227_, new_n51228_, new_n51229_, new_n51230_,
    new_n51231_, new_n51232_, new_n51233_, new_n51234_, new_n51235_,
    new_n51236_, new_n51237_, new_n51238_, new_n51239_, new_n51240_,
    new_n51241_, new_n51242_, new_n51243_, new_n51244_, new_n51245_,
    new_n51246_, new_n51247_, new_n51248_, new_n51249_, new_n51250_,
    new_n51251_, new_n51252_, new_n51253_, new_n51254_, new_n51255_,
    new_n51256_, new_n51257_, new_n51258_, new_n51259_, new_n51260_,
    new_n51261_, new_n51262_, new_n51263_, new_n51264_, new_n51265_,
    new_n51266_, new_n51267_, new_n51268_, new_n51269_, new_n51270_,
    new_n51271_, new_n51272_, new_n51273_, new_n51274_, new_n51275_,
    new_n51276_, new_n51277_, new_n51278_, new_n51279_, new_n51280_,
    new_n51281_, new_n51282_, new_n51283_, new_n51284_, new_n51285_,
    new_n51286_, new_n51287_, new_n51288_, new_n51289_, new_n51290_,
    new_n51291_, new_n51292_, new_n51293_, new_n51294_, new_n51295_,
    new_n51296_, new_n51297_, new_n51298_, new_n51299_, new_n51300_,
    new_n51301_, new_n51302_, new_n51303_, new_n51304_, new_n51305_,
    new_n51306_, new_n51307_, new_n51308_, new_n51309_, new_n51310_,
    new_n51311_, new_n51312_, new_n51313_, new_n51314_, new_n51315_,
    new_n51316_, new_n51317_, new_n51318_, new_n51319_, new_n51320_,
    new_n51321_, new_n51322_, new_n51323_, new_n51324_, new_n51325_,
    new_n51326_, new_n51327_, new_n51328_, new_n51329_, new_n51330_,
    new_n51331_, new_n51332_, new_n51333_, new_n51334_, new_n51335_,
    new_n51336_, new_n51337_, new_n51338_, new_n51339_, new_n51340_,
    new_n51341_, new_n51342_, new_n51343_, new_n51344_, new_n51345_,
    new_n51346_, new_n51347_, new_n51348_, new_n51349_, new_n51350_,
    new_n51351_, new_n51352_, new_n51353_, new_n51354_, new_n51355_,
    new_n51356_, new_n51357_, new_n51358_, new_n51359_, new_n51360_,
    new_n51361_, new_n51362_, new_n51363_, new_n51364_, new_n51365_,
    new_n51366_, new_n51367_, new_n51368_, new_n51369_, new_n51370_,
    new_n51371_, new_n51372_, new_n51373_, new_n51374_, new_n51375_,
    new_n51376_, new_n51377_, new_n51378_, new_n51379_, new_n51380_,
    new_n51381_, new_n51382_, new_n51383_, new_n51384_, new_n51385_,
    new_n51386_, new_n51387_, new_n51388_, new_n51389_, new_n51390_,
    new_n51391_, new_n51392_, new_n51393_, new_n51394_, new_n51395_,
    new_n51396_, new_n51397_, new_n51398_, new_n51399_, new_n51400_,
    new_n51401_, new_n51402_, new_n51403_, new_n51404_, new_n51405_,
    new_n51406_, new_n51407_, new_n51408_, new_n51409_, new_n51410_,
    new_n51411_, new_n51412_, new_n51413_, new_n51414_, new_n51415_,
    new_n51416_, new_n51417_, new_n51418_, new_n51419_, new_n51420_,
    new_n51421_, new_n51422_, new_n51423_, new_n51424_, new_n51425_,
    new_n51426_, new_n51427_, new_n51428_, new_n51429_, new_n51430_,
    new_n51431_, new_n51432_, new_n51433_, new_n51434_, new_n51435_,
    new_n51436_, new_n51437_, new_n51438_, new_n51439_, new_n51440_,
    new_n51441_, new_n51442_, new_n51443_, new_n51444_, new_n51445_,
    new_n51446_, new_n51447_, new_n51448_, new_n51449_, new_n51450_,
    new_n51451_, new_n51452_, new_n51453_, new_n51454_, new_n51455_,
    new_n51456_, new_n51457_, new_n51458_, new_n51459_, new_n51460_,
    new_n51461_, new_n51462_, new_n51463_, new_n51464_, new_n51465_,
    new_n51466_, new_n51467_, new_n51468_, new_n51469_, new_n51470_,
    new_n51471_, new_n51472_, new_n51473_, new_n51474_, new_n51475_,
    new_n51476_, new_n51477_, new_n51478_, new_n51479_, new_n51480_,
    new_n51481_, new_n51482_, new_n51483_, new_n51484_, new_n51485_,
    new_n51486_, new_n51487_, new_n51488_, new_n51489_, new_n51490_,
    new_n51491_, new_n51492_, new_n51493_, new_n51494_, new_n51495_,
    new_n51496_, new_n51497_, new_n51498_, new_n51499_, new_n51500_,
    new_n51501_, new_n51502_, new_n51503_, new_n51504_, new_n51505_,
    new_n51506_, new_n51507_, new_n51508_, new_n51509_, new_n51510_,
    new_n51511_, new_n51512_, new_n51513_, new_n51514_, new_n51515_,
    new_n51516_, new_n51517_, new_n51518_, new_n51519_, new_n51520_,
    new_n51521_, new_n51522_, new_n51523_, new_n51524_, new_n51525_,
    new_n51526_, new_n51527_, new_n51528_, new_n51529_, new_n51530_,
    new_n51531_, new_n51532_, new_n51533_, new_n51534_, new_n51535_,
    new_n51536_, new_n51537_, new_n51538_, new_n51539_, new_n51540_,
    new_n51541_, new_n51542_, new_n51543_, new_n51544_, new_n51545_,
    new_n51546_, new_n51547_, new_n51548_, new_n51549_, new_n51550_,
    new_n51551_, new_n51552_, new_n51553_, new_n51554_, new_n51555_,
    new_n51556_, new_n51557_, new_n51558_, new_n51559_, new_n51560_,
    new_n51561_, new_n51562_, new_n51563_, new_n51564_, new_n51565_,
    new_n51566_, new_n51567_, new_n51568_, new_n51569_, new_n51570_,
    new_n51571_, new_n51572_, new_n51573_, new_n51574_, new_n51575_,
    new_n51576_, new_n51577_, new_n51578_, new_n51579_, new_n51580_,
    new_n51581_, new_n51582_, new_n51583_, new_n51584_, new_n51585_,
    new_n51586_, new_n51587_, new_n51588_, new_n51589_, new_n51590_,
    new_n51591_, new_n51592_, new_n51593_, new_n51594_, new_n51595_,
    new_n51596_, new_n51597_, new_n51598_, new_n51599_, new_n51600_,
    new_n51601_, new_n51602_, new_n51603_, new_n51604_, new_n51605_,
    new_n51606_, new_n51607_, new_n51608_, new_n51609_, new_n51610_,
    new_n51611_, new_n51612_, new_n51613_, new_n51614_, new_n51615_,
    new_n51616_, new_n51617_, new_n51618_, new_n51619_, new_n51620_,
    new_n51621_, new_n51622_, new_n51623_, new_n51624_, new_n51625_,
    new_n51626_, new_n51627_, new_n51628_, new_n51629_, new_n51630_,
    new_n51631_, new_n51632_, new_n51633_, new_n51634_, new_n51635_,
    new_n51636_, new_n51637_, new_n51638_, new_n51639_, new_n51640_,
    new_n51641_, new_n51642_, new_n51643_, new_n51644_, new_n51645_,
    new_n51646_, new_n51647_, new_n51648_, new_n51649_, new_n51650_,
    new_n51651_, new_n51652_, new_n51653_, new_n51654_, new_n51655_,
    new_n51656_, new_n51657_, new_n51658_, new_n51659_, new_n51660_,
    new_n51661_, new_n51662_, new_n51663_, new_n51664_, new_n51665_,
    new_n51666_, new_n51667_, new_n51668_, new_n51669_, new_n51670_,
    new_n51671_, new_n51672_, new_n51673_, new_n51674_, new_n51675_,
    new_n51676_, new_n51677_, new_n51678_, new_n51679_, new_n51680_,
    new_n51681_, new_n51682_, new_n51683_, new_n51684_, new_n51685_,
    new_n51686_, new_n51687_, new_n51688_, new_n51689_, new_n51690_,
    new_n51691_, new_n51692_, new_n51693_, new_n51694_, new_n51695_,
    new_n51696_, new_n51697_, new_n51698_, new_n51699_, new_n51700_,
    new_n51701_, new_n51702_, new_n51703_, new_n51704_, new_n51705_,
    new_n51706_, new_n51707_, new_n51708_, new_n51709_, new_n51710_,
    new_n51711_, new_n51712_, new_n51713_, new_n51714_, new_n51715_,
    new_n51716_, new_n51717_, new_n51718_, new_n51719_, new_n51720_,
    new_n51721_, new_n51722_, new_n51723_, new_n51724_, new_n51725_,
    new_n51726_, new_n51727_, new_n51728_, new_n51729_, new_n51730_,
    new_n51731_, new_n51732_, new_n51733_, new_n51734_, new_n51735_,
    new_n51736_, new_n51737_, new_n51738_, new_n51739_, new_n51740_,
    new_n51741_, new_n51742_, new_n51743_, new_n51744_, new_n51745_,
    new_n51746_, new_n51747_, new_n51748_, new_n51749_, new_n51750_,
    new_n51751_, new_n51752_, new_n51753_, new_n51754_, new_n51755_,
    new_n51756_, new_n51757_, new_n51758_, new_n51759_, new_n51760_,
    new_n51761_, new_n51762_, new_n51763_, new_n51764_, new_n51765_,
    new_n51766_, new_n51767_, new_n51768_, new_n51769_, new_n51770_,
    new_n51771_, new_n51772_, new_n51773_, new_n51774_, new_n51775_,
    new_n51776_, new_n51777_, new_n51778_, new_n51779_, new_n51780_,
    new_n51781_, new_n51782_, new_n51783_, new_n51784_, new_n51785_,
    new_n51786_, new_n51787_, new_n51788_, new_n51789_, new_n51790_,
    new_n51791_, new_n51792_, new_n51793_, new_n51794_, new_n51795_,
    new_n51796_, new_n51797_, new_n51798_, new_n51799_, new_n51800_,
    new_n51801_, new_n51802_, new_n51803_, new_n51804_, new_n51805_,
    new_n51806_, new_n51807_, new_n51808_, new_n51809_, new_n51810_,
    new_n51811_, new_n51812_, new_n51813_, new_n51814_, new_n51815_,
    new_n51816_, new_n51817_, new_n51818_, new_n51819_, new_n51820_,
    new_n51821_, new_n51822_, new_n51823_, new_n51824_, new_n51825_,
    new_n51826_, new_n51827_, new_n51828_, new_n51829_, new_n51830_,
    new_n51831_, new_n51832_, new_n51833_, new_n51834_, new_n51835_,
    new_n51836_, new_n51837_, new_n51838_, new_n51839_, new_n51840_,
    new_n51841_, new_n51842_, new_n51843_, new_n51844_, new_n51845_,
    new_n51846_, new_n51847_, new_n51848_, new_n51849_, new_n51850_,
    new_n51851_, new_n51852_, new_n51853_, new_n51854_, new_n51855_,
    new_n51856_, new_n51857_, new_n51858_, new_n51859_, new_n51860_,
    new_n51861_, new_n51862_, new_n51863_, new_n51864_, new_n51865_,
    new_n51866_, new_n51867_, new_n51868_, new_n51869_, new_n51870_,
    new_n51871_, new_n51872_, new_n51873_, new_n51874_, new_n51875_,
    new_n51876_, new_n51877_, new_n51878_, new_n51879_, new_n51880_,
    new_n51881_, new_n51882_, new_n51883_, new_n51884_, new_n51885_,
    new_n51886_, new_n51887_, new_n51888_, new_n51889_, new_n51890_,
    new_n51891_, new_n51892_, new_n51893_, new_n51894_, new_n51895_,
    new_n51896_, new_n51897_, new_n51898_, new_n51899_, new_n51900_,
    new_n51901_, new_n51902_, new_n51903_, new_n51904_, new_n51905_,
    new_n51906_, new_n51907_, new_n51908_, new_n51909_, new_n51910_,
    new_n51911_, new_n51912_, new_n51913_, new_n51914_, new_n51915_,
    new_n51916_, new_n51917_, new_n51918_, new_n51919_, new_n51920_,
    new_n51921_, new_n51922_, new_n51923_, new_n51924_, new_n51925_,
    new_n51926_, new_n51927_, new_n51928_, new_n51929_, new_n51930_,
    new_n51931_, new_n51932_, new_n51933_, new_n51934_, new_n51935_,
    new_n51936_, new_n51937_, new_n51938_, new_n51939_, new_n51940_,
    new_n51941_, new_n51942_, new_n51943_, new_n51944_, new_n51945_,
    new_n51946_, new_n51947_, new_n51948_, new_n51949_, new_n51950_,
    new_n51951_, new_n51952_, new_n51953_, new_n51954_, new_n51955_,
    new_n51956_, new_n51957_, new_n51958_, new_n51959_, new_n51960_,
    new_n51961_, new_n51962_, new_n51963_, new_n51964_, new_n51965_,
    new_n51966_, new_n51967_, new_n51968_, new_n51969_, new_n51970_,
    new_n51971_, new_n51972_, new_n51973_, new_n51974_, new_n51975_,
    new_n51976_, new_n51977_, new_n51978_, new_n51979_, new_n51980_,
    new_n51981_, new_n51982_, new_n51983_, new_n51984_, new_n51985_,
    new_n51986_, new_n51987_, new_n51988_, new_n51989_, new_n51990_,
    new_n51991_, new_n51992_, new_n51993_, new_n51994_, new_n51995_,
    new_n51996_, new_n51997_, new_n51998_, new_n51999_, new_n52000_,
    new_n52001_, new_n52002_, new_n52003_, new_n52004_, new_n52005_,
    new_n52006_, new_n52007_, new_n52008_, new_n52009_, new_n52010_,
    new_n52011_, new_n52012_, new_n52013_, new_n52014_, new_n52015_,
    new_n52016_, new_n52017_, new_n52018_, new_n52019_, new_n52020_,
    new_n52021_, new_n52022_, new_n52023_, new_n52024_, new_n52025_,
    new_n52026_, new_n52027_, new_n52028_, new_n52029_, new_n52030_,
    new_n52031_, new_n52032_, new_n52033_, new_n52034_, new_n52035_,
    new_n52036_, new_n52037_, new_n52038_, new_n52039_, new_n52040_,
    new_n52041_, new_n52042_, new_n52043_, new_n52044_, new_n52045_,
    new_n52046_, new_n52047_, new_n52048_, new_n52049_, new_n52050_,
    new_n52051_, new_n52052_, new_n52053_, new_n52054_, new_n52055_,
    new_n52056_, new_n52057_, new_n52058_, new_n52059_, new_n52060_,
    new_n52061_, new_n52062_, new_n52063_, new_n52064_, new_n52065_,
    new_n52066_, new_n52067_, new_n52068_, new_n52069_, new_n52070_,
    new_n52071_, new_n52072_, new_n52073_, new_n52074_, new_n52075_,
    new_n52076_, new_n52077_, new_n52078_, new_n52079_, new_n52080_,
    new_n52081_, new_n52082_, new_n52083_, new_n52084_, new_n52085_,
    new_n52086_, new_n52087_, new_n52088_, new_n52089_, new_n52090_,
    new_n52091_, new_n52092_, new_n52093_, new_n52094_, new_n52095_,
    new_n52096_, new_n52097_, new_n52098_, new_n52099_, new_n52100_,
    new_n52101_, new_n52102_, new_n52103_, new_n52104_, new_n52105_,
    new_n52106_, new_n52107_, new_n52108_, new_n52109_, new_n52110_,
    new_n52111_, new_n52112_, new_n52113_, new_n52114_, new_n52115_,
    new_n52116_, new_n52117_, new_n52118_, new_n52119_, new_n52120_,
    new_n52121_, new_n52122_, new_n52123_, new_n52124_, new_n52125_,
    new_n52126_, new_n52127_, new_n52128_, new_n52129_, new_n52130_,
    new_n52131_, new_n52132_, new_n52133_, new_n52134_, new_n52135_,
    new_n52136_, new_n52137_, new_n52138_, new_n52139_, new_n52140_,
    new_n52141_, new_n52142_, new_n52143_, new_n52144_, new_n52145_,
    new_n52146_, new_n52147_, new_n52148_, new_n52149_, new_n52150_,
    new_n52151_, new_n52152_, new_n52153_, new_n52154_, new_n52155_,
    new_n52156_, new_n52157_, new_n52158_, new_n52159_, new_n52160_,
    new_n52161_, new_n52162_, new_n52163_, new_n52164_, new_n52165_,
    new_n52166_, new_n52167_, new_n52168_, new_n52169_, new_n52170_,
    new_n52171_, new_n52172_, new_n52173_, new_n52174_, new_n52175_,
    new_n52176_, new_n52177_, new_n52178_, new_n52179_, new_n52180_,
    new_n52181_, new_n52182_, new_n52183_, new_n52184_, new_n52185_,
    new_n52186_, new_n52187_, new_n52188_, new_n52189_, new_n52190_,
    new_n52191_, new_n52192_, new_n52193_, new_n52194_, new_n52195_,
    new_n52196_, new_n52197_, new_n52198_, new_n52199_, new_n52200_,
    new_n52201_, new_n52202_, new_n52203_, new_n52204_, new_n52205_,
    new_n52206_, new_n52207_, new_n52208_, new_n52209_, new_n52210_,
    new_n52211_, new_n52212_, new_n52213_, new_n52214_, new_n52215_,
    new_n52216_, new_n52217_, new_n52218_, new_n52219_, new_n52220_,
    new_n52221_, new_n52222_, new_n52223_, new_n52224_, new_n52225_,
    new_n52226_, new_n52227_, new_n52228_, new_n52229_, new_n52230_,
    new_n52231_, new_n52232_, new_n52233_, new_n52234_, new_n52235_,
    new_n52236_, new_n52237_, new_n52238_, new_n52239_, new_n52240_,
    new_n52241_, new_n52242_, new_n52243_, new_n52244_, new_n52245_,
    new_n52246_, new_n52247_, new_n52248_, new_n52249_, new_n52250_,
    new_n52251_, new_n52252_, new_n52253_, new_n52254_, new_n52255_,
    new_n52256_, new_n52257_, new_n52258_, new_n52259_, new_n52260_,
    new_n52261_, new_n52262_, new_n52263_, new_n52264_, new_n52265_,
    new_n52266_, new_n52267_, new_n52268_, new_n52269_, new_n52270_,
    new_n52271_, new_n52272_, new_n52273_, new_n52274_, new_n52275_,
    new_n52276_, new_n52277_, new_n52278_, new_n52279_, new_n52280_,
    new_n52281_, new_n52282_, new_n52283_, new_n52284_, new_n52285_,
    new_n52286_, new_n52287_, new_n52288_, new_n52289_, new_n52290_,
    new_n52291_, new_n52292_, new_n52293_, new_n52294_, new_n52295_,
    new_n52296_, new_n52297_, new_n52298_, new_n52299_, new_n52300_,
    new_n52301_, new_n52302_, new_n52303_, new_n52304_, new_n52305_,
    new_n52306_, new_n52307_, new_n52308_, new_n52309_, new_n52310_,
    new_n52311_, new_n52312_, new_n52313_, new_n52314_, new_n52315_,
    new_n52316_, new_n52317_, new_n52318_, new_n52319_, new_n52320_,
    new_n52321_, new_n52322_, new_n52323_, new_n52324_, new_n52325_,
    new_n52326_, new_n52327_, new_n52328_, new_n52329_, new_n52330_,
    new_n52331_, new_n52332_, new_n52333_, new_n52334_, new_n52335_,
    new_n52336_, new_n52337_, new_n52338_, new_n52339_, new_n52340_,
    new_n52341_, new_n52342_, new_n52343_, new_n52344_, new_n52345_,
    new_n52346_, new_n52347_, new_n52348_, new_n52349_, new_n52350_,
    new_n52351_, new_n52352_, new_n52353_, new_n52354_, new_n52355_,
    new_n52356_, new_n52357_, new_n52358_, new_n52359_, new_n52360_,
    new_n52361_, new_n52362_, new_n52363_, new_n52364_, new_n52365_,
    new_n52366_, new_n52367_, new_n52368_, new_n52369_, new_n52370_,
    new_n52371_, new_n52372_, new_n52373_, new_n52374_, new_n52375_,
    new_n52376_, new_n52377_, new_n52378_, new_n52379_, new_n52380_,
    new_n52381_, new_n52382_, new_n52383_, new_n52384_, new_n52385_,
    new_n52386_, new_n52387_, new_n52388_, new_n52389_, new_n52390_,
    new_n52391_, new_n52392_, new_n52393_, new_n52394_, new_n52395_,
    new_n52396_, new_n52397_, new_n52398_, new_n52399_, new_n52400_,
    new_n52401_, new_n52402_, new_n52403_, new_n52404_, new_n52405_,
    new_n52406_, new_n52407_, new_n52408_, new_n52409_, new_n52410_,
    new_n52411_, new_n52412_, new_n52413_, new_n52414_, new_n52415_,
    new_n52416_, new_n52417_, new_n52418_, new_n52419_, new_n52420_,
    new_n52421_, new_n52422_, new_n52423_, new_n52424_, new_n52425_,
    new_n52426_, new_n52427_, new_n52428_, new_n52429_, new_n52430_,
    new_n52431_, new_n52432_, new_n52433_, new_n52434_, new_n52435_,
    new_n52436_, new_n52437_, new_n52438_, new_n52439_, new_n52440_,
    new_n52441_, new_n52442_, new_n52443_, new_n52444_, new_n52445_,
    new_n52446_, new_n52447_, new_n52448_, new_n52449_, new_n52450_,
    new_n52451_, new_n52452_, new_n52453_, new_n52454_, new_n52455_,
    new_n52456_, new_n52457_, new_n52458_, new_n52459_, new_n52460_,
    new_n52461_, new_n52462_, new_n52463_, new_n52464_, new_n52465_,
    new_n52466_, new_n52467_, new_n52468_, new_n52469_, new_n52470_,
    new_n52471_, new_n52472_, new_n52473_, new_n52474_, new_n52475_,
    new_n52476_, new_n52477_, new_n52478_, new_n52479_, new_n52480_,
    new_n52481_, new_n52482_, new_n52483_, new_n52484_, new_n52485_,
    new_n52486_, new_n52487_, new_n52488_, new_n52489_, new_n52490_,
    new_n52491_, new_n52492_, new_n52493_, new_n52494_, new_n52495_,
    new_n52496_, new_n52497_, new_n52498_, new_n52499_, new_n52500_,
    new_n52501_, new_n52502_, new_n52503_, new_n52504_, new_n52505_,
    new_n52506_, new_n52507_, new_n52508_, new_n52509_, new_n52510_,
    new_n52511_, new_n52512_, new_n52513_, new_n52514_, new_n52515_,
    new_n52516_, new_n52517_, new_n52518_, new_n52519_, new_n52520_,
    new_n52521_, new_n52522_, new_n52523_, new_n52524_, new_n52525_,
    new_n52526_, new_n52527_, new_n52528_, new_n52529_, new_n52530_,
    new_n52531_, new_n52532_, new_n52533_, new_n52534_, new_n52535_,
    new_n52536_, new_n52537_, new_n52538_, new_n52539_, new_n52540_,
    new_n52541_, new_n52542_, new_n52543_, new_n52544_, new_n52545_,
    new_n52546_, new_n52547_, new_n52548_, new_n52549_, new_n52550_,
    new_n52551_, new_n52552_, new_n52553_, new_n52554_, new_n52555_,
    new_n52556_, new_n52557_, new_n52558_, new_n52559_, new_n52560_,
    new_n52561_, new_n52562_, new_n52563_, new_n52564_, new_n52565_,
    new_n52566_, new_n52567_, new_n52568_, new_n52569_, new_n52570_,
    new_n52571_, new_n52572_, new_n52573_, new_n52574_, new_n52575_,
    new_n52576_, new_n52577_, new_n52578_, new_n52579_, new_n52580_,
    new_n52581_, new_n52582_, new_n52583_, new_n52584_, new_n52585_,
    new_n52586_, new_n52587_, new_n52588_, new_n52589_, new_n52590_,
    new_n52591_, new_n52592_, new_n52593_, new_n52594_, new_n52595_,
    new_n52596_, new_n52597_, new_n52598_, new_n52599_, new_n52600_,
    new_n52601_, new_n52602_, new_n52603_, new_n52604_, new_n52605_,
    new_n52606_, new_n52607_, new_n52608_, new_n52609_, new_n52610_,
    new_n52611_, new_n52612_, new_n52613_, new_n52614_, new_n52615_,
    new_n52616_, new_n52617_, new_n52618_, new_n52619_, new_n52620_,
    new_n52621_, new_n52622_, new_n52623_, new_n52624_, new_n52625_,
    new_n52626_, new_n52627_, new_n52628_, new_n52629_, new_n52630_,
    new_n52631_, new_n52632_, new_n52633_, new_n52634_, new_n52635_,
    new_n52636_, new_n52637_, new_n52638_, new_n52639_, new_n52640_,
    new_n52641_, new_n52642_, new_n52643_, new_n52644_, new_n52645_,
    new_n52646_, new_n52647_, new_n52648_, new_n52649_, new_n52650_,
    new_n52651_, new_n52652_, new_n52653_, new_n52654_, new_n52655_,
    new_n52656_, new_n52657_, new_n52658_, new_n52659_, new_n52660_,
    new_n52661_, new_n52662_, new_n52663_, new_n52664_, new_n52665_,
    new_n52666_, new_n52667_, new_n52668_, new_n52669_, new_n52670_,
    new_n52671_, new_n52672_, new_n52673_, new_n52674_, new_n52675_,
    new_n52676_, new_n52677_, new_n52678_, new_n52679_, new_n52680_,
    new_n52681_, new_n52682_, new_n52683_, new_n52684_, new_n52685_,
    new_n52686_, new_n52687_, new_n52688_, new_n52689_, new_n52690_,
    new_n52691_, new_n52692_, new_n52693_, new_n52694_, new_n52695_,
    new_n52696_, new_n52697_, new_n52698_, new_n52699_, new_n52700_,
    new_n52701_, new_n52702_, new_n52703_, new_n52704_, new_n52705_,
    new_n52706_, new_n52707_, new_n52708_, new_n52709_, new_n52710_,
    new_n52711_, new_n52712_, new_n52713_, new_n52714_, new_n52715_,
    new_n52716_, new_n52717_, new_n52718_, new_n52719_, new_n52720_,
    new_n52721_, new_n52722_, new_n52723_, new_n52724_, new_n52725_,
    new_n52726_, new_n52727_, new_n52728_, new_n52729_, new_n52730_,
    new_n52731_, new_n52732_, new_n52733_, new_n52734_, new_n52735_,
    new_n52736_, new_n52737_, new_n52738_, new_n52739_, new_n52740_,
    new_n52741_, new_n52742_, new_n52743_, new_n52744_, new_n52745_,
    new_n52746_, new_n52747_, new_n52748_, new_n52749_, new_n52750_,
    new_n52751_, new_n52752_, new_n52753_, new_n52754_, new_n52755_,
    new_n52756_, new_n52757_, new_n52758_, new_n52759_, new_n52760_,
    new_n52761_, new_n52762_, new_n52763_, new_n52764_, new_n52765_,
    new_n52766_, new_n52767_, new_n52768_, new_n52769_, new_n52770_,
    new_n52771_, new_n52772_, new_n52773_, new_n52774_, new_n52775_,
    new_n52776_, new_n52777_, new_n52778_, new_n52779_, new_n52780_,
    new_n52781_, new_n52782_, new_n52783_, new_n52784_, new_n52785_,
    new_n52786_, new_n52787_, new_n52788_, new_n52789_, new_n52790_,
    new_n52791_, new_n52792_, new_n52793_, new_n52794_, new_n52795_,
    new_n52796_, new_n52797_, new_n52798_, new_n52799_, new_n52800_,
    new_n52801_, new_n52802_, new_n52803_, new_n52804_, new_n52805_,
    new_n52806_, new_n52807_, new_n52808_, new_n52809_, new_n52810_,
    new_n52811_, new_n52812_, new_n52813_, new_n52814_, new_n52815_,
    new_n52816_, new_n52817_, new_n52818_, new_n52819_, new_n52820_,
    new_n52821_, new_n52822_, new_n52823_, new_n52824_, new_n52825_,
    new_n52826_, new_n52827_, new_n52828_, new_n52829_, new_n52830_,
    new_n52831_, new_n52832_, new_n52833_, new_n52834_, new_n52835_,
    new_n52836_, new_n52837_, new_n52838_, new_n52839_, new_n52840_,
    new_n52841_, new_n52842_, new_n52843_, new_n52844_, new_n52845_,
    new_n52846_, new_n52847_, new_n52848_, new_n52849_, new_n52850_,
    new_n52851_, new_n52852_, new_n52853_, new_n52854_, new_n52855_,
    new_n52856_, new_n52857_, new_n52858_, new_n52859_, new_n52860_,
    new_n52861_, new_n52862_, new_n52863_, new_n52864_, new_n52865_,
    new_n52866_, new_n52867_, new_n52868_, new_n52869_, new_n52870_,
    new_n52871_, new_n52872_, new_n52873_, new_n52874_, new_n52875_,
    new_n52876_, new_n52877_, new_n52878_, new_n52879_, new_n52880_,
    new_n52881_, new_n52882_, new_n52883_, new_n52884_, new_n52885_,
    new_n52886_, new_n52887_, new_n52888_, new_n52889_, new_n52890_,
    new_n52891_, new_n52892_, new_n52893_, new_n52894_, new_n52895_,
    new_n52896_, new_n52897_, new_n52898_, new_n52899_, new_n52900_,
    new_n52901_, new_n52902_, new_n52903_, new_n52904_, new_n52905_,
    new_n52906_, new_n52907_, new_n52908_, new_n52909_, new_n52910_,
    new_n52911_, new_n52912_, new_n52913_, new_n52914_, new_n52915_,
    new_n52916_, new_n52917_, new_n52918_, new_n52919_, new_n52920_,
    new_n52921_, new_n52922_, new_n52923_, new_n52924_, new_n52925_,
    new_n52926_, new_n52927_, new_n52928_, new_n52929_, new_n52930_,
    new_n52931_, new_n52932_, new_n52933_, new_n52934_, new_n52935_,
    new_n52936_, new_n52937_, new_n52938_, new_n52939_, new_n52940_,
    new_n52941_, new_n52942_, new_n52943_, new_n52944_, new_n52945_,
    new_n52946_, new_n52947_, new_n52948_, new_n52949_, new_n52950_,
    new_n52951_, new_n52952_, new_n52953_, new_n52954_, new_n52955_,
    new_n52956_, new_n52957_, new_n52958_, new_n52959_, new_n52960_,
    new_n52961_, new_n52962_, new_n52963_, new_n52964_, new_n52965_,
    new_n52966_, new_n52967_, new_n52968_, new_n52969_, new_n52970_,
    new_n52971_, new_n52972_, new_n52973_, new_n52974_, new_n52975_,
    new_n52976_, new_n52977_, new_n52978_, new_n52979_, new_n52980_,
    new_n52981_, new_n52982_, new_n52983_, new_n52984_, new_n52985_,
    new_n52986_, new_n52987_, new_n52988_, new_n52989_, new_n52990_,
    new_n52991_, new_n52992_, new_n52993_, new_n52994_, new_n52995_,
    new_n52996_, new_n52997_, new_n52998_, new_n52999_, new_n53000_,
    new_n53001_, new_n53002_, new_n53003_, new_n53004_, new_n53005_,
    new_n53006_, new_n53007_, new_n53008_, new_n53009_, new_n53010_,
    new_n53011_, new_n53012_, new_n53013_, new_n53014_, new_n53015_,
    new_n53016_, new_n53017_, new_n53018_, new_n53019_, new_n53020_,
    new_n53021_, new_n53022_, new_n53023_, new_n53024_, new_n53025_,
    new_n53026_, new_n53027_, new_n53028_, new_n53029_, new_n53030_,
    new_n53031_, new_n53032_, new_n53033_, new_n53034_, new_n53035_,
    new_n53036_, new_n53037_, new_n53038_, new_n53039_, new_n53040_,
    new_n53041_, new_n53042_, new_n53043_, new_n53044_, new_n53045_,
    new_n53046_, new_n53047_, new_n53048_, new_n53049_, new_n53050_,
    new_n53051_, new_n53052_, new_n53053_, new_n53054_, new_n53055_,
    new_n53056_, new_n53057_, new_n53058_, new_n53059_, new_n53060_,
    new_n53061_, new_n53062_, new_n53063_, new_n53064_, new_n53065_,
    new_n53066_, new_n53067_, new_n53068_, new_n53069_, new_n53070_,
    new_n53071_, new_n53072_, new_n53073_, new_n53074_, new_n53075_,
    new_n53076_, new_n53077_, new_n53078_, new_n53079_, new_n53080_,
    new_n53081_, new_n53082_, new_n53083_, new_n53084_, new_n53085_,
    new_n53086_, new_n53087_, new_n53088_, new_n53089_, new_n53090_,
    new_n53091_, new_n53092_, new_n53093_, new_n53094_, new_n53095_,
    new_n53096_, new_n53097_, new_n53098_, new_n53099_, new_n53100_,
    new_n53101_, new_n53102_, new_n53103_, new_n53104_, new_n53105_,
    new_n53106_, new_n53107_, new_n53108_, new_n53109_, new_n53110_,
    new_n53111_, new_n53112_, new_n53113_, new_n53114_, new_n53115_,
    new_n53116_, new_n53117_, new_n53118_, new_n53119_, new_n53120_,
    new_n53121_, new_n53122_, new_n53123_, new_n53124_, new_n53125_,
    new_n53126_, new_n53127_, new_n53128_, new_n53129_, new_n53130_,
    new_n53131_, new_n53132_, new_n53133_, new_n53134_, new_n53135_,
    new_n53136_, new_n53137_, new_n53138_, new_n53139_, new_n53140_,
    new_n53141_, new_n53142_, new_n53143_, new_n53144_, new_n53145_,
    new_n53146_, new_n53147_, new_n53148_, new_n53149_, new_n53150_,
    new_n53151_, new_n53152_, new_n53153_, new_n53154_, new_n53155_,
    new_n53156_, new_n53157_, new_n53158_, new_n53159_, new_n53160_,
    new_n53161_, new_n53162_, new_n53163_, new_n53164_, new_n53165_,
    new_n53166_, new_n53167_, new_n53168_, new_n53169_, new_n53170_,
    new_n53171_, new_n53172_, new_n53173_, new_n53174_, new_n53175_,
    new_n53176_, new_n53177_, new_n53178_, new_n53179_, new_n53180_,
    new_n53181_, new_n53182_, new_n53183_, new_n53184_, new_n53185_,
    new_n53186_, new_n53187_, new_n53188_, new_n53189_, new_n53190_,
    new_n53191_, new_n53192_, new_n53193_, new_n53194_, new_n53195_,
    new_n53196_, new_n53197_, new_n53198_, new_n53199_, new_n53200_,
    new_n53201_, new_n53202_, new_n53203_, new_n53204_, new_n53205_,
    new_n53206_, new_n53207_, new_n53208_, new_n53209_, new_n53210_,
    new_n53211_, new_n53212_, new_n53213_, new_n53214_, new_n53215_,
    new_n53216_, new_n53217_, new_n53218_, new_n53219_, new_n53220_,
    new_n53221_, new_n53222_, new_n53223_, new_n53224_, new_n53225_,
    new_n53226_, new_n53227_, new_n53228_, new_n53229_, new_n53230_,
    new_n53231_, new_n53232_, new_n53233_, new_n53234_, new_n53235_,
    new_n53236_, new_n53237_, new_n53238_, new_n53239_, new_n53240_,
    new_n53241_, new_n53242_, new_n53243_, new_n53244_, new_n53245_,
    new_n53246_, new_n53247_, new_n53248_, new_n53249_, new_n53250_,
    new_n53251_, new_n53252_, new_n53253_, new_n53254_, new_n53255_,
    new_n53256_, new_n53257_, new_n53258_, new_n53259_, new_n53260_,
    new_n53261_, new_n53262_, new_n53263_, new_n53264_, new_n53265_,
    new_n53266_, new_n53267_, new_n53268_, new_n53269_, new_n53270_,
    new_n53271_, new_n53272_, new_n53273_, new_n53274_, new_n53275_,
    new_n53276_, new_n53277_, new_n53278_, new_n53279_, new_n53280_,
    new_n53281_, new_n53282_, new_n53283_, new_n53284_, new_n53285_,
    new_n53286_, new_n53287_, new_n53288_, new_n53289_, new_n53290_,
    new_n53291_, new_n53292_, new_n53293_, new_n53294_, new_n53295_,
    new_n53296_, new_n53297_, new_n53298_, new_n53299_, new_n53300_,
    new_n53301_, new_n53302_, new_n53303_, new_n53304_, new_n53305_,
    new_n53306_, new_n53307_, new_n53308_, new_n53309_, new_n53310_,
    new_n53311_, new_n53312_, new_n53313_, new_n53314_, new_n53315_,
    new_n53316_, new_n53317_, new_n53318_, new_n53319_, new_n53320_,
    new_n53321_, new_n53322_, new_n53323_, new_n53324_, new_n53325_,
    new_n53326_, new_n53327_, new_n53328_, new_n53329_, new_n53330_,
    new_n53331_, new_n53332_, new_n53333_, new_n53334_, new_n53335_,
    new_n53336_, new_n53337_, new_n53338_, new_n53339_, new_n53340_,
    new_n53341_, new_n53342_, new_n53343_, new_n53344_, new_n53345_,
    new_n53346_, new_n53347_, new_n53348_, new_n53349_, new_n53350_,
    new_n53351_, new_n53352_, new_n53353_, new_n53354_, new_n53355_,
    new_n53356_, new_n53357_, new_n53358_, new_n53359_, new_n53360_,
    new_n53361_, new_n53362_, new_n53363_, new_n53364_, new_n53365_,
    new_n53366_, new_n53367_, new_n53368_, new_n53369_, new_n53370_,
    new_n53371_, new_n53372_, new_n53373_, new_n53374_, new_n53375_,
    new_n53376_, new_n53377_, new_n53378_, new_n53379_, new_n53380_,
    new_n53381_, new_n53382_, new_n53383_, new_n53384_, new_n53385_,
    new_n53386_, new_n53387_, new_n53388_, new_n53389_, new_n53390_,
    new_n53391_, new_n53392_, new_n53393_, new_n53394_, new_n53395_,
    new_n53396_, new_n53397_, new_n53398_, new_n53399_, new_n53400_,
    new_n53401_, new_n53402_, new_n53403_, new_n53404_, new_n53405_,
    new_n53406_, new_n53407_, new_n53408_, new_n53409_, new_n53410_,
    new_n53411_, new_n53412_, new_n53413_, new_n53414_, new_n53415_,
    new_n53416_, new_n53417_, new_n53418_, new_n53419_, new_n53420_,
    new_n53421_, new_n53422_, new_n53423_, new_n53424_, new_n53425_,
    new_n53426_, new_n53427_, new_n53428_, new_n53429_, new_n53430_,
    new_n53431_, new_n53432_, new_n53433_, new_n53434_, new_n53435_,
    new_n53436_, new_n53437_, new_n53438_, new_n53439_, new_n53440_,
    new_n53441_, new_n53442_, new_n53443_, new_n53444_, new_n53445_,
    new_n53446_, new_n53447_, new_n53448_, new_n53449_, new_n53450_,
    new_n53451_, new_n53452_, new_n53453_, new_n53454_, new_n53455_,
    new_n53456_, new_n53457_, new_n53458_, new_n53459_, new_n53460_,
    new_n53461_, new_n53462_, new_n53463_, new_n53464_, new_n53465_,
    new_n53466_, new_n53467_, new_n53468_, new_n53469_, new_n53470_,
    new_n53471_, new_n53472_, new_n53473_, new_n53474_, new_n53475_,
    new_n53476_, new_n53477_, new_n53478_, new_n53479_, new_n53480_,
    new_n53481_, new_n53482_, new_n53483_, new_n53484_, new_n53485_,
    new_n53486_, new_n53487_, new_n53488_, new_n53489_, new_n53490_,
    new_n53491_, new_n53492_, new_n53493_, new_n53494_, new_n53495_,
    new_n53496_, new_n53497_, new_n53498_, new_n53499_, new_n53500_,
    new_n53501_, new_n53502_, new_n53503_, new_n53504_, new_n53505_,
    new_n53506_, new_n53507_, new_n53508_, new_n53509_, new_n53510_,
    new_n53511_, new_n53512_, new_n53513_, new_n53514_, new_n53515_,
    new_n53516_, new_n53517_, new_n53518_, new_n53519_, new_n53520_,
    new_n53521_, new_n53522_, new_n53523_, new_n53524_, new_n53525_,
    new_n53526_, new_n53527_, new_n53528_, new_n53529_, new_n53530_,
    new_n53531_, new_n53532_, new_n53533_, new_n53534_, new_n53535_,
    new_n53536_, new_n53537_, new_n53538_, new_n53539_, new_n53540_,
    new_n53541_, new_n53542_, new_n53543_, new_n53544_, new_n53545_,
    new_n53546_, new_n53547_, new_n53548_, new_n53549_, new_n53550_,
    new_n53551_, new_n53552_, new_n53553_, new_n53554_, new_n53555_,
    new_n53556_, new_n53557_, new_n53558_, new_n53559_, new_n53560_,
    new_n53561_, new_n53562_, new_n53563_, new_n53564_, new_n53565_,
    new_n53566_, new_n53567_, new_n53568_, new_n53569_, new_n53570_,
    new_n53571_, new_n53572_, new_n53573_, new_n53574_, new_n53575_,
    new_n53576_, new_n53577_, new_n53578_, new_n53579_, new_n53580_,
    new_n53581_, new_n53582_, new_n53583_, new_n53584_, new_n53585_,
    new_n53586_, new_n53587_, new_n53588_, new_n53589_, new_n53590_,
    new_n53591_, new_n53592_, new_n53593_, new_n53594_, new_n53595_,
    new_n53596_, new_n53597_, new_n53598_, new_n53599_, new_n53600_,
    new_n53601_, new_n53602_, new_n53603_, new_n53604_, new_n53605_,
    new_n53606_, new_n53607_, new_n53608_, new_n53609_, new_n53610_,
    new_n53611_, new_n53612_, new_n53613_, new_n53614_, new_n53615_,
    new_n53616_, new_n53617_, new_n53618_, new_n53619_, new_n53620_,
    new_n53621_, new_n53622_, new_n53623_, new_n53624_, new_n53625_,
    new_n53626_, new_n53627_, new_n53628_, new_n53629_, new_n53630_,
    new_n53631_, new_n53632_, new_n53633_, new_n53634_, new_n53635_,
    new_n53636_, new_n53637_, new_n53638_, new_n53639_, new_n53640_,
    new_n53641_, new_n53642_, new_n53643_, new_n53644_, new_n53645_,
    new_n53646_, new_n53647_, new_n53648_, new_n53649_, new_n53650_,
    new_n53651_, new_n53652_, new_n53653_, new_n53654_, new_n53655_,
    new_n53656_, new_n53657_, new_n53658_, new_n53659_, new_n53660_,
    new_n53661_, new_n53662_, new_n53663_, new_n53664_, new_n53665_,
    new_n53666_, new_n53667_, new_n53668_, new_n53669_, new_n53670_,
    new_n53671_, new_n53672_, new_n53673_, new_n53674_, new_n53675_,
    new_n53676_, new_n53677_, new_n53678_, new_n53679_, new_n53680_,
    new_n53681_, new_n53682_, new_n53683_, new_n53684_, new_n53685_,
    new_n53686_, new_n53687_, new_n53688_, new_n53689_, new_n53690_,
    new_n53691_, new_n53692_, new_n53693_, new_n53694_, new_n53695_,
    new_n53696_, new_n53697_, new_n53698_, new_n53699_, new_n53700_,
    new_n53701_, new_n53702_, new_n53703_, new_n53704_, new_n53705_,
    new_n53706_, new_n53707_, new_n53708_, new_n53709_, new_n53710_,
    new_n53711_, new_n53712_, new_n53713_, new_n53714_, new_n53715_,
    new_n53716_, new_n53717_, new_n53718_, new_n53719_, new_n53720_,
    new_n53721_, new_n53722_, new_n53723_, new_n53724_, new_n53725_,
    new_n53726_, new_n53727_, new_n53728_, new_n53729_, new_n53730_,
    new_n53731_, new_n53732_, new_n53733_, new_n53734_, new_n53735_,
    new_n53736_, new_n53737_, new_n53738_, new_n53739_, new_n53740_,
    new_n53741_, new_n53742_, new_n53743_, new_n53744_, new_n53745_,
    new_n53746_, new_n53747_, new_n53748_, new_n53749_, new_n53750_,
    new_n53751_, new_n53752_, new_n53753_, new_n53754_, new_n53755_,
    new_n53756_, new_n53757_, new_n53758_, new_n53759_, new_n53760_,
    new_n53761_, new_n53762_, new_n53763_, new_n53764_, new_n53765_,
    new_n53766_, new_n53767_, new_n53768_, new_n53769_, new_n53770_,
    new_n53771_, new_n53772_, new_n53773_, new_n53774_, new_n53775_,
    new_n53776_, new_n53777_, new_n53778_, new_n53779_, new_n53780_,
    new_n53781_, new_n53782_, new_n53783_, new_n53784_, new_n53785_,
    new_n53786_, new_n53787_, new_n53788_, new_n53789_, new_n53790_,
    new_n53791_, new_n53792_, new_n53793_, new_n53794_, new_n53795_,
    new_n53796_, new_n53797_, new_n53798_, new_n53799_, new_n53800_,
    new_n53801_, new_n53802_, new_n53803_, new_n53804_, new_n53805_,
    new_n53806_, new_n53807_, new_n53808_, new_n53809_, new_n53810_,
    new_n53811_, new_n53812_, new_n53813_, new_n53814_, new_n53815_,
    new_n53816_, new_n53817_, new_n53818_, new_n53819_, new_n53820_,
    new_n53821_, new_n53822_, new_n53823_, new_n53824_, new_n53825_,
    new_n53826_, new_n53827_, new_n53828_, new_n53829_, new_n53830_,
    new_n53831_, new_n53832_, new_n53833_, new_n53834_, new_n53835_,
    new_n53836_, new_n53837_, new_n53838_, new_n53839_, new_n53840_,
    new_n53841_, new_n53842_, new_n53843_, new_n53844_, new_n53845_,
    new_n53846_, new_n53847_, new_n53848_, new_n53849_, new_n53850_,
    new_n53851_, new_n53852_, new_n53853_, new_n53854_, new_n53855_,
    new_n53856_, new_n53857_, new_n53858_, new_n53859_, new_n53860_,
    new_n53861_, new_n53862_, new_n53863_, new_n53864_, new_n53865_,
    new_n53866_, new_n53867_, new_n53868_, new_n53869_, new_n53870_,
    new_n53871_, new_n53872_, new_n53873_, new_n53874_, new_n53875_,
    new_n53876_, new_n53877_, new_n53878_, new_n53879_, new_n53880_,
    new_n53881_, new_n53882_, new_n53883_, new_n53884_, new_n53885_,
    new_n53886_, new_n53887_, new_n53888_, new_n53889_, new_n53890_,
    new_n53891_, new_n53892_, new_n53893_, new_n53894_, new_n53895_,
    new_n53896_, new_n53897_, new_n53898_, new_n53899_, new_n53900_,
    new_n53901_, new_n53902_, new_n53903_, new_n53904_, new_n53905_,
    new_n53906_, new_n53907_, new_n53908_, new_n53909_, new_n53910_,
    new_n53911_, new_n53912_, new_n53913_, new_n53914_, new_n53915_,
    new_n53916_, new_n53917_, new_n53918_, new_n53919_, new_n53920_,
    new_n53921_, new_n53922_, new_n53923_, new_n53924_, new_n53925_,
    new_n53926_, new_n53927_, new_n53928_, new_n53929_, new_n53930_,
    new_n53931_, new_n53932_, new_n53933_, new_n53934_, new_n53935_,
    new_n53936_, new_n53937_, new_n53938_, new_n53939_, new_n53940_,
    new_n53941_, new_n53942_, new_n53943_, new_n53944_, new_n53945_,
    new_n53946_, new_n53947_, new_n53948_, new_n53949_, new_n53950_,
    new_n53951_, new_n53952_, new_n53953_, new_n53954_, new_n53955_,
    new_n53956_, new_n53957_, new_n53958_, new_n53959_, new_n53960_,
    new_n53961_, new_n53962_, new_n53963_, new_n53964_, new_n53965_,
    new_n53966_, new_n53967_, new_n53968_, new_n53969_, new_n53970_,
    new_n53971_, new_n53972_, new_n53973_, new_n53974_, new_n53975_,
    new_n53976_, new_n53977_, new_n53978_, new_n53979_, new_n53980_,
    new_n53981_, new_n53982_, new_n53983_, new_n53984_, new_n53985_,
    new_n53986_, new_n53987_, new_n53988_, new_n53989_, new_n53990_,
    new_n53991_, new_n53992_, new_n53993_, new_n53994_, new_n53995_,
    new_n53996_, new_n53997_, new_n53998_, new_n53999_, new_n54000_,
    new_n54001_, new_n54002_, new_n54003_, new_n54004_, new_n54005_,
    new_n54006_, new_n54007_, new_n54008_, new_n54009_, new_n54010_,
    new_n54011_, new_n54012_, new_n54013_, new_n54014_, new_n54015_,
    new_n54016_, new_n54017_, new_n54018_, new_n54019_, new_n54020_,
    new_n54021_, new_n54022_, new_n54023_, new_n54024_, new_n54025_,
    new_n54026_, new_n54027_, new_n54028_, new_n54029_, new_n54030_,
    new_n54031_, new_n54032_, new_n54033_, new_n54034_, new_n54035_,
    new_n54036_, new_n54037_, new_n54038_, new_n54039_, new_n54040_,
    new_n54041_, new_n54042_, new_n54043_, new_n54044_, new_n54045_,
    new_n54046_, new_n54047_, new_n54048_, new_n54049_, new_n54050_,
    new_n54051_, new_n54052_, new_n54053_, new_n54054_, new_n54055_,
    new_n54056_, new_n54057_, new_n54058_, new_n54059_, new_n54060_,
    new_n54061_, new_n54062_, new_n54063_, new_n54064_, new_n54065_,
    new_n54066_, new_n54067_, new_n54068_, new_n54069_, new_n54070_,
    new_n54071_, new_n54072_, new_n54073_, new_n54074_, new_n54075_,
    new_n54076_, new_n54077_, new_n54078_, new_n54079_, new_n54080_,
    new_n54081_, new_n54082_, new_n54083_, new_n54084_, new_n54085_,
    new_n54086_, new_n54087_, new_n54088_, new_n54089_, new_n54090_,
    new_n54091_, new_n54092_, new_n54093_, new_n54094_, new_n54095_,
    new_n54096_, new_n54097_, new_n54098_, new_n54099_, new_n54100_,
    new_n54101_, new_n54102_, new_n54103_, new_n54104_, new_n54105_,
    new_n54106_, new_n54107_, new_n54108_, new_n54109_, new_n54110_,
    new_n54111_, new_n54112_, new_n54113_, new_n54114_, new_n54115_,
    new_n54116_, new_n54117_, new_n54118_, new_n54119_, new_n54120_,
    new_n54121_, new_n54122_, new_n54123_, new_n54124_, new_n54125_,
    new_n54126_, new_n54127_, new_n54128_, new_n54129_, new_n54130_,
    new_n54131_, new_n54132_, new_n54133_, new_n54134_, new_n54135_,
    new_n54136_, new_n54137_, new_n54138_, new_n54139_, new_n54140_,
    new_n54141_, new_n54142_, new_n54143_, new_n54144_, new_n54145_,
    new_n54146_, new_n54147_, new_n54148_, new_n54149_, new_n54150_,
    new_n54151_, new_n54152_, new_n54153_, new_n54154_, new_n54155_,
    new_n54156_, new_n54157_, new_n54158_, new_n54159_, new_n54160_,
    new_n54161_, new_n54162_, new_n54163_, new_n54164_, new_n54165_,
    new_n54166_, new_n54167_, new_n54168_, new_n54169_, new_n54170_,
    new_n54171_, new_n54172_, new_n54173_, new_n54174_, new_n54175_,
    new_n54176_, new_n54177_, new_n54178_, new_n54179_, new_n54180_,
    new_n54181_, new_n54182_, new_n54183_, new_n54184_, new_n54185_,
    new_n54186_, new_n54187_, new_n54188_, new_n54189_, new_n54190_,
    new_n54191_, new_n54192_, new_n54193_, new_n54194_, new_n54195_,
    new_n54196_, new_n54197_, new_n54198_, new_n54199_, new_n54200_,
    new_n54201_, new_n54202_, new_n54203_, new_n54204_, new_n54205_,
    new_n54206_, new_n54207_, new_n54208_, new_n54209_, new_n54210_,
    new_n54211_, new_n54212_, new_n54213_, new_n54214_, new_n54215_,
    new_n54216_, new_n54217_, new_n54218_, new_n54219_, new_n54220_,
    new_n54221_, new_n54222_, new_n54223_, new_n54224_, new_n54225_,
    new_n54226_, new_n54227_, new_n54228_, new_n54229_, new_n54230_,
    new_n54231_, new_n54232_, new_n54233_, new_n54234_, new_n54235_,
    new_n54236_, new_n54237_, new_n54238_, new_n54239_, new_n54240_,
    new_n54241_, new_n54242_, new_n54243_, new_n54244_, new_n54245_,
    new_n54246_, new_n54247_, new_n54248_, new_n54249_, new_n54250_,
    new_n54251_, new_n54252_, new_n54253_, new_n54254_, new_n54255_,
    new_n54256_, new_n54257_, new_n54258_, new_n54259_, new_n54260_,
    new_n54261_, new_n54262_, new_n54263_, new_n54264_, new_n54265_,
    new_n54266_, new_n54267_, new_n54268_, new_n54269_, new_n54270_,
    new_n54271_, new_n54272_, new_n54273_, new_n54274_, new_n54275_,
    new_n54276_, new_n54277_, new_n54278_, new_n54279_, new_n54280_,
    new_n54281_, new_n54282_, new_n54283_, new_n54284_, new_n54285_,
    new_n54286_, new_n54287_, new_n54288_, new_n54289_, new_n54290_,
    new_n54291_, new_n54292_, new_n54293_, new_n54294_, new_n54295_,
    new_n54296_, new_n54297_, new_n54298_, new_n54299_, new_n54300_,
    new_n54301_, new_n54302_, new_n54303_, new_n54304_, new_n54305_,
    new_n54306_, new_n54307_, new_n54308_, new_n54309_, new_n54310_,
    new_n54311_, new_n54312_, new_n54313_, new_n54314_, new_n54315_,
    new_n54316_, new_n54317_, new_n54318_, new_n54319_, new_n54320_,
    new_n54321_, new_n54322_, new_n54323_, new_n54324_, new_n54325_,
    new_n54326_, new_n54327_, new_n54328_, new_n54329_, new_n54330_,
    new_n54331_, new_n54332_, new_n54333_, new_n54334_, new_n54335_,
    new_n54336_, new_n54337_, new_n54338_, new_n54339_, new_n54340_,
    new_n54341_, new_n54342_, new_n54343_, new_n54344_, new_n54345_,
    new_n54346_, new_n54347_, new_n54348_, new_n54349_, new_n54350_,
    new_n54351_, new_n54352_, new_n54353_, new_n54354_, new_n54355_,
    new_n54356_, new_n54357_, new_n54358_, new_n54359_, new_n54360_,
    new_n54361_, new_n54362_, new_n54363_, new_n54364_, new_n54365_,
    new_n54366_, new_n54367_, new_n54368_, new_n54369_, new_n54370_,
    new_n54371_, new_n54372_, new_n54373_, new_n54374_, new_n54375_,
    new_n54376_, new_n54377_, new_n54378_, new_n54379_, new_n54380_,
    new_n54381_, new_n54382_, new_n54383_, new_n54384_, new_n54385_,
    new_n54386_, new_n54387_, new_n54388_, new_n54389_, new_n54390_,
    new_n54391_, new_n54392_, new_n54393_, new_n54394_, new_n54395_,
    new_n54396_, new_n54397_, new_n54398_, new_n54399_, new_n54400_,
    new_n54401_, new_n54402_, new_n54403_, new_n54404_, new_n54405_,
    new_n54406_, new_n54407_, new_n54408_, new_n54409_, new_n54410_,
    new_n54411_, new_n54412_, new_n54413_, new_n54414_, new_n54415_,
    new_n54416_, new_n54417_, new_n54418_, new_n54419_, new_n54420_,
    new_n54421_, new_n54422_, new_n54423_, new_n54424_, new_n54425_,
    new_n54426_, new_n54427_, new_n54428_, new_n54429_, new_n54430_,
    new_n54431_, new_n54432_, new_n54433_, new_n54434_, new_n54435_,
    new_n54436_, new_n54437_, new_n54438_, new_n54439_, new_n54440_,
    new_n54441_, new_n54442_, new_n54443_, new_n54444_, new_n54445_,
    new_n54446_, new_n54447_, new_n54448_, new_n54449_, new_n54450_,
    new_n54451_, new_n54452_, new_n54453_, new_n54454_, new_n54455_,
    new_n54456_, new_n54457_, new_n54458_, new_n54459_, new_n54460_,
    new_n54461_, new_n54462_, new_n54463_, new_n54464_, new_n54465_,
    new_n54466_, new_n54467_, new_n54468_, new_n54469_, new_n54470_,
    new_n54471_, new_n54472_, new_n54473_, new_n54474_, new_n54475_,
    new_n54476_, new_n54477_, new_n54478_, new_n54479_, new_n54480_,
    new_n54481_, new_n54482_, new_n54483_, new_n54484_, new_n54485_,
    new_n54486_, new_n54487_, new_n54488_, new_n54489_, new_n54490_,
    new_n54491_, new_n54492_, new_n54493_, new_n54494_, new_n54495_,
    new_n54496_, new_n54497_, new_n54498_, new_n54499_, new_n54500_,
    new_n54501_, new_n54502_, new_n54503_, new_n54504_, new_n54505_,
    new_n54506_, new_n54507_, new_n54508_, new_n54509_, new_n54510_,
    new_n54511_, new_n54512_, new_n54513_, new_n54514_, new_n54515_,
    new_n54516_, new_n54517_, new_n54518_, new_n54519_, new_n54520_,
    new_n54521_, new_n54522_, new_n54523_, new_n54524_, new_n54525_,
    new_n54526_, new_n54527_, new_n54528_, new_n54529_, new_n54530_,
    new_n54531_, new_n54532_, new_n54533_, new_n54534_, new_n54535_,
    new_n54536_, new_n54537_, new_n54538_, new_n54539_, new_n54540_,
    new_n54541_, new_n54542_, new_n54543_, new_n54544_, new_n54545_,
    new_n54546_, new_n54547_, new_n54548_, new_n54549_, new_n54550_,
    new_n54551_, new_n54552_, new_n54553_, new_n54554_, new_n54555_,
    new_n54556_, new_n54557_, new_n54558_, new_n54559_, new_n54560_,
    new_n54561_, new_n54562_, new_n54563_, new_n54564_, new_n54565_,
    new_n54566_, new_n54567_, new_n54568_, new_n54569_, new_n54570_,
    new_n54571_, new_n54572_, new_n54573_, new_n54574_, new_n54575_,
    new_n54576_, new_n54577_, new_n54578_, new_n54579_, new_n54580_,
    new_n54581_, new_n54582_, new_n54583_, new_n54584_, new_n54585_,
    new_n54586_, new_n54587_, new_n54588_, new_n54589_, new_n54590_,
    new_n54591_, new_n54592_, new_n54593_, new_n54594_, new_n54595_,
    new_n54596_, new_n54597_, new_n54598_, new_n54599_, new_n54600_,
    new_n54601_, new_n54602_, new_n54603_, new_n54604_, new_n54605_,
    new_n54606_, new_n54607_, new_n54608_, new_n54609_, new_n54610_,
    new_n54611_, new_n54612_, new_n54613_, new_n54614_, new_n54615_,
    new_n54616_, new_n54617_, new_n54618_, new_n54619_, new_n54620_,
    new_n54621_, new_n54622_, new_n54623_, new_n54624_, new_n54625_,
    new_n54626_, new_n54627_, new_n54628_, new_n54629_, new_n54630_,
    new_n54631_, new_n54632_, new_n54633_, new_n54634_, new_n54635_,
    new_n54636_, new_n54637_, new_n54638_, new_n54639_, new_n54640_,
    new_n54641_, new_n54642_, new_n54643_, new_n54644_, new_n54645_,
    new_n54646_, new_n54647_, new_n54648_, new_n54649_, new_n54650_,
    new_n54651_, new_n54652_, new_n54653_, new_n54654_, new_n54655_,
    new_n54656_, new_n54657_, new_n54658_, new_n54659_, new_n54660_,
    new_n54661_, new_n54662_, new_n54663_, new_n54664_, new_n54665_,
    new_n54666_, new_n54667_, new_n54668_, new_n54669_, new_n54670_,
    new_n54671_, new_n54672_, new_n54673_, new_n54674_, new_n54675_,
    new_n54676_, new_n54677_, new_n54678_, new_n54679_, new_n54680_,
    new_n54681_, new_n54682_, new_n54683_, new_n54684_, new_n54685_,
    new_n54686_, new_n54687_, new_n54688_, new_n54689_, new_n54690_,
    new_n54691_, new_n54692_, new_n54693_, new_n54694_, new_n54695_,
    new_n54696_, new_n54697_, new_n54698_, new_n54699_, new_n54700_,
    new_n54701_, new_n54702_, new_n54703_, new_n54704_, new_n54705_,
    new_n54706_, new_n54707_, new_n54708_, new_n54709_, new_n54710_,
    new_n54711_, new_n54712_, new_n54713_, new_n54714_, new_n54715_,
    new_n54716_, new_n54717_, new_n54718_, new_n54719_, new_n54720_,
    new_n54721_, new_n54722_, new_n54723_, new_n54724_, new_n54725_,
    new_n54726_, new_n54727_, new_n54728_, new_n54729_, new_n54730_,
    new_n54731_, new_n54732_, new_n54733_, new_n54734_, new_n54735_,
    new_n54736_, new_n54737_, new_n54738_, new_n54739_, new_n54740_,
    new_n54741_, new_n54742_, new_n54743_, new_n54744_, new_n54745_,
    new_n54746_, new_n54747_, new_n54748_, new_n54749_, new_n54750_,
    new_n54751_, new_n54752_, new_n54753_, new_n54754_, new_n54755_,
    new_n54756_, new_n54757_, new_n54758_, new_n54759_, new_n54760_,
    new_n54761_, new_n54762_, new_n54763_, new_n54764_, new_n54765_,
    new_n54766_, new_n54767_, new_n54768_, new_n54769_, new_n54770_,
    new_n54771_, new_n54772_, new_n54773_, new_n54774_, new_n54775_,
    new_n54776_, new_n54777_, new_n54778_, new_n54779_, new_n54780_,
    new_n54781_, new_n54782_, new_n54783_, new_n54784_, new_n54785_,
    new_n54786_, new_n54787_, new_n54788_, new_n54789_, new_n54790_,
    new_n54791_, new_n54792_, new_n54793_, new_n54794_, new_n54795_,
    new_n54796_, new_n54797_, new_n54798_, new_n54799_, new_n54800_,
    new_n54801_, new_n54802_, new_n54803_, new_n54804_, new_n54805_,
    new_n54806_, new_n54807_, new_n54808_, new_n54809_, new_n54810_,
    new_n54811_, new_n54812_, new_n54813_, new_n54814_, new_n54815_,
    new_n54816_, new_n54817_, new_n54818_, new_n54819_, new_n54820_,
    new_n54821_, new_n54822_, new_n54823_, new_n54824_, new_n54825_,
    new_n54826_, new_n54827_, new_n54828_, new_n54829_, new_n54830_,
    new_n54831_, new_n54832_, new_n54833_, new_n54834_, new_n54835_,
    new_n54836_, new_n54837_, new_n54838_, new_n54839_, new_n54840_,
    new_n54841_, new_n54842_, new_n54843_, new_n54844_, new_n54845_,
    new_n54846_, new_n54847_, new_n54848_, new_n54849_, new_n54850_,
    new_n54851_, new_n54852_, new_n54853_, new_n54854_, new_n54855_,
    new_n54856_, new_n54857_, new_n54858_, new_n54859_, new_n54860_,
    new_n54861_, new_n54862_, new_n54863_, new_n54864_, new_n54865_,
    new_n54866_, new_n54867_, new_n54868_, new_n54869_, new_n54870_,
    new_n54871_, new_n54872_, new_n54873_, new_n54874_, new_n54875_,
    new_n54876_, new_n54877_, new_n54878_, new_n54879_, new_n54880_,
    new_n54881_, new_n54882_, new_n54883_, new_n54884_, new_n54885_,
    new_n54886_, new_n54887_, new_n54888_, new_n54889_, new_n54890_,
    new_n54891_, new_n54892_, new_n54893_, new_n54894_, new_n54895_,
    new_n54896_, new_n54897_, new_n54898_, new_n54899_, new_n54900_,
    new_n54901_, new_n54902_, new_n54903_, new_n54904_, new_n54905_,
    new_n54906_, new_n54907_, new_n54908_, new_n54909_, new_n54910_,
    new_n54911_, new_n54912_, new_n54913_, new_n54914_, new_n54915_,
    new_n54916_, new_n54917_, new_n54918_, new_n54919_, new_n54920_,
    new_n54921_, new_n54922_, new_n54923_, new_n54924_, new_n54925_,
    new_n54926_, new_n54927_, new_n54928_, new_n54929_, new_n54930_,
    new_n54931_, new_n54932_, new_n54933_, new_n54934_, new_n54935_,
    new_n54936_, new_n54937_, new_n54938_, new_n54939_, new_n54940_,
    new_n54941_, new_n54942_, new_n54943_, new_n54944_, new_n54945_,
    new_n54946_, new_n54947_, new_n54948_, new_n54949_, new_n54950_,
    new_n54951_, new_n54952_, new_n54953_, new_n54954_, new_n54955_,
    new_n54956_, new_n54957_, new_n54958_, new_n54959_, new_n54960_,
    new_n54961_, new_n54962_, new_n54963_, new_n54964_, new_n54965_,
    new_n54966_, new_n54967_, new_n54968_, new_n54969_, new_n54970_,
    new_n54971_, new_n54972_, new_n54973_, new_n54974_, new_n54975_,
    new_n54976_, new_n54977_, new_n54978_, new_n54979_, new_n54980_,
    new_n54981_, new_n54982_, new_n54983_, new_n54984_, new_n54985_,
    new_n54986_, new_n54987_, new_n54988_, new_n54989_, new_n54990_,
    new_n54991_, new_n54992_, new_n54993_, new_n54994_, new_n54995_,
    new_n54996_, new_n54997_, new_n54998_, new_n54999_, new_n55000_,
    new_n55001_, new_n55002_, new_n55003_, new_n55004_, new_n55005_,
    new_n55006_, new_n55007_, new_n55008_, new_n55009_, new_n55010_,
    new_n55011_, new_n55012_, new_n55013_, new_n55014_, new_n55015_,
    new_n55016_, new_n55017_, new_n55018_, new_n55019_, new_n55020_,
    new_n55021_, new_n55022_, new_n55023_, new_n55024_, new_n55025_,
    new_n55026_, new_n55027_, new_n55028_, new_n55029_, new_n55030_,
    new_n55031_, new_n55032_, new_n55033_, new_n55034_, new_n55035_,
    new_n55036_, new_n55037_, new_n55038_, new_n55039_, new_n55040_,
    new_n55041_, new_n55042_, new_n55043_, new_n55044_, new_n55045_,
    new_n55046_, new_n55047_, new_n55048_, new_n55049_, new_n55050_,
    new_n55051_, new_n55052_, new_n55053_, new_n55054_, new_n55055_,
    new_n55056_, new_n55057_, new_n55058_, new_n55059_, new_n55060_,
    new_n55061_, new_n55062_, new_n55063_, new_n55064_, new_n55065_,
    new_n55066_, new_n55067_, new_n55068_, new_n55069_, new_n55070_,
    new_n55071_, new_n55072_, new_n55073_, new_n55074_, new_n55075_,
    new_n55076_, new_n55077_, new_n55078_, new_n55079_, new_n55080_,
    new_n55081_, new_n55082_, new_n55083_, new_n55084_, new_n55085_,
    new_n55086_, new_n55087_, new_n55088_, new_n55089_, new_n55090_,
    new_n55091_, new_n55092_, new_n55093_, new_n55094_, new_n55095_,
    new_n55096_, new_n55097_, new_n55098_, new_n55099_, new_n55100_,
    new_n55101_, new_n55102_, new_n55103_, new_n55104_, new_n55105_,
    new_n55106_, new_n55107_, new_n55108_, new_n55109_, new_n55110_,
    new_n55111_, new_n55112_, new_n55113_, new_n55114_, new_n55115_,
    new_n55116_, new_n55117_, new_n55118_, new_n55119_, new_n55120_,
    new_n55121_, new_n55122_, new_n55123_, new_n55124_, new_n55125_,
    new_n55126_, new_n55127_, new_n55128_, new_n55129_, new_n55130_,
    new_n55131_, new_n55132_, new_n55133_, new_n55134_, new_n55135_,
    new_n55136_, new_n55137_, new_n55138_, new_n55139_, new_n55140_,
    new_n55141_, new_n55142_, new_n55143_, new_n55144_, new_n55145_,
    new_n55146_, new_n55147_, new_n55148_, new_n55149_, new_n55150_,
    new_n55151_, new_n55152_, new_n55153_, new_n55154_, new_n55155_,
    new_n55156_, new_n55157_, new_n55158_, new_n55159_, new_n55160_,
    new_n55161_, new_n55162_, new_n55163_, new_n55164_, new_n55165_,
    new_n55166_, new_n55167_, new_n55168_, new_n55169_, new_n55170_,
    new_n55171_, new_n55172_, new_n55173_, new_n55174_, new_n55175_,
    new_n55176_, new_n55177_, new_n55178_, new_n55179_, new_n55180_,
    new_n55181_, new_n55182_, new_n55183_, new_n55184_, new_n55185_,
    new_n55186_, new_n55187_, new_n55188_, new_n55189_, new_n55190_,
    new_n55191_, new_n55192_, new_n55193_, new_n55194_, new_n55195_,
    new_n55196_, new_n55197_, new_n55198_, new_n55199_, new_n55200_,
    new_n55201_, new_n55202_, new_n55203_, new_n55204_, new_n55205_,
    new_n55206_, new_n55207_, new_n55208_, new_n55209_, new_n55210_,
    new_n55211_, new_n55212_, new_n55213_, new_n55214_, new_n55215_,
    new_n55216_, new_n55217_, new_n55218_, new_n55219_, new_n55220_,
    new_n55221_, new_n55222_, new_n55223_, new_n55224_, new_n55225_,
    new_n55226_, new_n55227_, new_n55228_, new_n55229_, new_n55230_,
    new_n55231_, new_n55232_, new_n55233_, new_n55234_, new_n55235_,
    new_n55236_, new_n55237_, new_n55238_, new_n55239_, new_n55240_,
    new_n55241_, new_n55242_, new_n55243_, new_n55244_, new_n55245_,
    new_n55246_, new_n55247_, new_n55248_, new_n55249_, new_n55250_,
    new_n55251_, new_n55252_, new_n55253_, new_n55254_, new_n55255_,
    new_n55256_, new_n55257_, new_n55258_, new_n55259_, new_n55260_,
    new_n55261_, new_n55262_, new_n55263_, new_n55264_, new_n55265_,
    new_n55266_, new_n55267_, new_n55268_, new_n55269_, new_n55270_,
    new_n55271_, new_n55272_, new_n55273_, new_n55274_, new_n55275_,
    new_n55276_, new_n55277_, new_n55278_, new_n55279_, new_n55280_,
    new_n55281_, new_n55282_, new_n55283_, new_n55284_, new_n55285_,
    new_n55286_, new_n55287_, new_n55288_, new_n55289_, new_n55290_,
    new_n55291_, new_n55292_, new_n55293_, new_n55294_, new_n55295_,
    new_n55296_, new_n55297_, new_n55298_, new_n55299_, new_n55300_,
    new_n55301_, new_n55302_, new_n55303_, new_n55304_, new_n55305_,
    new_n55306_, new_n55307_, new_n55308_, new_n55309_, new_n55310_,
    new_n55311_, new_n55312_, new_n55313_, new_n55314_, new_n55315_,
    new_n55316_, new_n55317_, new_n55318_, new_n55319_, new_n55320_,
    new_n55321_, new_n55322_, new_n55323_, new_n55324_, new_n55325_,
    new_n55326_, new_n55327_, new_n55328_, new_n55329_, new_n55330_,
    new_n55331_, new_n55332_, new_n55333_, new_n55334_, new_n55335_,
    new_n55336_, new_n55337_, new_n55338_, new_n55339_, new_n55340_,
    new_n55341_, new_n55342_, new_n55343_, new_n55344_, new_n55345_,
    new_n55346_, new_n55347_, new_n55348_, new_n55349_, new_n55350_,
    new_n55351_, new_n55352_, new_n55353_, new_n55354_, new_n55355_,
    new_n55356_, new_n55357_, new_n55358_, new_n55359_, new_n55360_,
    new_n55361_, new_n55362_, new_n55363_, new_n55364_, new_n55365_,
    new_n55366_, new_n55367_, new_n55368_, new_n55369_, new_n55370_,
    new_n55371_, new_n55372_, new_n55373_, new_n55374_, new_n55375_,
    new_n55376_, new_n55377_, new_n55378_, new_n55379_, new_n55380_,
    new_n55381_, new_n55382_, new_n55383_, new_n55384_, new_n55385_,
    new_n55386_, new_n55387_, new_n55388_, new_n55389_, new_n55390_,
    new_n55391_, new_n55392_, new_n55393_, new_n55394_, new_n55395_,
    new_n55396_, new_n55397_, new_n55398_, new_n55399_, new_n55400_,
    new_n55401_, new_n55402_, new_n55403_, new_n55404_, new_n55405_,
    new_n55406_, new_n55407_, new_n55408_, new_n55409_, new_n55410_,
    new_n55411_, new_n55412_, new_n55413_, new_n55414_, new_n55415_,
    new_n55416_, new_n55417_, new_n55418_, new_n55419_, new_n55420_,
    new_n55421_, new_n55422_, new_n55423_, new_n55424_, new_n55425_,
    new_n55426_, new_n55427_, new_n55428_, new_n55429_, new_n55430_,
    new_n55431_, new_n55432_, new_n55433_, new_n55434_, new_n55435_,
    new_n55436_, new_n55437_, new_n55438_, new_n55439_, new_n55440_,
    new_n55441_, new_n55442_, new_n55443_, new_n55444_, new_n55445_,
    new_n55446_, new_n55447_, new_n55448_, new_n55449_, new_n55450_,
    new_n55451_, new_n55452_, new_n55453_, new_n55454_, new_n55455_,
    new_n55456_, new_n55457_, new_n55458_, new_n55459_, new_n55460_,
    new_n55461_, new_n55462_, new_n55463_, new_n55464_, new_n55465_,
    new_n55466_, new_n55467_, new_n55468_, new_n55469_, new_n55470_,
    new_n55471_, new_n55472_, new_n55473_, new_n55474_, new_n55475_,
    new_n55476_, new_n55477_, new_n55478_, new_n55479_, new_n55480_,
    new_n55481_, new_n55482_, new_n55483_, new_n55484_, new_n55485_,
    new_n55486_, new_n55487_, new_n55488_, new_n55489_, new_n55490_,
    new_n55491_, new_n55492_, new_n55493_, new_n55494_, new_n55495_,
    new_n55496_, new_n55497_, new_n55498_, new_n55499_, new_n55500_,
    new_n55501_, new_n55502_, new_n55503_, new_n55504_, new_n55505_,
    new_n55506_, new_n55507_, new_n55508_, new_n55509_, new_n55510_,
    new_n55511_, new_n55512_, new_n55513_, new_n55514_, new_n55515_,
    new_n55516_, new_n55517_, new_n55518_, new_n55519_, new_n55520_,
    new_n55521_, new_n55522_, new_n55523_, new_n55524_, new_n55525_,
    new_n55526_, new_n55527_, new_n55528_, new_n55529_, new_n55530_,
    new_n55531_, new_n55532_, new_n55533_, new_n55534_, new_n55535_,
    new_n55536_, new_n55537_, new_n55538_, new_n55539_, new_n55540_,
    new_n55541_, new_n55542_, new_n55543_, new_n55544_, new_n55545_,
    new_n55546_, new_n55547_, new_n55548_, new_n55549_, new_n55550_,
    new_n55551_, new_n55552_, new_n55553_, new_n55554_, new_n55555_,
    new_n55556_, new_n55557_, new_n55558_, new_n55559_, new_n55560_,
    new_n55561_, new_n55562_, new_n55563_, new_n55564_, new_n55565_,
    new_n55566_, new_n55567_, new_n55568_, new_n55569_, new_n55570_,
    new_n55571_, new_n55572_, new_n55573_, new_n55574_, new_n55575_,
    new_n55576_, new_n55577_, new_n55578_, new_n55579_, new_n55580_,
    new_n55581_, new_n55582_, new_n55583_, new_n55584_, new_n55585_,
    new_n55586_, new_n55587_, new_n55588_, new_n55589_, new_n55590_,
    new_n55591_, new_n55592_, new_n55593_, new_n55594_, new_n55595_,
    new_n55596_, new_n55597_, new_n55598_, new_n55599_, new_n55600_,
    new_n55601_, new_n55602_, new_n55603_, new_n55604_, new_n55605_,
    new_n55606_, new_n55607_, new_n55608_, new_n55609_, new_n55610_,
    new_n55611_, new_n55612_, new_n55613_, new_n55614_, new_n55615_,
    new_n55616_, new_n55617_, new_n55618_, new_n55619_, new_n55620_,
    new_n55621_, new_n55622_, new_n55623_, new_n55624_, new_n55625_,
    new_n55626_, new_n55627_, new_n55628_, new_n55629_, new_n55630_,
    new_n55631_, new_n55632_, new_n55633_, new_n55634_, new_n55635_,
    new_n55636_, new_n55637_, new_n55638_, new_n55639_, new_n55640_,
    new_n55641_, new_n55642_, new_n55643_, new_n55644_, new_n55645_,
    new_n55646_, new_n55647_, new_n55648_, new_n55649_, new_n55650_,
    new_n55651_, new_n55652_, new_n55653_, new_n55654_, new_n55655_,
    new_n55656_, new_n55657_, new_n55658_, new_n55659_, new_n55660_,
    new_n55661_, new_n55662_, new_n55663_, new_n55664_, new_n55665_,
    new_n55666_, new_n55667_, new_n55668_, new_n55669_, new_n55670_,
    new_n55671_, new_n55672_, new_n55673_, new_n55674_, new_n55675_,
    new_n55676_, new_n55677_, new_n55678_, new_n55679_, new_n55680_,
    new_n55681_, new_n55682_, new_n55683_, new_n55684_, new_n55685_,
    new_n55686_, new_n55687_, new_n55688_, new_n55689_, new_n55690_,
    new_n55691_, new_n55692_, new_n55693_, new_n55694_, new_n55695_,
    new_n55696_, new_n55697_, new_n55698_, new_n55699_, new_n55700_,
    new_n55701_, new_n55702_, new_n55703_, new_n55704_, new_n55705_,
    new_n55706_, new_n55707_, new_n55708_, new_n55709_, new_n55710_,
    new_n55711_, new_n55712_, new_n55713_, new_n55714_, new_n55715_,
    new_n55716_, new_n55717_, new_n55718_, new_n55719_, new_n55720_,
    new_n55721_, new_n55722_, new_n55723_, new_n55724_, new_n55725_,
    new_n55726_, new_n55727_, new_n55728_, new_n55729_, new_n55730_,
    new_n55731_, new_n55732_, new_n55733_, new_n55734_, new_n55735_,
    new_n55736_, new_n55737_, new_n55738_, new_n55739_, new_n55740_,
    new_n55741_, new_n55742_, new_n55743_, new_n55744_, new_n55745_,
    new_n55746_, new_n55747_, new_n55748_, new_n55749_, new_n55750_,
    new_n55751_, new_n55752_, new_n55753_, new_n55754_, new_n55755_,
    new_n55756_, new_n55757_, new_n55758_, new_n55759_, new_n55760_,
    new_n55761_, new_n55762_, new_n55763_, new_n55764_, new_n55765_,
    new_n55766_, new_n55767_, new_n55768_, new_n55769_, new_n55770_,
    new_n55771_, new_n55772_, new_n55773_, new_n55774_, new_n55775_,
    new_n55776_, new_n55777_, new_n55778_, new_n55779_, new_n55780_,
    new_n55781_, new_n55782_, new_n55783_, new_n55784_, new_n55785_,
    new_n55786_, new_n55787_, new_n55788_, new_n55789_, new_n55790_,
    new_n55791_, new_n55792_, new_n55793_, new_n55794_, new_n55795_,
    new_n55796_, new_n55797_, new_n55798_, new_n55799_, new_n55800_,
    new_n55801_, new_n55802_, new_n55803_, new_n55804_, new_n55805_,
    new_n55806_, new_n55807_, new_n55808_, new_n55809_, new_n55810_,
    new_n55811_, new_n55812_, new_n55813_, new_n55814_, new_n55815_,
    new_n55816_, new_n55817_, new_n55818_, new_n55819_, new_n55820_,
    new_n55821_, new_n55822_, new_n55823_, new_n55824_, new_n55825_,
    new_n55826_, new_n55827_, new_n55828_, new_n55829_, new_n55830_,
    new_n55831_, new_n55832_, new_n55833_, new_n55834_, new_n55835_,
    new_n55836_, new_n55837_, new_n55838_, new_n55839_, new_n55840_,
    new_n55841_, new_n55842_, new_n55843_, new_n55844_, new_n55845_,
    new_n55846_, new_n55847_, new_n55848_, new_n55849_, new_n55850_,
    new_n55851_, new_n55852_, new_n55853_, new_n55854_, new_n55855_,
    new_n55856_, new_n55857_, new_n55858_, new_n55859_, new_n55860_,
    new_n55861_, new_n55862_, new_n55863_, new_n55864_, new_n55865_,
    new_n55866_, new_n55867_, new_n55868_, new_n55869_, new_n55870_,
    new_n55871_, new_n55872_, new_n55873_, new_n55874_, new_n55875_,
    new_n55876_, new_n55877_, new_n55878_, new_n55879_, new_n55880_,
    new_n55881_, new_n55882_, new_n55883_, new_n55884_, new_n55885_,
    new_n55886_, new_n55887_, new_n55888_, new_n55889_, new_n55890_,
    new_n55891_, new_n55892_, new_n55893_, new_n55894_, new_n55895_,
    new_n55896_, new_n55897_, new_n55898_, new_n55899_, new_n55900_,
    new_n55901_, new_n55902_, new_n55903_, new_n55904_, new_n55905_,
    new_n55906_, new_n55907_, new_n55908_, new_n55909_, new_n55910_,
    new_n55911_, new_n55912_, new_n55913_, new_n55914_, new_n55915_,
    new_n55916_, new_n55917_, new_n55918_, new_n55919_, new_n55920_,
    new_n55921_, new_n55922_, new_n55923_, new_n55924_, new_n55925_,
    new_n55926_, new_n55927_, new_n55928_, new_n55929_, new_n55930_,
    new_n55931_, new_n55932_, new_n55933_, new_n55934_, new_n55935_,
    new_n55936_, new_n55937_, new_n55938_, new_n55939_, new_n55940_,
    new_n55941_, new_n55942_, new_n55943_, new_n55944_, new_n55945_,
    new_n55946_, new_n55947_, new_n55948_, new_n55949_, new_n55950_,
    new_n55951_, new_n55952_, new_n55953_, new_n55954_, new_n55955_,
    new_n55956_, new_n55957_, new_n55958_, new_n55959_, new_n55960_,
    new_n55961_, new_n55962_, new_n55963_, new_n55964_, new_n55965_,
    new_n55966_, new_n55967_, new_n55968_, new_n55969_, new_n55970_,
    new_n55971_, new_n55972_, new_n55973_, new_n55974_, new_n55975_,
    new_n55976_, new_n55977_, new_n55978_, new_n55979_, new_n55980_,
    new_n55981_, new_n55982_, new_n55983_, new_n55984_, new_n55985_,
    new_n55986_, new_n55987_, new_n55988_, new_n55989_, new_n55990_,
    new_n55991_, new_n55992_, new_n55993_, new_n55994_, new_n55995_,
    new_n55996_, new_n55997_, new_n55998_, new_n55999_, new_n56000_,
    new_n56001_, new_n56002_, new_n56003_, new_n56004_, new_n56005_,
    new_n56006_, new_n56007_, new_n56008_, new_n56009_, new_n56010_,
    new_n56011_, new_n56012_, new_n56013_, new_n56014_, new_n56015_,
    new_n56016_, new_n56017_, new_n56018_, new_n56019_, new_n56020_,
    new_n56021_, new_n56022_, new_n56023_, new_n56024_, new_n56025_,
    new_n56026_, new_n56027_, new_n56028_, new_n56029_, new_n56030_,
    new_n56031_, new_n56032_, new_n56033_, new_n56034_, new_n56035_,
    new_n56036_, new_n56037_, new_n56038_, new_n56039_, new_n56040_,
    new_n56041_, new_n56042_, new_n56043_, new_n56044_, new_n56045_,
    new_n56046_, new_n56047_, new_n56048_, new_n56049_, new_n56050_,
    new_n56051_, new_n56052_, new_n56053_, new_n56054_, new_n56055_,
    new_n56056_, new_n56057_, new_n56058_, new_n56059_, new_n56060_,
    new_n56061_, new_n56062_, new_n56063_, new_n56064_, new_n56065_,
    new_n56066_, new_n56067_, new_n56068_, new_n56069_, new_n56070_,
    new_n56071_, new_n56072_, new_n56073_, new_n56074_, new_n56075_,
    new_n56076_, new_n56077_, new_n56078_, new_n56079_, new_n56080_,
    new_n56081_, new_n56082_, new_n56083_, new_n56084_, new_n56085_,
    new_n56086_, new_n56087_, new_n56088_, new_n56089_, new_n56090_,
    new_n56091_, new_n56092_, new_n56093_, new_n56094_, new_n56095_,
    new_n56096_, new_n56097_, new_n56098_, new_n56099_, new_n56100_,
    new_n56101_, new_n56102_, new_n56103_, new_n56104_, new_n56105_,
    new_n56106_, new_n56107_, new_n56108_, new_n56109_, new_n56110_,
    new_n56111_, new_n56112_, new_n56113_, new_n56114_, new_n56115_,
    new_n56116_, new_n56117_, new_n56118_, new_n56119_, new_n56120_,
    new_n56121_, new_n56122_, new_n56123_, new_n56124_, new_n56125_,
    new_n56126_, new_n56127_, new_n56128_, new_n56129_, new_n56130_,
    new_n56131_, new_n56132_, new_n56133_, new_n56134_, new_n56135_,
    new_n56136_, new_n56137_, new_n56138_, new_n56139_, new_n56140_,
    new_n56141_, new_n56142_, new_n56143_, new_n56144_, new_n56145_,
    new_n56146_, new_n56147_, new_n56148_, new_n56149_, new_n56150_,
    new_n56151_, new_n56152_, new_n56153_, new_n56154_, new_n56155_,
    new_n56156_, new_n56157_, new_n56158_, new_n56159_, new_n56160_,
    new_n56161_, new_n56162_, new_n56163_, new_n56164_, new_n56165_,
    new_n56166_, new_n56167_, new_n56168_, new_n56169_, new_n56170_,
    new_n56171_, new_n56172_, new_n56173_, new_n56174_, new_n56175_,
    new_n56176_, new_n56177_, new_n56178_, new_n56179_, new_n56180_,
    new_n56181_, new_n56182_, new_n56183_, new_n56184_, new_n56185_,
    new_n56186_, new_n56187_, new_n56188_, new_n56189_, new_n56190_,
    new_n56191_, new_n56192_, new_n56193_, new_n56194_, new_n56195_,
    new_n56196_, new_n56197_, new_n56198_, new_n56199_, new_n56200_,
    new_n56201_, new_n56202_, new_n56203_, new_n56204_, new_n56205_,
    new_n56206_, new_n56207_, new_n56208_, new_n56209_, new_n56210_,
    new_n56211_, new_n56212_, new_n56213_, new_n56214_, new_n56215_,
    new_n56216_, new_n56217_, new_n56218_, new_n56219_, new_n56220_,
    new_n56221_, new_n56222_, new_n56223_, new_n56224_, new_n56225_,
    new_n56226_, new_n56227_, new_n56228_, new_n56229_, new_n56230_,
    new_n56231_, new_n56232_, new_n56233_, new_n56234_, new_n56235_,
    new_n56236_, new_n56237_, new_n56238_, new_n56239_, new_n56240_,
    new_n56241_, new_n56242_, new_n56243_, new_n56244_, new_n56245_,
    new_n56246_, new_n56247_, new_n56248_, new_n56249_, new_n56250_,
    new_n56251_, new_n56252_, new_n56253_, new_n56254_, new_n56255_,
    new_n56256_, new_n56257_, new_n56258_, new_n56259_, new_n56260_,
    new_n56261_, new_n56262_, new_n56263_, new_n56264_, new_n56265_,
    new_n56266_, new_n56267_, new_n56268_, new_n56269_, new_n56270_,
    new_n56271_, new_n56272_, new_n56273_, new_n56274_, new_n56275_,
    new_n56276_, new_n56277_, new_n56278_, new_n56279_, new_n56280_,
    new_n56281_, new_n56282_, new_n56283_, new_n56284_, new_n56285_,
    new_n56286_, new_n56287_, new_n56288_, new_n56289_, new_n56290_,
    new_n56291_, new_n56292_, new_n56293_, new_n56294_, new_n56295_,
    new_n56296_, new_n56297_, new_n56298_, new_n56299_, new_n56300_,
    new_n56301_, new_n56302_, new_n56303_, new_n56304_, new_n56305_,
    new_n56306_, new_n56307_, new_n56308_, new_n56309_, new_n56310_,
    new_n56311_, new_n56312_, new_n56313_, new_n56314_, new_n56315_,
    new_n56316_, new_n56317_, new_n56318_, new_n56319_, new_n56320_,
    new_n56321_, new_n56322_, new_n56323_, new_n56324_, new_n56325_,
    new_n56326_, new_n56327_, new_n56328_, new_n56329_, new_n56330_,
    new_n56331_, new_n56332_, new_n56333_, new_n56334_, new_n56335_,
    new_n56336_, new_n56337_, new_n56338_, new_n56339_, new_n56340_,
    new_n56341_, new_n56342_, new_n56343_, new_n56344_, new_n56345_,
    new_n56346_, new_n56347_, new_n56348_, new_n56349_, new_n56350_,
    new_n56351_, new_n56352_, new_n56353_, new_n56354_, new_n56355_,
    new_n56356_, new_n56357_, new_n56358_, new_n56359_, new_n56360_,
    new_n56361_, new_n56362_, new_n56363_, new_n56364_, new_n56365_,
    new_n56366_, new_n56367_, new_n56368_, new_n56369_, new_n56370_,
    new_n56371_, new_n56372_, new_n56373_, new_n56374_, new_n56375_,
    new_n56376_, new_n56377_, new_n56378_, new_n56379_, new_n56380_,
    new_n56381_, new_n56382_, new_n56383_, new_n56384_, new_n56385_,
    new_n56386_, new_n56387_, new_n56388_, new_n56389_, new_n56390_,
    new_n56391_, new_n56392_, new_n56393_, new_n56394_, new_n56395_,
    new_n56396_, new_n56397_, new_n56398_, new_n56399_, new_n56400_,
    new_n56401_, new_n56402_, new_n56403_, new_n56404_, new_n56405_,
    new_n56406_, new_n56407_, new_n56408_, new_n56409_, new_n56410_,
    new_n56411_, new_n56412_, new_n56413_, new_n56414_, new_n56415_,
    new_n56416_, new_n56417_, new_n56418_, new_n56419_, new_n56420_,
    new_n56421_, new_n56422_, new_n56423_, new_n56424_, new_n56425_,
    new_n56426_, new_n56427_, new_n56428_, new_n56429_, new_n56430_,
    new_n56431_, new_n56432_, new_n56433_, new_n56434_, new_n56435_,
    new_n56436_, new_n56437_, new_n56438_, new_n56439_, new_n56440_,
    new_n56441_, new_n56442_, new_n56443_, new_n56444_, new_n56445_,
    new_n56446_, new_n56447_, new_n56448_, new_n56449_, new_n56450_,
    new_n56451_, new_n56452_, new_n56453_, new_n56454_, new_n56455_,
    new_n56456_, new_n56457_, new_n56458_, new_n56459_, new_n56460_,
    new_n56461_, new_n56462_, new_n56463_, new_n56464_, new_n56465_,
    new_n56466_, new_n56467_, new_n56468_, new_n56469_, new_n56470_,
    new_n56471_, new_n56472_, new_n56473_, new_n56474_, new_n56475_,
    new_n56476_, new_n56477_, new_n56478_, new_n56479_, new_n56480_,
    new_n56481_, new_n56482_, new_n56483_, new_n56484_, new_n56485_,
    new_n56486_, new_n56487_, new_n56488_, new_n56489_, new_n56490_,
    new_n56491_, new_n56492_, new_n56493_, new_n56494_, new_n56495_,
    new_n56496_, new_n56497_, new_n56498_, new_n56499_, new_n56500_,
    new_n56501_, new_n56502_, new_n56503_, new_n56504_, new_n56505_,
    new_n56506_, new_n56507_, new_n56508_, new_n56509_, new_n56510_,
    new_n56511_, new_n56512_, new_n56513_, new_n56514_, new_n56515_,
    new_n56516_, new_n56517_, new_n56518_, new_n56519_, new_n56520_,
    new_n56521_, new_n56522_, new_n56523_, new_n56524_, new_n56525_,
    new_n56526_, new_n56527_, new_n56528_, new_n56529_, new_n56530_,
    new_n56531_, new_n56532_, new_n56533_, new_n56534_, new_n56535_,
    new_n56536_, new_n56537_, new_n56538_, new_n56539_, new_n56540_,
    new_n56541_, new_n56542_, new_n56543_, new_n56544_, new_n56545_,
    new_n56546_, new_n56547_, new_n56548_, new_n56549_, new_n56550_,
    new_n56551_, new_n56552_, new_n56553_, new_n56554_, new_n56555_,
    new_n56556_, new_n56557_, new_n56558_, new_n56559_, new_n56560_,
    new_n56561_, new_n56562_, new_n56563_, new_n56564_, new_n56565_,
    new_n56566_, new_n56567_, new_n56568_, new_n56569_, new_n56570_,
    new_n56571_, new_n56572_, new_n56573_, new_n56574_, new_n56575_,
    new_n56576_, new_n56577_, new_n56578_, new_n56579_, new_n56580_,
    new_n56581_, new_n56582_, new_n56583_, new_n56584_, new_n56585_,
    new_n56586_, new_n56587_, new_n56588_, new_n56589_, new_n56590_,
    new_n56591_, new_n56592_, new_n56593_, new_n56594_, new_n56595_,
    new_n56596_, new_n56597_, new_n56598_, new_n56599_, new_n56600_,
    new_n56601_, new_n56602_, new_n56603_, new_n56604_, new_n56605_,
    new_n56606_, new_n56607_, new_n56608_, new_n56609_, new_n56610_,
    new_n56611_, new_n56612_, new_n56613_, new_n56614_, new_n56615_,
    new_n56616_, new_n56617_, new_n56618_, new_n56619_, new_n56620_,
    new_n56621_, new_n56622_, new_n56623_, new_n56624_, new_n56625_,
    new_n56626_, new_n56627_, new_n56628_, new_n56629_, new_n56630_,
    new_n56631_, new_n56632_, new_n56633_, new_n56634_, new_n56635_,
    new_n56636_, new_n56637_, new_n56638_, new_n56639_, new_n56640_,
    new_n56641_, new_n56642_, new_n56643_, new_n56644_, new_n56645_,
    new_n56646_, new_n56647_, new_n56648_, new_n56649_, new_n56650_,
    new_n56651_, new_n56652_, new_n56653_, new_n56654_, new_n56655_,
    new_n56656_, new_n56657_, new_n56658_, new_n56659_, new_n56660_,
    new_n56661_, new_n56662_, new_n56663_, new_n56664_, new_n56665_,
    new_n56666_, new_n56667_, new_n56668_, new_n56669_, new_n56670_,
    new_n56671_, new_n56672_, new_n56673_, new_n56674_, new_n56675_,
    new_n56676_, new_n56677_, new_n56678_, new_n56679_, new_n56680_,
    new_n56681_, new_n56682_, new_n56683_, new_n56684_, new_n56685_,
    new_n56686_, new_n56687_, new_n56688_, new_n56689_, new_n56690_,
    new_n56691_, new_n56692_, new_n56693_, new_n56694_, new_n56695_,
    new_n56696_, new_n56697_, new_n56698_, new_n56699_, new_n56700_,
    new_n56701_, new_n56702_, new_n56703_, new_n56704_, new_n56705_,
    new_n56706_, new_n56707_, new_n56708_, new_n56709_, new_n56710_,
    new_n56711_, new_n56712_, new_n56713_, new_n56714_, new_n56715_,
    new_n56716_, new_n56717_, new_n56718_, new_n56719_, new_n56720_,
    new_n56721_, new_n56722_, new_n56723_, new_n56724_, new_n56725_,
    new_n56726_, new_n56727_, new_n56728_, new_n56729_, new_n56730_,
    new_n56731_, new_n56732_, new_n56733_, new_n56734_, new_n56735_,
    new_n56736_, new_n56737_, new_n56738_, new_n56739_, new_n56740_,
    new_n56741_, new_n56742_, new_n56743_, new_n56744_, new_n56745_,
    new_n56746_, new_n56747_, new_n56748_, new_n56749_, new_n56750_,
    new_n56751_, new_n56752_, new_n56753_, new_n56754_, new_n56755_,
    new_n56756_, new_n56757_, new_n56758_, new_n56759_, new_n56760_,
    new_n56761_, new_n56762_, new_n56763_, new_n56764_, new_n56765_,
    new_n56766_, new_n56767_, new_n56768_, new_n56769_, new_n56770_,
    new_n56771_, new_n56772_, new_n56773_, new_n56774_, new_n56775_,
    new_n56776_, new_n56777_, new_n56778_, new_n56779_, new_n56780_,
    new_n56781_, new_n56782_, new_n56783_, new_n56784_, new_n56785_,
    new_n56786_, new_n56787_, new_n56788_, new_n56789_, new_n56790_,
    new_n56791_, new_n56792_, new_n56793_, new_n56794_, new_n56795_,
    new_n56796_, new_n56797_, new_n56798_, new_n56799_, new_n56800_,
    new_n56801_, new_n56802_, new_n56803_, new_n56804_, new_n56805_,
    new_n56806_, new_n56807_, new_n56808_, new_n56809_, new_n56810_,
    new_n56811_, new_n56812_, new_n56813_, new_n56814_, new_n56815_,
    new_n56816_, new_n56817_, new_n56818_, new_n56819_, new_n56820_,
    new_n56821_, new_n56822_, new_n56823_, new_n56824_, new_n56825_,
    new_n56826_, new_n56827_, new_n56828_, new_n56829_, new_n56830_,
    new_n56831_, new_n56832_, new_n56833_, new_n56834_, new_n56835_,
    new_n56836_, new_n56837_, new_n56838_, new_n56839_, new_n56840_,
    new_n56841_, new_n56842_, new_n56843_, new_n56844_, new_n56845_,
    new_n56846_, new_n56847_, new_n56848_, new_n56849_, new_n56850_,
    new_n56851_, new_n56852_, new_n56853_, new_n56854_, new_n56855_,
    new_n56856_, new_n56857_, new_n56858_, new_n56859_, new_n56860_,
    new_n56861_, new_n56862_, new_n56863_, new_n56864_, new_n56865_,
    new_n56866_, new_n56867_, new_n56868_, new_n56869_, new_n56870_,
    new_n56871_, new_n56872_, new_n56873_, new_n56874_, new_n56875_,
    new_n56876_, new_n56877_, new_n56878_, new_n56879_, new_n56880_,
    new_n56881_, new_n56882_, new_n56883_, new_n56884_, new_n56885_,
    new_n56886_, new_n56887_, new_n56888_, new_n56889_, new_n56890_,
    new_n56891_, new_n56892_, new_n56893_, new_n56894_, new_n56895_,
    new_n56896_, new_n56897_, new_n56898_, new_n56899_, new_n56900_,
    new_n56901_, new_n56902_, new_n56903_, new_n56904_, new_n56905_,
    new_n56906_, new_n56907_, new_n56908_, new_n56909_, new_n56910_,
    new_n56911_, new_n56912_, new_n56913_, new_n56914_, new_n56915_,
    new_n56916_, new_n56917_, new_n56918_, new_n56919_, new_n56920_,
    new_n56921_, new_n56922_, new_n56923_, new_n56924_, new_n56925_,
    new_n56926_, new_n56927_, new_n56928_, new_n56929_, new_n56930_,
    new_n56931_, new_n56932_, new_n56933_, new_n56934_, new_n56935_,
    new_n56936_, new_n56937_, new_n56938_, new_n56939_, new_n56940_,
    new_n56941_, new_n56942_, new_n56943_, new_n56944_, new_n56945_,
    new_n56946_, new_n56947_, new_n56948_, new_n56949_, new_n56950_,
    new_n56951_, new_n56952_, new_n56953_, new_n56954_, new_n56955_,
    new_n56956_, new_n56957_, new_n56958_, new_n56959_, new_n56960_,
    new_n56961_, new_n56962_, new_n56963_, new_n56964_, new_n56965_,
    new_n56966_, new_n56967_, new_n56968_, new_n56969_, new_n56970_,
    new_n56971_, new_n56972_, new_n56973_, new_n56974_, new_n56975_,
    new_n56976_, new_n56977_, new_n56978_, new_n56979_, new_n56980_,
    new_n56981_, new_n56982_, new_n56983_, new_n56984_, new_n56985_,
    new_n56986_, new_n56987_, new_n56988_, new_n56989_, new_n56990_,
    new_n56991_, new_n56992_, new_n56993_, new_n56994_, new_n56995_,
    new_n56996_, new_n56997_, new_n56998_, new_n56999_, new_n57000_,
    new_n57001_, new_n57002_, new_n57003_, new_n57004_, new_n57005_,
    new_n57006_, new_n57007_, new_n57008_, new_n57009_, new_n57010_,
    new_n57011_, new_n57012_, new_n57013_, new_n57014_, new_n57015_,
    new_n57016_, new_n57017_, new_n57018_, new_n57019_, new_n57020_,
    new_n57021_, new_n57022_, new_n57023_, new_n57024_, new_n57025_,
    new_n57026_, new_n57027_, new_n57028_, new_n57029_, new_n57030_,
    new_n57031_, new_n57032_, new_n57033_, new_n57034_, new_n57035_,
    new_n57036_, new_n57037_, new_n57038_, new_n57039_, new_n57040_,
    new_n57041_, new_n57042_, new_n57043_, new_n57044_, new_n57045_,
    new_n57046_, new_n57047_, new_n57048_, new_n57049_, new_n57050_,
    new_n57051_, new_n57052_, new_n57053_, new_n57054_, new_n57055_,
    new_n57056_, new_n57057_, new_n57058_, new_n57059_, new_n57060_,
    new_n57061_, new_n57062_, new_n57063_, new_n57064_, new_n57065_,
    new_n57066_, new_n57067_, new_n57068_, new_n57069_, new_n57070_,
    new_n57071_, new_n57072_, new_n57073_, new_n57074_, new_n57075_,
    new_n57076_, new_n57077_, new_n57078_, new_n57079_, new_n57080_,
    new_n57081_, new_n57082_, new_n57083_, new_n57084_, new_n57085_,
    new_n57086_, new_n57087_, new_n57088_, new_n57089_, new_n57090_,
    new_n57091_, new_n57092_, new_n57093_, new_n57094_, new_n57095_,
    new_n57096_, new_n57097_, new_n57098_, new_n57099_, new_n57100_,
    new_n57101_, new_n57102_, new_n57103_, new_n57104_, new_n57105_,
    new_n57106_, new_n57107_, new_n57108_, new_n57109_, new_n57110_,
    new_n57111_, new_n57112_, new_n57113_, new_n57114_, new_n57115_,
    new_n57116_, new_n57117_, new_n57118_, new_n57119_, new_n57120_,
    new_n57121_, new_n57122_, new_n57123_, new_n57124_, new_n57125_,
    new_n57126_, new_n57127_, new_n57128_, new_n57129_, new_n57130_,
    new_n57131_, new_n57132_, new_n57133_, new_n57134_, new_n57135_,
    new_n57136_, new_n57137_, new_n57138_, new_n57139_, new_n57140_,
    new_n57141_, new_n57142_, new_n57143_, new_n57144_, new_n57145_,
    new_n57146_, new_n57147_, new_n57148_, new_n57149_, new_n57150_,
    new_n57151_, new_n57152_, new_n57153_, new_n57154_, new_n57155_,
    new_n57156_, new_n57157_, new_n57158_, new_n57159_, new_n57160_,
    new_n57161_, new_n57162_, new_n57163_, new_n57164_, new_n57165_,
    new_n57166_, new_n57167_, new_n57168_, new_n57169_, new_n57170_,
    new_n57171_, new_n57172_, new_n57173_, new_n57174_, new_n57175_,
    new_n57176_, new_n57177_, new_n57178_, new_n57179_, new_n57180_,
    new_n57181_, new_n57182_, new_n57183_, new_n57184_, new_n57185_,
    new_n57186_, new_n57187_, new_n57188_, new_n57189_, new_n57190_,
    new_n57191_, new_n57192_, new_n57193_, new_n57194_, new_n57195_,
    new_n57196_, new_n57197_, new_n57198_, new_n57199_, new_n57200_,
    new_n57201_, new_n57202_, new_n57203_, new_n57204_, new_n57205_,
    new_n57206_, new_n57207_, new_n57208_, new_n57209_, new_n57210_,
    new_n57211_, new_n57212_, new_n57213_, new_n57214_, new_n57215_,
    new_n57216_, new_n57217_, new_n57218_, new_n57219_, new_n57220_,
    new_n57221_, new_n57222_, new_n57223_, new_n57224_, new_n57225_,
    new_n57226_, new_n57227_, new_n57228_, new_n57229_, new_n57230_,
    new_n57231_, new_n57232_, new_n57233_, new_n57234_, new_n57235_,
    new_n57236_, new_n57237_, new_n57238_, new_n57239_, new_n57240_,
    new_n57241_, new_n57242_, new_n57243_, new_n57244_, new_n57245_,
    new_n57246_, new_n57247_, new_n57248_, new_n57249_, new_n57250_,
    new_n57251_, new_n57252_, new_n57253_, new_n57254_, new_n57255_,
    new_n57256_, new_n57257_, new_n57258_, new_n57259_, new_n57260_,
    new_n57261_, new_n57262_, new_n57263_, new_n57264_, new_n57265_,
    new_n57266_, new_n57267_, new_n57268_, new_n57269_, new_n57270_,
    new_n57271_, new_n57272_, new_n57273_, new_n57274_, new_n57275_,
    new_n57276_, new_n57277_, new_n57278_, new_n57279_, new_n57280_,
    new_n57281_, new_n57282_, new_n57283_, new_n57284_, new_n57285_,
    new_n57286_, new_n57287_, new_n57288_, new_n57289_, new_n57290_,
    new_n57291_, new_n57292_, new_n57293_, new_n57294_, new_n57295_,
    new_n57296_, new_n57297_, new_n57298_, new_n57299_, new_n57300_,
    new_n57301_, new_n57302_, new_n57303_, new_n57304_, new_n57305_,
    new_n57306_, new_n57307_, new_n57308_, new_n57309_, new_n57310_,
    new_n57311_, new_n57312_, new_n57313_, new_n57314_, new_n57315_,
    new_n57316_, new_n57317_, new_n57318_, new_n57319_, new_n57320_,
    new_n57321_, new_n57322_, new_n57323_, new_n57324_, new_n57325_,
    new_n57326_, new_n57327_, new_n57328_, new_n57329_, new_n57330_,
    new_n57331_, new_n57332_, new_n57333_, new_n57334_, new_n57335_,
    new_n57336_, new_n57337_, new_n57338_, new_n57339_, new_n57340_,
    new_n57341_, new_n57342_, new_n57343_, new_n57344_, new_n57345_,
    new_n57346_, new_n57347_, new_n57348_, new_n57349_, new_n57350_,
    new_n57351_, new_n57352_, new_n57353_, new_n57354_, new_n57355_,
    new_n57356_, new_n57357_, new_n57358_, new_n57359_, new_n57360_,
    new_n57361_, new_n57362_, new_n57363_, new_n57364_, new_n57365_,
    new_n57366_, new_n57367_, new_n57368_, new_n57369_, new_n57370_,
    new_n57371_, new_n57372_, new_n57373_, new_n57374_, new_n57375_,
    new_n57376_, new_n57377_, new_n57378_, new_n57379_, new_n57380_,
    new_n57381_, new_n57382_, new_n57383_, new_n57384_, new_n57385_,
    new_n57386_, new_n57387_, new_n57388_, new_n57389_, new_n57390_,
    new_n57391_, new_n57392_, new_n57393_, new_n57394_, new_n57395_,
    new_n57396_, new_n57397_, new_n57398_, new_n57399_, new_n57400_,
    new_n57401_, new_n57402_, new_n57403_, new_n57404_, new_n57405_,
    new_n57406_, new_n57407_, new_n57408_, new_n57409_, new_n57410_,
    new_n57411_, new_n57412_, new_n57413_, new_n57414_, new_n57415_,
    new_n57416_, new_n57417_, new_n57418_, new_n57419_, new_n57420_,
    new_n57421_, new_n57422_, new_n57423_, new_n57424_, new_n57425_,
    new_n57426_, new_n57427_, new_n57428_, new_n57429_, new_n57430_,
    new_n57431_, new_n57432_, new_n57433_, new_n57434_, new_n57435_,
    new_n57436_, new_n57437_, new_n57438_, new_n57439_, new_n57440_,
    new_n57441_, new_n57442_, new_n57443_, new_n57444_, new_n57445_,
    new_n57446_, new_n57447_, new_n57448_, new_n57449_, new_n57450_,
    new_n57451_, new_n57452_, new_n57453_, new_n57454_, new_n57455_,
    new_n57456_, new_n57457_, new_n57458_, new_n57459_, new_n57460_,
    new_n57461_, new_n57462_, new_n57463_, new_n57464_, new_n57465_,
    new_n57466_, new_n57467_, new_n57468_, new_n57469_, new_n57470_,
    new_n57471_, new_n57472_, new_n57473_, new_n57474_, new_n57475_,
    new_n57476_, new_n57477_, new_n57478_, new_n57479_, new_n57480_,
    new_n57481_, new_n57482_, new_n57483_, new_n57484_, new_n57485_,
    new_n57486_, new_n57487_, new_n57488_, new_n57489_, new_n57490_,
    new_n57491_, new_n57492_, new_n57493_, new_n57494_, new_n57495_,
    new_n57496_, new_n57497_, new_n57498_, new_n57499_, new_n57500_,
    new_n57501_, new_n57502_, new_n57503_, new_n57504_, new_n57505_,
    new_n57506_, new_n57507_, new_n57508_, new_n57509_, new_n57510_,
    new_n57511_, new_n57512_, new_n57513_, new_n57514_, new_n57515_,
    new_n57516_, new_n57517_, new_n57518_, new_n57519_, new_n57520_,
    new_n57521_, new_n57522_, new_n57523_, new_n57524_, new_n57525_,
    new_n57526_, new_n57527_, new_n57528_, new_n57529_, new_n57530_,
    new_n57531_, new_n57532_, new_n57533_, new_n57534_, new_n57535_,
    new_n57536_, new_n57537_, new_n57538_, new_n57539_, new_n57540_,
    new_n57541_, new_n57542_, new_n57543_, new_n57544_, new_n57545_,
    new_n57546_, new_n57547_, new_n57548_, new_n57549_, new_n57550_,
    new_n57551_, new_n57552_, new_n57553_, new_n57554_, new_n57555_,
    new_n57556_, new_n57557_, new_n57558_, new_n57559_, new_n57560_,
    new_n57561_, new_n57562_, new_n57563_, new_n57564_, new_n57565_,
    new_n57566_, new_n57567_, new_n57568_, new_n57569_, new_n57570_,
    new_n57571_, new_n57572_, new_n57573_, new_n57574_, new_n57575_,
    new_n57576_, new_n57577_, new_n57578_, new_n57579_, new_n57580_,
    new_n57581_, new_n57582_, new_n57583_, new_n57584_, new_n57585_,
    new_n57586_, new_n57587_, new_n57588_, new_n57589_, new_n57590_,
    new_n57591_, new_n57592_, new_n57593_, new_n57594_, new_n57595_,
    new_n57596_, new_n57597_, new_n57598_, new_n57599_, new_n57600_,
    new_n57601_, new_n57602_, new_n57603_, new_n57604_, new_n57605_,
    new_n57606_, new_n57607_, new_n57608_, new_n57609_, new_n57610_,
    new_n57611_, new_n57612_, new_n57613_, new_n57614_, new_n57615_,
    new_n57616_, new_n57617_, new_n57618_, new_n57619_, new_n57620_,
    new_n57621_, new_n57622_, new_n57623_, new_n57624_, new_n57625_,
    new_n57626_, new_n57627_, new_n57628_, new_n57629_, new_n57630_,
    new_n57631_, new_n57632_, new_n57633_, new_n57634_, new_n57635_,
    new_n57636_, new_n57637_, new_n57638_, new_n57639_, new_n57640_,
    new_n57641_, new_n57642_, new_n57643_, new_n57644_, new_n57645_,
    new_n57646_, new_n57647_, new_n57648_, new_n57649_, new_n57650_,
    new_n57651_, new_n57652_, new_n57653_, new_n57654_, new_n57655_,
    new_n57656_, new_n57657_, new_n57658_, new_n57659_, new_n57660_,
    new_n57661_, new_n57662_, new_n57663_, new_n57664_, new_n57665_,
    new_n57666_, new_n57667_, new_n57668_, new_n57669_, new_n57670_,
    new_n57671_, new_n57672_, new_n57673_, new_n57674_, new_n57675_,
    new_n57676_, new_n57677_, new_n57678_, new_n57679_, new_n57680_,
    new_n57681_, new_n57682_, new_n57683_, new_n57684_, new_n57685_,
    new_n57686_, new_n57687_, new_n57688_, new_n57689_, new_n57690_,
    new_n57691_, new_n57692_, new_n57693_, new_n57694_, new_n57695_,
    new_n57696_, new_n57697_, new_n57698_, new_n57699_, new_n57700_,
    new_n57701_, new_n57702_, new_n57703_, new_n57704_, new_n57705_,
    new_n57706_, new_n57707_, new_n57708_, new_n57709_, new_n57710_,
    new_n57711_, new_n57712_, new_n57713_, new_n57714_, new_n57715_,
    new_n57716_, new_n57717_, new_n57718_, new_n57719_, new_n57720_,
    new_n57721_, new_n57722_, new_n57723_, new_n57724_, new_n57725_,
    new_n57726_, new_n57727_, new_n57728_, new_n57729_, new_n57730_,
    new_n57731_, new_n57732_, new_n57733_, new_n57734_, new_n57735_,
    new_n57736_, new_n57737_, new_n57738_, new_n57739_, new_n57740_,
    new_n57741_, new_n57742_, new_n57743_, new_n57744_, new_n57745_,
    new_n57746_, new_n57747_, new_n57748_, new_n57749_, new_n57750_,
    new_n57751_, new_n57752_, new_n57753_, new_n57754_, new_n57755_,
    new_n57756_, new_n57757_, new_n57758_, new_n57759_, new_n57760_,
    new_n57761_, new_n57762_, new_n57763_, new_n57764_, new_n57765_,
    new_n57766_, new_n57767_, new_n57768_, new_n57769_, new_n57770_,
    new_n57771_, new_n57772_, new_n57773_, new_n57774_, new_n57775_,
    new_n57776_, new_n57777_, new_n57778_, new_n57779_, new_n57780_,
    new_n57781_, new_n57782_, new_n57783_, new_n57784_, new_n57785_,
    new_n57786_, new_n57787_, new_n57788_, new_n57789_, new_n57790_,
    new_n57791_, new_n57792_, new_n57793_, new_n57794_, new_n57795_,
    new_n57796_, new_n57797_, new_n57798_, new_n57799_, new_n57800_,
    new_n57801_, new_n57802_, new_n57803_, new_n57804_, new_n57805_,
    new_n57806_, new_n57807_, new_n57808_, new_n57809_, new_n57810_,
    new_n57811_, new_n57812_, new_n57813_, new_n57814_, new_n57815_,
    new_n57816_, new_n57817_, new_n57818_, new_n57819_, new_n57820_,
    new_n57821_, new_n57822_, new_n57823_, new_n57824_, new_n57825_,
    new_n57826_, new_n57827_, new_n57828_, new_n57829_, new_n57830_,
    new_n57831_, new_n57832_, new_n57833_, new_n57834_, new_n57835_,
    new_n57836_, new_n57837_, new_n57838_, new_n57839_, new_n57840_,
    new_n57841_, new_n57842_, new_n57843_, new_n57844_, new_n57845_,
    new_n57846_, new_n57847_, new_n57848_, new_n57849_, new_n57850_,
    new_n57851_, new_n57852_, new_n57853_, new_n57854_, new_n57855_,
    new_n57856_, new_n57857_, new_n57858_, new_n57859_, new_n57860_,
    new_n57861_, new_n57862_, new_n57863_, new_n57864_, new_n57865_,
    new_n57866_, new_n57867_, new_n57868_, new_n57869_, new_n57870_,
    new_n57871_, new_n57872_, new_n57873_, new_n57874_, new_n57875_,
    new_n57876_, new_n57877_, new_n57878_, new_n57879_, new_n57880_,
    new_n57881_, new_n57882_, new_n57883_, new_n57884_, new_n57885_,
    new_n57886_, new_n57887_, new_n57888_, new_n57889_, new_n57890_,
    new_n57891_, new_n57892_, new_n57893_, new_n57894_, new_n57895_,
    new_n57896_, new_n57897_, new_n57898_, new_n57899_, new_n57900_,
    new_n57901_, new_n57902_, new_n57903_, new_n57904_, new_n57905_,
    new_n57906_, new_n57907_, new_n57908_, new_n57909_, new_n57910_,
    new_n57911_, new_n57912_, new_n57913_, new_n57914_, new_n57915_,
    new_n57916_, new_n57917_, new_n57918_, new_n57919_, new_n57920_,
    new_n57921_, new_n57922_, new_n57923_, new_n57924_, new_n57925_,
    new_n57926_, new_n57927_, new_n57928_, new_n57929_, new_n57930_,
    new_n57931_, new_n57932_, new_n57933_, new_n57934_, new_n57935_,
    new_n57936_, new_n57937_, new_n57938_, new_n57939_, new_n57940_,
    new_n57941_, new_n57942_, new_n57943_, new_n57944_, new_n57945_,
    new_n57946_, new_n57947_, new_n57948_, new_n57949_, new_n57950_,
    new_n57951_, new_n57952_, new_n57953_, new_n57954_, new_n57955_,
    new_n57956_, new_n57957_, new_n57958_, new_n57959_, new_n57960_,
    new_n57961_, new_n57962_, new_n57963_, new_n57964_, new_n57965_,
    new_n57966_, new_n57967_, new_n57968_, new_n57969_, new_n57970_,
    new_n57971_, new_n57972_, new_n57973_, new_n57974_, new_n57975_,
    new_n57976_, new_n57977_, new_n57978_, new_n57979_, new_n57980_,
    new_n57981_, new_n57982_, new_n57983_, new_n57984_, new_n57985_,
    new_n57986_, new_n57987_, new_n57988_, new_n57989_, new_n57990_,
    new_n57991_, new_n57992_, new_n57993_, new_n57994_, new_n57995_,
    new_n57996_, new_n57997_, new_n57998_, new_n57999_, new_n58000_,
    new_n58001_, new_n58002_, new_n58003_, new_n58004_, new_n58005_,
    new_n58006_, new_n58007_, new_n58008_, new_n58009_, new_n58010_,
    new_n58011_, new_n58012_, new_n58013_, new_n58014_, new_n58015_,
    new_n58016_, new_n58017_, new_n58018_, new_n58019_, new_n58020_,
    new_n58021_, new_n58022_, new_n58023_, new_n58024_, new_n58025_,
    new_n58026_, new_n58027_, new_n58028_, new_n58029_, new_n58030_,
    new_n58031_, new_n58032_, new_n58033_, new_n58034_, new_n58035_,
    new_n58036_, new_n58037_, new_n58038_, new_n58039_, new_n58040_,
    new_n58041_, new_n58042_, new_n58043_, new_n58044_, new_n58045_,
    new_n58046_, new_n58047_, new_n58048_, new_n58049_, new_n58050_,
    new_n58051_, new_n58052_, new_n58053_, new_n58054_, new_n58055_,
    new_n58056_, new_n58057_, new_n58058_, new_n58059_, new_n58060_,
    new_n58061_, new_n58062_, new_n58063_, new_n58064_, new_n58065_,
    new_n58066_, new_n58067_, new_n58068_, new_n58069_, new_n58070_,
    new_n58071_, new_n58072_, new_n58073_, new_n58074_, new_n58075_,
    new_n58076_, new_n58077_, new_n58078_, new_n58079_, new_n58080_,
    new_n58081_, new_n58082_, new_n58083_, new_n58084_, new_n58085_,
    new_n58086_, new_n58087_, new_n58088_, new_n58089_, new_n58090_,
    new_n58091_, new_n58092_, new_n58093_, new_n58094_, new_n58095_,
    new_n58096_, new_n58097_, new_n58098_, new_n58099_, new_n58100_,
    new_n58101_, new_n58102_, new_n58103_, new_n58104_, new_n58105_,
    new_n58106_, new_n58107_, new_n58108_, new_n58109_, new_n58110_,
    new_n58111_, new_n58112_, new_n58113_, new_n58114_, new_n58115_,
    new_n58116_, new_n58117_, new_n58118_, new_n58119_, new_n58120_,
    new_n58121_, new_n58122_, new_n58123_, new_n58124_, new_n58125_,
    new_n58126_, new_n58127_, new_n58128_, new_n58129_, new_n58130_,
    new_n58131_, new_n58132_, new_n58133_, new_n58134_, new_n58135_,
    new_n58136_, new_n58137_, new_n58138_, new_n58139_, new_n58140_,
    new_n58141_, new_n58142_, new_n58143_, new_n58144_, new_n58145_,
    new_n58146_, new_n58147_, new_n58148_, new_n58149_, new_n58150_,
    new_n58151_, new_n58152_, new_n58153_, new_n58154_, new_n58155_,
    new_n58156_, new_n58157_, new_n58158_, new_n58159_, new_n58160_,
    new_n58161_, new_n58162_, new_n58163_, new_n58164_, new_n58165_,
    new_n58166_, new_n58167_, new_n58168_, new_n58169_, new_n58170_,
    new_n58171_, new_n58172_, new_n58173_, new_n58174_, new_n58175_,
    new_n58176_, new_n58177_, new_n58178_, new_n58179_, new_n58180_,
    new_n58181_, new_n58182_, new_n58183_, new_n58184_, new_n58185_,
    new_n58186_, new_n58187_, new_n58188_, new_n58189_, new_n58190_,
    new_n58191_, new_n58192_, new_n58193_, new_n58194_, new_n58195_,
    new_n58196_, new_n58197_, new_n58198_, new_n58199_, new_n58200_,
    new_n58201_, new_n58202_, new_n58203_, new_n58204_, new_n58205_,
    new_n58206_, new_n58207_, new_n58208_, new_n58209_, new_n58210_,
    new_n58211_, new_n58212_, new_n58213_, new_n58214_, new_n58215_,
    new_n58216_, new_n58217_, new_n58218_, new_n58219_, new_n58220_,
    new_n58221_, new_n58222_, new_n58223_, new_n58224_, new_n58225_,
    new_n58226_, new_n58227_, new_n58228_, new_n58229_, new_n58230_,
    new_n58231_, new_n58232_, new_n58233_, new_n58234_, new_n58235_,
    new_n58236_, new_n58237_, new_n58238_, new_n58239_, new_n58240_,
    new_n58241_, new_n58242_, new_n58243_, new_n58244_, new_n58245_,
    new_n58246_, new_n58247_, new_n58248_, new_n58249_, new_n58250_,
    new_n58251_, new_n58252_, new_n58253_, new_n58254_, new_n58255_,
    new_n58256_, new_n58257_, new_n58258_, new_n58259_, new_n58260_,
    new_n58261_, new_n58262_, new_n58263_, new_n58264_, new_n58265_,
    new_n58266_, new_n58267_, new_n58268_, new_n58269_, new_n58270_,
    new_n58271_, new_n58272_, new_n58273_, new_n58274_, new_n58275_,
    new_n58276_, new_n58277_, new_n58278_, new_n58279_, new_n58280_,
    new_n58281_, new_n58282_, new_n58283_, new_n58284_, new_n58285_,
    new_n58286_, new_n58287_, new_n58288_, new_n58289_, new_n58290_,
    new_n58291_, new_n58292_, new_n58293_, new_n58294_, new_n58295_,
    new_n58296_, new_n58297_, new_n58298_, new_n58299_, new_n58300_,
    new_n58301_, new_n58302_, new_n58303_, new_n58304_, new_n58305_,
    new_n58306_, new_n58307_, new_n58308_, new_n58309_, new_n58310_,
    new_n58311_, new_n58312_, new_n58313_, new_n58314_, new_n58315_,
    new_n58316_, new_n58317_, new_n58318_, new_n58319_, new_n58320_,
    new_n58321_, new_n58322_, new_n58323_, new_n58324_, new_n58325_,
    new_n58326_, new_n58327_, new_n58328_, new_n58329_, new_n58330_,
    new_n58331_, new_n58332_, new_n58333_, new_n58334_, new_n58335_,
    new_n58336_, new_n58337_, new_n58338_, new_n58339_, new_n58340_,
    new_n58341_, new_n58342_, new_n58343_, new_n58344_, new_n58345_,
    new_n58346_, new_n58347_, new_n58348_, new_n58349_, new_n58350_,
    new_n58351_, new_n58352_, new_n58353_, new_n58354_, new_n58355_,
    new_n58356_, new_n58357_, new_n58358_, new_n58359_, new_n58360_,
    new_n58361_, new_n58362_, new_n58363_, new_n58364_, new_n58365_,
    new_n58366_, new_n58367_, new_n58368_, new_n58369_, new_n58370_,
    new_n58371_, new_n58372_, new_n58373_, new_n58374_, new_n58375_,
    new_n58376_, new_n58377_, new_n58378_, new_n58379_, new_n58380_,
    new_n58381_, new_n58382_, new_n58383_, new_n58384_, new_n58385_,
    new_n58386_, new_n58387_, new_n58388_, new_n58389_, new_n58390_,
    new_n58391_, new_n58392_, new_n58393_, new_n58394_, new_n58395_,
    new_n58396_, new_n58397_, new_n58398_, new_n58399_, new_n58400_,
    new_n58401_, new_n58402_, new_n58403_, new_n58404_, new_n58405_,
    new_n58406_, new_n58407_, new_n58408_, new_n58409_, new_n58410_,
    new_n58411_, new_n58412_, new_n58413_, new_n58414_, new_n58415_,
    new_n58416_, new_n58417_, new_n58418_, new_n58419_, new_n58420_,
    new_n58421_, new_n58422_, new_n58423_, new_n58424_, new_n58425_,
    new_n58426_, new_n58427_, new_n58428_, new_n58429_, new_n58430_,
    new_n58431_, new_n58432_, new_n58433_, new_n58434_, new_n58435_,
    new_n58436_, new_n58437_, new_n58438_, new_n58439_, new_n58440_,
    new_n58441_, new_n58442_, new_n58443_, new_n58444_, new_n58445_,
    new_n58446_, new_n58447_, new_n58448_, new_n58449_, new_n58450_,
    new_n58451_, new_n58452_, new_n58453_, new_n58454_, new_n58455_,
    new_n58456_, new_n58457_, new_n58458_, new_n58459_, new_n58460_,
    new_n58461_, new_n58462_, new_n58463_, new_n58464_, new_n58465_,
    new_n58466_, new_n58467_, new_n58468_, new_n58469_, new_n58470_,
    new_n58471_, new_n58472_, new_n58473_, new_n58474_, new_n58475_,
    new_n58476_, new_n58477_, new_n58478_, new_n58479_, new_n58480_,
    new_n58481_, new_n58482_, new_n58483_, new_n58484_, new_n58485_,
    new_n58486_, new_n58487_, new_n58488_, new_n58489_, new_n58490_,
    new_n58491_, new_n58492_, new_n58493_, new_n58494_, new_n58495_,
    new_n58496_, new_n58497_, new_n58498_, new_n58499_, new_n58500_,
    new_n58501_, new_n58502_, new_n58503_, new_n58504_, new_n58505_,
    new_n58506_, new_n58507_, new_n58508_, new_n58509_, new_n58510_,
    new_n58511_, new_n58512_, new_n58513_, new_n58514_, new_n58515_,
    new_n58516_, new_n58517_, new_n58518_, new_n58519_, new_n58520_,
    new_n58521_, new_n58522_, new_n58523_, new_n58524_, new_n58525_,
    new_n58526_, new_n58527_, new_n58528_, new_n58529_, new_n58530_,
    new_n58531_, new_n58532_, new_n58533_, new_n58534_, new_n58535_,
    new_n58536_, new_n58537_, new_n58538_, new_n58539_, new_n58540_,
    new_n58541_, new_n58542_, new_n58543_, new_n58544_, new_n58545_,
    new_n58546_, new_n58547_, new_n58548_, new_n58549_, new_n58550_,
    new_n58551_, new_n58552_, new_n58553_, new_n58554_, new_n58555_,
    new_n58556_, new_n58557_, new_n58558_, new_n58559_, new_n58560_,
    new_n58561_, new_n58562_, new_n58563_, new_n58564_, new_n58565_,
    new_n58566_, new_n58567_, new_n58568_, new_n58569_, new_n58570_,
    new_n58571_, new_n58572_, new_n58573_, new_n58574_, new_n58575_,
    new_n58576_, new_n58577_, new_n58578_, new_n58579_, new_n58580_,
    new_n58581_, new_n58582_, new_n58583_, new_n58584_, new_n58585_,
    new_n58586_, new_n58587_, new_n58588_, new_n58589_, new_n58590_,
    new_n58591_, new_n58592_, new_n58593_, new_n58594_, new_n58595_,
    new_n58596_, new_n58597_, new_n58598_, new_n58599_, new_n58600_,
    new_n58601_, new_n58602_, new_n58603_, new_n58604_, new_n58605_,
    new_n58606_, new_n58607_, new_n58608_, new_n58609_, new_n58610_,
    new_n58611_, new_n58612_, new_n58613_, new_n58614_, new_n58615_,
    new_n58616_, new_n58617_, new_n58618_, new_n58619_, new_n58620_,
    new_n58621_, new_n58622_, new_n58623_, new_n58624_, new_n58625_,
    new_n58626_, new_n58627_, new_n58628_, new_n58629_, new_n58630_,
    new_n58631_, new_n58632_, new_n58633_, new_n58634_, new_n58635_,
    new_n58636_, new_n58637_, new_n58638_, new_n58639_, new_n58640_,
    new_n58641_, new_n58642_, new_n58643_, new_n58644_, new_n58645_,
    new_n58646_, new_n58647_, new_n58648_, new_n58649_, new_n58650_,
    new_n58651_, new_n58652_, new_n58653_, new_n58654_, new_n58655_,
    new_n58656_, new_n58657_, new_n58658_, new_n58659_, new_n58660_,
    new_n58661_, new_n58662_, new_n58663_, new_n58664_, new_n58665_,
    new_n58666_, new_n58667_, new_n58668_, new_n58669_, new_n58670_,
    new_n58671_, new_n58672_, new_n58673_, new_n58674_, new_n58675_,
    new_n58676_, new_n58677_, new_n58678_, new_n58679_, new_n58680_,
    new_n58681_, new_n58682_, new_n58683_, new_n58684_, new_n58685_,
    new_n58686_, new_n58687_, new_n58688_, new_n58689_, new_n58690_,
    new_n58691_, new_n58692_, new_n58693_, new_n58694_, new_n58695_,
    new_n58696_, new_n58697_, new_n58698_, new_n58699_, new_n58700_,
    new_n58701_, new_n58702_, new_n58703_, new_n58704_, new_n58705_,
    new_n58706_, new_n58707_, new_n58708_, new_n58709_, new_n58710_,
    new_n58711_, new_n58712_, new_n58713_, new_n58714_, new_n58715_,
    new_n58716_, new_n58717_, new_n58718_, new_n58719_, new_n58720_,
    new_n58721_, new_n58722_, new_n58723_, new_n58724_, new_n58725_,
    new_n58726_, new_n58727_, new_n58728_, new_n58729_, new_n58730_,
    new_n58731_, new_n58732_, new_n58733_, new_n58734_, new_n58735_,
    new_n58736_, new_n58737_, new_n58738_, new_n58739_, new_n58740_,
    new_n58741_, new_n58742_, new_n58743_, new_n58744_, new_n58745_,
    new_n58746_, new_n58747_, new_n58748_, new_n58749_, new_n58750_,
    new_n58751_, new_n58752_, new_n58753_, new_n58754_, new_n58755_,
    new_n58756_, new_n58757_, new_n58758_, new_n58759_, new_n58760_,
    new_n58761_, new_n58762_, new_n58763_, new_n58764_, new_n58765_,
    new_n58766_, new_n58767_, new_n58768_, new_n58769_, new_n58770_,
    new_n58771_, new_n58772_, new_n58773_, new_n58774_, new_n58775_,
    new_n58776_, new_n58777_, new_n58778_, new_n58779_, new_n58780_,
    new_n58781_, new_n58782_, new_n58783_, new_n58784_, new_n58785_,
    new_n58786_, new_n58787_, new_n58788_, new_n58789_, new_n58790_,
    new_n58791_, new_n58792_, new_n58793_, new_n58794_, new_n58795_,
    new_n58796_, new_n58797_, new_n58798_, new_n58799_, new_n58800_,
    new_n58801_, new_n58802_, new_n58803_, new_n58804_, new_n58805_,
    new_n58806_, new_n58807_, new_n58808_, new_n58809_, new_n58810_,
    new_n58811_, new_n58812_, new_n58813_, new_n58814_, new_n58815_,
    new_n58816_, new_n58817_, new_n58818_, new_n58819_, new_n58820_,
    new_n58821_, new_n58822_, new_n58823_, new_n58824_, new_n58825_,
    new_n58826_, new_n58827_, new_n58828_, new_n58829_, new_n58830_,
    new_n58831_, new_n58832_, new_n58833_, new_n58834_, new_n58835_,
    new_n58836_, new_n58837_, new_n58838_, new_n58839_, new_n58840_,
    new_n58841_, new_n58842_, new_n58843_, new_n58844_, new_n58845_,
    new_n58846_, new_n58847_, new_n58848_, new_n58849_, new_n58850_,
    new_n58851_, new_n58852_, new_n58853_, new_n58854_, new_n58855_,
    new_n58856_, new_n58857_, new_n58858_, new_n58859_, new_n58860_,
    new_n58861_, new_n58862_, new_n58863_, new_n58864_, new_n58865_,
    new_n58866_, new_n58867_, new_n58868_, new_n58869_, new_n58870_,
    new_n58871_, new_n58872_, new_n58873_, new_n58874_, new_n58875_,
    new_n58876_, new_n58877_, new_n58878_, new_n58879_, new_n58880_,
    new_n58881_, new_n58882_, new_n58883_, new_n58884_, new_n58885_,
    new_n58886_, new_n58887_, new_n58888_, new_n58889_, new_n58890_,
    new_n58891_, new_n58892_, new_n58893_, new_n58894_, new_n58895_,
    new_n58896_, new_n58897_, new_n58898_, new_n58899_, new_n58900_,
    new_n58901_, new_n58902_, new_n58903_, new_n58904_, new_n58905_,
    new_n58906_, new_n58907_, new_n58908_, new_n58909_, new_n58910_,
    new_n58911_, new_n58912_, new_n58913_, new_n58914_, new_n58915_,
    new_n58916_, new_n58917_, new_n58918_, new_n58919_, new_n58920_,
    new_n58921_, new_n58922_, new_n58923_, new_n58924_, new_n58925_,
    new_n58926_, new_n58927_, new_n58928_, new_n58929_, new_n58930_,
    new_n58931_, new_n58932_, new_n58933_, new_n58934_, new_n58935_,
    new_n58936_, new_n58937_, new_n58938_, new_n58939_, new_n58940_,
    new_n58941_, new_n58942_, new_n58943_, new_n58944_, new_n58945_,
    new_n58946_, new_n58947_, new_n58948_, new_n58949_, new_n58950_,
    new_n58951_, new_n58952_, new_n58953_, new_n58954_, new_n58955_,
    new_n58956_, new_n58957_, new_n58958_, new_n58959_, new_n58960_,
    new_n58961_, new_n58962_, new_n58963_, new_n58964_, new_n58965_,
    new_n58966_, new_n58967_, new_n58968_, new_n58969_, new_n58970_,
    new_n58971_, new_n58972_, new_n58973_, new_n58974_, new_n58975_,
    new_n58976_, new_n58977_, new_n58978_, new_n58979_, new_n58980_,
    new_n58981_, new_n58982_, new_n58983_, new_n58984_, new_n58985_,
    new_n58986_, new_n58987_, new_n58988_, new_n58989_, new_n58990_,
    new_n58991_, new_n58992_, new_n58993_, new_n58994_, new_n58995_,
    new_n58996_, new_n58997_, new_n58998_, new_n58999_, new_n59000_,
    new_n59001_, new_n59002_, new_n59003_, new_n59004_, new_n59005_,
    new_n59006_, new_n59007_, new_n59008_, new_n59009_, new_n59010_,
    new_n59011_, new_n59012_, new_n59013_, new_n59014_, new_n59015_,
    new_n59016_, new_n59017_, new_n59018_, new_n59019_, new_n59020_,
    new_n59021_, new_n59022_, new_n59023_, new_n59024_, new_n59025_,
    new_n59026_, new_n59027_, new_n59028_, new_n59029_, new_n59030_,
    new_n59031_, new_n59032_, new_n59033_, new_n59034_, new_n59035_,
    new_n59036_, new_n59037_, new_n59038_, new_n59039_, new_n59040_,
    new_n59041_, new_n59042_, new_n59043_, new_n59044_, new_n59045_,
    new_n59046_, new_n59047_, new_n59048_, new_n59049_, new_n59050_,
    new_n59051_, new_n59052_, new_n59053_, new_n59054_, new_n59055_,
    new_n59056_, new_n59057_, new_n59058_, new_n59059_, new_n59060_,
    new_n59061_, new_n59062_, new_n59063_, new_n59064_, new_n59065_,
    new_n59066_, new_n59067_, new_n59068_, new_n59069_, new_n59070_,
    new_n59071_, new_n59072_, new_n59073_, new_n59074_, new_n59075_,
    new_n59076_, new_n59077_, new_n59078_, new_n59079_, new_n59080_,
    new_n59081_, new_n59082_, new_n59083_, new_n59084_, new_n59085_,
    new_n59086_, new_n59087_, new_n59088_, new_n59089_, new_n59090_,
    new_n59091_, new_n59092_, new_n59093_, new_n59094_, new_n59095_,
    new_n59096_, new_n59097_, new_n59098_, new_n59099_, new_n59100_,
    new_n59101_, new_n59102_, new_n59103_, new_n59104_, new_n59105_,
    new_n59106_, new_n59107_, new_n59108_, new_n59109_, new_n59110_,
    new_n59111_, new_n59112_, new_n59113_, new_n59114_, new_n59115_,
    new_n59116_, new_n59117_, new_n59118_, new_n59119_, new_n59120_,
    new_n59121_, new_n59122_, new_n59123_, new_n59124_, new_n59125_,
    new_n59126_, new_n59127_, new_n59128_, new_n59129_, new_n59130_,
    new_n59131_, new_n59132_, new_n59133_, new_n59134_, new_n59135_,
    new_n59136_, new_n59137_, new_n59138_, new_n59139_, new_n59140_,
    new_n59141_, new_n59142_, new_n59143_, new_n59144_, new_n59145_,
    new_n59146_, new_n59147_, new_n59148_, new_n59149_, new_n59150_,
    new_n59151_, new_n59152_, new_n59153_, new_n59154_, new_n59155_,
    new_n59156_, new_n59157_, new_n59158_, new_n59159_, new_n59160_,
    new_n59161_, new_n59162_, new_n59163_, new_n59164_, new_n59165_,
    new_n59166_, new_n59167_, new_n59168_, new_n59169_, new_n59170_,
    new_n59171_, new_n59172_, new_n59173_, new_n59174_, new_n59175_,
    new_n59176_, new_n59177_, new_n59178_, new_n59179_, new_n59180_,
    new_n59181_, new_n59182_, new_n59183_, new_n59184_, new_n59185_,
    new_n59186_, new_n59187_, new_n59188_, new_n59189_, new_n59190_,
    new_n59191_, new_n59192_, new_n59193_, new_n59194_, new_n59195_,
    new_n59196_, new_n59197_, new_n59198_, new_n59199_, new_n59200_,
    new_n59201_, new_n59202_, new_n59203_, new_n59204_, new_n59205_,
    new_n59206_, new_n59207_, new_n59208_, new_n59209_, new_n59210_,
    new_n59211_, new_n59212_, new_n59213_, new_n59214_, new_n59215_,
    new_n59216_, new_n59217_, new_n59218_, new_n59219_, new_n59220_,
    new_n59221_, new_n59222_, new_n59223_, new_n59224_, new_n59225_,
    new_n59226_, new_n59227_, new_n59228_, new_n59229_, new_n59230_,
    new_n59231_, new_n59232_, new_n59233_, new_n59234_, new_n59235_,
    new_n59236_, new_n59237_, new_n59238_, new_n59239_, new_n59240_,
    new_n59241_, new_n59242_, new_n59243_, new_n59244_, new_n59245_,
    new_n59246_, new_n59247_, new_n59248_, new_n59249_, new_n59250_,
    new_n59251_, new_n59252_, new_n59253_, new_n59254_, new_n59255_,
    new_n59256_, new_n59257_, new_n59258_, new_n59259_, new_n59260_,
    new_n59261_, new_n59262_, new_n59263_, new_n59264_, new_n59265_,
    new_n59266_, new_n59267_, new_n59268_, new_n59269_, new_n59270_,
    new_n59271_, new_n59272_, new_n59273_, new_n59274_, new_n59275_,
    new_n59276_, new_n59277_, new_n59278_, new_n59279_, new_n59280_,
    new_n59281_, new_n59282_, new_n59283_, new_n59284_, new_n59285_,
    new_n59286_, new_n59287_, new_n59288_, new_n59289_, new_n59290_,
    new_n59291_, new_n59292_, new_n59293_, new_n59294_, new_n59295_,
    new_n59296_, new_n59297_, new_n59298_, new_n59299_, new_n59300_,
    new_n59301_, new_n59302_, new_n59303_, new_n59304_, new_n59305_,
    new_n59306_, new_n59307_, new_n59308_, new_n59309_, new_n59310_,
    new_n59311_, new_n59312_, new_n59313_, new_n59314_, new_n59315_,
    new_n59316_, new_n59317_, new_n59318_, new_n59319_, new_n59320_,
    new_n59321_, new_n59322_, new_n59323_, new_n59324_, new_n59325_,
    new_n59326_, new_n59327_, new_n59328_, new_n59329_, new_n59330_,
    new_n59331_, new_n59332_, new_n59333_, new_n59334_, new_n59335_,
    new_n59336_, new_n59337_, new_n59338_, new_n59339_, new_n59340_,
    new_n59341_, new_n59342_, new_n59343_, new_n59344_, new_n59345_,
    new_n59346_, new_n59347_, new_n59348_, new_n59349_, new_n59350_,
    new_n59351_, new_n59352_, new_n59353_, new_n59354_, new_n59355_,
    new_n59356_, new_n59357_, new_n59358_, new_n59359_, new_n59360_,
    new_n59361_, new_n59362_, new_n59363_, new_n59364_, new_n59365_,
    new_n59366_, new_n59367_, new_n59368_, new_n59369_, new_n59370_,
    new_n59371_, new_n59372_, new_n59373_, new_n59374_, new_n59375_,
    new_n59376_, new_n59377_, new_n59378_, new_n59379_, new_n59380_,
    new_n59381_, new_n59382_, new_n59383_, new_n59384_, new_n59385_,
    new_n59386_, new_n59387_, new_n59388_, new_n59389_, new_n59390_,
    new_n59391_, new_n59392_, new_n59393_, new_n59394_, new_n59395_,
    new_n59396_, new_n59397_, new_n59398_, new_n59399_, new_n59400_,
    new_n59401_, new_n59402_, new_n59403_, new_n59404_, new_n59405_,
    new_n59406_, new_n59407_, new_n59408_, new_n59409_, new_n59410_,
    new_n59411_, new_n59412_, new_n59413_, new_n59414_, new_n59415_,
    new_n59416_, new_n59417_, new_n59418_, new_n59419_, new_n59420_,
    new_n59421_, new_n59422_, new_n59423_, new_n59424_, new_n59425_,
    new_n59426_, new_n59427_, new_n59428_, new_n59429_, new_n59430_,
    new_n59431_, new_n59432_, new_n59433_, new_n59434_, new_n59435_,
    new_n59436_, new_n59437_, new_n59438_, new_n59439_, new_n59440_,
    new_n59441_, new_n59442_, new_n59443_, new_n59444_, new_n59445_,
    new_n59446_, new_n59447_, new_n59448_, new_n59449_, new_n59450_,
    new_n59451_, new_n59452_, new_n59453_, new_n59454_, new_n59455_,
    new_n59456_, new_n59457_, new_n59458_, new_n59459_, new_n59460_,
    new_n59461_, new_n59462_, new_n59463_, new_n59464_, new_n59465_,
    new_n59466_, new_n59467_, new_n59468_, new_n59469_, new_n59470_,
    new_n59471_, new_n59472_, new_n59473_, new_n59474_, new_n59475_,
    new_n59476_, new_n59477_, new_n59478_, new_n59479_, new_n59480_,
    new_n59481_, new_n59482_, new_n59483_, new_n59484_, new_n59485_,
    new_n59486_, new_n59487_, new_n59488_, new_n59489_, new_n59490_,
    new_n59491_, new_n59492_, new_n59493_, new_n59494_, new_n59495_,
    new_n59496_, new_n59497_, new_n59498_, new_n59499_, new_n59500_,
    new_n59501_, new_n59502_, new_n59503_, new_n59504_, new_n59505_,
    new_n59506_, new_n59507_, new_n59508_, new_n59509_, new_n59510_,
    new_n59511_, new_n59512_, new_n59513_, new_n59514_, new_n59515_,
    new_n59516_, new_n59517_, new_n59518_, new_n59519_, new_n59520_,
    new_n59521_, new_n59522_, new_n59523_, new_n59524_, new_n59525_,
    new_n59526_, new_n59527_, new_n59528_, new_n59529_, new_n59530_,
    new_n59531_, new_n59532_, new_n59533_, new_n59534_, new_n59535_,
    new_n59536_, new_n59537_, new_n59538_, new_n59539_, new_n59540_,
    new_n59541_, new_n59542_, new_n59543_, new_n59544_, new_n59545_,
    new_n59546_, new_n59547_, new_n59548_, new_n59549_, new_n59550_,
    new_n59551_, new_n59552_, new_n59553_, new_n59554_, new_n59555_,
    new_n59556_, new_n59557_, new_n59558_, new_n59559_, new_n59560_,
    new_n59561_, new_n59562_, new_n59563_, new_n59564_, new_n59565_,
    new_n59566_, new_n59567_, new_n59568_, new_n59569_, new_n59570_,
    new_n59571_, new_n59572_, new_n59573_, new_n59574_, new_n59575_,
    new_n59576_, new_n59577_, new_n59578_, new_n59579_, new_n59580_,
    new_n59581_, new_n59582_, new_n59583_, new_n59584_, new_n59585_,
    new_n59586_, new_n59587_, new_n59588_, new_n59589_, new_n59590_,
    new_n59591_, new_n59592_, new_n59593_, new_n59594_, new_n59595_,
    new_n59596_, new_n59597_, new_n59598_, new_n59599_, new_n59600_,
    new_n59601_, new_n59602_, new_n59603_, new_n59604_, new_n59605_,
    new_n59606_, new_n59607_, new_n59608_, new_n59609_, new_n59610_,
    new_n59611_, new_n59612_, new_n59613_, new_n59614_, new_n59615_,
    new_n59616_, new_n59617_, new_n59618_, new_n59619_, new_n59620_,
    new_n59621_, new_n59622_, new_n59623_, new_n59624_, new_n59625_,
    new_n59626_, new_n59627_, new_n59628_, new_n59629_, new_n59630_,
    new_n59631_, new_n59632_, new_n59633_, new_n59634_, new_n59635_,
    new_n59636_, new_n59637_, new_n59638_, new_n59639_, new_n59640_,
    new_n59641_, new_n59642_, new_n59643_, new_n59644_, new_n59645_,
    new_n59646_, new_n59647_, new_n59648_, new_n59649_, new_n59650_,
    new_n59651_, new_n59652_, new_n59653_, new_n59654_, new_n59655_,
    new_n59656_, new_n59657_, new_n59658_, new_n59659_, new_n59660_,
    new_n59661_, new_n59662_, new_n59663_, new_n59664_, new_n59665_,
    new_n59666_, new_n59667_, new_n59668_, new_n59669_, new_n59670_,
    new_n59671_, new_n59672_, new_n59673_, new_n59674_, new_n59675_,
    new_n59676_, new_n59677_, new_n59678_, new_n59679_, new_n59680_,
    new_n59681_, new_n59682_, new_n59683_, new_n59684_, new_n59685_,
    new_n59686_, new_n59687_, new_n59688_, new_n59689_, new_n59690_,
    new_n59691_, new_n59692_, new_n59693_, new_n59694_, new_n59695_,
    new_n59696_, new_n59697_, new_n59698_, new_n59699_, new_n59700_,
    new_n59701_, new_n59702_, new_n59703_, new_n59704_, new_n59705_,
    new_n59706_, new_n59707_, new_n59708_, new_n59709_, new_n59710_,
    new_n59711_, new_n59712_, new_n59713_, new_n59714_, new_n59715_,
    new_n59716_, new_n59717_, new_n59718_, new_n59719_, new_n59720_,
    new_n59721_, new_n59722_, new_n59723_, new_n59724_, new_n59725_,
    new_n59726_, new_n59727_, new_n59728_, new_n59729_, new_n59730_,
    new_n59731_, new_n59732_, new_n59733_, new_n59734_, new_n59735_,
    new_n59736_, new_n59737_, new_n59738_, new_n59739_, new_n59740_,
    new_n59741_, new_n59742_, new_n59743_, new_n59744_, new_n59745_,
    new_n59746_, new_n59747_, new_n59748_, new_n59749_, new_n59750_,
    new_n59751_, new_n59752_, new_n59753_, new_n59754_, new_n59755_,
    new_n59756_, new_n59757_, new_n59758_, new_n59759_, new_n59760_,
    new_n59761_, new_n59762_, new_n59763_, new_n59764_, new_n59765_,
    new_n59766_, new_n59767_, new_n59768_, new_n59769_, new_n59770_,
    new_n59771_, new_n59772_, new_n59773_, new_n59774_, new_n59775_,
    new_n59776_, new_n59777_, new_n59778_, new_n59779_, new_n59780_,
    new_n59781_, new_n59782_, new_n59783_, new_n59784_, new_n59785_,
    new_n59786_, new_n59787_, new_n59788_, new_n59789_, new_n59790_,
    new_n59791_, new_n59792_, new_n59793_, new_n59794_, new_n59795_,
    new_n59796_, new_n59797_, new_n59798_, new_n59799_, new_n59800_,
    new_n59801_, new_n59802_, new_n59803_, new_n59804_, new_n59805_,
    new_n59806_, new_n59807_, new_n59808_, new_n59809_, new_n59810_,
    new_n59811_, new_n59812_, new_n59813_, new_n59814_, new_n59815_,
    new_n59816_, new_n59817_, new_n59818_, new_n59819_, new_n59820_,
    new_n59821_, new_n59822_, new_n59823_, new_n59824_, new_n59825_,
    new_n59826_, new_n59827_, new_n59828_, new_n59829_, new_n59830_,
    new_n59831_, new_n59832_, new_n59833_, new_n59834_, new_n59835_,
    new_n59836_, new_n59837_, new_n59838_, new_n59839_, new_n59840_,
    new_n59841_, new_n59842_, new_n59843_, new_n59844_, new_n59845_,
    new_n59846_, new_n59847_, new_n59848_, new_n59849_, new_n59850_,
    new_n59851_, new_n59852_, new_n59853_, new_n59854_, new_n59855_,
    new_n59856_, new_n59857_, new_n59858_, new_n59859_, new_n59860_,
    new_n59861_, new_n59862_, new_n59863_, new_n59864_, new_n59865_,
    new_n59866_, new_n59867_, new_n59868_, new_n59869_, new_n59870_,
    new_n59871_, new_n59872_, new_n59873_, new_n59874_, new_n59875_,
    new_n59876_, new_n59877_, new_n59878_, new_n59879_, new_n59880_,
    new_n59881_, new_n59882_, new_n59883_, new_n59884_, new_n59885_,
    new_n59886_, new_n59887_, new_n59888_, new_n59889_, new_n59890_,
    new_n59891_, new_n59892_, new_n59893_, new_n59894_, new_n59895_,
    new_n59896_, new_n59897_, new_n59898_, new_n59899_, new_n59900_,
    new_n59901_, new_n59902_, new_n59903_, new_n59904_, new_n59905_,
    new_n59906_, new_n59907_, new_n59908_, new_n59909_, new_n59910_,
    new_n59911_, new_n59912_, new_n59913_, new_n59914_, new_n59915_,
    new_n59916_, new_n59917_, new_n59918_, new_n59919_, new_n59920_,
    new_n59921_, new_n59922_, new_n59923_, new_n59924_, new_n59925_,
    new_n59926_, new_n59927_, new_n59928_, new_n59929_, new_n59930_,
    new_n59931_, new_n59932_, new_n59933_, new_n59934_, new_n59935_,
    new_n59936_, new_n59937_, new_n59938_, new_n59939_, new_n59940_,
    new_n59941_, new_n59942_, new_n59943_, new_n59944_, new_n59945_,
    new_n59946_, new_n59947_, new_n59948_, new_n59949_, new_n59950_,
    new_n59951_, new_n59952_, new_n59953_, new_n59954_, new_n59955_,
    new_n59956_, new_n59957_, new_n59958_, new_n59959_, new_n59960_,
    new_n59961_, new_n59962_, new_n59963_, new_n59964_, new_n59965_,
    new_n59966_, new_n59967_, new_n59968_, new_n59969_, new_n59970_,
    new_n59971_, new_n59972_, new_n59973_, new_n59974_, new_n59975_,
    new_n59976_, new_n59977_, new_n59978_, new_n59979_, new_n59980_,
    new_n59981_, new_n59982_, new_n59983_, new_n59984_, new_n59985_,
    new_n59986_, new_n59987_, new_n59988_, new_n59989_, new_n59990_,
    new_n59991_, new_n59992_, new_n59993_, new_n59994_, new_n59995_,
    new_n59996_, new_n59997_, new_n59998_, new_n59999_, new_n60000_,
    new_n60001_, new_n60002_, new_n60003_, new_n60004_, new_n60005_,
    new_n60006_, new_n60007_, new_n60008_, new_n60009_, new_n60010_,
    new_n60011_, new_n60012_, new_n60013_, new_n60014_, new_n60015_,
    new_n60016_, new_n60017_, new_n60018_, new_n60019_, new_n60020_,
    new_n60021_, new_n60022_, new_n60023_, new_n60024_, new_n60025_,
    new_n60026_, new_n60027_, new_n60028_, new_n60029_, new_n60030_,
    new_n60031_, new_n60032_, new_n60033_, new_n60034_, new_n60035_,
    new_n60036_, new_n60037_, new_n60038_, new_n60039_, new_n60040_,
    new_n60041_, new_n60042_, new_n60043_, new_n60044_, new_n60045_,
    new_n60046_, new_n60047_, new_n60048_, new_n60049_, new_n60050_,
    new_n60051_, new_n60052_, new_n60053_, new_n60054_, new_n60055_,
    new_n60056_, new_n60057_, new_n60058_, new_n60059_, new_n60060_,
    new_n60061_, new_n60062_, new_n60063_, new_n60064_, new_n60065_,
    new_n60066_, new_n60067_, new_n60068_, new_n60069_, new_n60070_,
    new_n60071_, new_n60072_, new_n60073_, new_n60074_, new_n60075_,
    new_n60076_, new_n60077_, new_n60078_, new_n60079_, new_n60080_,
    new_n60081_, new_n60082_, new_n60083_, new_n60084_, new_n60085_,
    new_n60086_, new_n60087_, new_n60088_, new_n60089_, new_n60090_,
    new_n60091_, new_n60092_, new_n60093_, new_n60094_, new_n60095_,
    new_n60096_, new_n60097_, new_n60098_, new_n60099_, new_n60100_,
    new_n60101_, new_n60102_, new_n60103_, new_n60104_, new_n60105_,
    new_n60106_, new_n60107_, new_n60108_, new_n60109_, new_n60110_,
    new_n60111_, new_n60112_, new_n60113_, new_n60114_, new_n60115_,
    new_n60116_, new_n60117_, new_n60118_, new_n60119_, new_n60120_,
    new_n60121_, new_n60122_, new_n60123_, new_n60124_, new_n60125_,
    new_n60126_, new_n60127_, new_n60128_, new_n60129_, new_n60130_,
    new_n60131_, new_n60132_, new_n60133_, new_n60134_, new_n60135_,
    new_n60136_, new_n60137_, new_n60138_, new_n60139_, new_n60140_,
    new_n60141_, new_n60142_, new_n60143_, new_n60144_, new_n60145_,
    new_n60146_, new_n60147_, new_n60148_, new_n60149_, new_n60150_,
    new_n60151_, new_n60152_, new_n60153_, new_n60154_, new_n60155_,
    new_n60156_, new_n60157_, new_n60158_, new_n60159_, new_n60160_,
    new_n60161_, new_n60162_, new_n60163_, new_n60164_, new_n60165_,
    new_n60166_, new_n60167_, new_n60168_, new_n60169_, new_n60170_,
    new_n60171_, new_n60172_, new_n60173_, new_n60174_, new_n60175_,
    new_n60176_, new_n60177_, new_n60178_, new_n60179_, new_n60180_,
    new_n60181_, new_n60182_, new_n60183_, new_n60184_, new_n60185_,
    new_n60186_, new_n60187_, new_n60188_, new_n60189_, new_n60190_,
    new_n60191_, new_n60192_, new_n60193_, new_n60194_, new_n60195_,
    new_n60196_, new_n60197_, new_n60198_, new_n60199_, new_n60200_,
    new_n60201_, new_n60202_, new_n60203_, new_n60204_, new_n60205_,
    new_n60206_, new_n60207_, new_n60208_, new_n60209_, new_n60210_,
    new_n60211_, new_n60212_, new_n60213_, new_n60214_, new_n60215_,
    new_n60216_, new_n60217_, new_n60218_, new_n60219_, new_n60220_,
    new_n60221_, new_n60222_, new_n60223_, new_n60224_, new_n60225_,
    new_n60226_, new_n60227_, new_n60228_, new_n60229_, new_n60230_,
    new_n60231_, new_n60232_, new_n60233_, new_n60234_, new_n60235_,
    new_n60236_, new_n60237_, new_n60238_, new_n60239_, new_n60240_,
    new_n60241_, new_n60242_, new_n60243_, new_n60244_, new_n60245_,
    new_n60246_, new_n60247_, new_n60248_, new_n60249_, new_n60250_,
    new_n60251_, new_n60252_, new_n60253_, new_n60254_, new_n60255_,
    new_n60256_, new_n60257_, new_n60258_, new_n60259_, new_n60260_,
    new_n60261_, new_n60262_, new_n60263_, new_n60264_, new_n60265_,
    new_n60266_, new_n60267_, new_n60268_, new_n60269_, new_n60270_,
    new_n60271_, new_n60272_, new_n60273_, new_n60274_, new_n60275_,
    new_n60276_, new_n60277_, new_n60278_, new_n60279_, new_n60280_,
    new_n60281_, new_n60282_, new_n60283_, new_n60284_, new_n60285_,
    new_n60286_, new_n60287_, new_n60288_, new_n60289_, new_n60290_,
    new_n60291_, new_n60292_, new_n60293_, new_n60294_, new_n60295_,
    new_n60296_, new_n60297_, new_n60298_, new_n60299_, new_n60300_,
    new_n60301_, new_n60302_, new_n60303_, new_n60304_, new_n60305_,
    new_n60306_, new_n60307_, new_n60308_, new_n60309_, new_n60310_,
    new_n60311_, new_n60312_, new_n60313_, new_n60314_, new_n60315_,
    new_n60316_, new_n60317_, new_n60318_, new_n60319_, new_n60320_,
    new_n60321_, new_n60322_, new_n60323_, new_n60324_, new_n60325_,
    new_n60326_, new_n60327_, new_n60328_, new_n60329_, new_n60330_,
    new_n60331_, new_n60332_, new_n60333_, new_n60334_, new_n60335_,
    new_n60336_, new_n60337_, new_n60338_, new_n60339_, new_n60340_,
    new_n60341_, new_n60342_, new_n60343_, new_n60344_, new_n60345_,
    new_n60346_, new_n60347_, new_n60348_, new_n60349_, new_n60350_,
    new_n60351_, new_n60352_, new_n60353_, new_n60354_, new_n60355_,
    new_n60356_, new_n60357_, new_n60358_, new_n60359_, new_n60360_,
    new_n60361_, new_n60362_, new_n60363_, new_n60364_, new_n60365_,
    new_n60366_, new_n60367_, new_n60368_, new_n60369_, new_n60370_,
    new_n60371_, new_n60372_, new_n60373_, new_n60374_, new_n60375_,
    new_n60376_, new_n60377_, new_n60378_, new_n60379_, new_n60380_,
    new_n60381_, new_n60382_, new_n60383_, new_n60384_, new_n60385_,
    new_n60386_, new_n60387_, new_n60388_, new_n60389_, new_n60390_,
    new_n60391_, new_n60392_, new_n60393_, new_n60394_, new_n60395_,
    new_n60396_, new_n60397_, new_n60398_, new_n60399_, new_n60400_,
    new_n60401_, new_n60402_, new_n60403_, new_n60404_, new_n60405_,
    new_n60406_, new_n60407_, new_n60408_, new_n60409_, new_n60410_,
    new_n60411_, new_n60412_, new_n60413_, new_n60414_, new_n60415_,
    new_n60416_, new_n60417_, new_n60418_, new_n60419_, new_n60420_,
    new_n60421_, new_n60422_, new_n60423_, new_n60424_, new_n60425_,
    new_n60426_, new_n60427_, new_n60428_, new_n60429_, new_n60430_,
    new_n60431_, new_n60432_, new_n60433_, new_n60434_, new_n60435_,
    new_n60436_, new_n60437_, new_n60438_, new_n60439_, new_n60440_,
    new_n60441_, new_n60442_, new_n60443_, new_n60444_, new_n60445_,
    new_n60446_, new_n60447_, new_n60448_, new_n60449_, new_n60450_,
    new_n60451_, new_n60452_, new_n60453_, new_n60454_, new_n60455_,
    new_n60456_, new_n60457_, new_n60458_, new_n60459_, new_n60460_,
    new_n60461_, new_n60462_, new_n60463_, new_n60464_, new_n60465_,
    new_n60466_, new_n60467_, new_n60468_, new_n60469_, new_n60470_,
    new_n60471_, new_n60472_, new_n60473_, new_n60474_, new_n60475_,
    new_n60476_, new_n60477_, new_n60478_, new_n60479_, new_n60480_,
    new_n60481_, new_n60482_, new_n60483_, new_n60484_, new_n60485_,
    new_n60486_, new_n60487_, new_n60488_, new_n60489_, new_n60490_,
    new_n60491_, new_n60492_, new_n60493_, new_n60494_, new_n60495_,
    new_n60496_, new_n60497_, new_n60498_, new_n60499_, new_n60500_,
    new_n60501_, new_n60502_, new_n60503_, new_n60504_, new_n60505_,
    new_n60506_, new_n60507_, new_n60508_, new_n60509_, new_n60510_,
    new_n60511_, new_n60512_, new_n60513_, new_n60514_, new_n60515_,
    new_n60516_, new_n60517_, new_n60518_, new_n60519_, new_n60520_,
    new_n60521_, new_n60522_, new_n60523_, new_n60524_, new_n60525_,
    new_n60526_, new_n60527_, new_n60528_, new_n60529_, new_n60530_,
    new_n60531_, new_n60532_, new_n60533_, new_n60534_, new_n60535_,
    new_n60536_, new_n60537_, new_n60538_, new_n60539_, new_n60540_,
    new_n60541_, new_n60542_, new_n60543_, new_n60544_, new_n60545_,
    new_n60546_, new_n60547_, new_n60548_, new_n60549_, new_n60550_,
    new_n60551_, new_n60552_, new_n60553_, new_n60554_, new_n60555_,
    new_n60556_, new_n60557_, new_n60558_, new_n60559_, new_n60560_,
    new_n60561_, new_n60562_, new_n60563_, new_n60564_, new_n60565_,
    new_n60566_, new_n60567_, new_n60568_, new_n60569_, new_n60570_,
    new_n60571_, new_n60572_, new_n60573_, new_n60574_, new_n60575_,
    new_n60576_, new_n60577_, new_n60578_, new_n60579_, new_n60580_,
    new_n60581_, new_n60582_, new_n60583_, new_n60584_, new_n60585_,
    new_n60586_, new_n60587_, new_n60588_, new_n60589_, new_n60590_,
    new_n60591_, new_n60592_, new_n60593_, new_n60594_, new_n60595_,
    new_n60596_, new_n60597_, new_n60598_, new_n60599_, new_n60600_,
    new_n60601_, new_n60602_, new_n60603_, new_n60604_, new_n60605_,
    new_n60606_, new_n60607_, new_n60608_, new_n60609_, new_n60610_,
    new_n60611_, new_n60612_, new_n60613_, new_n60614_, new_n60615_,
    new_n60616_, new_n60617_, new_n60618_, new_n60619_, new_n60620_,
    new_n60621_, new_n60622_, new_n60623_, new_n60624_, new_n60625_,
    new_n60626_, new_n60627_, new_n60628_, new_n60629_, new_n60630_,
    new_n60631_, new_n60632_, new_n60633_, new_n60634_, new_n60635_,
    new_n60636_, new_n60637_, new_n60638_, new_n60639_, new_n60640_,
    new_n60641_, new_n60642_, new_n60643_, new_n60644_, new_n60645_,
    new_n60646_, new_n60647_, new_n60648_, new_n60649_, new_n60650_,
    new_n60651_, new_n60652_, new_n60653_, new_n60654_, new_n60655_,
    new_n60656_, new_n60657_, new_n60658_, new_n60659_, new_n60660_,
    new_n60661_, new_n60662_, new_n60663_, new_n60664_, new_n60665_,
    new_n60666_, new_n60667_, new_n60668_, new_n60669_, new_n60670_,
    new_n60671_, new_n60672_, new_n60673_, new_n60674_, new_n60675_,
    new_n60676_, new_n60677_, new_n60678_, new_n60679_, new_n60680_,
    new_n60681_, new_n60682_, new_n60683_, new_n60684_, new_n60685_,
    new_n60686_, new_n60687_, new_n60688_, new_n60689_, new_n60690_,
    new_n60691_, new_n60692_, new_n60693_, new_n60694_, new_n60695_,
    new_n60696_, new_n60697_, new_n60698_, new_n60699_, new_n60700_,
    new_n60701_, new_n60702_, new_n60703_, new_n60704_, new_n60705_,
    new_n60706_, new_n60707_, new_n60708_, new_n60709_, new_n60710_,
    new_n60711_, new_n60712_, new_n60713_, new_n60714_, new_n60715_,
    new_n60716_, new_n60717_, new_n60718_, new_n60719_, new_n60720_,
    new_n60721_, new_n60722_, new_n60723_, new_n60724_, new_n60725_,
    new_n60726_, new_n60727_, new_n60728_, new_n60729_, new_n60730_,
    new_n60731_, new_n60732_, new_n60733_, new_n60734_, new_n60735_,
    new_n60736_, new_n60737_, new_n60738_, new_n60739_, new_n60740_,
    new_n60741_, new_n60742_, new_n60743_, new_n60744_, new_n60745_,
    new_n60746_, new_n60747_, new_n60748_, new_n60749_, new_n60750_,
    new_n60751_, new_n60752_, new_n60753_, new_n60754_, new_n60755_,
    new_n60756_, new_n60757_, new_n60758_, new_n60759_, new_n60760_,
    new_n60761_, new_n60762_, new_n60763_, new_n60764_, new_n60765_,
    new_n60766_, new_n60767_, new_n60768_, new_n60769_, new_n60770_,
    new_n60771_, new_n60772_, new_n60773_, new_n60774_, new_n60775_,
    new_n60776_, new_n60777_, new_n60778_, new_n60779_, new_n60780_,
    new_n60781_, new_n60782_, new_n60783_, new_n60784_, new_n60785_,
    new_n60786_, new_n60787_, new_n60788_, new_n60789_, new_n60790_,
    new_n60791_, new_n60792_, new_n60793_, new_n60794_, new_n60795_,
    new_n60796_, new_n60797_, new_n60798_, new_n60799_, new_n60800_,
    new_n60801_, new_n60802_, new_n60803_, new_n60804_, new_n60805_,
    new_n60806_, new_n60807_, new_n60808_, new_n60809_, new_n60810_,
    new_n60811_, new_n60812_, new_n60813_, new_n60814_, new_n60815_,
    new_n60816_, new_n60817_, new_n60818_, new_n60819_, new_n60820_,
    new_n60821_, new_n60822_, new_n60823_, new_n60824_, new_n60825_,
    new_n60826_, new_n60827_, new_n60828_, new_n60829_, new_n60830_,
    new_n60831_, new_n60832_, new_n60833_, new_n60834_, new_n60835_,
    new_n60836_, new_n60837_, new_n60838_, new_n60839_, new_n60840_,
    new_n60841_, new_n60842_, new_n60843_, new_n60844_, new_n60845_,
    new_n60846_, new_n60847_, new_n60848_, new_n60849_, new_n60850_,
    new_n60851_, new_n60852_, new_n60853_, new_n60854_, new_n60855_,
    new_n60856_, new_n60857_, new_n60858_, new_n60859_, new_n60860_,
    new_n60861_, new_n60862_, new_n60863_, new_n60864_, new_n60865_,
    new_n60866_, new_n60867_, new_n60868_, new_n60869_, new_n60870_,
    new_n60871_, new_n60872_, new_n60873_, new_n60874_, new_n60875_,
    new_n60876_, new_n60877_, new_n60878_, new_n60879_, new_n60880_,
    new_n60881_, new_n60882_, new_n60883_, new_n60884_, new_n60885_,
    new_n60886_, new_n60887_, new_n60888_, new_n60889_, new_n60890_,
    new_n60891_, new_n60892_, new_n60893_, new_n60894_, new_n60895_,
    new_n60896_, new_n60897_, new_n60898_, new_n60899_, new_n60900_,
    new_n60901_, new_n60902_, new_n60903_, new_n60904_, new_n60905_,
    new_n60906_, new_n60907_, new_n60908_, new_n60909_, new_n60910_,
    new_n60911_, new_n60912_, new_n60913_, new_n60914_, new_n60915_,
    new_n60916_, new_n60917_, new_n60918_, new_n60919_, new_n60920_,
    new_n60921_, new_n60922_, new_n60923_, new_n60924_, new_n60925_,
    new_n60926_, new_n60927_, new_n60928_, new_n60929_, new_n60930_,
    new_n60931_, new_n60932_, new_n60933_, new_n60934_, new_n60935_,
    new_n60936_, new_n60937_, new_n60938_, new_n60939_, new_n60940_,
    new_n60941_, new_n60942_, new_n60943_, new_n60944_, new_n60945_,
    new_n60946_, new_n60947_, new_n60948_, new_n60949_, new_n60950_,
    new_n60951_, new_n60952_, new_n60953_, new_n60954_, new_n60955_,
    new_n60956_, new_n60957_, new_n60958_, new_n60959_, new_n60960_,
    new_n60961_, new_n60962_, new_n60963_, new_n60964_, new_n60965_,
    new_n60966_, new_n60967_, new_n60968_, new_n60969_, new_n60970_,
    new_n60971_, new_n60972_, new_n60973_, new_n60974_, new_n60975_,
    new_n60976_, new_n60977_, new_n60978_, new_n60979_, new_n60980_,
    new_n60981_, new_n60982_, new_n60983_, new_n60984_, new_n60985_,
    new_n60986_, new_n60987_, new_n60988_, new_n60989_, new_n60990_,
    new_n60991_, new_n60992_, new_n60993_, new_n60994_, new_n60995_,
    new_n60996_, new_n60997_, new_n60998_, new_n60999_, new_n61000_,
    new_n61001_, new_n61002_, new_n61003_, new_n61004_, new_n61005_,
    new_n61006_, new_n61007_, new_n61008_, new_n61009_, new_n61010_,
    new_n61011_, new_n61012_, new_n61013_, new_n61014_, new_n61015_,
    new_n61016_, new_n61017_, new_n61018_, new_n61019_, new_n61020_,
    new_n61021_, new_n61022_, new_n61023_, new_n61024_, new_n61025_,
    new_n61026_, new_n61027_, new_n61028_, new_n61029_, new_n61030_,
    new_n61031_, new_n61032_, new_n61033_, new_n61034_, new_n61035_,
    new_n61036_, new_n61037_, new_n61038_, new_n61039_, new_n61040_,
    new_n61041_, new_n61042_, new_n61043_, new_n61044_, new_n61045_,
    new_n61046_, new_n61047_, new_n61048_, new_n61049_, new_n61050_,
    new_n61051_, new_n61052_, new_n61053_, new_n61054_, new_n61055_,
    new_n61056_, new_n61057_, new_n61058_, new_n61059_, new_n61060_,
    new_n61061_, new_n61062_, new_n61063_, new_n61064_, new_n61065_,
    new_n61066_, new_n61067_, new_n61068_, new_n61069_, new_n61070_,
    new_n61071_, new_n61072_, new_n61073_, new_n61074_, new_n61075_,
    new_n61076_, new_n61077_, new_n61078_, new_n61079_, new_n61080_,
    new_n61081_, new_n61082_, new_n61083_, new_n61084_, new_n61085_,
    new_n61086_, new_n61087_, new_n61088_, new_n61089_, new_n61090_,
    new_n61091_, new_n61092_, new_n61093_, new_n61094_, new_n61095_,
    new_n61096_, new_n61097_, new_n61098_, new_n61099_, new_n61100_,
    new_n61101_, new_n61102_, new_n61103_, new_n61104_, new_n61105_,
    new_n61106_, new_n61107_, new_n61108_, new_n61109_, new_n61110_,
    new_n61111_, new_n61112_, new_n61113_, new_n61114_, new_n61115_,
    new_n61116_, new_n61117_, new_n61118_, new_n61119_, new_n61120_,
    new_n61121_, new_n61122_, new_n61123_, new_n61124_, new_n61125_,
    new_n61126_, new_n61127_, new_n61128_, new_n61129_, new_n61130_,
    new_n61131_, new_n61132_, new_n61133_, new_n61134_, new_n61135_,
    new_n61136_, new_n61137_, new_n61138_, new_n61139_, new_n61140_,
    new_n61141_, new_n61142_, new_n61143_, new_n61144_, new_n61145_,
    new_n61146_, new_n61147_, new_n61148_, new_n61149_, new_n61150_,
    new_n61151_, new_n61152_, new_n61153_, new_n61154_, new_n61155_,
    new_n61156_, new_n61157_, new_n61158_, new_n61159_, new_n61160_,
    new_n61161_, new_n61162_, new_n61163_, new_n61164_, new_n61165_,
    new_n61166_, new_n61167_, new_n61168_, new_n61169_, new_n61170_,
    new_n61171_, new_n61172_, new_n61173_, new_n61174_, new_n61175_,
    new_n61176_, new_n61177_, new_n61178_, new_n61179_, new_n61180_,
    new_n61181_, new_n61182_, new_n61183_, new_n61184_, new_n61185_,
    new_n61186_, new_n61187_, new_n61188_, new_n61189_, new_n61190_,
    new_n61191_, new_n61192_, new_n61193_, new_n61194_, new_n61195_,
    new_n61196_, new_n61197_, new_n61198_, new_n61199_, new_n61200_,
    new_n61201_, new_n61202_, new_n61203_, new_n61204_, new_n61205_,
    new_n61206_, new_n61207_, new_n61208_, new_n61209_, new_n61210_,
    new_n61211_, new_n61212_, new_n61213_, new_n61214_, new_n61215_,
    new_n61216_, new_n61217_, new_n61218_, new_n61219_, new_n61220_,
    new_n61221_, new_n61222_, new_n61223_, new_n61224_, new_n61225_,
    new_n61226_, new_n61227_, new_n61228_, new_n61229_, new_n61230_,
    new_n61231_, new_n61232_, new_n61233_, new_n61234_, new_n61235_,
    new_n61236_, new_n61237_, new_n61238_, new_n61239_, new_n61240_,
    new_n61241_, new_n61242_, new_n61243_, new_n61244_, new_n61245_,
    new_n61246_, new_n61247_, new_n61248_, new_n61249_, new_n61250_,
    new_n61251_, new_n61252_, new_n61253_, new_n61254_, new_n61255_,
    new_n61256_, new_n61257_, new_n61258_, new_n61259_, new_n61260_,
    new_n61261_, new_n61262_, new_n61263_, new_n61264_, new_n61265_,
    new_n61266_, new_n61267_, new_n61268_, new_n61269_, new_n61270_,
    new_n61271_, new_n61272_, new_n61273_, new_n61274_, new_n61275_,
    new_n61276_, new_n61277_, new_n61278_, new_n61279_, new_n61280_,
    new_n61281_, new_n61282_, new_n61283_, new_n61284_, new_n61285_,
    new_n61286_, new_n61287_, new_n61288_, new_n61289_, new_n61290_,
    new_n61291_, new_n61292_, new_n61293_, new_n61294_, new_n61295_,
    new_n61296_, new_n61297_, new_n61298_, new_n61299_, new_n61300_,
    new_n61301_, new_n61302_, new_n61303_, new_n61304_, new_n61305_,
    new_n61306_, new_n61307_, new_n61308_, new_n61309_, new_n61310_,
    new_n61311_, new_n61312_, new_n61313_, new_n61314_, new_n61315_,
    new_n61316_, new_n61317_, new_n61318_, new_n61319_, new_n61320_,
    new_n61321_, new_n61322_, new_n61323_, new_n61324_, new_n61325_,
    new_n61326_, new_n61327_, new_n61328_, new_n61329_, new_n61330_,
    new_n61331_, new_n61332_, new_n61333_, new_n61334_, new_n61335_,
    new_n61336_, new_n61337_, new_n61338_, new_n61339_, new_n61340_,
    new_n61341_, new_n61342_, new_n61343_, new_n61344_, new_n61345_,
    new_n61346_, new_n61347_, new_n61348_, new_n61349_, new_n61350_,
    new_n61351_, new_n61352_, new_n61353_, new_n61354_, new_n61355_,
    new_n61356_, new_n61357_, new_n61358_, new_n61359_, new_n61360_,
    new_n61361_, new_n61362_, new_n61363_, new_n61364_, new_n61365_,
    new_n61366_, new_n61367_, new_n61368_, new_n61369_, new_n61370_,
    new_n61371_, new_n61372_, new_n61373_, new_n61374_, new_n61375_,
    new_n61376_, new_n61377_, new_n61378_, new_n61379_, new_n61380_,
    new_n61381_, new_n61382_, new_n61383_, new_n61384_, new_n61385_,
    new_n61386_, new_n61387_, new_n61388_, new_n61389_, new_n61390_,
    new_n61391_, new_n61392_, new_n61393_, new_n61394_, new_n61395_,
    new_n61396_, new_n61397_, new_n61398_, new_n61399_, new_n61400_,
    new_n61401_, new_n61402_, new_n61403_, new_n61404_, new_n61405_,
    new_n61406_, new_n61407_, new_n61408_, new_n61409_, new_n61410_,
    new_n61411_, new_n61412_, new_n61413_, new_n61414_, new_n61415_,
    new_n61416_, new_n61417_, new_n61418_, new_n61419_, new_n61420_,
    new_n61421_, new_n61422_, new_n61423_, new_n61424_, new_n61425_,
    new_n61426_, new_n61427_, new_n61428_, new_n61429_, new_n61430_,
    new_n61431_, new_n61432_, new_n61433_, new_n61434_, new_n61435_,
    new_n61436_, new_n61437_, new_n61438_, new_n61439_, new_n61440_,
    new_n61441_, new_n61442_, new_n61443_, new_n61444_, new_n61445_,
    new_n61446_, new_n61447_, new_n61448_, new_n61449_, new_n61450_,
    new_n61451_, new_n61452_, new_n61453_, new_n61454_, new_n61455_,
    new_n61456_, new_n61457_, new_n61458_, new_n61459_, new_n61460_,
    new_n61461_, new_n61462_, new_n61463_, new_n61464_, new_n61465_,
    new_n61466_, new_n61467_, new_n61468_, new_n61469_, new_n61470_,
    new_n61471_, new_n61472_, new_n61473_, new_n61474_, new_n61475_,
    new_n61476_, new_n61477_, new_n61478_, new_n61479_, new_n61480_,
    new_n61481_, new_n61482_, new_n61483_, new_n61484_, new_n61485_,
    new_n61486_, new_n61487_, new_n61488_, new_n61489_, new_n61490_,
    new_n61491_, new_n61492_, new_n61493_, new_n61494_, new_n61495_,
    new_n61496_, new_n61497_, new_n61498_, new_n61499_, new_n61500_,
    new_n61501_, new_n61502_, new_n61503_, new_n61504_, new_n61505_,
    new_n61506_, new_n61507_, new_n61508_, new_n61509_, new_n61510_,
    new_n61511_, new_n61512_, new_n61513_, new_n61514_, new_n61515_,
    new_n61516_, new_n61517_, new_n61518_, new_n61519_, new_n61520_,
    new_n61521_, new_n61522_, new_n61523_, new_n61524_, new_n61525_,
    new_n61526_, new_n61527_, new_n61528_, new_n61529_, new_n61530_,
    new_n61531_, new_n61532_, new_n61533_, new_n61534_, new_n61535_,
    new_n61536_, new_n61537_, new_n61538_, new_n61539_, new_n61540_,
    new_n61541_, new_n61542_, new_n61543_, new_n61544_, new_n61545_,
    new_n61546_, new_n61547_, new_n61548_, new_n61549_, new_n61550_,
    new_n61551_, new_n61552_, new_n61553_, new_n61554_, new_n61555_,
    new_n61556_, new_n61557_, new_n61558_, new_n61559_, new_n61560_,
    new_n61561_, new_n61562_, new_n61563_, new_n61564_, new_n61565_,
    new_n61566_, new_n61567_, new_n61568_, new_n61569_, new_n61570_,
    new_n61571_, new_n61572_, new_n61573_, new_n61574_, new_n61575_,
    new_n61576_, new_n61577_, new_n61578_, new_n61579_, new_n61580_,
    new_n61581_, new_n61582_, new_n61583_, new_n61584_, new_n61585_,
    new_n61586_, new_n61587_, new_n61588_, new_n61589_, new_n61590_,
    new_n61591_, new_n61592_, new_n61593_, new_n61594_, new_n61595_,
    new_n61596_, new_n61597_, new_n61598_, new_n61599_, new_n61600_,
    new_n61601_, new_n61602_, new_n61603_, new_n61604_, new_n61605_,
    new_n61606_, new_n61607_, new_n61608_, new_n61609_, new_n61610_,
    new_n61611_, new_n61612_, new_n61613_, new_n61614_, new_n61615_,
    new_n61616_, new_n61617_, new_n61618_, new_n61619_, new_n61620_,
    new_n61621_, new_n61622_, new_n61623_, new_n61624_, new_n61625_,
    new_n61626_, new_n61627_, new_n61628_, new_n61629_, new_n61630_,
    new_n61631_, new_n61632_, new_n61633_, new_n61634_, new_n61635_,
    new_n61636_, new_n61637_, new_n61638_, new_n61639_, new_n61640_,
    new_n61641_, new_n61642_, new_n61643_, new_n61644_, new_n61645_,
    new_n61646_, new_n61647_, new_n61648_, new_n61649_, new_n61650_,
    new_n61651_, new_n61652_, new_n61653_, new_n61654_, new_n61655_,
    new_n61656_, new_n61657_, new_n61658_, new_n61659_, new_n61660_,
    new_n61661_, new_n61662_, new_n61663_, new_n61664_, new_n61665_,
    new_n61666_, new_n61667_, new_n61668_, new_n61669_, new_n61670_,
    new_n61671_, new_n61672_, new_n61673_, new_n61674_, new_n61675_,
    new_n61676_, new_n61677_, new_n61678_, new_n61679_, new_n61680_,
    new_n61681_, new_n61682_, new_n61683_, new_n61684_, new_n61685_,
    new_n61686_, new_n61687_, new_n61688_, new_n61689_, new_n61690_,
    new_n61691_, new_n61692_, new_n61693_, new_n61694_, new_n61695_,
    new_n61696_, new_n61697_, new_n61698_, new_n61699_, new_n61700_,
    new_n61701_, new_n61702_, new_n61703_, new_n61704_, new_n61705_,
    new_n61706_, new_n61707_, new_n61708_, new_n61709_, new_n61710_,
    new_n61711_, new_n61712_, new_n61713_, new_n61714_, new_n61715_,
    new_n61716_, new_n61717_, new_n61718_, new_n61719_, new_n61720_,
    new_n61721_, new_n61722_, new_n61723_, new_n61724_, new_n61725_,
    new_n61726_, new_n61727_, new_n61728_, new_n61729_, new_n61730_,
    new_n61731_, new_n61732_, new_n61733_, new_n61734_, new_n61735_,
    new_n61736_, new_n61737_, new_n61738_, new_n61739_, new_n61740_,
    new_n61741_, new_n61742_, new_n61743_, new_n61744_, new_n61745_,
    new_n61746_, new_n61747_, new_n61748_, new_n61749_, new_n61750_,
    new_n61751_, new_n61752_, new_n61753_, new_n61754_, new_n61755_,
    new_n61756_, new_n61757_, new_n61758_, new_n61759_, new_n61760_,
    new_n61761_, new_n61762_, new_n61763_, new_n61764_, new_n61765_,
    new_n61766_, new_n61767_, new_n61768_, new_n61769_, new_n61770_,
    new_n61771_, new_n61772_, new_n61773_, new_n61774_, new_n61775_,
    new_n61776_, new_n61777_, new_n61778_, new_n61779_, new_n61780_,
    new_n61781_, new_n61782_, new_n61783_, new_n61784_, new_n61785_,
    new_n61786_, new_n61787_, new_n61788_, new_n61789_, new_n61790_,
    new_n61791_, new_n61792_, new_n61793_, new_n61794_, new_n61795_,
    new_n61796_, new_n61797_, new_n61798_, new_n61799_, new_n61800_,
    new_n61801_, new_n61802_, new_n61803_, new_n61804_, new_n61805_,
    new_n61806_, new_n61807_, new_n61808_, new_n61809_, new_n61810_,
    new_n61811_, new_n61812_, new_n61813_, new_n61814_, new_n61815_,
    new_n61816_, new_n61817_, new_n61818_, new_n61819_, new_n61820_,
    new_n61821_, new_n61822_, new_n61823_, new_n61824_, new_n61825_,
    new_n61826_, new_n61827_, new_n61828_, new_n61829_, new_n61830_,
    new_n61831_, new_n61832_, new_n61833_, new_n61834_, new_n61835_,
    new_n61836_, new_n61837_, new_n61838_, new_n61839_, new_n61840_,
    new_n61841_, new_n61842_, new_n61843_, new_n61844_, new_n61845_,
    new_n61846_, new_n61847_, new_n61848_, new_n61849_, new_n61850_,
    new_n61851_, new_n61852_, new_n61853_, new_n61854_, new_n61855_,
    new_n61856_, new_n61857_, new_n61858_, new_n61859_, new_n61860_,
    new_n61861_, new_n61862_, new_n61863_, new_n61864_, new_n61865_,
    new_n61866_, new_n61867_, new_n61868_, new_n61869_, new_n61870_,
    new_n61871_, new_n61872_, new_n61873_, new_n61874_, new_n61875_,
    new_n61876_, new_n61877_, new_n61878_, new_n61879_, new_n61880_,
    new_n61881_, new_n61882_, new_n61883_, new_n61884_, new_n61885_,
    new_n61886_, new_n61887_, new_n61888_, new_n61889_, new_n61890_,
    new_n61891_, new_n61892_, new_n61893_, new_n61894_, new_n61895_,
    new_n61896_, new_n61897_, new_n61898_, new_n61899_, new_n61900_,
    new_n61901_, new_n61902_, new_n61903_, new_n61904_, new_n61905_,
    new_n61906_, new_n61907_, new_n61908_, new_n61909_, new_n61910_,
    new_n61911_, new_n61912_, new_n61913_, new_n61914_, new_n61915_,
    new_n61916_, new_n61917_, new_n61918_, new_n61919_, new_n61920_,
    new_n61921_, new_n61922_, new_n61923_, new_n61924_, new_n61925_,
    new_n61926_, new_n61927_, new_n61928_, new_n61929_, new_n61930_,
    new_n61931_, new_n61932_, new_n61933_, new_n61934_, new_n61935_,
    new_n61936_, new_n61937_, new_n61938_, new_n61939_, new_n61940_,
    new_n61941_, new_n61942_, new_n61943_, new_n61944_, new_n61945_,
    new_n61946_, new_n61947_, new_n61948_, new_n61949_, new_n61950_,
    new_n61951_, new_n61952_, new_n61953_, new_n61954_, new_n61955_,
    new_n61956_, new_n61957_, new_n61958_, new_n61959_, new_n61960_,
    new_n61961_, new_n61962_, new_n61963_, new_n61964_, new_n61965_,
    new_n61966_, new_n61967_, new_n61968_, new_n61969_, new_n61970_,
    new_n61971_, new_n61972_, new_n61973_, new_n61974_, new_n61975_,
    new_n61976_, new_n61977_, new_n61978_, new_n61979_, new_n61980_,
    new_n61981_, new_n61982_, new_n61983_, new_n61984_, new_n61985_,
    new_n61986_, new_n61987_, new_n61988_, new_n61989_, new_n61990_,
    new_n61991_, new_n61992_, new_n61993_, new_n61994_, new_n61995_,
    new_n61996_, new_n61997_, new_n61998_, new_n61999_, new_n62000_,
    new_n62001_, new_n62002_, new_n62003_, new_n62004_, new_n62005_,
    new_n62006_, new_n62007_, new_n62008_, new_n62009_, new_n62010_,
    new_n62011_, new_n62012_, new_n62013_, new_n62014_, new_n62015_,
    new_n62016_, new_n62017_, new_n62018_, new_n62019_, new_n62020_,
    new_n62021_, new_n62022_, new_n62023_, new_n62024_, new_n62025_,
    new_n62026_, new_n62027_, new_n62028_, new_n62029_, new_n62030_,
    new_n62031_, new_n62032_, new_n62033_, new_n62034_, new_n62035_,
    new_n62036_, new_n62037_, new_n62038_, new_n62039_, new_n62040_,
    new_n62041_, new_n62042_, new_n62043_, new_n62044_, new_n62045_,
    new_n62046_, new_n62047_, new_n62048_, new_n62049_, new_n62050_,
    new_n62051_, new_n62052_, new_n62053_, new_n62054_, new_n62055_,
    new_n62056_, new_n62057_, new_n62058_, new_n62059_, new_n62060_,
    new_n62061_, new_n62062_, new_n62063_, new_n62064_, new_n62065_,
    new_n62066_, new_n62067_, new_n62068_, new_n62069_, new_n62070_,
    new_n62071_, new_n62072_, new_n62073_, new_n62074_, new_n62075_,
    new_n62076_, new_n62077_, new_n62078_, new_n62079_, new_n62080_,
    new_n62081_, new_n62082_, new_n62083_, new_n62084_, new_n62085_,
    new_n62086_, new_n62087_, new_n62088_, new_n62089_, new_n62090_,
    new_n62091_, new_n62092_, new_n62093_, new_n62094_, new_n62095_,
    new_n62096_, new_n62097_, new_n62098_, new_n62099_, new_n62100_,
    new_n62101_, new_n62102_, new_n62103_, new_n62104_, new_n62105_,
    new_n62106_, new_n62107_, new_n62108_, new_n62109_, new_n62110_,
    new_n62111_, new_n62112_, new_n62113_, new_n62114_, new_n62115_,
    new_n62116_, new_n62117_, new_n62118_, new_n62119_, new_n62120_,
    new_n62121_, new_n62122_, new_n62123_, new_n62124_, new_n62125_,
    new_n62126_, new_n62127_, new_n62128_, new_n62129_, new_n62130_,
    new_n62131_, new_n62132_, new_n62133_, new_n62134_, new_n62135_,
    new_n62136_, new_n62137_, new_n62138_, new_n62139_, new_n62140_,
    new_n62141_, new_n62142_, new_n62143_, new_n62144_, new_n62145_,
    new_n62146_, new_n62147_, new_n62148_, new_n62149_, new_n62150_,
    new_n62151_, new_n62152_, new_n62153_, new_n62154_, new_n62155_,
    new_n62156_, new_n62157_, new_n62158_, new_n62159_, new_n62160_,
    new_n62161_, new_n62162_, new_n62163_, new_n62164_, new_n62165_,
    new_n62166_, new_n62167_, new_n62168_, new_n62169_, new_n62170_,
    new_n62171_, new_n62172_, new_n62173_, new_n62174_, new_n62175_,
    new_n62176_, new_n62177_, new_n62178_, new_n62179_, new_n62180_,
    new_n62181_, new_n62182_, new_n62183_, new_n62184_, new_n62185_,
    new_n62186_, new_n62187_, new_n62188_, new_n62189_, new_n62190_,
    new_n62191_, new_n62192_, new_n62193_, new_n62194_, new_n62195_,
    new_n62196_, new_n62197_, new_n62198_, new_n62199_, new_n62200_,
    new_n62201_, new_n62202_, new_n62203_, new_n62204_, new_n62205_,
    new_n62206_, new_n62207_, new_n62208_, new_n62209_, new_n62210_,
    new_n62211_, new_n62212_, new_n62213_, new_n62214_, new_n62215_,
    new_n62216_, new_n62217_, new_n62218_, new_n62219_, new_n62220_,
    new_n62221_, new_n62222_, new_n62223_, new_n62224_, new_n62225_,
    new_n62226_, new_n62227_, new_n62228_, new_n62229_, new_n62230_,
    new_n62231_, new_n62232_, new_n62233_, new_n62234_, new_n62235_,
    new_n62236_, new_n62237_, new_n62238_, new_n62239_, new_n62240_,
    new_n62241_, new_n62242_, new_n62243_, new_n62244_, new_n62245_,
    new_n62246_, new_n62247_, new_n62248_, new_n62249_, new_n62250_,
    new_n62251_, new_n62252_, new_n62253_, new_n62254_, new_n62255_,
    new_n62256_, new_n62257_, new_n62258_, new_n62259_, new_n62260_,
    new_n62261_, new_n62262_, new_n62263_, new_n62264_, new_n62265_,
    new_n62266_, new_n62267_, new_n62268_, new_n62269_, new_n62270_,
    new_n62271_, new_n62272_, new_n62273_, new_n62274_, new_n62275_,
    new_n62276_, new_n62277_, new_n62278_, new_n62279_, new_n62280_,
    new_n62281_, new_n62282_, new_n62283_, new_n62284_, new_n62285_,
    new_n62286_, new_n62287_, new_n62288_, new_n62289_, new_n62290_,
    new_n62291_, new_n62292_, new_n62293_, new_n62294_, new_n62295_,
    new_n62296_, new_n62297_, new_n62298_, new_n62299_, new_n62300_,
    new_n62301_, new_n62302_, new_n62303_, new_n62304_, new_n62305_,
    new_n62306_, new_n62307_, new_n62308_, new_n62309_, new_n62310_,
    new_n62311_, new_n62312_, new_n62313_, new_n62314_, new_n62315_,
    new_n62316_, new_n62317_, new_n62318_, new_n62319_, new_n62320_,
    new_n62321_, new_n62322_, new_n62323_, new_n62324_, new_n62325_,
    new_n62326_, new_n62327_, new_n62328_, new_n62329_, new_n62330_,
    new_n62331_, new_n62332_, new_n62333_, new_n62334_, new_n62335_,
    new_n62336_, new_n62337_, new_n62338_, new_n62339_, new_n62340_,
    new_n62341_, new_n62342_, new_n62343_, new_n62344_, new_n62345_,
    new_n62346_, new_n62347_, new_n62348_, new_n62349_, new_n62350_,
    new_n62351_, new_n62352_, new_n62353_, new_n62354_, new_n62355_,
    new_n62356_, new_n62357_, new_n62358_, new_n62359_, new_n62360_,
    new_n62361_, new_n62362_, new_n62363_, new_n62364_, new_n62365_,
    new_n62366_, new_n62367_, new_n62368_, new_n62369_, new_n62370_,
    new_n62371_, new_n62372_, new_n62373_, new_n62374_, new_n62375_,
    new_n62376_, new_n62377_, new_n62378_, new_n62379_, new_n62380_,
    new_n62381_, new_n62382_, new_n62383_, new_n62384_, new_n62385_,
    new_n62386_, new_n62387_, new_n62388_, new_n62389_, new_n62390_,
    new_n62391_, new_n62392_, new_n62393_, new_n62394_, new_n62395_,
    new_n62396_, new_n62397_, new_n62398_, new_n62399_, new_n62400_,
    new_n62401_, new_n62402_, new_n62403_, new_n62404_, new_n62405_,
    new_n62406_, new_n62407_, new_n62408_, new_n62409_, new_n62410_,
    new_n62411_, new_n62412_, new_n62413_, new_n62414_, new_n62415_,
    new_n62416_, new_n62417_, new_n62418_, new_n62419_, new_n62420_,
    new_n62421_, new_n62422_, new_n62423_, new_n62424_, new_n62425_,
    new_n62426_, new_n62427_, new_n62428_, new_n62429_, new_n62430_,
    new_n62431_, new_n62432_, new_n62433_, new_n62434_, new_n62435_,
    new_n62436_, new_n62437_, new_n62438_, new_n62439_, new_n62440_,
    new_n62441_, new_n62442_, new_n62443_, new_n62444_, new_n62445_,
    new_n62446_, new_n62447_, new_n62448_, new_n62449_, new_n62450_,
    new_n62451_, new_n62452_, new_n62453_, new_n62454_, new_n62455_,
    new_n62456_, new_n62457_, new_n62458_, new_n62459_, new_n62460_,
    new_n62461_, new_n62462_, new_n62463_, new_n62464_, new_n62465_,
    new_n62466_, new_n62467_, new_n62468_, new_n62469_, new_n62470_,
    new_n62471_, new_n62472_, new_n62473_, new_n62474_, new_n62475_,
    new_n62476_, new_n62477_, new_n62478_, new_n62479_, new_n62480_,
    new_n62481_, new_n62482_, new_n62483_, new_n62484_, new_n62485_,
    new_n62486_, new_n62487_, new_n62488_, new_n62489_, new_n62490_,
    new_n62491_, new_n62492_, new_n62493_, new_n62494_, new_n62495_,
    new_n62496_, new_n62497_, new_n62498_, new_n62499_, new_n62500_,
    new_n62501_, new_n62502_, new_n62503_, new_n62504_, new_n62505_,
    new_n62506_, new_n62507_, new_n62508_, new_n62509_, new_n62510_,
    new_n62511_, new_n62512_, new_n62513_, new_n62514_, new_n62515_,
    new_n62516_, new_n62517_, new_n62518_, new_n62519_, new_n62520_,
    new_n62521_, new_n62522_, new_n62523_, new_n62524_, new_n62525_,
    new_n62526_, new_n62527_, new_n62528_, new_n62529_, new_n62530_,
    new_n62531_, new_n62532_, new_n62533_, new_n62534_, new_n62535_,
    new_n62536_, new_n62537_, new_n62538_, new_n62539_, new_n62540_,
    new_n62541_, new_n62542_, new_n62543_, new_n62544_, new_n62545_,
    new_n62546_, new_n62547_, new_n62548_, new_n62549_, new_n62550_,
    new_n62551_, new_n62552_, new_n62553_, new_n62554_, new_n62555_,
    new_n62556_, new_n62557_, new_n62558_, new_n62559_, new_n62560_,
    new_n62561_, new_n62562_, new_n62563_, new_n62564_, new_n62565_,
    new_n62566_, new_n62567_, new_n62568_, new_n62569_, new_n62570_,
    new_n62571_, new_n62572_, new_n62573_, new_n62574_, new_n62575_,
    new_n62576_, new_n62577_, new_n62578_, new_n62579_, new_n62580_,
    new_n62581_, new_n62582_, new_n62583_, new_n62584_, new_n62585_,
    new_n62586_, new_n62587_, new_n62588_, new_n62589_, new_n62590_,
    new_n62591_, new_n62592_, new_n62593_, new_n62594_, new_n62595_,
    new_n62596_, new_n62597_, new_n62598_, new_n62599_, new_n62600_,
    new_n62601_, new_n62602_, new_n62603_, new_n62604_, new_n62605_,
    new_n62606_, new_n62607_, new_n62608_, new_n62609_, new_n62610_,
    new_n62611_, new_n62612_, new_n62613_, new_n62614_, new_n62615_,
    new_n62616_, new_n62617_, new_n62618_, new_n62619_, new_n62620_,
    new_n62621_, new_n62622_, new_n62623_, new_n62624_, new_n62625_,
    new_n62626_, new_n62627_, new_n62628_, new_n62629_, new_n62630_,
    new_n62631_, new_n62632_, new_n62633_, new_n62634_, new_n62635_,
    new_n62636_, new_n62637_, new_n62638_, new_n62639_, new_n62640_,
    new_n62641_, new_n62642_, new_n62643_, new_n62644_, new_n62645_,
    new_n62646_, new_n62647_, new_n62648_, new_n62649_, new_n62650_,
    new_n62651_, new_n62652_, new_n62653_, new_n62654_, new_n62655_,
    new_n62656_, new_n62657_, new_n62658_, new_n62659_, new_n62660_,
    new_n62661_, new_n62662_, new_n62663_, new_n62664_, new_n62665_,
    new_n62666_, new_n62667_, new_n62668_, new_n62669_, new_n62670_,
    new_n62671_, new_n62672_, new_n62673_, new_n62674_, new_n62675_,
    new_n62676_, new_n62677_, new_n62678_, new_n62679_, new_n62680_,
    new_n62681_, new_n62682_, new_n62683_, new_n62684_, new_n62685_,
    new_n62686_, new_n62687_, new_n62688_, new_n62689_, new_n62690_,
    new_n62691_, new_n62692_, new_n62693_, new_n62694_, new_n62695_,
    new_n62696_, new_n62697_, new_n62698_, new_n62699_, new_n62700_,
    new_n62701_, new_n62702_, new_n62703_, new_n62704_, new_n62705_,
    new_n62706_, new_n62707_, new_n62708_, new_n62709_, new_n62710_,
    new_n62711_, new_n62712_, new_n62713_, new_n62714_, new_n62715_,
    new_n62716_, new_n62717_, new_n62718_, new_n62719_, new_n62720_,
    new_n62721_, new_n62722_, new_n62723_, new_n62724_, new_n62725_,
    new_n62726_, new_n62727_, new_n62728_, new_n62729_, new_n62730_,
    new_n62731_, new_n62732_, new_n62733_, new_n62734_, new_n62735_,
    new_n62736_, new_n62737_, new_n62738_, new_n62739_, new_n62740_,
    new_n62741_, new_n62742_, new_n62743_, new_n62744_, new_n62745_,
    new_n62746_, new_n62747_, new_n62748_, new_n62749_, new_n62750_,
    new_n62751_, new_n62752_, new_n62753_, new_n62754_, new_n62755_,
    new_n62756_, new_n62757_, new_n62758_, new_n62759_, new_n62760_,
    new_n62761_, new_n62762_, new_n62763_, new_n62764_, new_n62765_,
    new_n62766_, new_n62767_, new_n62768_, new_n62769_, new_n62770_,
    new_n62771_, new_n62772_, new_n62773_, new_n62774_, new_n62775_,
    new_n62776_, new_n62777_, new_n62778_, new_n62779_, new_n62780_,
    new_n62781_, new_n62782_, new_n62783_, new_n62784_, new_n62785_,
    new_n62786_, new_n62787_, new_n62788_, new_n62789_, new_n62790_,
    new_n62791_, new_n62792_, new_n62793_, new_n62794_, new_n62795_,
    new_n62796_, new_n62797_, new_n62798_, new_n62799_, new_n62800_,
    new_n62801_, new_n62802_, new_n62803_, new_n62804_, new_n62805_,
    new_n62806_, new_n62807_, new_n62808_, new_n62809_, new_n62810_,
    new_n62811_, new_n62812_, new_n62813_, new_n62814_, new_n62815_,
    new_n62816_, new_n62817_, new_n62818_, new_n62819_, new_n62820_,
    new_n62821_, new_n62822_, new_n62823_, new_n62824_, new_n62825_,
    new_n62826_, new_n62827_, new_n62828_, new_n62829_, new_n62830_,
    new_n62831_, new_n62832_, new_n62833_, new_n62834_, new_n62835_,
    new_n62836_, new_n62837_, new_n62838_, new_n62839_, new_n62840_,
    new_n62841_, new_n62842_, new_n62843_, new_n62844_, new_n62845_,
    new_n62846_, new_n62847_, new_n62848_, new_n62849_, new_n62850_,
    new_n62851_, new_n62852_, new_n62853_, new_n62854_, new_n62855_,
    new_n62856_, new_n62857_, new_n62858_, new_n62859_, new_n62860_,
    new_n62861_, new_n62862_, new_n62863_, new_n62864_, new_n62865_,
    new_n62866_, new_n62867_, new_n62868_, new_n62869_, new_n62870_,
    new_n62871_, new_n62872_, new_n62873_, new_n62874_, new_n62875_,
    new_n62876_, new_n62877_, new_n62878_, new_n62879_, new_n62880_,
    new_n62881_, new_n62882_, new_n62883_, new_n62884_, new_n62885_,
    new_n62886_, new_n62887_, new_n62888_, new_n62889_, new_n62890_,
    new_n62891_, new_n62892_, new_n62893_, new_n62894_, new_n62895_,
    new_n62896_, new_n62897_, new_n62898_, new_n62899_, new_n62900_,
    new_n62901_, new_n62902_, new_n62903_, new_n62904_, new_n62905_,
    new_n62906_, new_n62907_, new_n62908_, new_n62909_, new_n62910_,
    new_n62911_, new_n62912_, new_n62913_, new_n62914_, new_n62915_,
    new_n62916_, new_n62917_, new_n62918_, new_n62919_, new_n62920_,
    new_n62921_, new_n62922_, new_n62923_, new_n62924_, new_n62925_,
    new_n62926_, new_n62927_, new_n62928_, new_n62929_, new_n62930_,
    new_n62931_, new_n62932_, new_n62933_, new_n62934_, new_n62935_,
    new_n62936_, new_n62937_, new_n62938_, new_n62939_, new_n62940_,
    new_n62941_, new_n62942_, new_n62943_, new_n62944_, new_n62945_,
    new_n62946_, new_n62947_, new_n62948_, new_n62949_, new_n62950_,
    new_n62951_, new_n62952_, new_n62953_, new_n62954_, new_n62955_,
    new_n62956_, new_n62957_, new_n62958_, new_n62959_, new_n62960_,
    new_n62961_, new_n62962_, new_n62963_, new_n62964_, new_n62965_,
    new_n62966_, new_n62967_, new_n62968_, new_n62969_, new_n62970_,
    new_n62971_, new_n62972_, new_n62973_, new_n62974_, new_n62975_,
    new_n62976_, new_n62977_, new_n62978_, new_n62979_, new_n62980_,
    new_n62981_, new_n62982_, new_n62983_, new_n62984_, new_n62985_,
    new_n62986_, new_n62987_, new_n62988_, new_n62989_, new_n62990_,
    new_n62991_, new_n62992_, new_n62993_, new_n62994_, new_n62995_,
    new_n62996_, new_n62997_, new_n62998_, new_n62999_, new_n63000_,
    new_n63001_, new_n63002_, new_n63003_, new_n63004_, new_n63005_,
    new_n63006_, new_n63007_, new_n63008_, new_n63009_, new_n63010_,
    new_n63011_, new_n63012_, new_n63013_, new_n63014_, new_n63015_,
    new_n63016_, new_n63017_, new_n63018_, new_n63019_, new_n63020_,
    new_n63021_, new_n63022_, new_n63023_, new_n63024_, new_n63025_,
    new_n63026_, new_n63027_, new_n63028_, new_n63029_, new_n63030_,
    new_n63031_, new_n63032_, new_n63033_, new_n63034_, new_n63035_,
    new_n63036_, new_n63037_, new_n63038_, new_n63039_, new_n63040_,
    new_n63041_, new_n63042_, new_n63043_, new_n63044_, new_n63045_,
    new_n63046_, new_n63047_, new_n63048_, new_n63049_, new_n63050_,
    new_n63051_, new_n63052_, new_n63053_, new_n63054_, new_n63055_,
    new_n63056_, new_n63057_, new_n63058_, new_n63059_, new_n63060_,
    new_n63061_, new_n63062_, new_n63063_, new_n63064_, new_n63065_,
    new_n63066_, new_n63067_, new_n63068_, new_n63069_, new_n63070_,
    new_n63071_, new_n63072_, new_n63073_, new_n63074_, new_n63075_,
    new_n63076_, new_n63077_, new_n63078_, new_n63079_, new_n63080_,
    new_n63081_, new_n63082_, new_n63083_, new_n63084_, new_n63085_,
    new_n63086_, new_n63087_, new_n63088_, new_n63089_, new_n63090_,
    new_n63091_, new_n63092_, new_n63093_, new_n63094_, new_n63095_,
    new_n63096_, new_n63097_, new_n63098_, new_n63099_, new_n63100_,
    new_n63101_, new_n63102_, new_n63103_, new_n63104_, new_n63105_,
    new_n63106_, new_n63107_, new_n63108_, new_n63109_, new_n63110_,
    new_n63111_, new_n63112_, new_n63113_, new_n63114_, new_n63115_,
    new_n63116_, new_n63117_, new_n63118_, new_n63119_, new_n63120_,
    new_n63121_, new_n63122_, new_n63123_, new_n63124_, new_n63125_,
    new_n63126_, new_n63127_, new_n63128_, new_n63129_, new_n63130_,
    new_n63131_, new_n63132_, new_n63133_, new_n63134_, new_n63135_,
    new_n63136_, new_n63137_, new_n63138_, new_n63139_, new_n63140_,
    new_n63141_, new_n63142_, new_n63143_, new_n63144_, new_n63145_,
    new_n63146_, new_n63147_, new_n63148_, new_n63149_, new_n63150_,
    new_n63151_, new_n63152_, new_n63153_, new_n63154_, new_n63155_,
    new_n63156_, new_n63157_, new_n63158_, new_n63159_, new_n63160_,
    new_n63161_, new_n63162_, new_n63163_, new_n63164_, new_n63165_,
    new_n63166_, new_n63167_, new_n63168_, new_n63169_, new_n63170_,
    new_n63171_, new_n63172_, new_n63173_, new_n63174_, new_n63175_,
    new_n63176_, new_n63177_, new_n63178_, new_n63179_, new_n63180_,
    new_n63181_, new_n63182_, new_n63183_, new_n63184_, new_n63185_,
    new_n63186_, new_n63187_, new_n63188_, new_n63189_, new_n63190_,
    new_n63191_, new_n63192_, new_n63193_, new_n63194_, new_n63195_,
    new_n63196_, new_n63197_, new_n63198_, new_n63199_, new_n63200_,
    new_n63201_, new_n63202_, new_n63203_, new_n63204_, new_n63205_,
    new_n63206_, new_n63207_, new_n63208_, new_n63209_, new_n63210_,
    new_n63211_, new_n63212_, new_n63213_, new_n63214_, new_n63215_,
    new_n63216_, new_n63217_, new_n63218_, new_n63219_, new_n63220_,
    new_n63221_, new_n63222_, new_n63223_, new_n63224_, new_n63225_,
    new_n63226_, new_n63227_, new_n63228_, new_n63229_, new_n63230_,
    new_n63231_, new_n63232_, new_n63233_, new_n63234_, new_n63235_,
    new_n63236_, new_n63237_, new_n63238_, new_n63239_, new_n63240_,
    new_n63241_, new_n63242_, new_n63243_, new_n63244_, new_n63245_,
    new_n63246_, new_n63247_, new_n63248_, new_n63249_, new_n63250_,
    new_n63251_, new_n63252_, new_n63253_, new_n63254_, new_n63255_,
    new_n63256_, new_n63257_, new_n63258_, new_n63259_, new_n63260_,
    new_n63261_, new_n63262_, new_n63263_, new_n63264_, new_n63265_,
    new_n63266_, new_n63267_, new_n63268_, new_n63269_, new_n63270_,
    new_n63271_, new_n63272_, new_n63273_, new_n63274_, new_n63275_,
    new_n63276_, new_n63277_, new_n63278_, new_n63279_, new_n63280_,
    new_n63281_, new_n63282_, new_n63283_, new_n63284_, new_n63285_,
    new_n63286_, new_n63287_, new_n63288_, new_n63289_, new_n63290_,
    new_n63291_, new_n63292_, new_n63293_, new_n63294_, new_n63295_,
    new_n63296_, new_n63297_, new_n63298_, new_n63299_, new_n63300_,
    new_n63301_, new_n63302_, new_n63303_, new_n63304_, new_n63305_,
    new_n63306_, new_n63307_, new_n63308_, new_n63309_, new_n63310_,
    new_n63311_, new_n63312_, new_n63313_, new_n63314_, new_n63315_,
    new_n63316_, new_n63317_, new_n63318_, new_n63319_, new_n63320_,
    new_n63321_, new_n63322_, new_n63323_, new_n63324_, new_n63325_,
    new_n63326_, new_n63327_, new_n63328_, new_n63329_, new_n63330_,
    new_n63331_, new_n63332_, new_n63333_, new_n63334_, new_n63335_,
    new_n63336_, new_n63337_, new_n63338_, new_n63339_, new_n63340_,
    new_n63341_, new_n63342_, new_n63343_, new_n63344_, new_n63345_,
    new_n63346_, new_n63347_, new_n63348_, new_n63349_, new_n63350_,
    new_n63351_, new_n63352_, new_n63353_, new_n63354_, new_n63355_,
    new_n63356_, new_n63357_, new_n63358_, new_n63359_, new_n63360_,
    new_n63361_, new_n63362_, new_n63363_, new_n63364_, new_n63365_,
    new_n63366_, new_n63367_, new_n63368_, new_n63369_, new_n63370_,
    new_n63371_, new_n63372_, new_n63373_, new_n63374_, new_n63375_,
    new_n63376_, new_n63377_, new_n63378_, new_n63379_, new_n63380_,
    new_n63381_, new_n63382_, new_n63383_, new_n63384_, new_n63385_,
    new_n63386_, new_n63387_, new_n63388_, new_n63389_, new_n63390_,
    new_n63391_, new_n63392_, new_n63393_, new_n63394_, new_n63395_,
    new_n63396_, new_n63397_, new_n63398_, new_n63399_, new_n63400_,
    new_n63401_, new_n63402_, new_n63403_, new_n63404_, new_n63405_,
    new_n63406_, new_n63407_, new_n63408_, new_n63409_, new_n63410_,
    new_n63411_, new_n63412_, new_n63413_, new_n63414_, new_n63415_,
    new_n63416_, new_n63417_, new_n63418_, new_n63419_, new_n63420_,
    new_n63421_, new_n63422_, new_n63423_, new_n63424_, new_n63425_,
    new_n63426_, new_n63427_, new_n63428_, new_n63429_, new_n63430_,
    new_n63431_, new_n63432_, new_n63433_, new_n63434_, new_n63435_,
    new_n63436_, new_n63437_, new_n63438_, new_n63439_, new_n63440_,
    new_n63441_, new_n63442_, new_n63443_, new_n63444_, new_n63445_,
    new_n63446_, new_n63447_, new_n63448_, new_n63449_, new_n63450_,
    new_n63451_, new_n63452_, new_n63453_, new_n63454_, new_n63455_,
    new_n63456_, new_n63457_, new_n63458_, new_n63459_, new_n63460_,
    new_n63461_, new_n63462_, new_n63463_, new_n63464_, new_n63465_,
    new_n63466_, new_n63467_, new_n63468_, new_n63469_, new_n63470_,
    new_n63471_, new_n63472_, new_n63473_, new_n63474_, new_n63475_,
    new_n63476_, new_n63477_, new_n63478_, new_n63479_, new_n63480_,
    new_n63481_, new_n63482_, new_n63483_, new_n63484_, new_n63485_,
    new_n63486_, new_n63487_, new_n63488_, new_n63489_, new_n63490_,
    new_n63491_, new_n63492_, new_n63493_, new_n63494_, new_n63495_,
    new_n63496_, new_n63497_, new_n63498_, new_n63499_, new_n63500_,
    new_n63501_, new_n63502_, new_n63503_, new_n63504_, new_n63505_,
    new_n63506_, new_n63507_, new_n63508_, new_n63509_, new_n63510_,
    new_n63511_, new_n63512_, new_n63513_, new_n63514_, new_n63515_,
    new_n63516_, new_n63517_, new_n63518_, new_n63519_, new_n63520_,
    new_n63521_, new_n63522_, new_n63523_, new_n63524_, new_n63525_,
    new_n63526_, new_n63527_, new_n63528_, new_n63529_, new_n63530_,
    new_n63531_, new_n63532_, new_n63533_, new_n63534_, new_n63535_,
    new_n63536_, new_n63537_, new_n63538_, new_n63539_, new_n63540_,
    new_n63541_, new_n63542_, new_n63543_, new_n63544_, new_n63545_,
    new_n63546_, new_n63547_, new_n63548_, new_n63549_, new_n63550_,
    new_n63551_, new_n63552_, new_n63553_, new_n63554_, new_n63555_,
    new_n63556_, new_n63557_, new_n63558_, new_n63559_, new_n63560_,
    new_n63561_, new_n63562_, new_n63563_, new_n63564_, new_n63565_,
    new_n63566_, new_n63567_, new_n63568_, new_n63569_, new_n63570_,
    new_n63571_, new_n63572_, new_n63573_, new_n63574_, new_n63575_,
    new_n63576_, new_n63577_, new_n63578_, new_n63579_, new_n63580_,
    new_n63581_, new_n63582_, new_n63583_, new_n63584_, new_n63585_,
    new_n63586_, new_n63587_, new_n63588_, new_n63589_, new_n63590_,
    new_n63591_, new_n63592_, new_n63593_, new_n63594_, new_n63595_,
    new_n63596_, new_n63597_, new_n63598_, new_n63599_, new_n63600_,
    new_n63601_, new_n63602_, new_n63603_, new_n63604_, new_n63605_,
    new_n63606_, new_n63607_, new_n63608_, new_n63609_, new_n63610_,
    new_n63611_, new_n63612_, new_n63613_, new_n63614_, new_n63615_,
    new_n63616_, new_n63617_, new_n63618_, new_n63619_, new_n63620_,
    new_n63621_, new_n63622_, new_n63623_, new_n63624_, new_n63625_,
    new_n63626_, new_n63627_, new_n63628_, new_n63629_, new_n63630_,
    new_n63631_, new_n63632_, new_n63633_, new_n63634_, new_n63635_,
    new_n63636_, new_n63637_, new_n63638_, new_n63639_, new_n63640_,
    new_n63641_, new_n63642_, new_n63643_, new_n63644_, new_n63645_,
    new_n63646_, new_n63647_, new_n63648_, new_n63649_, new_n63650_,
    new_n63651_, new_n63652_, new_n63653_, new_n63654_, new_n63655_,
    new_n63656_, new_n63657_, new_n63658_, new_n63659_, new_n63660_,
    new_n63661_, new_n63662_, new_n63663_, new_n63664_, new_n63665_,
    new_n63666_, new_n63667_, new_n63668_, new_n63669_, new_n63670_,
    new_n63671_, new_n63672_, new_n63673_, new_n63674_, new_n63675_,
    new_n63676_, new_n63677_, new_n63678_, new_n63679_, new_n63680_,
    new_n63681_, new_n63682_, new_n63683_, new_n63684_, new_n63685_,
    new_n63686_, new_n63687_, new_n63688_, new_n63689_, new_n63690_,
    new_n63691_, new_n63692_, new_n63693_, new_n63694_, new_n63695_,
    new_n63696_, new_n63697_, new_n63698_, new_n63699_, new_n63700_,
    new_n63701_, new_n63702_, new_n63703_, new_n63704_, new_n63705_,
    new_n63706_, new_n63707_, new_n63708_, new_n63709_, new_n63710_,
    new_n63711_, new_n63712_, new_n63713_, new_n63714_, new_n63715_,
    new_n63716_, new_n63717_, new_n63718_, new_n63719_, new_n63720_,
    new_n63721_, new_n63722_, new_n63723_, new_n63724_, new_n63725_,
    new_n63726_, new_n63727_, new_n63728_, new_n63729_, new_n63730_,
    new_n63731_, new_n63732_, new_n63733_, new_n63734_, new_n63735_,
    new_n63736_, new_n63737_, new_n63738_, new_n63739_, new_n63740_,
    new_n63741_, new_n63742_, new_n63743_, new_n63744_, new_n63745_,
    new_n63746_, new_n63747_, new_n63748_, new_n63749_, new_n63750_,
    new_n63751_, new_n63752_, new_n63753_, new_n63754_, new_n63755_,
    new_n63756_, new_n63757_, new_n63758_, new_n63759_, new_n63760_,
    new_n63761_, new_n63762_, new_n63763_, new_n63764_, new_n63765_,
    new_n63766_, new_n63767_, new_n63768_, new_n63769_, new_n63770_,
    new_n63771_, new_n63772_, new_n63773_, new_n63774_, new_n63775_,
    new_n63776_, new_n63777_, new_n63778_, new_n63779_, new_n63780_,
    new_n63781_, new_n63782_, new_n63783_, new_n63784_, new_n63785_,
    new_n63786_, new_n63787_, new_n63788_, new_n63789_, new_n63790_,
    new_n63791_, new_n63792_, new_n63793_, new_n63794_, new_n63795_,
    new_n63796_, new_n63797_, new_n63798_, new_n63799_, new_n63800_,
    new_n63801_, new_n63802_, new_n63803_, new_n63804_, new_n63805_,
    new_n63806_, new_n63807_, new_n63808_, new_n63809_, new_n63810_,
    new_n63811_, new_n63812_, new_n63813_, new_n63814_, new_n63815_,
    new_n63816_, new_n63817_, new_n63818_, new_n63819_, new_n63820_,
    new_n63821_, new_n63822_, new_n63823_, new_n63824_, new_n63825_,
    new_n63826_, new_n63827_, new_n63828_, new_n63829_, new_n63830_,
    new_n63831_, new_n63832_, new_n63833_, new_n63834_, new_n63835_,
    new_n63836_, new_n63837_, new_n63838_, new_n63839_, new_n63840_,
    new_n63841_, new_n63842_, new_n63843_, new_n63844_, new_n63845_,
    new_n63846_, new_n63847_, new_n63848_, new_n63849_, new_n63850_,
    new_n63851_, new_n63852_, new_n63853_, new_n63854_, new_n63855_,
    new_n63856_, new_n63857_, new_n63858_, new_n63859_, new_n63860_,
    new_n63861_, new_n63862_, new_n63863_, new_n63864_, new_n63865_,
    new_n63866_, new_n63867_, new_n63868_, new_n63869_, new_n63870_,
    new_n63871_, new_n63872_, new_n63873_, new_n63874_, new_n63875_,
    new_n63876_, new_n63877_, new_n63878_, new_n63879_, new_n63880_,
    new_n63881_, new_n63882_, new_n63883_, new_n63884_, new_n63885_,
    new_n63886_, new_n63887_, new_n63888_, new_n63889_, new_n63890_,
    new_n63891_, new_n63892_, new_n63893_, new_n63894_, new_n63895_,
    new_n63896_, new_n63897_, new_n63898_, new_n63899_, new_n63900_,
    new_n63901_, new_n63902_, new_n63903_, new_n63904_, new_n63905_,
    new_n63906_, new_n63907_, new_n63908_, new_n63909_, new_n63910_,
    new_n63911_, new_n63912_, new_n63913_, new_n63914_, new_n63915_,
    new_n63916_, new_n63917_, new_n63918_, new_n63919_, new_n63920_,
    new_n63921_, new_n63922_, new_n63923_, new_n63924_, new_n63925_,
    new_n63926_, new_n63927_, new_n63928_, new_n63929_, new_n63930_,
    new_n63931_, new_n63932_, new_n63933_, new_n63934_, new_n63935_,
    new_n63936_, new_n63937_, new_n63938_, new_n63939_, new_n63940_,
    new_n63941_, new_n63942_, new_n63943_, new_n63944_, new_n63945_,
    new_n63946_, new_n63947_, new_n63948_, new_n63949_, new_n63950_,
    new_n63951_, new_n63952_, new_n63953_, new_n63954_, new_n63955_,
    new_n63956_, new_n63957_, new_n63958_, new_n63959_, new_n63960_,
    new_n63961_, new_n63962_, new_n63963_, new_n63964_, new_n63965_,
    new_n63966_, new_n63967_, new_n63968_, new_n63969_, new_n63970_,
    new_n63971_, new_n63972_, new_n63973_, new_n63974_, new_n63975_,
    new_n63976_, new_n63977_, new_n63978_, new_n63979_, new_n63980_,
    new_n63981_, new_n63982_, new_n63983_, new_n63984_, new_n63985_,
    new_n63986_, new_n63987_, new_n63988_, new_n63989_, new_n63990_,
    new_n63991_, new_n63992_, new_n63993_, new_n63994_, new_n63995_,
    new_n63996_, new_n63997_, new_n63998_, new_n63999_, new_n64000_,
    new_n64001_, new_n64002_, new_n64003_, new_n64004_, new_n64005_,
    new_n64006_, new_n64007_, new_n64008_, new_n64009_, new_n64010_,
    new_n64011_, new_n64012_, new_n64013_, new_n64014_, new_n64015_,
    new_n64016_, new_n64017_, new_n64018_, new_n64019_, new_n64020_,
    new_n64021_, new_n64022_, new_n64023_, new_n64024_, new_n64025_,
    new_n64026_, new_n64027_, new_n64028_, new_n64029_, new_n64030_,
    new_n64031_, new_n64032_, new_n64033_, new_n64034_, new_n64035_,
    new_n64036_, new_n64037_, new_n64038_, new_n64039_, new_n64040_,
    new_n64041_, new_n64042_, new_n64043_, new_n64044_, new_n64045_,
    new_n64046_, new_n64047_, new_n64048_, new_n64049_, new_n64050_,
    new_n64051_, new_n64052_, new_n64053_, new_n64054_, new_n64055_,
    new_n64056_, new_n64057_, new_n64058_, new_n64059_, new_n64060_,
    new_n64061_, new_n64062_, new_n64063_, new_n64064_, new_n64065_,
    new_n64066_, new_n64067_, new_n64068_, new_n64069_, new_n64070_,
    new_n64071_, new_n64072_, new_n64073_, new_n64074_, new_n64075_,
    new_n64076_, new_n64077_, new_n64078_, new_n64079_, new_n64080_,
    new_n64081_, new_n64082_, new_n64083_, new_n64084_, new_n64085_,
    new_n64086_, new_n64087_, new_n64088_, new_n64089_, new_n64090_,
    new_n64091_, new_n64092_, new_n64093_, new_n64094_, new_n64095_,
    new_n64096_, new_n64097_, new_n64098_, new_n64099_, new_n64100_,
    new_n64101_, new_n64102_, new_n64103_, new_n64104_, new_n64105_,
    new_n64106_, new_n64107_, new_n64108_, new_n64109_, new_n64110_,
    new_n64111_, new_n64112_, new_n64113_, new_n64114_, new_n64115_,
    new_n64116_, new_n64117_, new_n64118_, new_n64119_, new_n64120_,
    new_n64121_, new_n64122_, new_n64123_, new_n64124_, new_n64125_,
    new_n64126_, new_n64127_, new_n64128_, new_n64129_, new_n64130_,
    new_n64131_, new_n64132_, new_n64133_, new_n64134_, new_n64135_,
    new_n64136_, new_n64137_, new_n64138_, new_n64139_, new_n64140_,
    new_n64141_, new_n64142_, new_n64143_, new_n64144_, new_n64145_,
    new_n64146_, new_n64147_, new_n64148_, new_n64149_, new_n64150_,
    new_n64151_, new_n64152_, new_n64153_, new_n64154_, new_n64155_,
    new_n64156_, new_n64157_, new_n64158_, new_n64159_, new_n64160_,
    new_n64161_, new_n64162_, new_n64163_, new_n64164_, new_n64165_,
    new_n64166_, new_n64167_, new_n64168_, new_n64169_, new_n64170_,
    new_n64171_, new_n64172_, new_n64173_, new_n64174_, new_n64175_,
    new_n64176_, new_n64177_, new_n64178_, new_n64179_, new_n64180_,
    new_n64181_, new_n64182_, new_n64183_, new_n64184_, new_n64185_,
    new_n64186_, new_n64187_, new_n64188_, new_n64189_, new_n64190_,
    new_n64191_, new_n64192_, new_n64193_, new_n64194_, new_n64195_,
    new_n64196_, new_n64197_, new_n64198_, new_n64199_, new_n64200_,
    new_n64201_, new_n64202_, new_n64203_, new_n64204_, new_n64205_,
    new_n64206_, new_n64207_, new_n64208_, new_n64209_, new_n64210_,
    new_n64211_, new_n64212_, new_n64213_, new_n64214_, new_n64215_,
    new_n64216_, new_n64217_, new_n64218_, new_n64219_, new_n64220_,
    new_n64221_, new_n64222_, new_n64223_, new_n64224_, new_n64225_,
    new_n64226_, new_n64227_, new_n64228_, new_n64229_, new_n64230_,
    new_n64231_, new_n64232_, new_n64233_, new_n64234_, new_n64235_,
    new_n64236_, new_n64237_, new_n64238_, new_n64239_, new_n64240_,
    new_n64241_, new_n64242_, new_n64243_, new_n64244_, new_n64245_,
    new_n64246_, new_n64247_, new_n64248_, new_n64249_, new_n64250_,
    new_n64251_, new_n64252_, new_n64253_, new_n64254_, new_n64255_,
    new_n64256_, new_n64257_, new_n64258_, new_n64259_, new_n64260_,
    new_n64261_, new_n64262_, new_n64263_, new_n64264_, new_n64265_,
    new_n64266_, new_n64267_, new_n64268_, new_n64269_, new_n64270_,
    new_n64271_, new_n64272_, new_n64273_, new_n64274_, new_n64275_,
    new_n64276_, new_n64277_, new_n64278_, new_n64279_, new_n64280_,
    new_n64281_, new_n64282_, new_n64283_, new_n64284_, new_n64285_,
    new_n64286_, new_n64287_, new_n64288_, new_n64289_, new_n64290_,
    new_n64291_, new_n64292_, new_n64293_, new_n64294_, new_n64295_,
    new_n64296_, new_n64297_, new_n64298_, new_n64299_, new_n64300_,
    new_n64301_, new_n64302_, new_n64303_, new_n64304_, new_n64305_,
    new_n64306_, new_n64307_, new_n64308_, new_n64309_, new_n64310_,
    new_n64311_, new_n64312_, new_n64313_, new_n64314_, new_n64315_,
    new_n64316_, new_n64317_, new_n64318_, new_n64319_, new_n64320_,
    new_n64321_, new_n64322_, new_n64323_, new_n64324_, new_n64325_,
    new_n64326_, new_n64327_, new_n64328_, new_n64329_, new_n64330_,
    new_n64331_, new_n64332_, new_n64333_, new_n64334_, new_n64335_,
    new_n64336_, new_n64337_, new_n64338_, new_n64339_, new_n64340_,
    new_n64341_, new_n64342_, new_n64343_, new_n64344_, new_n64345_,
    new_n64346_, new_n64347_, new_n64348_, new_n64349_, new_n64350_,
    new_n64351_, new_n64352_, new_n64353_, new_n64354_, new_n64355_,
    new_n64356_, new_n64357_, new_n64358_, new_n64359_, new_n64360_,
    new_n64361_, new_n64362_, new_n64363_, new_n64364_, new_n64365_,
    new_n64366_, new_n64367_, new_n64368_, new_n64369_, new_n64370_,
    new_n64371_, new_n64372_, new_n64373_, new_n64374_, new_n64375_,
    new_n64376_, new_n64377_, new_n64378_, new_n64379_, new_n64380_,
    new_n64381_, new_n64382_, new_n64383_, new_n64384_, new_n64385_,
    new_n64386_, new_n64387_, new_n64388_, new_n64389_, new_n64390_,
    new_n64391_, new_n64392_, new_n64393_, new_n64394_, new_n64395_,
    new_n64396_, new_n64397_, new_n64398_, new_n64399_, new_n64400_,
    new_n64401_, new_n64402_, new_n64403_, new_n64404_, new_n64405_,
    new_n64406_, new_n64407_, new_n64408_, new_n64409_, new_n64410_,
    new_n64411_, new_n64412_, new_n64413_, new_n64414_, new_n64415_,
    new_n64416_, new_n64417_, new_n64418_, new_n64419_, new_n64420_,
    new_n64421_, new_n64422_, new_n64423_, new_n64424_, new_n64425_,
    new_n64426_, new_n64427_, new_n64428_, new_n64429_, new_n64430_,
    new_n64431_, new_n64432_, new_n64433_, new_n64434_, new_n64435_,
    new_n64436_, new_n64437_, new_n64438_, new_n64439_, new_n64440_,
    new_n64441_, new_n64442_, new_n64443_, new_n64444_, new_n64445_,
    new_n64446_, new_n64447_, new_n64448_, new_n64449_, new_n64450_,
    new_n64451_, new_n64452_, new_n64453_, new_n64454_, new_n64455_,
    new_n64456_, new_n64457_, new_n64458_, new_n64459_, new_n64460_,
    new_n64461_, new_n64462_, new_n64463_, new_n64464_, new_n64465_,
    new_n64466_, new_n64467_, new_n64468_, new_n64469_, new_n64470_,
    new_n64471_, new_n64472_, new_n64473_, new_n64474_, new_n64475_,
    new_n64476_, new_n64477_, new_n64478_, new_n64479_, new_n64480_,
    new_n64481_, new_n64482_, new_n64483_, new_n64484_, new_n64485_,
    new_n64486_, new_n64487_, new_n64488_, new_n64489_, new_n64490_,
    new_n64491_, new_n64492_, new_n64493_, new_n64494_, new_n64495_,
    new_n64496_, new_n64497_, new_n64498_, new_n64499_, new_n64500_,
    new_n64501_, new_n64502_, new_n64503_, new_n64504_, new_n64505_,
    new_n64506_, new_n64507_, new_n64508_, new_n64509_, new_n64510_,
    new_n64511_, new_n64512_, new_n64513_, new_n64514_, new_n64515_,
    new_n64516_, new_n64517_, new_n64518_, new_n64519_, new_n64520_,
    new_n64521_, new_n64522_, new_n64523_, new_n64524_, new_n64525_,
    new_n64526_, new_n64527_, new_n64528_, new_n64529_, new_n64530_,
    new_n64531_, new_n64532_, new_n64533_, new_n64534_, new_n64535_,
    new_n64536_, new_n64537_, new_n64538_, new_n64539_, new_n64540_,
    new_n64541_, new_n64542_, new_n64543_, new_n64544_, new_n64545_,
    new_n64546_, new_n64547_, new_n64548_, new_n64549_, new_n64550_,
    new_n64551_, new_n64552_, new_n64553_, new_n64554_, new_n64555_,
    new_n64556_, new_n64557_, new_n64558_, new_n64559_, new_n64560_,
    new_n64561_, new_n64562_, new_n64563_, new_n64564_, new_n64565_,
    new_n64566_, new_n64567_, new_n64568_, new_n64569_, new_n64570_,
    new_n64571_, new_n64572_, new_n64573_, new_n64574_, new_n64575_,
    new_n64576_, new_n64577_, new_n64578_, new_n64579_, new_n64580_,
    new_n64581_, new_n64582_, new_n64583_, new_n64584_, new_n64585_,
    new_n64586_, new_n64587_, new_n64588_, new_n64589_, new_n64590_,
    new_n64591_, new_n64592_, new_n64593_, new_n64594_, new_n64595_,
    new_n64596_, new_n64597_, new_n64598_, new_n64599_, new_n64600_,
    new_n64601_, new_n64602_, new_n64603_, new_n64604_, new_n64605_,
    new_n64606_, new_n64607_, new_n64608_, new_n64609_, new_n64610_,
    new_n64611_, new_n64612_, new_n64613_, new_n64614_, new_n64615_,
    new_n64616_, new_n64617_, new_n64618_, new_n64619_, new_n64620_,
    new_n64621_, new_n64622_, new_n64623_, new_n64624_, new_n64625_,
    new_n64626_, new_n64627_, new_n64628_, new_n64629_, new_n64630_,
    new_n64631_, new_n64632_, new_n64633_, new_n64634_, new_n64635_,
    new_n64636_, new_n64637_, new_n64638_, new_n64639_, new_n64640_,
    new_n64641_, new_n64642_, new_n64643_, new_n64644_, new_n64645_,
    new_n64646_, new_n64647_, new_n64648_, new_n64649_, new_n64650_,
    new_n64651_, new_n64652_, new_n64653_, new_n64654_, new_n64655_,
    new_n64656_, new_n64657_, new_n64658_, new_n64659_, new_n64660_,
    new_n64661_, new_n64662_, new_n64663_, new_n64664_, new_n64665_,
    new_n64666_, new_n64667_, new_n64668_, new_n64669_, new_n64670_,
    new_n64671_, new_n64672_, new_n64673_, new_n64674_, new_n64675_,
    new_n64676_, new_n64677_, new_n64678_, new_n64679_, new_n64680_,
    new_n64681_, new_n64682_, new_n64683_, new_n64684_, new_n64685_,
    new_n64686_, new_n64687_, new_n64688_, new_n64689_, new_n64690_,
    new_n64691_, new_n64692_, new_n64693_, new_n64694_, new_n64695_,
    new_n64696_, new_n64697_, new_n64698_, new_n64699_, new_n64700_,
    new_n64701_, new_n64702_, new_n64703_, new_n64704_, new_n64705_,
    new_n64706_, new_n64707_, new_n64708_, new_n64709_, new_n64710_,
    new_n64711_, new_n64712_, new_n64713_, new_n64714_, new_n64715_,
    new_n64716_, new_n64717_, new_n64718_, new_n64719_, new_n64720_,
    new_n64721_, new_n64722_, new_n64723_, new_n64724_, new_n64725_,
    new_n64726_, new_n64727_, new_n64728_, new_n64729_, new_n64730_,
    new_n64731_, new_n64732_, new_n64733_, new_n64734_, new_n64735_,
    new_n64736_, new_n64737_, new_n64738_, new_n64739_, new_n64740_,
    new_n64741_, new_n64742_, new_n64743_, new_n64744_, new_n64745_,
    new_n64746_, new_n64747_, new_n64748_, new_n64749_, new_n64750_,
    new_n64751_, new_n64752_, new_n64753_, new_n64754_, new_n64755_,
    new_n64756_, new_n64757_, new_n64758_, new_n64759_, new_n64760_,
    new_n64761_, new_n64762_, new_n64763_, new_n64764_, new_n64765_,
    new_n64766_, new_n64767_, new_n64768_, new_n64769_, new_n64770_,
    new_n64771_, new_n64772_, new_n64773_, new_n64774_, new_n64775_,
    new_n64776_, new_n64777_, new_n64778_, new_n64779_, new_n64780_,
    new_n64781_, new_n64782_, new_n64783_, new_n64784_, new_n64785_,
    new_n64786_, new_n64787_, new_n64788_, new_n64789_, new_n64790_,
    new_n64791_, new_n64792_, new_n64793_, new_n64794_, new_n64795_,
    new_n64796_, new_n64797_, new_n64798_, new_n64799_, new_n64800_,
    new_n64801_, new_n64802_, new_n64803_, new_n64804_, new_n64805_,
    new_n64806_, new_n64807_, new_n64808_, new_n64809_, new_n64810_,
    new_n64811_, new_n64812_, new_n64813_, new_n64814_, new_n64815_,
    new_n64816_, new_n64817_, new_n64818_, new_n64819_, new_n64820_,
    new_n64821_, new_n64822_, new_n64823_, new_n64824_, new_n64825_,
    new_n64826_, new_n64827_, new_n64828_, new_n64829_, new_n64830_,
    new_n64831_, new_n64832_, new_n64833_, new_n64834_, new_n64835_,
    new_n64836_, new_n64837_, new_n64838_, new_n64839_, new_n64840_,
    new_n64841_, new_n64842_, new_n64843_, new_n64844_, new_n64845_,
    new_n64846_, new_n64847_, new_n64848_, new_n64849_, new_n64850_,
    new_n64851_, new_n64852_, new_n64853_, new_n64854_, new_n64855_,
    new_n64856_, new_n64857_, new_n64858_, new_n64859_, new_n64860_,
    new_n64861_, new_n64862_, new_n64863_, new_n64864_, new_n64865_,
    new_n64866_, new_n64867_, new_n64868_, new_n64869_, new_n64870_,
    new_n64871_, new_n64872_, new_n64873_, new_n64874_, new_n64875_,
    new_n64876_, new_n64877_, new_n64878_, new_n64879_, new_n64880_,
    new_n64881_, new_n64882_, new_n64883_, new_n64884_, new_n64885_,
    new_n64886_, new_n64887_, new_n64888_, new_n64889_, new_n64890_,
    new_n64891_, new_n64892_, new_n64893_, new_n64894_, new_n64895_,
    new_n64896_, new_n64897_, new_n64898_, new_n64899_, new_n64900_,
    new_n64901_, new_n64902_, new_n64903_, new_n64904_, new_n64905_,
    new_n64906_, new_n64907_, new_n64908_, new_n64909_, new_n64910_,
    new_n64911_, new_n64912_, new_n64913_, new_n64914_, new_n64915_,
    new_n64916_, new_n64917_, new_n64918_, new_n64919_, new_n64920_,
    new_n64921_, new_n64922_, new_n64923_, new_n64924_, new_n64925_,
    new_n64926_, new_n64927_, new_n64928_, new_n64929_, new_n64930_,
    new_n64931_, new_n64932_, new_n64933_, new_n64934_, new_n64935_,
    new_n64936_, new_n64937_, new_n64938_, new_n64939_, new_n64940_,
    new_n64941_, new_n64942_, new_n64943_, new_n64944_, new_n64945_,
    new_n64946_, new_n64947_, new_n64948_, new_n64949_, new_n64950_,
    new_n64951_, new_n64952_, new_n64953_, new_n64954_, new_n64955_,
    new_n64956_, new_n64957_, new_n64958_, new_n64959_, new_n64960_,
    new_n64961_, new_n64962_, new_n64963_, new_n64964_, new_n64965_,
    new_n64966_, new_n64967_, new_n64968_, new_n64969_, new_n64970_,
    new_n64971_, new_n64972_, new_n64973_, new_n64974_, new_n64975_,
    new_n64976_, new_n64977_, new_n64978_, new_n64979_, new_n64980_,
    new_n64981_, new_n64982_, new_n64983_, new_n64984_, new_n64985_,
    new_n64986_, new_n64987_, new_n64988_, new_n64989_, new_n64990_,
    new_n64991_, new_n64992_, new_n64993_, new_n64994_, new_n64995_,
    new_n64996_, new_n64997_, new_n64998_, new_n64999_, new_n65000_,
    new_n65001_, new_n65002_, new_n65003_, new_n65004_, new_n65005_,
    new_n65006_, new_n65007_, new_n65008_, new_n65009_, new_n65010_,
    new_n65011_, new_n65012_, new_n65013_, new_n65014_, new_n65015_,
    new_n65016_, new_n65017_, new_n65018_, new_n65019_, new_n65020_,
    new_n65021_, new_n65022_, new_n65023_, new_n65024_, new_n65025_,
    new_n65026_, new_n65027_, new_n65028_, new_n65029_, new_n65030_,
    new_n65031_, new_n65032_, new_n65033_, new_n65034_, new_n65035_,
    new_n65036_, new_n65037_, new_n65038_, new_n65039_, new_n65040_,
    new_n65041_, new_n65042_, new_n65043_, new_n65044_, new_n65045_,
    new_n65046_, new_n65047_, new_n65048_, new_n65049_, new_n65050_,
    new_n65051_, new_n65052_, new_n65053_, new_n65054_, new_n65055_,
    new_n65056_, new_n65057_, new_n65058_, new_n65059_, new_n65060_,
    new_n65061_, new_n65062_, new_n65063_, new_n65064_, new_n65065_,
    new_n65066_, new_n65067_, new_n65068_, new_n65069_, new_n65070_,
    new_n65071_, new_n65072_, new_n65073_, new_n65074_, new_n65075_,
    new_n65076_, new_n65077_, new_n65078_, new_n65079_, new_n65080_,
    new_n65081_, new_n65082_, new_n65083_, new_n65084_, new_n65085_,
    new_n65086_, new_n65087_, new_n65088_, new_n65089_, new_n65090_,
    new_n65091_, new_n65092_, new_n65093_, new_n65094_, new_n65095_,
    new_n65096_, new_n65097_, new_n65098_, new_n65099_, new_n65100_,
    new_n65101_, new_n65102_, new_n65103_, new_n65104_, new_n65105_,
    new_n65106_, new_n65107_, new_n65108_, new_n65109_, new_n65110_,
    new_n65111_, new_n65112_, new_n65113_, new_n65114_, new_n65115_,
    new_n65116_, new_n65117_, new_n65118_, new_n65119_, new_n65120_,
    new_n65121_, new_n65122_, new_n65123_, new_n65124_, new_n65125_,
    new_n65126_, new_n65127_, new_n65128_, new_n65129_, new_n65130_,
    new_n65131_, new_n65132_, new_n65133_, new_n65134_, new_n65135_,
    new_n65136_, new_n65137_, new_n65138_, new_n65139_, new_n65140_,
    new_n65141_, new_n65142_, new_n65143_, new_n65144_, new_n65145_,
    new_n65146_, new_n65147_, new_n65148_, new_n65149_, new_n65150_,
    new_n65151_, new_n65152_, new_n65153_, new_n65154_, new_n65155_,
    new_n65156_, new_n65157_, new_n65158_, new_n65159_, new_n65160_,
    new_n65161_, new_n65162_, new_n65163_, new_n65164_, new_n65165_,
    new_n65166_, new_n65167_, new_n65168_, new_n65169_, new_n65170_,
    new_n65171_, new_n65172_, new_n65173_, new_n65174_, new_n65175_,
    new_n65176_, new_n65177_, new_n65178_, new_n65179_, new_n65180_,
    new_n65181_, new_n65182_, new_n65183_, new_n65184_, new_n65185_,
    new_n65186_, new_n65187_, new_n65188_, new_n65189_, new_n65190_,
    new_n65191_, new_n65192_, new_n65193_, new_n65194_, new_n65195_,
    new_n65196_, new_n65197_, new_n65198_, new_n65199_, new_n65200_,
    new_n65201_, new_n65202_, new_n65203_, new_n65204_, new_n65205_,
    new_n65206_, new_n65207_, new_n65208_, new_n65209_, new_n65210_,
    new_n65211_, new_n65212_, new_n65213_, new_n65214_, new_n65215_,
    new_n65216_, new_n65217_, new_n65218_, new_n65219_, new_n65220_,
    new_n65221_, new_n65222_, new_n65223_, new_n65224_, new_n65225_,
    new_n65226_, new_n65227_, new_n65228_, new_n65229_, new_n65230_,
    new_n65231_, new_n65232_, new_n65233_, new_n65234_, new_n65235_,
    new_n65236_, new_n65237_, new_n65238_, new_n65239_, new_n65240_,
    new_n65241_, new_n65242_, new_n65243_, new_n65244_, new_n65245_,
    new_n65246_, new_n65247_, new_n65248_, new_n65249_, new_n65250_,
    new_n65251_, new_n65252_, new_n65253_, new_n65254_, new_n65255_,
    new_n65256_, new_n65257_, new_n65258_, new_n65259_, new_n65260_,
    new_n65261_, new_n65262_, new_n65263_, new_n65264_, new_n65265_,
    new_n65266_, new_n65267_, new_n65268_, new_n65269_, new_n65270_,
    new_n65271_, new_n65272_, new_n65273_, new_n65274_, new_n65275_,
    new_n65276_, new_n65277_, new_n65278_, new_n65279_, new_n65280_,
    new_n65281_, new_n65282_, new_n65283_, new_n65284_, new_n65285_,
    new_n65286_, new_n65287_, new_n65288_, new_n65289_, new_n65290_,
    new_n65291_, new_n65292_, new_n65293_, new_n65294_, new_n65295_,
    new_n65296_, new_n65297_, new_n65298_, new_n65299_, new_n65300_,
    new_n65301_, new_n65302_, new_n65303_, new_n65304_, new_n65305_,
    new_n65306_, new_n65307_, new_n65308_, new_n65309_, new_n65310_,
    new_n65311_, new_n65312_, new_n65313_, new_n65314_, new_n65315_,
    new_n65316_, new_n65317_, new_n65318_, new_n65319_, new_n65320_,
    new_n65321_, new_n65322_, new_n65323_, new_n65324_, new_n65325_,
    new_n65326_, new_n65327_, new_n65328_, new_n65329_, new_n65330_,
    new_n65331_, new_n65332_, new_n65333_, new_n65334_, new_n65335_,
    new_n65336_, new_n65337_, new_n65338_, new_n65339_, new_n65340_,
    new_n65341_, new_n65342_, new_n65343_, new_n65344_, new_n65345_,
    new_n65346_, new_n65347_, new_n65348_, new_n65349_, new_n65350_,
    new_n65351_, new_n65352_, new_n65353_, new_n65354_, new_n65355_,
    new_n65356_, new_n65357_, new_n65358_, new_n65359_, new_n65360_,
    new_n65361_, new_n65362_, new_n65363_, new_n65364_, new_n65365_,
    new_n65366_, new_n65367_, new_n65368_, new_n65369_, new_n65370_,
    new_n65371_, new_n65372_, new_n65373_, new_n65374_, new_n65375_,
    new_n65376_, new_n65377_, new_n65378_, new_n65379_, new_n65380_,
    new_n65381_, new_n65382_, new_n65383_, new_n65384_, new_n65385_,
    new_n65386_, new_n65387_, new_n65388_, new_n65389_, new_n65390_,
    new_n65391_, new_n65392_, new_n65393_, new_n65394_, new_n65395_,
    new_n65396_, new_n65397_, new_n65398_, new_n65399_, new_n65400_,
    new_n65401_, new_n65402_, new_n65403_, new_n65404_, new_n65405_,
    new_n65406_, new_n65407_, new_n65408_, new_n65409_, new_n65410_,
    new_n65411_, new_n65412_, new_n65413_, new_n65414_, new_n65415_,
    new_n65416_, new_n65417_, new_n65418_, new_n65419_, new_n65420_,
    new_n65421_, new_n65422_, new_n65423_, new_n65424_, new_n65425_,
    new_n65426_, new_n65427_, new_n65428_, new_n65429_, new_n65430_,
    new_n65431_, new_n65432_, new_n65433_, new_n65434_, new_n65435_,
    new_n65436_, new_n65437_, new_n65438_, new_n65439_, new_n65440_,
    new_n65441_, new_n65442_, new_n65443_, new_n65444_, new_n65445_,
    new_n65446_, new_n65447_, new_n65448_, new_n65449_, new_n65450_,
    new_n65451_, new_n65452_, new_n65453_, new_n65454_, new_n65455_,
    new_n65456_, new_n65457_, new_n65458_, new_n65459_, new_n65460_,
    new_n65461_, new_n65462_, new_n65463_, new_n65464_, new_n65465_,
    new_n65466_, new_n65467_, new_n65468_, new_n65469_, new_n65470_,
    new_n65471_, new_n65472_, new_n65473_, new_n65474_, new_n65475_,
    new_n65476_, new_n65477_, new_n65478_, new_n65479_, new_n65480_,
    new_n65481_, new_n65482_, new_n65483_, new_n65484_, new_n65485_,
    new_n65486_, new_n65487_, new_n65488_, new_n65489_, new_n65490_,
    new_n65491_, new_n65492_, new_n65493_, new_n65494_, new_n65495_,
    new_n65496_, new_n65497_, new_n65498_, new_n65499_, new_n65500_,
    new_n65501_, new_n65502_, new_n65503_, new_n65504_, new_n65505_,
    new_n65506_, new_n65507_, new_n65508_, new_n65509_, new_n65510_,
    new_n65511_, new_n65512_, new_n65513_, new_n65514_, new_n65515_,
    new_n65516_, new_n65517_, new_n65518_, new_n65519_, new_n65520_,
    new_n65521_, new_n65522_, new_n65523_, new_n65524_, new_n65525_,
    new_n65526_, new_n65527_, new_n65528_, new_n65529_, new_n65530_,
    new_n65531_, new_n65532_, new_n65533_, new_n65534_, new_n65535_,
    new_n65536_, new_n65537_, new_n65538_, new_n65539_, new_n65540_,
    new_n65541_, new_n65542_, new_n65543_, new_n65544_, new_n65545_,
    new_n65546_, new_n65547_, new_n65548_, new_n65549_, new_n65550_,
    new_n65551_, new_n65552_, new_n65553_, new_n65554_, new_n65555_,
    new_n65556_, new_n65557_, new_n65558_, new_n65559_, new_n65560_,
    new_n65561_, new_n65562_, new_n65563_, new_n65564_, new_n65565_,
    new_n65566_, new_n65567_, new_n65568_, new_n65569_, new_n65570_,
    new_n65571_, new_n65572_, new_n65573_, new_n65574_, new_n65575_,
    new_n65576_, new_n65577_, new_n65578_, new_n65579_, new_n65580_,
    new_n65581_, new_n65582_, new_n65583_, new_n65584_, new_n65585_,
    new_n65586_, new_n65587_, new_n65588_, new_n65589_, new_n65590_,
    new_n65591_, new_n65592_, new_n65593_, new_n65594_, new_n65595_,
    new_n65596_, new_n65597_, new_n65598_, new_n65599_, new_n65600_,
    new_n65601_, new_n65602_, new_n65603_, new_n65604_, new_n65605_,
    new_n65606_, new_n65607_, new_n65608_, new_n65609_, new_n65610_,
    new_n65611_, new_n65612_, new_n65613_, new_n65614_, new_n65615_,
    new_n65616_, new_n65617_, new_n65618_, new_n65619_, new_n65620_,
    new_n65621_, new_n65622_, new_n65623_, new_n65624_, new_n65625_,
    new_n65626_, new_n65627_, new_n65628_, new_n65629_, new_n65630_,
    new_n65631_, new_n65632_, new_n65633_, new_n65634_, new_n65635_,
    new_n65636_, new_n65637_, new_n65638_, new_n65639_, new_n65640_,
    new_n65641_, new_n65642_, new_n65643_, new_n65644_, new_n65645_,
    new_n65646_, new_n65647_, new_n65648_, new_n65649_, new_n65650_,
    new_n65651_, new_n65652_, new_n65653_, new_n65654_, new_n65655_,
    new_n65656_, new_n65657_, new_n65658_, new_n65659_, new_n65660_,
    new_n65661_, new_n65662_, new_n65663_, new_n65664_, new_n65665_,
    new_n65666_, new_n65667_, new_n65668_, new_n65669_, new_n65670_,
    new_n65671_, new_n65672_, new_n65673_, new_n65674_, new_n65675_,
    new_n65676_, new_n65677_, new_n65678_, new_n65679_, new_n65680_,
    new_n65681_, new_n65682_, new_n65683_, new_n65684_, new_n65685_,
    new_n65686_, new_n65687_, new_n65688_, new_n65689_, new_n65690_,
    new_n65691_, new_n65692_, new_n65693_, new_n65694_, new_n65695_,
    new_n65696_, new_n65697_, new_n65698_, new_n65699_, new_n65700_,
    new_n65701_, new_n65702_, new_n65703_, new_n65704_, new_n65705_,
    new_n65706_, new_n65707_, new_n65708_, new_n65709_, new_n65710_,
    new_n65711_, new_n65712_, new_n65713_, new_n65714_, new_n65715_,
    new_n65716_, new_n65717_, new_n65718_, new_n65719_, new_n65720_,
    new_n65721_, new_n65722_, new_n65723_, new_n65724_, new_n65725_,
    new_n65726_, new_n65727_, new_n65728_, new_n65729_, new_n65730_,
    new_n65731_, new_n65732_, new_n65733_, new_n65734_, new_n65735_,
    new_n65736_, new_n65737_, new_n65738_, new_n65739_, new_n65740_,
    new_n65741_, new_n65742_, new_n65743_, new_n65744_, new_n65745_,
    new_n65746_, new_n65747_, new_n65748_, new_n65749_, new_n65750_,
    new_n65751_, new_n65752_, new_n65753_, new_n65754_, new_n65755_,
    new_n65756_, new_n65757_, new_n65758_, new_n65759_, new_n65760_,
    new_n65761_, new_n65762_, new_n65763_, new_n65764_, new_n65765_,
    new_n65766_, new_n65767_, new_n65768_, new_n65769_, new_n65770_,
    new_n65771_, new_n65772_, new_n65773_, new_n65774_, new_n65775_,
    new_n65776_, new_n65777_, new_n65778_, new_n65779_, new_n65780_,
    new_n65781_, new_n65782_, new_n65783_, new_n65784_, new_n65785_,
    new_n65786_, new_n65787_, new_n65788_, new_n65789_, new_n65790_,
    new_n65791_, new_n65792_, new_n65793_, new_n65794_, new_n65795_,
    new_n65796_, new_n65797_, new_n65798_, new_n65799_, new_n65800_,
    new_n65801_, new_n65802_, new_n65803_, new_n65804_, new_n65805_,
    new_n65806_, new_n65807_, new_n65808_, new_n65809_, new_n65810_,
    new_n65811_, new_n65812_, new_n65813_, new_n65814_, new_n65815_,
    new_n65816_, new_n65817_, new_n65818_, new_n65819_, new_n65820_,
    new_n65821_, new_n65822_, new_n65823_, new_n65824_, new_n65825_,
    new_n65826_, new_n65827_, new_n65828_, new_n65829_, new_n65830_,
    new_n65831_, new_n65832_, new_n65833_, new_n65834_, new_n65835_,
    new_n65836_, new_n65837_, new_n65838_, new_n65839_, new_n65840_,
    new_n65841_, new_n65842_, new_n65843_, new_n65844_, new_n65845_,
    new_n65846_, new_n65847_, new_n65848_, new_n65849_, new_n65850_,
    new_n65851_, new_n65852_, new_n65853_, new_n65854_, new_n65855_,
    new_n65856_, new_n65857_, new_n65858_, new_n65859_, new_n65860_,
    new_n65861_, new_n65862_, new_n65863_, new_n65864_, new_n65865_,
    new_n65866_, new_n65867_, new_n65868_, new_n65869_, new_n65870_,
    new_n65871_, new_n65872_, new_n65873_, new_n65874_, new_n65875_,
    new_n65876_, new_n65877_, new_n65878_, new_n65879_, new_n65880_,
    new_n65881_, new_n65882_, new_n65883_, new_n65884_, new_n65885_,
    new_n65886_, new_n65887_, new_n65888_, new_n65889_, new_n65890_,
    new_n65891_, new_n65892_, new_n65893_, new_n65894_, new_n65895_,
    new_n65896_, new_n65897_, new_n65898_, new_n65899_, new_n65900_,
    new_n65901_, new_n65902_, new_n65903_, new_n65904_, new_n65905_,
    new_n65906_, new_n65907_, new_n65908_, new_n65909_, new_n65910_,
    new_n65911_, new_n65912_, new_n65913_, new_n65914_, new_n65915_,
    new_n65916_, new_n65917_, new_n65918_, new_n65919_, new_n65920_,
    new_n65921_, new_n65922_, new_n65923_, new_n65924_, new_n65925_,
    new_n65926_, new_n65927_, new_n65928_, new_n65929_, new_n65930_,
    new_n65931_, new_n65932_, new_n65933_, new_n65934_, new_n65935_,
    new_n65936_, new_n65937_, new_n65938_, new_n65939_, new_n65940_,
    new_n65941_, new_n65942_, new_n65943_, new_n65944_, new_n65945_,
    new_n65946_, new_n65947_, new_n65948_, new_n65949_, new_n65950_,
    new_n65951_, new_n65952_, new_n65953_, new_n65954_, new_n65955_,
    new_n65956_, new_n65957_, new_n65958_, new_n65959_, new_n65960_,
    new_n65961_, new_n65962_, new_n65963_, new_n65964_, new_n65965_,
    new_n65966_, new_n65967_, new_n65968_, new_n65969_, new_n65970_,
    new_n65971_, new_n65972_, new_n65973_, new_n65974_, new_n65975_,
    new_n65976_, new_n65977_, new_n65978_, new_n65979_, new_n65980_,
    new_n65981_, new_n65982_, new_n65983_, new_n65984_, new_n65985_,
    new_n65986_, new_n65987_, new_n65988_, new_n65989_, new_n65990_,
    new_n65991_, new_n65992_, new_n65993_, new_n65994_, new_n65995_,
    new_n65996_, new_n65997_, new_n65998_, new_n65999_, new_n66000_,
    new_n66001_, new_n66002_, new_n66003_, new_n66004_, new_n66005_,
    new_n66006_, new_n66007_, new_n66008_, new_n66009_, new_n66010_,
    new_n66011_, new_n66012_, new_n66013_, new_n66014_, new_n66015_,
    new_n66016_, new_n66017_, new_n66018_, new_n66019_, new_n66020_,
    new_n66021_, new_n66022_, new_n66023_, new_n66024_, new_n66025_,
    new_n66026_, new_n66027_, new_n66028_, new_n66029_, new_n66030_,
    new_n66031_, new_n66032_, new_n66033_, new_n66034_, new_n66035_,
    new_n66036_, new_n66037_, new_n66038_, new_n66039_, new_n66040_,
    new_n66041_, new_n66042_, new_n66043_, new_n66044_, new_n66045_,
    new_n66046_, new_n66047_, new_n66048_, new_n66049_, new_n66050_,
    new_n66051_, new_n66052_, new_n66053_, new_n66054_, new_n66055_,
    new_n66056_, new_n66057_, new_n66058_, new_n66059_, new_n66060_,
    new_n66061_, new_n66062_, new_n66063_, new_n66064_, new_n66065_,
    new_n66066_, new_n66067_, new_n66068_, new_n66069_, new_n66070_,
    new_n66071_, new_n66072_, new_n66073_, new_n66074_, new_n66075_,
    new_n66076_, new_n66077_, new_n66078_, new_n66079_, new_n66080_,
    new_n66081_, new_n66082_, new_n66083_, new_n66084_, new_n66085_,
    new_n66086_, new_n66087_, new_n66088_, new_n66089_, new_n66090_,
    new_n66091_, new_n66092_, new_n66093_, new_n66094_, new_n66095_,
    new_n66096_, new_n66097_, new_n66098_, new_n66099_, new_n66100_,
    new_n66101_, new_n66102_, new_n66103_, new_n66104_, new_n66105_,
    new_n66106_, new_n66107_, new_n66108_, new_n66109_, new_n66110_,
    new_n66111_, new_n66112_, new_n66113_, new_n66114_, new_n66115_,
    new_n66116_, new_n66117_, new_n66118_, new_n66119_, new_n66120_,
    new_n66121_, new_n66122_, new_n66123_, new_n66124_, new_n66125_,
    new_n66126_, new_n66127_, new_n66128_, new_n66129_, new_n66130_,
    new_n66131_, new_n66132_, new_n66133_, new_n66134_, new_n66135_,
    new_n66136_, new_n66137_, new_n66138_, new_n66139_, new_n66140_,
    new_n66141_, new_n66142_, new_n66143_, new_n66144_, new_n66145_,
    new_n66146_, new_n66147_, new_n66148_, new_n66149_, new_n66150_,
    new_n66151_, new_n66152_, new_n66153_, new_n66154_, new_n66155_,
    new_n66156_, new_n66157_, new_n66158_, new_n66159_, new_n66160_,
    new_n66161_, new_n66162_, new_n66163_, new_n66164_, new_n66165_,
    new_n66166_, new_n66167_, new_n66168_, new_n66169_, new_n66170_,
    new_n66171_, new_n66172_, new_n66173_, new_n66174_, new_n66175_,
    new_n66176_, new_n66177_, new_n66178_, new_n66179_, new_n66180_,
    new_n66181_, new_n66182_, new_n66183_, new_n66184_, new_n66185_,
    new_n66186_, new_n66187_, new_n66188_, new_n66189_, new_n66190_,
    new_n66191_, new_n66192_, new_n66193_, new_n66194_, new_n66195_,
    new_n66196_, new_n66197_, new_n66198_, new_n66199_, new_n66200_,
    new_n66201_, new_n66202_, new_n66203_, new_n66204_, new_n66205_,
    new_n66206_, new_n66207_, new_n66208_, new_n66209_, new_n66210_,
    new_n66211_, new_n66212_, new_n66213_, new_n66214_, new_n66215_,
    new_n66216_, new_n66217_, new_n66218_, new_n66219_, new_n66220_,
    new_n66221_, new_n66222_, new_n66223_, new_n66224_, new_n66225_,
    new_n66226_, new_n66227_, new_n66228_, new_n66229_, new_n66230_,
    new_n66231_, new_n66232_, new_n66233_, new_n66234_, new_n66235_,
    new_n66236_, new_n66237_, new_n66238_, new_n66239_, new_n66240_,
    new_n66241_, new_n66242_, new_n66243_, new_n66244_, new_n66245_,
    new_n66246_, new_n66247_, new_n66248_, new_n66249_, new_n66250_,
    new_n66251_, new_n66252_, new_n66253_, new_n66254_, new_n66255_,
    new_n66256_, new_n66257_, new_n66258_, new_n66259_, new_n66260_,
    new_n66261_, new_n66262_, new_n66263_, new_n66264_, new_n66265_,
    new_n66266_, new_n66267_, new_n66268_, new_n66269_, new_n66270_,
    new_n66271_, new_n66272_, new_n66273_, new_n66274_, new_n66275_,
    new_n66276_, new_n66277_, new_n66278_, new_n66279_, new_n66280_,
    new_n66281_, new_n66282_, new_n66283_, new_n66284_, new_n66285_,
    new_n66286_, new_n66287_;
and  ( new_n258_, RIbb2d360_75, RIbb2f610_1 );
not  ( new_n259_, new_n258_ );
not  ( new_n260_, RIbb2f610_1 );
and  ( new_n261_, RIbb2f598_2, RIbb2f520_3 );
nor  ( new_n262_, new_n261_, new_n260_ );
not  ( new_n263_, new_n262_ );
not  ( new_n264_, RIbb2d3d8_74 );
xor  ( new_n265_, RIbb2f598_2, RIbb2f520_3 );
xor  ( new_n266_, RIbb2f598_2, new_n260_ );
nor  ( new_n267_, new_n266_, new_n265_ );
not  ( new_n268_, new_n267_ );
or   ( new_n269_, new_n268_, new_n264_ );
not  ( new_n270_, RIbb2d450_73 );
not  ( new_n271_, new_n265_ );
or   ( new_n272_, new_n271_, new_n270_ );
and  ( new_n273_, new_n272_, new_n269_ );
xor  ( new_n274_, new_n273_, new_n263_ );
not  ( new_n275_, RIbb2f430_5 );
and  ( new_n276_, RIbb2f3b8_6, RIbb2f340_7 );
nor  ( new_n277_, new_n276_, new_n275_ );
not  ( new_n278_, new_n277_ );
not  ( new_n279_, RIbb2d5b8_70 );
xor  ( new_n280_, RIbb2f3b8_6, RIbb2f340_7 );
xor  ( new_n281_, RIbb2f3b8_6, new_n275_ );
nor  ( new_n282_, new_n281_, new_n280_ );
not  ( new_n283_, new_n282_ );
or   ( new_n284_, new_n283_, new_n279_ );
not  ( new_n285_, RIbb2d630_69 );
not  ( new_n286_, new_n280_ );
or   ( new_n287_, new_n286_, new_n285_ );
and  ( new_n288_, new_n287_, new_n284_ );
xor  ( new_n289_, new_n288_, new_n278_ );
and  ( new_n290_, RIbb2f4a8_4, RIbb2f430_5 );
not  ( new_n291_, new_n290_ );
and  ( new_n292_, new_n291_, RIbb2f520_3 );
not  ( new_n293_, new_n292_ );
not  ( new_n294_, RIbb2d4c8_72 );
xor  ( new_n295_, RIbb2f4a8_4, RIbb2f430_5 );
not  ( new_n296_, RIbb2f520_3 );
xor  ( new_n297_, RIbb2f4a8_4, new_n296_ );
nor  ( new_n298_, new_n297_, new_n295_ );
not  ( new_n299_, new_n298_ );
or   ( new_n300_, new_n299_, new_n294_ );
not  ( new_n301_, RIbb2d540_71 );
not  ( new_n302_, new_n295_ );
or   ( new_n303_, new_n302_, new_n301_ );
and  ( new_n304_, new_n303_, new_n300_ );
xor  ( new_n305_, new_n304_, new_n293_ );
xnor ( new_n306_, new_n305_, new_n289_ );
xor  ( new_n307_, new_n306_, new_n274_ );
xor  ( new_n308_, new_n307_, new_n259_ );
not  ( new_n309_, RIbb2f340_7 );
and  ( new_n310_, RIbb2f2c8_8, RIbb2f250_9 );
nor  ( new_n311_, new_n310_, new_n309_ );
not  ( new_n312_, new_n311_ );
not  ( new_n313_, RIbb2d6a8_68 );
xor  ( new_n314_, RIbb2f2c8_8, RIbb2f250_9 );
xor  ( new_n315_, RIbb2f2c8_8, new_n309_ );
nor  ( new_n316_, new_n315_, new_n314_ );
not  ( new_n317_, new_n316_ );
or   ( new_n318_, new_n317_, new_n313_ );
not  ( new_n319_, RIbb2d720_67 );
not  ( new_n320_, new_n314_ );
or   ( new_n321_, new_n320_, new_n319_ );
and  ( new_n322_, new_n321_, new_n318_ );
xor  ( new_n323_, new_n322_, new_n312_ );
not  ( new_n324_, new_n323_ );
not  ( new_n325_, RIbb2f160_11 );
and  ( new_n326_, RIbb2f0e8_12, RIbb2f070_13 );
nor  ( new_n327_, new_n326_, new_n325_ );
not  ( new_n328_, new_n327_ );
not  ( new_n329_, RIbb2f250_9 );
and  ( new_n330_, RIbb2f1d8_10, RIbb2f160_11 );
nor  ( new_n331_, new_n330_, new_n329_ );
not  ( new_n332_, new_n331_ );
not  ( new_n333_, RIbb2d798_66 );
xor  ( new_n334_, RIbb2f1d8_10, RIbb2f160_11 );
xor  ( new_n335_, RIbb2f1d8_10, new_n329_ );
nor  ( new_n336_, new_n335_, new_n334_ );
not  ( new_n337_, new_n336_ );
or   ( new_n338_, new_n337_, new_n333_ );
not  ( new_n339_, RIbb2d810_65 );
not  ( new_n340_, new_n334_ );
or   ( new_n341_, new_n340_, new_n339_ );
and  ( new_n342_, new_n341_, new_n338_ );
xor  ( new_n343_, new_n342_, new_n332_ );
xor  ( new_n344_, new_n343_, new_n328_ );
xor  ( new_n345_, new_n344_, new_n324_ );
xnor ( new_n346_, new_n345_, new_n308_ );
not  ( new_n347_, new_n346_ );
not  ( new_n348_, RIbb2d360_75 );
or   ( new_n349_, new_n268_, new_n348_ );
or   ( new_n350_, new_n271_, new_n264_ );
and  ( new_n351_, new_n350_, new_n349_ );
xor  ( new_n352_, new_n351_, new_n263_ );
or   ( new_n353_, new_n283_, new_n301_ );
or   ( new_n354_, new_n286_, new_n279_ );
and  ( new_n355_, new_n354_, new_n353_ );
xor  ( new_n356_, new_n355_, new_n278_ );
or   ( new_n357_, new_n299_, new_n270_ );
or   ( new_n358_, new_n302_, new_n294_ );
and  ( new_n359_, new_n358_, new_n357_ );
xor  ( new_n360_, new_n359_, new_n293_ );
xor  ( new_n361_, new_n360_, new_n356_ );
xor  ( new_n362_, new_n361_, new_n352_ );
or   ( new_n363_, new_n317_, new_n285_ );
or   ( new_n364_, new_n320_, new_n313_ );
and  ( new_n365_, new_n364_, new_n363_ );
xor  ( new_n366_, new_n365_, new_n312_ );
or   ( new_n367_, new_n337_, new_n319_ );
or   ( new_n368_, new_n340_, new_n333_ );
and  ( new_n369_, new_n368_, new_n367_ );
xor  ( new_n370_, new_n369_, new_n331_ );
xor  ( new_n371_, RIbb2f0e8_12, RIbb2f070_13 );
xor  ( new_n372_, RIbb2f0e8_12, new_n325_ );
nor  ( new_n373_, new_n372_, new_n371_ );
and  ( new_n374_, new_n373_, RIbb2d810_65 );
xor  ( new_n375_, new_n374_, new_n328_ );
xor  ( new_n376_, new_n375_, new_n370_ );
xor  ( new_n377_, new_n376_, new_n366_ );
nand ( new_n378_, new_n377_, new_n362_ );
and  ( new_n379_, RIbb2f610_1, RIbb2d2e8_76 );
nor  ( new_n380_, new_n377_, new_n362_ );
or   ( new_n381_, new_n380_, new_n379_ );
and  ( new_n382_, new_n381_, new_n378_ );
xor  ( new_n383_, new_n382_, new_n347_ );
or   ( new_n384_, new_n317_, new_n279_ );
or   ( new_n385_, new_n320_, new_n285_ );
and  ( new_n386_, new_n385_, new_n384_ );
xor  ( new_n387_, new_n386_, new_n312_ );
or   ( new_n388_, new_n283_, new_n294_ );
or   ( new_n389_, new_n286_, new_n301_ );
and  ( new_n390_, new_n389_, new_n388_ );
xor  ( new_n391_, new_n390_, new_n278_ );
nand ( new_n392_, new_n391_, new_n387_ );
or   ( new_n393_, new_n299_, new_n264_ );
or   ( new_n394_, new_n302_, new_n270_ );
and  ( new_n395_, new_n394_, new_n393_ );
xor  ( new_n396_, new_n395_, new_n293_ );
or   ( new_n397_, new_n391_, new_n387_ );
nand ( new_n398_, new_n397_, new_n396_ );
and  ( new_n399_, new_n398_, new_n392_ );
not  ( new_n400_, RIbb2f070_13 );
and  ( new_n401_, RIbb2ef80_15, RIbb2eff8_14 );
nor  ( new_n402_, new_n401_, new_n400_ );
not  ( new_n403_, new_n402_ );
or   ( new_n404_, new_n337_, new_n313_ );
or   ( new_n405_, new_n340_, new_n319_ );
and  ( new_n406_, new_n405_, new_n404_ );
xor  ( new_n407_, new_n406_, new_n332_ );
nand ( new_n408_, new_n407_, new_n403_ );
not  ( new_n409_, new_n373_ );
or   ( new_n410_, new_n409_, new_n333_ );
not  ( new_n411_, new_n371_ );
or   ( new_n412_, new_n411_, new_n339_ );
and  ( new_n413_, new_n412_, new_n410_ );
xor  ( new_n414_, new_n413_, new_n328_ );
or   ( new_n415_, new_n407_, new_n403_ );
nand ( new_n416_, new_n415_, new_n414_ );
and  ( new_n417_, new_n416_, new_n408_ );
or   ( new_n418_, new_n417_, new_n399_ );
not  ( new_n419_, RIbb2d2e8_76 );
or   ( new_n420_, new_n268_, new_n419_ );
or   ( new_n421_, new_n271_, new_n348_ );
and  ( new_n422_, new_n421_, new_n420_ );
xor  ( new_n423_, new_n422_, new_n263_ );
and  ( new_n424_, RIbb2d270_77, RIbb2f610_1 );
nand ( new_n425_, new_n424_, new_n423_ );
and  ( new_n426_, new_n417_, new_n399_ );
or   ( new_n427_, new_n426_, new_n425_ );
and  ( new_n428_, new_n427_, new_n418_ );
xor  ( new_n429_, new_n428_, new_n383_ );
nor  ( new_n430_, new_n360_, new_n356_ );
and  ( new_n431_, new_n360_, new_n356_ );
nor  ( new_n432_, new_n431_, new_n352_ );
or   ( new_n433_, new_n432_, new_n430_ );
nand ( new_n434_, new_n375_, new_n370_ );
nor  ( new_n435_, new_n375_, new_n370_ );
or   ( new_n436_, new_n435_, new_n366_ );
and  ( new_n437_, new_n436_, new_n434_ );
xor  ( new_n438_, new_n437_, new_n379_ );
xor  ( new_n439_, new_n438_, new_n433_ );
xnor ( new_n440_, new_n439_, new_n429_ );
xor  ( new_n441_, new_n377_, new_n362_ );
xnor ( new_n442_, new_n441_, new_n379_ );
not  ( new_n443_, RIbb2d270_77 );
or   ( new_n444_, new_n268_, new_n443_ );
or   ( new_n445_, new_n271_, new_n419_ );
and  ( new_n446_, new_n445_, new_n444_ );
xor  ( new_n447_, new_n446_, new_n263_ );
and  ( new_n448_, RIbb2d1f8_78, RIbb2f610_1 );
or   ( new_n449_, new_n448_, new_n447_ );
or   ( new_n450_, new_n409_, new_n319_ );
or   ( new_n451_, new_n411_, new_n333_ );
and  ( new_n452_, new_n451_, new_n450_ );
xor  ( new_n453_, new_n452_, new_n327_ );
xor  ( new_n454_, RIbb2ef80_15, RIbb2eff8_14 );
xor  ( new_n455_, RIbb2eff8_14, new_n400_ );
nor  ( new_n456_, new_n455_, new_n454_ );
and  ( new_n457_, new_n456_, RIbb2d810_65 );
xor  ( new_n458_, new_n457_, new_n403_ );
nand ( new_n459_, new_n458_, new_n453_ );
or   ( new_n460_, new_n337_, new_n285_ );
or   ( new_n461_, new_n340_, new_n313_ );
and  ( new_n462_, new_n461_, new_n460_ );
xor  ( new_n463_, new_n462_, new_n332_ );
nor  ( new_n464_, new_n458_, new_n453_ );
or   ( new_n465_, new_n464_, new_n463_ );
and  ( new_n466_, new_n465_, new_n459_ );
or   ( new_n467_, new_n466_, new_n449_ );
and  ( new_n468_, new_n466_, new_n449_ );
or   ( new_n469_, new_n317_, new_n301_ );
or   ( new_n470_, new_n320_, new_n279_ );
and  ( new_n471_, new_n470_, new_n469_ );
xor  ( new_n472_, new_n471_, new_n312_ );
or   ( new_n473_, new_n283_, new_n270_ );
or   ( new_n474_, new_n286_, new_n294_ );
and  ( new_n475_, new_n474_, new_n473_ );
xor  ( new_n476_, new_n475_, new_n278_ );
nor  ( new_n477_, new_n476_, new_n472_ );
or   ( new_n478_, new_n299_, new_n348_ );
or   ( new_n479_, new_n302_, new_n264_ );
and  ( new_n480_, new_n479_, new_n478_ );
xor  ( new_n481_, new_n480_, new_n293_ );
and  ( new_n482_, new_n476_, new_n472_ );
nor  ( new_n483_, new_n482_, new_n481_ );
nor  ( new_n484_, new_n483_, new_n477_ );
or   ( new_n485_, new_n484_, new_n468_ );
and  ( new_n486_, new_n485_, new_n467_ );
or   ( new_n487_, new_n486_, new_n442_ );
and  ( new_n488_, new_n486_, new_n442_ );
xor  ( new_n489_, new_n391_, new_n387_ );
xor  ( new_n490_, new_n489_, new_n396_ );
xor  ( new_n491_, new_n407_, new_n403_ );
xor  ( new_n492_, new_n491_, new_n414_ );
nor  ( new_n493_, new_n492_, new_n490_ );
xor  ( new_n494_, new_n424_, new_n423_ );
and  ( new_n495_, new_n492_, new_n490_ );
nor  ( new_n496_, new_n495_, new_n494_ );
nor  ( new_n497_, new_n496_, new_n493_ );
or   ( new_n498_, new_n497_, new_n488_ );
and  ( new_n499_, new_n498_, new_n487_ );
xor  ( new_n500_, new_n499_, new_n440_ );
xor  ( new_n501_, new_n417_, new_n399_ );
xor  ( new_n502_, new_n501_, new_n425_ );
xnor ( new_n503_, new_n492_, new_n490_ );
xor  ( new_n504_, new_n503_, new_n494_ );
or   ( new_n505_, new_n299_, new_n419_ );
or   ( new_n506_, new_n302_, new_n348_ );
and  ( new_n507_, new_n506_, new_n505_ );
xor  ( new_n508_, new_n507_, new_n293_ );
not  ( new_n509_, RIbb2d1f8_78 );
or   ( new_n510_, new_n268_, new_n509_ );
or   ( new_n511_, new_n271_, new_n443_ );
and  ( new_n512_, new_n511_, new_n510_ );
xor  ( new_n513_, new_n512_, new_n263_ );
nor  ( new_n514_, new_n513_, new_n508_ );
not  ( new_n515_, RIbb2d180_79 );
or   ( new_n516_, new_n515_, new_n260_ );
nand ( new_n517_, new_n513_, new_n508_ );
and  ( new_n518_, new_n517_, new_n516_ );
or   ( new_n519_, new_n518_, new_n514_ );
not  ( new_n520_, RIbb2ef80_15 );
and  ( new_n521_, RIbb2ee90_17, RIbb2ef08_16 );
nor  ( new_n522_, new_n521_, new_n520_ );
not  ( new_n523_, new_n522_ );
not  ( new_n524_, new_n456_ );
or   ( new_n525_, new_n524_, new_n333_ );
not  ( new_n526_, new_n454_ );
or   ( new_n527_, new_n526_, new_n339_ );
and  ( new_n528_, new_n527_, new_n525_ );
xor  ( new_n529_, new_n528_, new_n403_ );
nand ( new_n530_, new_n529_, new_n523_ );
or   ( new_n531_, new_n409_, new_n313_ );
or   ( new_n532_, new_n411_, new_n319_ );
and  ( new_n533_, new_n532_, new_n531_ );
xor  ( new_n534_, new_n533_, new_n327_ );
nor  ( new_n535_, new_n529_, new_n523_ );
or   ( new_n536_, new_n535_, new_n534_ );
and  ( new_n537_, new_n536_, new_n530_ );
or   ( new_n538_, new_n537_, new_n519_ );
and  ( new_n539_, new_n537_, new_n519_ );
or   ( new_n540_, new_n337_, new_n279_ );
or   ( new_n541_, new_n340_, new_n285_ );
and  ( new_n542_, new_n541_, new_n540_ );
xor  ( new_n543_, new_n542_, new_n332_ );
or   ( new_n544_, new_n317_, new_n294_ );
or   ( new_n545_, new_n320_, new_n301_ );
and  ( new_n546_, new_n545_, new_n544_ );
xor  ( new_n547_, new_n546_, new_n312_ );
nor  ( new_n548_, new_n547_, new_n543_ );
or   ( new_n549_, new_n283_, new_n264_ );
or   ( new_n550_, new_n286_, new_n270_ );
and  ( new_n551_, new_n550_, new_n549_ );
xor  ( new_n552_, new_n551_, new_n278_ );
not  ( new_n553_, new_n552_ );
nand ( new_n554_, new_n547_, new_n543_ );
and  ( new_n555_, new_n554_, new_n553_ );
or   ( new_n556_, new_n555_, new_n548_ );
or   ( new_n557_, new_n556_, new_n539_ );
and  ( new_n558_, new_n557_, new_n538_ );
or   ( new_n559_, new_n558_, new_n504_ );
and  ( new_n560_, new_n558_, new_n504_ );
xnor ( new_n561_, new_n458_, new_n453_ );
xor  ( new_n562_, new_n561_, new_n463_ );
xnor ( new_n563_, new_n476_, new_n472_ );
xor  ( new_n564_, new_n563_, new_n481_ );
or   ( new_n565_, new_n564_, new_n562_ );
xor  ( new_n566_, new_n448_, new_n447_ );
and  ( new_n567_, new_n564_, new_n562_ );
or   ( new_n568_, new_n567_, new_n566_ );
and  ( new_n569_, new_n568_, new_n565_ );
or   ( new_n570_, new_n569_, new_n560_ );
and  ( new_n571_, new_n570_, new_n559_ );
or   ( new_n572_, new_n571_, new_n502_ );
and  ( new_n573_, new_n571_, new_n502_ );
xnor ( new_n574_, new_n486_, new_n442_ );
xor  ( new_n575_, new_n574_, new_n497_ );
or   ( new_n576_, new_n575_, new_n573_ );
and  ( new_n577_, new_n576_, new_n572_ );
nor  ( new_n578_, new_n577_, new_n500_ );
and  ( new_n579_, new_n439_, new_n429_ );
nor  ( new_n580_, new_n439_, new_n429_ );
nor  ( new_n581_, new_n499_, new_n580_ );
or   ( new_n582_, new_n581_, new_n579_ );
nor  ( new_n583_, new_n305_, new_n289_ );
and  ( new_n584_, new_n305_, new_n289_ );
nor  ( new_n585_, new_n584_, new_n274_ );
nor  ( new_n586_, new_n585_, new_n583_ );
not  ( new_n587_, new_n586_ );
and  ( new_n588_, new_n343_, new_n328_ );
nor  ( new_n589_, new_n343_, new_n328_ );
nor  ( new_n590_, new_n589_, new_n324_ );
nor  ( new_n591_, new_n590_, new_n588_ );
xor  ( new_n592_, new_n591_, new_n587_ );
not  ( new_n593_, new_n592_ );
or   ( new_n594_, new_n283_, new_n285_ );
or   ( new_n595_, new_n286_, new_n313_ );
and  ( new_n596_, new_n595_, new_n594_ );
xor  ( new_n597_, new_n596_, new_n278_ );
or   ( new_n598_, new_n317_, new_n319_ );
or   ( new_n599_, new_n320_, new_n333_ );
and  ( new_n600_, new_n599_, new_n598_ );
xor  ( new_n601_, new_n600_, new_n312_ );
and  ( new_n602_, new_n336_, RIbb2d810_65 );
xor  ( new_n603_, new_n602_, new_n332_ );
not  ( new_n604_, new_n603_ );
xor  ( new_n605_, new_n604_, new_n601_ );
xor  ( new_n606_, new_n605_, new_n597_ );
xor  ( new_n607_, new_n606_, new_n593_ );
nor  ( new_n608_, new_n437_, new_n379_ );
nand ( new_n609_, new_n437_, new_n379_ );
and  ( new_n610_, new_n609_, new_n433_ );
or   ( new_n611_, new_n610_, new_n608_ );
and  ( new_n612_, new_n307_, new_n259_ );
or   ( new_n613_, new_n307_, new_n259_ );
and  ( new_n614_, new_n345_, new_n613_ );
nor  ( new_n615_, new_n614_, new_n612_ );
not  ( new_n616_, new_n615_ );
xor  ( new_n617_, new_n616_, new_n611_ );
or   ( new_n618_, new_n260_, new_n264_ );
or   ( new_n619_, new_n299_, new_n301_ );
or   ( new_n620_, new_n302_, new_n279_ );
and  ( new_n621_, new_n620_, new_n619_ );
xor  ( new_n622_, new_n621_, new_n293_ );
or   ( new_n623_, new_n268_, new_n270_ );
or   ( new_n624_, new_n271_, new_n294_ );
and  ( new_n625_, new_n624_, new_n623_ );
xor  ( new_n626_, new_n625_, new_n263_ );
xor  ( new_n627_, new_n626_, new_n622_ );
xor  ( new_n628_, new_n627_, new_n618_ );
xor  ( new_n629_, new_n628_, new_n617_ );
not  ( new_n630_, new_n629_ );
xor  ( new_n631_, new_n630_, new_n607_ );
nor  ( new_n632_, new_n382_, new_n347_ );
and  ( new_n633_, new_n382_, new_n347_ );
nor  ( new_n634_, new_n428_, new_n633_ );
nor  ( new_n635_, new_n634_, new_n632_ );
xor  ( new_n636_, new_n635_, new_n631_ );
xor  ( new_n637_, new_n636_, new_n582_ );
and  ( new_n638_, new_n637_, new_n578_ );
xor  ( new_n639_, new_n571_, new_n502_ );
xor  ( new_n640_, new_n639_, new_n575_ );
xnor ( new_n641_, new_n564_, new_n562_ );
xor  ( new_n642_, new_n641_, new_n566_ );
or   ( new_n643_, new_n299_, new_n443_ );
or   ( new_n644_, new_n302_, new_n419_ );
and  ( new_n645_, new_n644_, new_n643_ );
xor  ( new_n646_, new_n645_, new_n293_ );
or   ( new_n647_, new_n268_, new_n515_ );
or   ( new_n648_, new_n271_, new_n509_ );
and  ( new_n649_, new_n648_, new_n647_ );
xor  ( new_n650_, new_n649_, new_n263_ );
or   ( new_n651_, new_n650_, new_n646_ );
and  ( new_n652_, RIbb2d108_80, RIbb2f610_1 );
and  ( new_n653_, new_n650_, new_n646_ );
or   ( new_n654_, new_n653_, new_n652_ );
and  ( new_n655_, new_n654_, new_n651_ );
or   ( new_n656_, new_n524_, new_n319_ );
or   ( new_n657_, new_n526_, new_n333_ );
and  ( new_n658_, new_n657_, new_n656_ );
xor  ( new_n659_, new_n658_, new_n402_ );
xor  ( new_n660_, RIbb2ee90_17, RIbb2ef08_16 );
xor  ( new_n661_, RIbb2ef08_16, new_n520_ );
nor  ( new_n662_, new_n661_, new_n660_ );
and  ( new_n663_, new_n662_, RIbb2d810_65 );
xor  ( new_n664_, new_n663_, new_n523_ );
nand ( new_n665_, new_n664_, new_n659_ );
nor  ( new_n666_, new_n664_, new_n659_ );
or   ( new_n667_, new_n409_, new_n285_ );
or   ( new_n668_, new_n411_, new_n313_ );
and  ( new_n669_, new_n668_, new_n667_ );
xor  ( new_n670_, new_n669_, new_n328_ );
or   ( new_n671_, new_n670_, new_n666_ );
and  ( new_n672_, new_n671_, new_n665_ );
or   ( new_n673_, new_n672_, new_n655_ );
and  ( new_n674_, new_n672_, new_n655_ );
or   ( new_n675_, new_n337_, new_n301_ );
or   ( new_n676_, new_n340_, new_n279_ );
and  ( new_n677_, new_n676_, new_n675_ );
xor  ( new_n678_, new_n677_, new_n332_ );
or   ( new_n679_, new_n317_, new_n270_ );
or   ( new_n680_, new_n320_, new_n294_ );
and  ( new_n681_, new_n680_, new_n679_ );
xor  ( new_n682_, new_n681_, new_n312_ );
nor  ( new_n683_, new_n682_, new_n678_ );
and  ( new_n684_, new_n682_, new_n678_ );
or   ( new_n685_, new_n283_, new_n348_ );
or   ( new_n686_, new_n286_, new_n264_ );
and  ( new_n687_, new_n686_, new_n685_ );
xor  ( new_n688_, new_n687_, new_n278_ );
nor  ( new_n689_, new_n688_, new_n684_ );
nor  ( new_n690_, new_n689_, new_n683_ );
or   ( new_n691_, new_n690_, new_n674_ );
and  ( new_n692_, new_n691_, new_n673_ );
nor  ( new_n693_, new_n692_, new_n642_ );
nand ( new_n694_, new_n692_, new_n642_ );
xor  ( new_n695_, new_n529_, new_n523_ );
xor  ( new_n696_, new_n695_, new_n534_ );
xor  ( new_n697_, new_n513_, new_n508_ );
xor  ( new_n698_, new_n697_, new_n516_ );
or   ( new_n699_, new_n698_, new_n696_ );
and  ( new_n700_, new_n698_, new_n696_ );
xor  ( new_n701_, new_n547_, new_n543_ );
xor  ( new_n702_, new_n701_, new_n553_ );
or   ( new_n703_, new_n702_, new_n700_ );
and  ( new_n704_, new_n703_, new_n699_ );
and  ( new_n705_, new_n704_, new_n694_ );
or   ( new_n706_, new_n705_, new_n693_ );
xnor ( new_n707_, new_n466_, new_n449_ );
xor  ( new_n708_, new_n707_, new_n484_ );
or   ( new_n709_, new_n708_, new_n706_ );
and  ( new_n710_, new_n708_, new_n706_ );
xor  ( new_n711_, new_n558_, new_n504_ );
xor  ( new_n712_, new_n711_, new_n569_ );
or   ( new_n713_, new_n712_, new_n710_ );
and  ( new_n714_, new_n713_, new_n709_ );
nor  ( new_n715_, new_n714_, new_n640_ );
xor  ( new_n716_, new_n577_, new_n500_ );
and  ( new_n717_, new_n716_, new_n715_ );
xor  ( new_n718_, new_n692_, new_n642_ );
xor  ( new_n719_, new_n718_, new_n704_ );
xor  ( new_n720_, new_n537_, new_n519_ );
xor  ( new_n721_, new_n720_, new_n556_ );
nor  ( new_n722_, new_n721_, new_n719_ );
and  ( new_n723_, new_n721_, new_n719_ );
xor  ( new_n724_, new_n650_, new_n646_ );
xnor ( new_n725_, new_n724_, new_n652_ );
xnor ( new_n726_, new_n682_, new_n678_ );
xor  ( new_n727_, new_n726_, new_n688_ );
nand ( new_n728_, new_n727_, new_n725_ );
or   ( new_n729_, new_n409_, new_n279_ );
or   ( new_n730_, new_n411_, new_n285_ );
and  ( new_n731_, new_n730_, new_n729_ );
xor  ( new_n732_, new_n731_, new_n328_ );
or   ( new_n733_, new_n337_, new_n294_ );
or   ( new_n734_, new_n340_, new_n301_ );
and  ( new_n735_, new_n734_, new_n733_ );
xor  ( new_n736_, new_n735_, new_n332_ );
nor  ( new_n737_, new_n736_, new_n732_ );
nand ( new_n738_, new_n736_, new_n732_ );
or   ( new_n739_, new_n317_, new_n264_ );
or   ( new_n740_, new_n320_, new_n270_ );
and  ( new_n741_, new_n740_, new_n739_ );
xor  ( new_n742_, new_n741_, new_n311_ );
and  ( new_n743_, new_n742_, new_n738_ );
or   ( new_n744_, new_n743_, new_n737_ );
not  ( new_n745_, RIbb2ee90_17 );
and  ( new_n746_, RIbb2eda0_19, RIbb2ee18_18 );
nor  ( new_n747_, new_n746_, new_n745_ );
not  ( new_n748_, new_n747_ );
or   ( new_n749_, new_n524_, new_n313_ );
or   ( new_n750_, new_n526_, new_n319_ );
and  ( new_n751_, new_n750_, new_n749_ );
xor  ( new_n752_, new_n751_, new_n403_ );
nand ( new_n753_, new_n752_, new_n748_ );
or   ( new_n754_, new_n752_, new_n748_ );
not  ( new_n755_, new_n662_ );
or   ( new_n756_, new_n755_, new_n333_ );
not  ( new_n757_, new_n660_ );
or   ( new_n758_, new_n757_, new_n339_ );
and  ( new_n759_, new_n758_, new_n756_ );
xor  ( new_n760_, new_n759_, new_n523_ );
nand ( new_n761_, new_n760_, new_n754_ );
and  ( new_n762_, new_n761_, new_n753_ );
nand ( new_n763_, new_n762_, new_n744_ );
nor  ( new_n764_, new_n762_, new_n744_ );
or   ( new_n765_, new_n283_, new_n419_ );
or   ( new_n766_, new_n286_, new_n348_ );
and  ( new_n767_, new_n766_, new_n765_ );
xor  ( new_n768_, new_n767_, new_n278_ );
or   ( new_n769_, new_n299_, new_n509_ );
or   ( new_n770_, new_n302_, new_n443_ );
and  ( new_n771_, new_n770_, new_n769_ );
xor  ( new_n772_, new_n771_, new_n293_ );
nor  ( new_n773_, new_n772_, new_n768_ );
and  ( new_n774_, new_n772_, new_n768_ );
not  ( new_n775_, RIbb2d108_80 );
or   ( new_n776_, new_n268_, new_n775_ );
or   ( new_n777_, new_n271_, new_n515_ );
and  ( new_n778_, new_n777_, new_n776_ );
xor  ( new_n779_, new_n778_, new_n263_ );
nor  ( new_n780_, new_n779_, new_n774_ );
nor  ( new_n781_, new_n780_, new_n773_ );
or   ( new_n782_, new_n781_, new_n764_ );
and  ( new_n783_, new_n782_, new_n763_ );
nor  ( new_n784_, new_n783_, new_n728_ );
and  ( new_n785_, new_n783_, new_n728_ );
xor  ( new_n786_, new_n698_, new_n696_ );
xnor ( new_n787_, new_n786_, new_n702_ );
nor  ( new_n788_, new_n787_, new_n785_ );
nor  ( new_n789_, new_n788_, new_n784_ );
not  ( new_n790_, new_n789_ );
nor  ( new_n791_, new_n790_, new_n723_ );
nor  ( new_n792_, new_n791_, new_n722_ );
xor  ( new_n793_, new_n708_, new_n706_ );
xor  ( new_n794_, new_n793_, new_n712_ );
nor  ( new_n795_, new_n794_, new_n792_ );
xor  ( new_n796_, new_n714_, new_n640_ );
and  ( new_n797_, new_n796_, new_n795_ );
xnor ( new_n798_, new_n794_, new_n792_ );
xor  ( new_n799_, new_n721_, new_n719_ );
xor  ( new_n800_, new_n799_, new_n790_ );
xor  ( new_n801_, new_n762_, new_n744_ );
xnor ( new_n802_, new_n801_, new_n781_ );
xor  ( new_n803_, new_n664_, new_n659_ );
xnor ( new_n804_, new_n803_, new_n670_ );
not  ( new_n805_, RIbb2d090_81 );
or   ( new_n806_, new_n805_, new_n260_ );
xor  ( new_n807_, new_n736_, new_n732_ );
xor  ( new_n808_, new_n807_, new_n742_ );
nand ( new_n809_, new_n808_, new_n806_ );
nor  ( new_n810_, new_n808_, new_n806_ );
xor  ( new_n811_, new_n772_, new_n768_ );
xor  ( new_n812_, new_n811_, new_n779_ );
or   ( new_n813_, new_n812_, new_n810_ );
and  ( new_n814_, new_n813_, new_n809_ );
xor  ( new_n815_, new_n814_, new_n804_ );
or   ( new_n816_, new_n755_, new_n319_ );
or   ( new_n817_, new_n757_, new_n333_ );
and  ( new_n818_, new_n817_, new_n816_ );
xor  ( new_n819_, new_n818_, new_n522_ );
xor  ( new_n820_, RIbb2eda0_19, RIbb2ee18_18 );
xor  ( new_n821_, RIbb2ee18_18, new_n745_ );
nor  ( new_n822_, new_n821_, new_n820_ );
and  ( new_n823_, new_n822_, RIbb2d810_65 );
xor  ( new_n824_, new_n823_, new_n748_ );
nand ( new_n825_, new_n824_, new_n819_ );
nor  ( new_n826_, new_n824_, new_n819_ );
or   ( new_n827_, new_n524_, new_n285_ );
or   ( new_n828_, new_n526_, new_n313_ );
and  ( new_n829_, new_n828_, new_n827_ );
xor  ( new_n830_, new_n829_, new_n403_ );
or   ( new_n831_, new_n830_, new_n826_ );
and  ( new_n832_, new_n831_, new_n825_ );
or   ( new_n833_, new_n409_, new_n301_ );
or   ( new_n834_, new_n411_, new_n279_ );
and  ( new_n835_, new_n834_, new_n833_ );
xor  ( new_n836_, new_n835_, new_n328_ );
or   ( new_n837_, new_n337_, new_n270_ );
or   ( new_n838_, new_n340_, new_n294_ );
and  ( new_n839_, new_n838_, new_n837_ );
xor  ( new_n840_, new_n839_, new_n332_ );
or   ( new_n841_, new_n840_, new_n836_ );
and  ( new_n842_, new_n840_, new_n836_ );
or   ( new_n843_, new_n317_, new_n348_ );
or   ( new_n844_, new_n320_, new_n264_ );
and  ( new_n845_, new_n844_, new_n843_ );
xor  ( new_n846_, new_n845_, new_n312_ );
or   ( new_n847_, new_n846_, new_n842_ );
and  ( new_n848_, new_n847_, new_n841_ );
or   ( new_n849_, new_n848_, new_n832_ );
and  ( new_n850_, new_n848_, new_n832_ );
or   ( new_n851_, new_n283_, new_n443_ );
or   ( new_n852_, new_n286_, new_n419_ );
and  ( new_n853_, new_n852_, new_n851_ );
xor  ( new_n854_, new_n853_, new_n278_ );
or   ( new_n855_, new_n299_, new_n515_ );
or   ( new_n856_, new_n302_, new_n509_ );
and  ( new_n857_, new_n856_, new_n855_ );
xor  ( new_n858_, new_n857_, new_n293_ );
nor  ( new_n859_, new_n858_, new_n854_ );
and  ( new_n860_, new_n858_, new_n854_ );
or   ( new_n861_, new_n268_, new_n805_ );
or   ( new_n862_, new_n271_, new_n775_ );
and  ( new_n863_, new_n862_, new_n861_ );
xor  ( new_n864_, new_n863_, new_n263_ );
nor  ( new_n865_, new_n864_, new_n860_ );
nor  ( new_n866_, new_n865_, new_n859_ );
or   ( new_n867_, new_n866_, new_n850_ );
and  ( new_n868_, new_n867_, new_n849_ );
xor  ( new_n869_, new_n868_, new_n815_ );
nor  ( new_n870_, new_n869_, new_n802_ );
xor  ( new_n871_, new_n808_, new_n806_ );
xor  ( new_n872_, new_n871_, new_n812_ );
xor  ( new_n873_, new_n752_, new_n748_ );
xor  ( new_n874_, new_n873_, new_n760_ );
or   ( new_n875_, new_n874_, new_n872_ );
nand ( new_n876_, new_n874_, new_n872_ );
xor  ( new_n877_, new_n848_, new_n832_ );
xnor ( new_n878_, new_n877_, new_n866_ );
nand ( new_n879_, new_n878_, new_n876_ );
and  ( new_n880_, new_n879_, new_n875_ );
xor  ( new_n881_, new_n840_, new_n836_ );
xnor ( new_n882_, new_n881_, new_n846_ );
xnor ( new_n883_, new_n824_, new_n819_ );
xor  ( new_n884_, new_n883_, new_n830_ );
or   ( new_n885_, new_n884_, new_n882_ );
not  ( new_n886_, RIbb2d018_82 );
or   ( new_n887_, new_n886_, new_n260_ );
xnor ( new_n888_, new_n858_, new_n854_ );
xor  ( new_n889_, new_n888_, new_n864_ );
and  ( new_n890_, new_n889_, new_n887_ );
nand ( new_n891_, new_n890_, new_n885_ );
nor  ( new_n892_, new_n890_, new_n885_ );
not  ( new_n893_, RIbb2eda0_19 );
and  ( new_n894_, RIbb2ecb0_21, RIbb2ed28_20 );
nor  ( new_n895_, new_n894_, new_n893_ );
not  ( new_n896_, new_n895_ );
not  ( new_n897_, new_n822_ );
or   ( new_n898_, new_n897_, new_n333_ );
not  ( new_n899_, new_n820_ );
or   ( new_n900_, new_n899_, new_n339_ );
and  ( new_n901_, new_n900_, new_n898_ );
xor  ( new_n902_, new_n901_, new_n748_ );
and  ( new_n903_, new_n902_, new_n896_ );
or   ( new_n904_, new_n902_, new_n896_ );
or   ( new_n905_, new_n755_, new_n313_ );
or   ( new_n906_, new_n757_, new_n319_ );
and  ( new_n907_, new_n906_, new_n905_ );
xor  ( new_n908_, new_n907_, new_n523_ );
and  ( new_n909_, new_n908_, new_n904_ );
or   ( new_n910_, new_n909_, new_n903_ );
or   ( new_n911_, new_n524_, new_n279_ );
or   ( new_n912_, new_n526_, new_n285_ );
and  ( new_n913_, new_n912_, new_n911_ );
xor  ( new_n914_, new_n913_, new_n403_ );
or   ( new_n915_, new_n409_, new_n294_ );
or   ( new_n916_, new_n411_, new_n301_ );
and  ( new_n917_, new_n916_, new_n915_ );
xor  ( new_n918_, new_n917_, new_n328_ );
or   ( new_n919_, new_n918_, new_n914_ );
and  ( new_n920_, new_n918_, new_n914_ );
or   ( new_n921_, new_n337_, new_n264_ );
or   ( new_n922_, new_n340_, new_n270_ );
and  ( new_n923_, new_n922_, new_n921_ );
xor  ( new_n924_, new_n923_, new_n332_ );
or   ( new_n925_, new_n924_, new_n920_ );
and  ( new_n926_, new_n925_, new_n919_ );
nor  ( new_n927_, new_n926_, new_n910_ );
and  ( new_n928_, new_n926_, new_n910_ );
or   ( new_n929_, new_n317_, new_n419_ );
or   ( new_n930_, new_n320_, new_n348_ );
and  ( new_n931_, new_n930_, new_n929_ );
xor  ( new_n932_, new_n931_, new_n312_ );
or   ( new_n933_, new_n283_, new_n509_ );
or   ( new_n934_, new_n286_, new_n443_ );
and  ( new_n935_, new_n934_, new_n933_ );
xor  ( new_n936_, new_n935_, new_n278_ );
nor  ( new_n937_, new_n936_, new_n932_ );
and  ( new_n938_, new_n936_, new_n932_ );
or   ( new_n939_, new_n299_, new_n775_ );
or   ( new_n940_, new_n302_, new_n515_ );
and  ( new_n941_, new_n940_, new_n939_ );
xor  ( new_n942_, new_n941_, new_n293_ );
nor  ( new_n943_, new_n942_, new_n938_ );
nor  ( new_n944_, new_n943_, new_n937_ );
nor  ( new_n945_, new_n944_, new_n928_ );
nor  ( new_n946_, new_n945_, new_n927_ );
or   ( new_n947_, new_n946_, new_n892_ );
and  ( new_n948_, new_n947_, new_n891_ );
or   ( new_n949_, new_n948_, new_n880_ );
and  ( new_n950_, new_n948_, new_n880_ );
xnor ( new_n951_, new_n727_, new_n725_ );
or   ( new_n952_, new_n951_, new_n950_ );
and  ( new_n953_, new_n952_, new_n949_ );
nand ( new_n954_, new_n953_, new_n870_ );
nor  ( new_n955_, new_n953_, new_n870_ );
not  ( new_n956_, new_n804_ );
and  ( new_n957_, new_n814_, new_n956_ );
or   ( new_n958_, new_n814_, new_n956_ );
and  ( new_n959_, new_n868_, new_n958_ );
nor  ( new_n960_, new_n959_, new_n957_ );
xnor ( new_n961_, new_n672_, new_n655_ );
xor  ( new_n962_, new_n961_, new_n690_ );
xor  ( new_n963_, new_n962_, new_n960_ );
xnor ( new_n964_, new_n783_, new_n728_ );
xor  ( new_n965_, new_n964_, new_n787_ );
xor  ( new_n966_, new_n965_, new_n963_ );
or   ( new_n967_, new_n966_, new_n955_ );
and  ( new_n968_, new_n967_, new_n954_ );
or   ( new_n969_, new_n968_, new_n800_ );
and  ( new_n970_, new_n968_, new_n800_ );
or   ( new_n971_, new_n962_, new_n960_ );
and  ( new_n972_, new_n962_, new_n960_ );
or   ( new_n973_, new_n965_, new_n972_ );
and  ( new_n974_, new_n973_, new_n971_ );
or   ( new_n975_, new_n974_, new_n970_ );
and  ( new_n976_, new_n975_, new_n969_ );
nor  ( new_n977_, new_n976_, new_n798_ );
xor  ( new_n978_, new_n889_, new_n887_ );
xnor ( new_n979_, new_n926_, new_n910_ );
xor  ( new_n980_, new_n979_, new_n944_ );
nor  ( new_n981_, new_n980_, new_n978_ );
nand ( new_n982_, new_n980_, new_n978_ );
xor  ( new_n983_, new_n884_, new_n882_ );
and  ( new_n984_, new_n983_, new_n982_ );
or   ( new_n985_, new_n984_, new_n981_ );
not  ( new_n986_, RIbb2cfa0_83 );
or   ( new_n987_, new_n268_, new_n986_ );
or   ( new_n988_, new_n271_, new_n886_ );
and  ( new_n989_, new_n988_, new_n987_ );
xor  ( new_n990_, new_n989_, new_n263_ );
and  ( new_n991_, RIbb2cf28_84, RIbb2f610_1 );
or   ( new_n992_, new_n991_, new_n990_ );
or   ( new_n993_, new_n268_, new_n886_ );
or   ( new_n994_, new_n271_, new_n805_ );
and  ( new_n995_, new_n994_, new_n993_ );
xor  ( new_n996_, new_n995_, new_n263_ );
or   ( new_n997_, new_n996_, new_n992_ );
and  ( new_n998_, new_n996_, new_n992_ );
and  ( new_n999_, RIbb2cfa0_83, RIbb2f610_1 );
or   ( new_n1000_, new_n999_, new_n998_ );
and  ( new_n1001_, new_n1000_, new_n997_ );
or   ( new_n1002_, new_n524_, new_n301_ );
or   ( new_n1003_, new_n526_, new_n279_ );
and  ( new_n1004_, new_n1003_, new_n1002_ );
xor  ( new_n1005_, new_n1004_, new_n403_ );
or   ( new_n1006_, new_n409_, new_n270_ );
or   ( new_n1007_, new_n411_, new_n294_ );
and  ( new_n1008_, new_n1007_, new_n1006_ );
xor  ( new_n1009_, new_n1008_, new_n328_ );
or   ( new_n1010_, new_n1009_, new_n1005_ );
and  ( new_n1011_, new_n1009_, new_n1005_ );
or   ( new_n1012_, new_n337_, new_n348_ );
or   ( new_n1013_, new_n340_, new_n264_ );
and  ( new_n1014_, new_n1013_, new_n1012_ );
xor  ( new_n1015_, new_n1014_, new_n332_ );
or   ( new_n1016_, new_n1015_, new_n1011_ );
and  ( new_n1017_, new_n1016_, new_n1010_ );
or   ( new_n1018_, new_n317_, new_n443_ );
or   ( new_n1019_, new_n320_, new_n419_ );
and  ( new_n1020_, new_n1019_, new_n1018_ );
xor  ( new_n1021_, new_n1020_, new_n312_ );
or   ( new_n1022_, new_n283_, new_n515_ );
or   ( new_n1023_, new_n286_, new_n509_ );
and  ( new_n1024_, new_n1023_, new_n1022_ );
xor  ( new_n1025_, new_n1024_, new_n278_ );
or   ( new_n1026_, new_n1025_, new_n1021_ );
and  ( new_n1027_, new_n1025_, new_n1021_ );
or   ( new_n1028_, new_n299_, new_n805_ );
or   ( new_n1029_, new_n302_, new_n775_ );
and  ( new_n1030_, new_n1029_, new_n1028_ );
xor  ( new_n1031_, new_n1030_, new_n293_ );
or   ( new_n1032_, new_n1031_, new_n1027_ );
and  ( new_n1033_, new_n1032_, new_n1026_ );
or   ( new_n1034_, new_n1033_, new_n1017_ );
and  ( new_n1035_, new_n1033_, new_n1017_ );
or   ( new_n1036_, new_n897_, new_n319_ );
or   ( new_n1037_, new_n899_, new_n333_ );
and  ( new_n1038_, new_n1037_, new_n1036_ );
xor  ( new_n1039_, new_n1038_, new_n747_ );
xor  ( new_n1040_, RIbb2ecb0_21, RIbb2ed28_20 );
xor  ( new_n1041_, RIbb2ed28_20, new_n893_ );
nor  ( new_n1042_, new_n1041_, new_n1040_ );
and  ( new_n1043_, new_n1042_, RIbb2d810_65 );
xor  ( new_n1044_, new_n1043_, new_n896_ );
and  ( new_n1045_, new_n1044_, new_n1039_ );
nor  ( new_n1046_, new_n1044_, new_n1039_ );
or   ( new_n1047_, new_n755_, new_n285_ );
or   ( new_n1048_, new_n757_, new_n313_ );
and  ( new_n1049_, new_n1048_, new_n1047_ );
xor  ( new_n1050_, new_n1049_, new_n523_ );
nor  ( new_n1051_, new_n1050_, new_n1046_ );
nor  ( new_n1052_, new_n1051_, new_n1045_ );
or   ( new_n1053_, new_n1052_, new_n1035_ );
and  ( new_n1054_, new_n1053_, new_n1034_ );
or   ( new_n1055_, new_n1054_, new_n1001_ );
and  ( new_n1056_, new_n1054_, new_n1001_ );
xor  ( new_n1057_, new_n902_, new_n895_ );
xor  ( new_n1058_, new_n1057_, new_n908_ );
xnor ( new_n1059_, new_n918_, new_n914_ );
xor  ( new_n1060_, new_n1059_, new_n924_ );
nor  ( new_n1061_, new_n1060_, new_n1058_ );
nand ( new_n1062_, new_n1060_, new_n1058_ );
xor  ( new_n1063_, new_n936_, new_n932_ );
xnor ( new_n1064_, new_n1063_, new_n942_ );
not  ( new_n1065_, new_n1064_ );
and  ( new_n1066_, new_n1065_, new_n1062_ );
or   ( new_n1067_, new_n1066_, new_n1061_ );
or   ( new_n1068_, new_n1067_, new_n1056_ );
and  ( new_n1069_, new_n1068_, new_n1055_ );
or   ( new_n1070_, new_n1069_, new_n985_ );
nand ( new_n1071_, new_n1069_, new_n985_ );
xor  ( new_n1072_, new_n874_, new_n872_ );
xor  ( new_n1073_, new_n1072_, new_n878_ );
nand ( new_n1074_, new_n1073_, new_n1071_ );
and  ( new_n1075_, new_n1074_, new_n1070_ );
xor  ( new_n1076_, new_n948_, new_n880_ );
xor  ( new_n1077_, new_n1076_, new_n951_ );
or   ( new_n1078_, new_n1077_, new_n1075_ );
and  ( new_n1079_, new_n1077_, new_n1075_ );
xor  ( new_n1080_, new_n869_, new_n802_ );
or   ( new_n1081_, new_n1080_, new_n1079_ );
and  ( new_n1082_, new_n1081_, new_n1078_ );
xnor ( new_n1083_, new_n953_, new_n870_ );
xor  ( new_n1084_, new_n1083_, new_n966_ );
nand ( new_n1085_, new_n1084_, new_n1082_ );
xor  ( new_n1086_, new_n968_, new_n800_ );
xor  ( new_n1087_, new_n1086_, new_n974_ );
nor  ( new_n1088_, new_n1087_, new_n1085_ );
xnor ( new_n1089_, new_n1077_, new_n1075_ );
xor  ( new_n1090_, new_n1089_, new_n1080_ );
xnor ( new_n1091_, new_n980_, new_n978_ );
xor  ( new_n1092_, new_n1091_, new_n983_ );
xnor ( new_n1093_, new_n1033_, new_n1017_ );
xor  ( new_n1094_, new_n1093_, new_n1052_ );
xnor ( new_n1095_, new_n996_, new_n992_ );
xor  ( new_n1096_, new_n1095_, new_n999_ );
or   ( new_n1097_, new_n1096_, new_n1094_ );
nand ( new_n1098_, new_n1096_, new_n1094_ );
xor  ( new_n1099_, new_n1060_, new_n1058_ );
xor  ( new_n1100_, new_n1099_, new_n1065_ );
nand ( new_n1101_, new_n1100_, new_n1098_ );
and  ( new_n1102_, new_n1101_, new_n1097_ );
or   ( new_n1103_, new_n1102_, new_n1092_ );
and  ( new_n1104_, new_n1102_, new_n1092_ );
xor  ( new_n1105_, new_n1009_, new_n1005_ );
xnor ( new_n1106_, new_n1105_, new_n1015_ );
xnor ( new_n1107_, new_n1044_, new_n1039_ );
xor  ( new_n1108_, new_n1107_, new_n1050_ );
nor  ( new_n1109_, new_n1108_, new_n1106_ );
or   ( new_n1110_, new_n409_, new_n264_ );
or   ( new_n1111_, new_n411_, new_n270_ );
and  ( new_n1112_, new_n1111_, new_n1110_ );
xor  ( new_n1113_, new_n1112_, new_n328_ );
or   ( new_n1114_, new_n524_, new_n294_ );
or   ( new_n1115_, new_n526_, new_n301_ );
and  ( new_n1116_, new_n1115_, new_n1114_ );
xor  ( new_n1117_, new_n1116_, new_n403_ );
and  ( new_n1118_, new_n1117_, new_n1113_ );
or   ( new_n1119_, new_n1117_, new_n1113_ );
or   ( new_n1120_, new_n755_, new_n279_ );
or   ( new_n1121_, new_n757_, new_n285_ );
and  ( new_n1122_, new_n1121_, new_n1120_ );
xor  ( new_n1123_, new_n1122_, new_n523_ );
and  ( new_n1124_, new_n1123_, new_n1119_ );
or   ( new_n1125_, new_n1124_, new_n1118_ );
not  ( new_n1126_, RIbb2ecb0_21 );
and  ( new_n1127_, RIbb2ebc0_23, RIbb2ec38_22 );
nor  ( new_n1128_, new_n1127_, new_n1126_ );
not  ( new_n1129_, new_n1128_ );
or   ( new_n1130_, new_n897_, new_n313_ );
or   ( new_n1131_, new_n899_, new_n319_ );
and  ( new_n1132_, new_n1131_, new_n1130_ );
xor  ( new_n1133_, new_n1132_, new_n748_ );
or   ( new_n1134_, new_n1133_, new_n1129_ );
not  ( new_n1135_, new_n1042_ );
or   ( new_n1136_, new_n1135_, new_n333_ );
not  ( new_n1137_, new_n1040_ );
or   ( new_n1138_, new_n1137_, new_n339_ );
and  ( new_n1139_, new_n1138_, new_n1136_ );
xor  ( new_n1140_, new_n1139_, new_n896_ );
and  ( new_n1141_, new_n1133_, new_n1129_ );
or   ( new_n1142_, new_n1141_, new_n1140_ );
and  ( new_n1143_, new_n1142_, new_n1134_ );
or   ( new_n1144_, new_n1143_, new_n1125_ );
nand ( new_n1145_, new_n1143_, new_n1125_ );
or   ( new_n1146_, new_n283_, new_n775_ );
or   ( new_n1147_, new_n286_, new_n515_ );
and  ( new_n1148_, new_n1147_, new_n1146_ );
xor  ( new_n1149_, new_n1148_, new_n278_ );
or   ( new_n1150_, new_n317_, new_n509_ );
or   ( new_n1151_, new_n320_, new_n443_ );
and  ( new_n1152_, new_n1151_, new_n1150_ );
xor  ( new_n1153_, new_n1152_, new_n312_ );
and  ( new_n1154_, new_n1153_, new_n1149_ );
nor  ( new_n1155_, new_n1153_, new_n1149_ );
or   ( new_n1156_, new_n337_, new_n419_ );
or   ( new_n1157_, new_n340_, new_n348_ );
and  ( new_n1158_, new_n1157_, new_n1156_ );
xor  ( new_n1159_, new_n1158_, new_n332_ );
not  ( new_n1160_, new_n1159_ );
nor  ( new_n1161_, new_n1160_, new_n1155_ );
nor  ( new_n1162_, new_n1161_, new_n1154_ );
nand ( new_n1163_, new_n1162_, new_n1145_ );
and  ( new_n1164_, new_n1163_, new_n1144_ );
nand ( new_n1165_, new_n1164_, new_n1109_ );
nor  ( new_n1166_, new_n1164_, new_n1109_ );
and  ( new_n1167_, RIbb2ceb0_85, RIbb2f610_1 );
not  ( new_n1168_, RIbb2cf28_84 );
or   ( new_n1169_, new_n268_, new_n1168_ );
or   ( new_n1170_, new_n271_, new_n986_ );
and  ( new_n1171_, new_n1170_, new_n1169_ );
xor  ( new_n1172_, new_n1171_, new_n263_ );
nand ( new_n1173_, new_n1172_, new_n1167_ );
or   ( new_n1174_, new_n1172_, new_n1167_ );
or   ( new_n1175_, new_n299_, new_n886_ );
or   ( new_n1176_, new_n302_, new_n805_ );
and  ( new_n1177_, new_n1176_, new_n1175_ );
xor  ( new_n1178_, new_n1177_, new_n293_ );
nand ( new_n1179_, new_n1178_, new_n1174_ );
and  ( new_n1180_, new_n1179_, new_n1173_ );
xnor ( new_n1181_, new_n1025_, new_n1021_ );
xor  ( new_n1182_, new_n1181_, new_n1031_ );
nor  ( new_n1183_, new_n1182_, new_n1180_ );
and  ( new_n1184_, new_n1182_, new_n1180_ );
xor  ( new_n1185_, new_n991_, new_n990_ );
nor  ( new_n1186_, new_n1185_, new_n1184_ );
nor  ( new_n1187_, new_n1186_, new_n1183_ );
or   ( new_n1188_, new_n1187_, new_n1166_ );
and  ( new_n1189_, new_n1188_, new_n1165_ );
or   ( new_n1190_, new_n1189_, new_n1104_ );
and  ( new_n1191_, new_n1190_, new_n1103_ );
xnor ( new_n1192_, new_n890_, new_n885_ );
xor  ( new_n1193_, new_n1192_, new_n946_ );
or   ( new_n1194_, new_n1193_, new_n1191_ );
and  ( new_n1195_, new_n1193_, new_n1191_ );
xor  ( new_n1196_, new_n1069_, new_n985_ );
xor  ( new_n1197_, new_n1196_, new_n1073_ );
or   ( new_n1198_, new_n1197_, new_n1195_ );
and  ( new_n1199_, new_n1198_, new_n1194_ );
nor  ( new_n1200_, new_n1199_, new_n1090_ );
xor  ( new_n1201_, new_n1084_, new_n1082_ );
and  ( new_n1202_, new_n1201_, new_n1200_ );
xor  ( new_n1203_, new_n1193_, new_n1191_ );
xor  ( new_n1204_, new_n1203_, new_n1197_ );
xor  ( new_n1205_, new_n1054_, new_n1001_ );
xor  ( new_n1206_, new_n1205_, new_n1067_ );
xor  ( new_n1207_, new_n1096_, new_n1094_ );
xor  ( new_n1208_, new_n1207_, new_n1100_ );
or   ( new_n1209_, new_n299_, new_n986_ );
or   ( new_n1210_, new_n302_, new_n886_ );
and  ( new_n1211_, new_n1210_, new_n1209_ );
xor  ( new_n1212_, new_n1211_, new_n293_ );
not  ( new_n1213_, RIbb2ceb0_85 );
or   ( new_n1214_, new_n268_, new_n1213_ );
or   ( new_n1215_, new_n271_, new_n1168_ );
and  ( new_n1216_, new_n1215_, new_n1214_ );
xor  ( new_n1217_, new_n1216_, new_n263_ );
or   ( new_n1218_, new_n1217_, new_n1212_ );
and  ( new_n1219_, RIbb2ce38_86, RIbb2f610_1 );
and  ( new_n1220_, new_n1217_, new_n1212_ );
or   ( new_n1221_, new_n1220_, new_n1219_ );
and  ( new_n1222_, new_n1221_, new_n1218_ );
xor  ( new_n1223_, new_n1172_, new_n1167_ );
xor  ( new_n1224_, new_n1223_, new_n1178_ );
or   ( new_n1225_, new_n1224_, new_n1222_ );
and  ( new_n1226_, new_n1224_, new_n1222_ );
xor  ( new_n1227_, new_n1153_, new_n1149_ );
xor  ( new_n1228_, new_n1227_, new_n1159_ );
or   ( new_n1229_, new_n1228_, new_n1226_ );
and  ( new_n1230_, new_n1229_, new_n1225_ );
or   ( new_n1231_, new_n337_, new_n443_ );
or   ( new_n1232_, new_n340_, new_n419_ );
and  ( new_n1233_, new_n1232_, new_n1231_ );
xor  ( new_n1234_, new_n1233_, new_n332_ );
or   ( new_n1235_, new_n317_, new_n515_ );
or   ( new_n1236_, new_n320_, new_n509_ );
and  ( new_n1237_, new_n1236_, new_n1235_ );
xor  ( new_n1238_, new_n1237_, new_n312_ );
or   ( new_n1239_, new_n1238_, new_n1234_ );
and  ( new_n1240_, new_n1238_, new_n1234_ );
or   ( new_n1241_, new_n283_, new_n805_ );
or   ( new_n1242_, new_n286_, new_n775_ );
and  ( new_n1243_, new_n1242_, new_n1241_ );
xor  ( new_n1244_, new_n1243_, new_n278_ );
or   ( new_n1245_, new_n1244_, new_n1240_ );
and  ( new_n1246_, new_n1245_, new_n1239_ );
or   ( new_n1247_, new_n1135_, new_n319_ );
or   ( new_n1248_, new_n1137_, new_n333_ );
and  ( new_n1249_, new_n1248_, new_n1247_ );
xor  ( new_n1250_, new_n1249_, new_n895_ );
xor  ( new_n1251_, RIbb2ebc0_23, RIbb2ec38_22 );
xor  ( new_n1252_, RIbb2ec38_22, new_n1126_ );
nor  ( new_n1253_, new_n1252_, new_n1251_ );
and  ( new_n1254_, new_n1253_, RIbb2d810_65 );
xor  ( new_n1255_, new_n1254_, new_n1129_ );
nand ( new_n1256_, new_n1255_, new_n1250_ );
nor  ( new_n1257_, new_n1255_, new_n1250_ );
or   ( new_n1258_, new_n897_, new_n285_ );
or   ( new_n1259_, new_n899_, new_n313_ );
and  ( new_n1260_, new_n1259_, new_n1258_ );
xor  ( new_n1261_, new_n1260_, new_n748_ );
or   ( new_n1262_, new_n1261_, new_n1257_ );
and  ( new_n1263_, new_n1262_, new_n1256_ );
nor  ( new_n1264_, new_n1263_, new_n1246_ );
and  ( new_n1265_, new_n1263_, new_n1246_ );
or   ( new_n1266_, new_n755_, new_n301_ );
or   ( new_n1267_, new_n757_, new_n279_ );
and  ( new_n1268_, new_n1267_, new_n1266_ );
xor  ( new_n1269_, new_n1268_, new_n523_ );
or   ( new_n1270_, new_n524_, new_n270_ );
or   ( new_n1271_, new_n526_, new_n294_ );
and  ( new_n1272_, new_n1271_, new_n1270_ );
xor  ( new_n1273_, new_n1272_, new_n403_ );
nor  ( new_n1274_, new_n1273_, new_n1269_ );
and  ( new_n1275_, new_n1273_, new_n1269_ );
or   ( new_n1276_, new_n409_, new_n348_ );
or   ( new_n1277_, new_n411_, new_n264_ );
and  ( new_n1278_, new_n1277_, new_n1276_ );
xor  ( new_n1279_, new_n1278_, new_n328_ );
nor  ( new_n1280_, new_n1279_, new_n1275_ );
nor  ( new_n1281_, new_n1280_, new_n1274_ );
nor  ( new_n1282_, new_n1281_, new_n1265_ );
nor  ( new_n1283_, new_n1282_, new_n1264_ );
xor  ( new_n1284_, new_n1133_, new_n1129_ );
xnor ( new_n1285_, new_n1284_, new_n1140_ );
xor  ( new_n1286_, new_n1117_, new_n1113_ );
xnor ( new_n1287_, new_n1286_, new_n1123_ );
nor  ( new_n1288_, new_n1287_, new_n1285_ );
and  ( new_n1289_, new_n1288_, new_n1283_ );
or   ( new_n1290_, new_n1289_, new_n1230_ );
or   ( new_n1291_, new_n1288_, new_n1283_ );
and  ( new_n1292_, new_n1291_, new_n1290_ );
or   ( new_n1293_, new_n1292_, new_n1208_ );
nand ( new_n1294_, new_n1292_, new_n1208_ );
xor  ( new_n1295_, new_n1143_, new_n1125_ );
xor  ( new_n1296_, new_n1295_, new_n1162_ );
xor  ( new_n1297_, new_n1182_, new_n1180_ );
xor  ( new_n1298_, new_n1297_, new_n1185_ );
nor  ( new_n1299_, new_n1298_, new_n1296_ );
and  ( new_n1300_, new_n1298_, new_n1296_ );
xor  ( new_n1301_, new_n1108_, new_n1106_ );
not  ( new_n1302_, new_n1301_ );
nor  ( new_n1303_, new_n1302_, new_n1300_ );
nor  ( new_n1304_, new_n1303_, new_n1299_ );
nand ( new_n1305_, new_n1304_, new_n1294_ );
and  ( new_n1306_, new_n1305_, new_n1293_ );
nand ( new_n1307_, new_n1306_, new_n1206_ );
nor  ( new_n1308_, new_n1306_, new_n1206_ );
xor  ( new_n1309_, new_n1102_, new_n1092_ );
xor  ( new_n1310_, new_n1309_, new_n1189_ );
or   ( new_n1311_, new_n1310_, new_n1308_ );
and  ( new_n1312_, new_n1311_, new_n1307_ );
nor  ( new_n1313_, new_n1312_, new_n1204_ );
xor  ( new_n1314_, new_n1199_, new_n1090_ );
and  ( new_n1315_, new_n1314_, new_n1313_ );
xor  ( new_n1316_, new_n1298_, new_n1296_ );
xor  ( new_n1317_, new_n1316_, new_n1302_ );
not  ( new_n1318_, RIbb2ce38_86 );
or   ( new_n1319_, new_n268_, new_n1318_ );
or   ( new_n1320_, new_n271_, new_n1213_ );
and  ( new_n1321_, new_n1320_, new_n1319_ );
xor  ( new_n1322_, new_n1321_, new_n263_ );
or   ( new_n1323_, new_n299_, new_n1168_ );
or   ( new_n1324_, new_n302_, new_n986_ );
and  ( new_n1325_, new_n1324_, new_n1323_ );
xor  ( new_n1326_, new_n1325_, new_n293_ );
and  ( new_n1327_, new_n1326_, new_n1322_ );
nor  ( new_n1328_, new_n1326_, new_n1322_ );
not  ( new_n1329_, new_n1328_ );
or   ( new_n1330_, new_n283_, new_n886_ );
or   ( new_n1331_, new_n286_, new_n805_ );
and  ( new_n1332_, new_n1331_, new_n1330_ );
xor  ( new_n1333_, new_n1332_, new_n278_ );
and  ( new_n1334_, new_n1333_, new_n1329_ );
nor  ( new_n1335_, new_n1334_, new_n1327_ );
xnor ( new_n1336_, new_n1217_, new_n1212_ );
xor  ( new_n1337_, new_n1336_, new_n1219_ );
nand ( new_n1338_, new_n1337_, new_n1335_ );
or   ( new_n1339_, new_n317_, new_n775_ );
or   ( new_n1340_, new_n320_, new_n515_ );
and  ( new_n1341_, new_n1340_, new_n1339_ );
xor  ( new_n1342_, new_n1341_, new_n312_ );
or   ( new_n1343_, new_n337_, new_n509_ );
or   ( new_n1344_, new_n340_, new_n443_ );
and  ( new_n1345_, new_n1344_, new_n1343_ );
xor  ( new_n1346_, new_n1345_, new_n332_ );
and  ( new_n1347_, new_n1346_, new_n1342_ );
or   ( new_n1348_, new_n1346_, new_n1342_ );
or   ( new_n1349_, new_n409_, new_n419_ );
or   ( new_n1350_, new_n411_, new_n348_ );
and  ( new_n1351_, new_n1350_, new_n1349_ );
xor  ( new_n1352_, new_n1351_, new_n328_ );
and  ( new_n1353_, new_n1352_, new_n1348_ );
or   ( new_n1354_, new_n1353_, new_n1347_ );
not  ( new_n1355_, RIbb2ebc0_23 );
and  ( new_n1356_, RIbb2ead0_25, RIbb2eb48_24 );
nor  ( new_n1357_, new_n1356_, new_n1355_ );
not  ( new_n1358_, new_n1357_ );
or   ( new_n1359_, new_n1135_, new_n313_ );
or   ( new_n1360_, new_n1137_, new_n319_ );
and  ( new_n1361_, new_n1360_, new_n1359_ );
xor  ( new_n1362_, new_n1361_, new_n896_ );
or   ( new_n1363_, new_n1362_, new_n1358_ );
not  ( new_n1364_, new_n1253_ );
or   ( new_n1365_, new_n1364_, new_n333_ );
not  ( new_n1366_, new_n1251_ );
or   ( new_n1367_, new_n1366_, new_n339_ );
and  ( new_n1368_, new_n1367_, new_n1365_ );
xor  ( new_n1369_, new_n1368_, new_n1129_ );
and  ( new_n1370_, new_n1362_, new_n1358_ );
or   ( new_n1371_, new_n1370_, new_n1369_ );
and  ( new_n1372_, new_n1371_, new_n1363_ );
or   ( new_n1373_, new_n1372_, new_n1354_ );
nand ( new_n1374_, new_n1372_, new_n1354_ );
or   ( new_n1375_, new_n524_, new_n264_ );
or   ( new_n1376_, new_n526_, new_n270_ );
and  ( new_n1377_, new_n1376_, new_n1375_ );
xor  ( new_n1378_, new_n1377_, new_n403_ );
or   ( new_n1379_, new_n755_, new_n294_ );
or   ( new_n1380_, new_n757_, new_n301_ );
and  ( new_n1381_, new_n1380_, new_n1379_ );
xor  ( new_n1382_, new_n1381_, new_n523_ );
and  ( new_n1383_, new_n1382_, new_n1378_ );
nor  ( new_n1384_, new_n1382_, new_n1378_ );
not  ( new_n1385_, new_n1384_ );
or   ( new_n1386_, new_n897_, new_n279_ );
or   ( new_n1387_, new_n899_, new_n285_ );
and  ( new_n1388_, new_n1387_, new_n1386_ );
xor  ( new_n1389_, new_n1388_, new_n748_ );
and  ( new_n1390_, new_n1389_, new_n1385_ );
nor  ( new_n1391_, new_n1390_, new_n1383_ );
nand ( new_n1392_, new_n1391_, new_n1374_ );
and  ( new_n1393_, new_n1392_, new_n1373_ );
nand ( new_n1394_, new_n1393_, new_n1338_ );
nor  ( new_n1395_, new_n1393_, new_n1338_ );
xnor ( new_n1396_, new_n1273_, new_n1269_ );
xor  ( new_n1397_, new_n1396_, new_n1279_ );
xnor ( new_n1398_, new_n1238_, new_n1234_ );
xor  ( new_n1399_, new_n1398_, new_n1244_ );
or   ( new_n1400_, new_n1399_, new_n1397_ );
and  ( new_n1401_, new_n1399_, new_n1397_ );
xor  ( new_n1402_, new_n1255_, new_n1250_ );
xnor ( new_n1403_, new_n1402_, new_n1261_ );
or   ( new_n1404_, new_n1403_, new_n1401_ );
and  ( new_n1405_, new_n1404_, new_n1400_ );
or   ( new_n1406_, new_n1405_, new_n1395_ );
and  ( new_n1407_, new_n1406_, new_n1394_ );
and  ( new_n1408_, new_n1407_, new_n1317_ );
xnor ( new_n1409_, new_n1287_, new_n1285_ );
xnor ( new_n1410_, new_n1224_, new_n1222_ );
xor  ( new_n1411_, new_n1410_, new_n1228_ );
nor  ( new_n1412_, new_n1411_, new_n1409_ );
and  ( new_n1413_, new_n1411_, new_n1409_ );
xor  ( new_n1414_, new_n1263_, new_n1246_ );
xnor ( new_n1415_, new_n1414_, new_n1281_ );
nor  ( new_n1416_, new_n1415_, new_n1413_ );
nor  ( new_n1417_, new_n1416_, new_n1412_ );
nor  ( new_n1418_, new_n1417_, new_n1408_ );
nor  ( new_n1419_, new_n1407_, new_n1317_ );
or   ( new_n1420_, new_n1419_, new_n1418_ );
xnor ( new_n1421_, new_n1164_, new_n1109_ );
xor  ( new_n1422_, new_n1421_, new_n1187_ );
nor  ( new_n1423_, new_n1422_, new_n1420_ );
nand ( new_n1424_, new_n1422_, new_n1420_ );
xor  ( new_n1425_, new_n1292_, new_n1208_ );
xor  ( new_n1426_, new_n1425_, new_n1304_ );
and  ( new_n1427_, new_n1426_, new_n1424_ );
or   ( new_n1428_, new_n1427_, new_n1423_ );
xor  ( new_n1429_, new_n1306_, new_n1206_ );
xor  ( new_n1430_, new_n1429_, new_n1310_ );
nor  ( new_n1431_, new_n1430_, new_n1428_ );
xor  ( new_n1432_, new_n1312_, new_n1204_ );
and  ( new_n1433_, new_n1432_, new_n1431_ );
xor  ( new_n1434_, new_n1407_, new_n1317_ );
xor  ( new_n1435_, new_n1434_, new_n1417_ );
xnor ( new_n1436_, new_n1288_, new_n1283_ );
xor  ( new_n1437_, new_n1436_, new_n1230_ );
or   ( new_n1438_, new_n1437_, new_n1435_ );
and  ( new_n1439_, new_n1437_, new_n1435_ );
xnor ( new_n1440_, new_n1411_, new_n1409_ );
xor  ( new_n1441_, new_n1440_, new_n1415_ );
xnor ( new_n1442_, new_n1337_, new_n1335_ );
xnor ( new_n1443_, new_n1399_, new_n1397_ );
xor  ( new_n1444_, new_n1443_, new_n1403_ );
or   ( new_n1445_, new_n1444_, new_n1442_ );
and  ( new_n1446_, new_n1444_, new_n1442_ );
xor  ( new_n1447_, new_n1372_, new_n1354_ );
xor  ( new_n1448_, new_n1447_, new_n1391_ );
not  ( new_n1449_, new_n1448_ );
or   ( new_n1450_, new_n1449_, new_n1446_ );
and  ( new_n1451_, new_n1450_, new_n1445_ );
and  ( new_n1452_, new_n1451_, new_n1441_ );
nor  ( new_n1453_, new_n1451_, new_n1441_ );
xor  ( new_n1454_, new_n1326_, new_n1322_ );
xor  ( new_n1455_, new_n1454_, new_n1333_ );
xor  ( new_n1456_, new_n1382_, new_n1378_ );
xor  ( new_n1457_, new_n1456_, new_n1389_ );
nor  ( new_n1458_, new_n1457_, new_n1455_ );
and  ( new_n1459_, new_n1457_, new_n1455_ );
xor  ( new_n1460_, new_n1346_, new_n1342_ );
xor  ( new_n1461_, new_n1460_, new_n1352_ );
nor  ( new_n1462_, new_n1461_, new_n1459_ );
or   ( new_n1463_, new_n1462_, new_n1458_ );
or   ( new_n1464_, new_n1135_, new_n285_ );
or   ( new_n1465_, new_n1137_, new_n313_ );
and  ( new_n1466_, new_n1465_, new_n1464_ );
xor  ( new_n1467_, new_n1466_, new_n896_ );
or   ( new_n1468_, new_n1364_, new_n319_ );
or   ( new_n1469_, new_n1366_, new_n333_ );
and  ( new_n1470_, new_n1469_, new_n1468_ );
xor  ( new_n1471_, new_n1470_, new_n1129_ );
and  ( new_n1472_, new_n1471_, new_n1467_ );
nor  ( new_n1473_, new_n1471_, new_n1467_ );
xor  ( new_n1474_, RIbb2ead0_25, RIbb2eb48_24 );
xor  ( new_n1475_, RIbb2eb48_24, new_n1355_ );
nor  ( new_n1476_, new_n1475_, new_n1474_ );
and  ( new_n1477_, new_n1476_, RIbb2d810_65 );
xor  ( new_n1478_, new_n1477_, new_n1358_ );
nor  ( new_n1479_, new_n1478_, new_n1473_ );
nor  ( new_n1480_, new_n1479_, new_n1472_ );
not  ( new_n1481_, new_n1480_ );
or   ( new_n1482_, new_n524_, new_n348_ );
or   ( new_n1483_, new_n526_, new_n264_ );
and  ( new_n1484_, new_n1483_, new_n1482_ );
xor  ( new_n1485_, new_n1484_, new_n403_ );
or   ( new_n1486_, new_n755_, new_n270_ );
or   ( new_n1487_, new_n757_, new_n294_ );
and  ( new_n1488_, new_n1487_, new_n1486_ );
xor  ( new_n1489_, new_n1488_, new_n523_ );
and  ( new_n1490_, new_n1489_, new_n1485_ );
nor  ( new_n1491_, new_n1489_, new_n1485_ );
not  ( new_n1492_, new_n1491_ );
or   ( new_n1493_, new_n897_, new_n301_ );
or   ( new_n1494_, new_n899_, new_n279_ );
and  ( new_n1495_, new_n1494_, new_n1493_ );
xor  ( new_n1496_, new_n1495_, new_n748_ );
and  ( new_n1497_, new_n1496_, new_n1492_ );
nor  ( new_n1498_, new_n1497_, new_n1490_ );
not  ( new_n1499_, new_n1498_ );
and  ( new_n1500_, new_n1499_, new_n1481_ );
and  ( new_n1501_, new_n1498_, new_n1480_ );
or   ( new_n1502_, new_n317_, new_n805_ );
or   ( new_n1503_, new_n320_, new_n775_ );
and  ( new_n1504_, new_n1503_, new_n1502_ );
xor  ( new_n1505_, new_n1504_, new_n312_ );
or   ( new_n1506_, new_n337_, new_n515_ );
or   ( new_n1507_, new_n340_, new_n509_ );
and  ( new_n1508_, new_n1507_, new_n1506_ );
xor  ( new_n1509_, new_n1508_, new_n332_ );
and  ( new_n1510_, new_n1509_, new_n1505_ );
nor  ( new_n1511_, new_n1509_, new_n1505_ );
or   ( new_n1512_, new_n409_, new_n443_ );
or   ( new_n1513_, new_n411_, new_n419_ );
and  ( new_n1514_, new_n1513_, new_n1512_ );
xor  ( new_n1515_, new_n1514_, new_n328_ );
not  ( new_n1516_, new_n1515_ );
nor  ( new_n1517_, new_n1516_, new_n1511_ );
nor  ( new_n1518_, new_n1517_, new_n1510_ );
nor  ( new_n1519_, new_n1518_, new_n1501_ );
nor  ( new_n1520_, new_n1519_, new_n1500_ );
nor  ( new_n1521_, new_n1520_, new_n1463_ );
and  ( new_n1522_, new_n1520_, new_n1463_ );
not  ( new_n1523_, RIbb2cd48_88 );
or   ( new_n1524_, new_n1523_, new_n260_ );
not  ( new_n1525_, RIbb2cdc0_87 );
or   ( new_n1526_, new_n268_, new_n1525_ );
or   ( new_n1527_, new_n271_, new_n1318_ );
and  ( new_n1528_, new_n1527_, new_n1526_ );
xor  ( new_n1529_, new_n1528_, new_n263_ );
or   ( new_n1530_, new_n299_, new_n1213_ );
or   ( new_n1531_, new_n302_, new_n1168_ );
and  ( new_n1532_, new_n1531_, new_n1530_ );
xor  ( new_n1533_, new_n1532_, new_n293_ );
nand ( new_n1534_, new_n1533_, new_n1529_ );
or   ( new_n1535_, new_n1533_, new_n1529_ );
or   ( new_n1536_, new_n283_, new_n986_ );
or   ( new_n1537_, new_n286_, new_n886_ );
and  ( new_n1538_, new_n1537_, new_n1536_ );
xor  ( new_n1539_, new_n1538_, new_n278_ );
nand ( new_n1540_, new_n1539_, new_n1535_ );
and  ( new_n1541_, new_n1540_, new_n1534_ );
nor  ( new_n1542_, new_n1541_, new_n1524_ );
and  ( new_n1543_, new_n1541_, new_n1524_ );
not  ( new_n1544_, new_n1543_ );
and  ( new_n1545_, RIbb2cdc0_87, RIbb2f610_1 );
and  ( new_n1546_, new_n1545_, new_n1544_ );
nor  ( new_n1547_, new_n1546_, new_n1542_ );
nor  ( new_n1548_, new_n1547_, new_n1522_ );
nor  ( new_n1549_, new_n1548_, new_n1521_ );
nor  ( new_n1550_, new_n1549_, new_n1453_ );
nor  ( new_n1551_, new_n1550_, new_n1452_ );
or   ( new_n1552_, new_n1551_, new_n1439_ );
and  ( new_n1553_, new_n1552_, new_n1438_ );
xor  ( new_n1554_, new_n1422_, new_n1420_ );
xor  ( new_n1555_, new_n1554_, new_n1426_ );
nor  ( new_n1556_, new_n1555_, new_n1553_ );
xor  ( new_n1557_, new_n1430_, new_n1428_ );
and  ( new_n1558_, new_n1557_, new_n1556_ );
xor  ( new_n1559_, new_n1393_, new_n1338_ );
xor  ( new_n1560_, new_n1559_, new_n1405_ );
xor  ( new_n1561_, new_n1533_, new_n1529_ );
xor  ( new_n1562_, new_n1561_, new_n1539_ );
or   ( new_n1563_, new_n1562_, new_n1524_ );
and  ( new_n1564_, new_n1562_, new_n1524_ );
or   ( new_n1565_, new_n317_, new_n886_ );
or   ( new_n1566_, new_n320_, new_n805_ );
and  ( new_n1567_, new_n1566_, new_n1565_ );
xor  ( new_n1568_, new_n1567_, new_n312_ );
or   ( new_n1569_, new_n283_, new_n1168_ );
or   ( new_n1570_, new_n286_, new_n986_ );
and  ( new_n1571_, new_n1570_, new_n1569_ );
xor  ( new_n1572_, new_n1571_, new_n278_ );
nor  ( new_n1573_, new_n1572_, new_n1568_ );
and  ( new_n1574_, new_n1572_, new_n1568_ );
or   ( new_n1575_, new_n299_, new_n1318_ );
or   ( new_n1576_, new_n302_, new_n1213_ );
and  ( new_n1577_, new_n1576_, new_n1575_ );
xor  ( new_n1578_, new_n1577_, new_n293_ );
nor  ( new_n1579_, new_n1578_, new_n1574_ );
nor  ( new_n1580_, new_n1579_, new_n1573_ );
or   ( new_n1581_, new_n1580_, new_n1564_ );
and  ( new_n1582_, new_n1581_, new_n1563_ );
not  ( new_n1583_, RIbb2ead0_25 );
and  ( new_n1584_, RIbb2e9e0_27, RIbb2ea58_26 );
nor  ( new_n1585_, new_n1584_, new_n1583_ );
not  ( new_n1586_, new_n1585_ );
or   ( new_n1587_, new_n1364_, new_n313_ );
or   ( new_n1588_, new_n1366_, new_n319_ );
and  ( new_n1589_, new_n1588_, new_n1587_ );
xor  ( new_n1590_, new_n1589_, new_n1129_ );
and  ( new_n1591_, new_n1590_, new_n1586_ );
or   ( new_n1592_, new_n1590_, new_n1586_ );
not  ( new_n1593_, new_n1476_ );
or   ( new_n1594_, new_n1593_, new_n333_ );
not  ( new_n1595_, new_n1474_ );
or   ( new_n1596_, new_n1595_, new_n339_ );
and  ( new_n1597_, new_n1596_, new_n1594_ );
xor  ( new_n1598_, new_n1597_, new_n1358_ );
and  ( new_n1599_, new_n1598_, new_n1592_ );
or   ( new_n1600_, new_n1599_, new_n1591_ );
or   ( new_n1601_, new_n1135_, new_n279_ );
or   ( new_n1602_, new_n1137_, new_n285_ );
and  ( new_n1603_, new_n1602_, new_n1601_ );
xor  ( new_n1604_, new_n1603_, new_n896_ );
or   ( new_n1605_, new_n897_, new_n294_ );
or   ( new_n1606_, new_n899_, new_n301_ );
and  ( new_n1607_, new_n1606_, new_n1605_ );
xor  ( new_n1608_, new_n1607_, new_n748_ );
or   ( new_n1609_, new_n1608_, new_n1604_ );
and  ( new_n1610_, new_n1608_, new_n1604_ );
or   ( new_n1611_, new_n755_, new_n264_ );
or   ( new_n1612_, new_n757_, new_n270_ );
and  ( new_n1613_, new_n1612_, new_n1611_ );
xor  ( new_n1614_, new_n1613_, new_n523_ );
or   ( new_n1615_, new_n1614_, new_n1610_ );
and  ( new_n1616_, new_n1615_, new_n1609_ );
or   ( new_n1617_, new_n1616_, new_n1600_ );
and  ( new_n1618_, new_n1616_, new_n1600_ );
or   ( new_n1619_, new_n524_, new_n419_ );
or   ( new_n1620_, new_n526_, new_n348_ );
and  ( new_n1621_, new_n1620_, new_n1619_ );
xor  ( new_n1622_, new_n1621_, new_n403_ );
or   ( new_n1623_, new_n409_, new_n509_ );
or   ( new_n1624_, new_n411_, new_n443_ );
and  ( new_n1625_, new_n1624_, new_n1623_ );
xor  ( new_n1626_, new_n1625_, new_n328_ );
nor  ( new_n1627_, new_n1626_, new_n1622_ );
and  ( new_n1628_, new_n1626_, new_n1622_ );
or   ( new_n1629_, new_n337_, new_n775_ );
or   ( new_n1630_, new_n340_, new_n515_ );
and  ( new_n1631_, new_n1630_, new_n1629_ );
xor  ( new_n1632_, new_n1631_, new_n332_ );
nor  ( new_n1633_, new_n1632_, new_n1628_ );
nor  ( new_n1634_, new_n1633_, new_n1627_ );
or   ( new_n1635_, new_n1634_, new_n1618_ );
and  ( new_n1636_, new_n1635_, new_n1617_ );
nor  ( new_n1637_, new_n1636_, new_n1582_ );
and  ( new_n1638_, new_n1636_, new_n1582_ );
xnor ( new_n1639_, new_n1471_, new_n1467_ );
xor  ( new_n1640_, new_n1639_, new_n1478_ );
xor  ( new_n1641_, new_n1489_, new_n1485_ );
xor  ( new_n1642_, new_n1641_, new_n1496_ );
nor  ( new_n1643_, new_n1642_, new_n1640_ );
and  ( new_n1644_, new_n1642_, new_n1640_ );
xor  ( new_n1645_, new_n1509_, new_n1505_ );
xor  ( new_n1646_, new_n1645_, new_n1515_ );
nor  ( new_n1647_, new_n1646_, new_n1644_ );
nor  ( new_n1648_, new_n1647_, new_n1643_ );
nor  ( new_n1649_, new_n1648_, new_n1638_ );
or   ( new_n1650_, new_n1649_, new_n1637_ );
xor  ( new_n1651_, new_n1444_, new_n1442_ );
xor  ( new_n1652_, new_n1651_, new_n1449_ );
not  ( new_n1653_, new_n1652_ );
or   ( new_n1654_, new_n1653_, new_n1650_ );
and  ( new_n1655_, new_n1653_, new_n1650_ );
xor  ( new_n1656_, new_n1457_, new_n1455_ );
xor  ( new_n1657_, new_n1656_, new_n1461_ );
xor  ( new_n1658_, new_n1541_, new_n1524_ );
xor  ( new_n1659_, new_n1658_, new_n1545_ );
nand ( new_n1660_, new_n1659_, new_n1657_ );
nor  ( new_n1661_, new_n1659_, new_n1657_ );
xor  ( new_n1662_, new_n1362_, new_n1358_ );
xnor ( new_n1663_, new_n1662_, new_n1369_ );
or   ( new_n1664_, new_n1663_, new_n1661_ );
and  ( new_n1665_, new_n1664_, new_n1660_ );
or   ( new_n1666_, new_n1665_, new_n1655_ );
and  ( new_n1667_, new_n1666_, new_n1654_ );
nand ( new_n1668_, new_n1667_, new_n1560_ );
xor  ( new_n1669_, new_n1451_, new_n1441_ );
xnor ( new_n1670_, new_n1669_, new_n1549_ );
and  ( new_n1671_, new_n1670_, new_n1668_ );
nor  ( new_n1672_, new_n1667_, new_n1560_ );
or   ( new_n1673_, new_n1672_, new_n1671_ );
xnor ( new_n1674_, new_n1437_, new_n1435_ );
xor  ( new_n1675_, new_n1674_, new_n1551_ );
and  ( new_n1676_, new_n1675_, new_n1673_ );
xor  ( new_n1677_, new_n1555_, new_n1553_ );
and  ( new_n1678_, new_n1677_, new_n1676_ );
xor  ( new_n1679_, new_n1636_, new_n1582_ );
xor  ( new_n1680_, new_n1679_, new_n1648_ );
xnor ( new_n1681_, new_n1659_, new_n1657_ );
xor  ( new_n1682_, new_n1681_, new_n1663_ );
nand ( new_n1683_, new_n1682_, new_n1680_ );
xor  ( new_n1684_, new_n1498_, new_n1481_ );
and  ( new_n1685_, new_n1684_, new_n1518_ );
not  ( new_n1686_, new_n1500_ );
and  ( new_n1687_, new_n1519_, new_n1686_ );
or   ( new_n1688_, new_n1687_, new_n1685_ );
xnor ( new_n1689_, new_n1642_, new_n1640_ );
xor  ( new_n1690_, new_n1689_, new_n1646_ );
xnor ( new_n1691_, new_n1562_, new_n1524_ );
xor  ( new_n1692_, new_n1691_, new_n1580_ );
or   ( new_n1693_, new_n1692_, new_n1690_ );
and  ( new_n1694_, new_n1692_, new_n1690_ );
xor  ( new_n1695_, new_n1616_, new_n1600_ );
xnor ( new_n1696_, new_n1695_, new_n1634_ );
or   ( new_n1697_, new_n1696_, new_n1694_ );
and  ( new_n1698_, new_n1697_, new_n1693_ );
or   ( new_n1699_, new_n1698_, new_n1688_ );
and  ( new_n1700_, new_n1698_, new_n1688_ );
or   ( new_n1701_, new_n1135_, new_n301_ );
or   ( new_n1702_, new_n1137_, new_n279_ );
and  ( new_n1703_, new_n1702_, new_n1701_ );
xor  ( new_n1704_, new_n1703_, new_n896_ );
or   ( new_n1705_, new_n897_, new_n270_ );
or   ( new_n1706_, new_n899_, new_n294_ );
and  ( new_n1707_, new_n1706_, new_n1705_ );
xor  ( new_n1708_, new_n1707_, new_n748_ );
or   ( new_n1709_, new_n1708_, new_n1704_ );
and  ( new_n1710_, new_n1708_, new_n1704_ );
or   ( new_n1711_, new_n755_, new_n348_ );
or   ( new_n1712_, new_n757_, new_n264_ );
and  ( new_n1713_, new_n1712_, new_n1711_ );
xor  ( new_n1714_, new_n1713_, new_n523_ );
or   ( new_n1715_, new_n1714_, new_n1710_ );
and  ( new_n1716_, new_n1715_, new_n1709_ );
or   ( new_n1717_, new_n524_, new_n443_ );
or   ( new_n1718_, new_n526_, new_n419_ );
and  ( new_n1719_, new_n1718_, new_n1717_ );
xor  ( new_n1720_, new_n1719_, new_n403_ );
or   ( new_n1721_, new_n409_, new_n515_ );
or   ( new_n1722_, new_n411_, new_n509_ );
and  ( new_n1723_, new_n1722_, new_n1721_ );
xor  ( new_n1724_, new_n1723_, new_n328_ );
or   ( new_n1725_, new_n1724_, new_n1720_ );
and  ( new_n1726_, new_n1724_, new_n1720_ );
or   ( new_n1727_, new_n337_, new_n805_ );
or   ( new_n1728_, new_n340_, new_n775_ );
and  ( new_n1729_, new_n1728_, new_n1727_ );
xor  ( new_n1730_, new_n1729_, new_n332_ );
or   ( new_n1731_, new_n1730_, new_n1726_ );
and  ( new_n1732_, new_n1731_, new_n1725_ );
or   ( new_n1733_, new_n1732_, new_n1716_ );
and  ( new_n1734_, new_n1732_, new_n1716_ );
or   ( new_n1735_, new_n1593_, new_n319_ );
or   ( new_n1736_, new_n1595_, new_n333_ );
and  ( new_n1737_, new_n1736_, new_n1735_ );
xor  ( new_n1738_, new_n1737_, new_n1357_ );
xor  ( new_n1739_, RIbb2e9e0_27, RIbb2ea58_26 );
xor  ( new_n1740_, RIbb2ea58_26, new_n1583_ );
nor  ( new_n1741_, new_n1740_, new_n1739_ );
and  ( new_n1742_, new_n1741_, RIbb2d810_65 );
xor  ( new_n1743_, new_n1742_, new_n1586_ );
nand ( new_n1744_, new_n1743_, new_n1738_ );
nor  ( new_n1745_, new_n1743_, new_n1738_ );
or   ( new_n1746_, new_n1364_, new_n285_ );
or   ( new_n1747_, new_n1366_, new_n313_ );
and  ( new_n1748_, new_n1747_, new_n1746_ );
xor  ( new_n1749_, new_n1748_, new_n1129_ );
or   ( new_n1750_, new_n1749_, new_n1745_ );
and  ( new_n1751_, new_n1750_, new_n1744_ );
or   ( new_n1752_, new_n1751_, new_n1734_ );
and  ( new_n1753_, new_n1752_, new_n1733_ );
not  ( new_n1754_, RIbb2ccd0_89 );
or   ( new_n1755_, new_n1754_, new_n260_ );
xnor ( new_n1756_, new_n1626_, new_n1622_ );
xor  ( new_n1757_, new_n1756_, new_n1632_ );
nand ( new_n1758_, new_n1757_, new_n1755_ );
nor  ( new_n1759_, new_n1757_, new_n1755_ );
xor  ( new_n1760_, new_n1572_, new_n1568_ );
xor  ( new_n1761_, new_n1760_, new_n1578_ );
or   ( new_n1762_, new_n1761_, new_n1759_ );
and  ( new_n1763_, new_n1762_, new_n1758_ );
and  ( new_n1764_, new_n1763_, new_n1753_ );
nor  ( new_n1765_, new_n1763_, new_n1753_ );
or   ( new_n1766_, new_n268_, new_n1754_ );
or   ( new_n1767_, new_n271_, new_n1523_ );
and  ( new_n1768_, new_n1767_, new_n1766_ );
xor  ( new_n1769_, new_n1768_, new_n263_ );
and  ( new_n1770_, RIbb2cc58_90, RIbb2f610_1 );
or   ( new_n1771_, new_n1770_, new_n1769_ );
or   ( new_n1772_, new_n317_, new_n986_ );
or   ( new_n1773_, new_n320_, new_n886_ );
and  ( new_n1774_, new_n1773_, new_n1772_ );
xor  ( new_n1775_, new_n1774_, new_n312_ );
or   ( new_n1776_, new_n283_, new_n1213_ );
or   ( new_n1777_, new_n286_, new_n1168_ );
and  ( new_n1778_, new_n1777_, new_n1776_ );
xor  ( new_n1779_, new_n1778_, new_n278_ );
or   ( new_n1780_, new_n1779_, new_n1775_ );
and  ( new_n1781_, new_n1779_, new_n1775_ );
or   ( new_n1782_, new_n299_, new_n1525_ );
or   ( new_n1783_, new_n302_, new_n1318_ );
and  ( new_n1784_, new_n1783_, new_n1782_ );
xor  ( new_n1785_, new_n1784_, new_n293_ );
or   ( new_n1786_, new_n1785_, new_n1781_ );
and  ( new_n1787_, new_n1786_, new_n1780_ );
and  ( new_n1788_, new_n1787_, new_n1771_ );
nor  ( new_n1789_, new_n1787_, new_n1771_ );
or   ( new_n1790_, new_n268_, new_n1523_ );
or   ( new_n1791_, new_n271_, new_n1525_ );
and  ( new_n1792_, new_n1791_, new_n1790_ );
xor  ( new_n1793_, new_n1792_, new_n263_ );
not  ( new_n1794_, new_n1793_ );
nor  ( new_n1795_, new_n1794_, new_n1789_ );
nor  ( new_n1796_, new_n1795_, new_n1788_ );
nor  ( new_n1797_, new_n1796_, new_n1765_ );
nor  ( new_n1798_, new_n1797_, new_n1764_ );
or   ( new_n1799_, new_n1798_, new_n1700_ );
and  ( new_n1800_, new_n1799_, new_n1699_ );
nor  ( new_n1801_, new_n1800_, new_n1683_ );
and  ( new_n1802_, new_n1800_, new_n1683_ );
not  ( new_n1803_, new_n1802_ );
xor  ( new_n1804_, new_n1520_, new_n1463_ );
xnor ( new_n1805_, new_n1804_, new_n1547_ );
and  ( new_n1806_, new_n1805_, new_n1803_ );
nor  ( new_n1807_, new_n1806_, new_n1801_ );
xnor ( new_n1808_, new_n1667_, new_n1560_ );
xor  ( new_n1809_, new_n1808_, new_n1670_ );
nor  ( new_n1810_, new_n1809_, new_n1807_ );
xor  ( new_n1811_, new_n1675_, new_n1673_ );
and  ( new_n1812_, new_n1811_, new_n1810_ );
xnor ( new_n1813_, new_n1809_, new_n1807_ );
xor  ( new_n1814_, new_n1652_, new_n1650_ );
xor  ( new_n1815_, new_n1814_, new_n1665_ );
xor  ( new_n1816_, new_n1800_, new_n1683_ );
xor  ( new_n1817_, new_n1816_, new_n1805_ );
nand ( new_n1818_, new_n1817_, new_n1815_ );
nor  ( new_n1819_, new_n1817_, new_n1815_ );
xor  ( new_n1820_, new_n1682_, new_n1680_ );
xnor ( new_n1821_, new_n1698_, new_n1688_ );
xor  ( new_n1822_, new_n1821_, new_n1798_ );
nand ( new_n1823_, new_n1822_, new_n1820_ );
nor  ( new_n1824_, new_n1822_, new_n1820_ );
xor  ( new_n1825_, new_n1757_, new_n1755_ );
xor  ( new_n1826_, new_n1825_, new_n1761_ );
xor  ( new_n1827_, new_n1590_, new_n1586_ );
xor  ( new_n1828_, new_n1827_, new_n1598_ );
and  ( new_n1829_, new_n1828_, new_n1826_ );
or   ( new_n1830_, new_n1828_, new_n1826_ );
xor  ( new_n1831_, new_n1608_, new_n1604_ );
xnor ( new_n1832_, new_n1831_, new_n1614_ );
not  ( new_n1833_, new_n1832_ );
and  ( new_n1834_, new_n1833_, new_n1830_ );
or   ( new_n1835_, new_n1834_, new_n1829_ );
xnor ( new_n1836_, new_n1692_, new_n1690_ );
xor  ( new_n1837_, new_n1836_, new_n1696_ );
and  ( new_n1838_, new_n1837_, new_n1835_ );
nor  ( new_n1839_, new_n1837_, new_n1835_ );
not  ( new_n1840_, RIbb2e9e0_27 );
and  ( new_n1841_, RIbb2e8f0_29, RIbb2e968_28 );
nor  ( new_n1842_, new_n1841_, new_n1840_ );
not  ( new_n1843_, new_n1842_ );
not  ( new_n1844_, new_n1741_ );
or   ( new_n1845_, new_n1844_, new_n333_ );
not  ( new_n1846_, new_n1739_ );
or   ( new_n1847_, new_n1846_, new_n339_ );
and  ( new_n1848_, new_n1847_, new_n1845_ );
xor  ( new_n1849_, new_n1848_, new_n1586_ );
and  ( new_n1850_, new_n1849_, new_n1843_ );
or   ( new_n1851_, new_n1849_, new_n1843_ );
or   ( new_n1852_, new_n1593_, new_n313_ );
or   ( new_n1853_, new_n1595_, new_n319_ );
and  ( new_n1854_, new_n1853_, new_n1852_ );
xor  ( new_n1855_, new_n1854_, new_n1358_ );
and  ( new_n1856_, new_n1855_, new_n1851_ );
or   ( new_n1857_, new_n1856_, new_n1850_ );
or   ( new_n1858_, new_n1364_, new_n279_ );
or   ( new_n1859_, new_n1366_, new_n285_ );
and  ( new_n1860_, new_n1859_, new_n1858_ );
xor  ( new_n1861_, new_n1860_, new_n1129_ );
or   ( new_n1862_, new_n1135_, new_n294_ );
or   ( new_n1863_, new_n1137_, new_n301_ );
and  ( new_n1864_, new_n1863_, new_n1862_ );
xor  ( new_n1865_, new_n1864_, new_n896_ );
or   ( new_n1866_, new_n1865_, new_n1861_ );
and  ( new_n1867_, new_n1865_, new_n1861_ );
or   ( new_n1868_, new_n897_, new_n264_ );
or   ( new_n1869_, new_n899_, new_n270_ );
and  ( new_n1870_, new_n1869_, new_n1868_ );
xor  ( new_n1871_, new_n1870_, new_n748_ );
or   ( new_n1872_, new_n1871_, new_n1867_ );
and  ( new_n1873_, new_n1872_, new_n1866_ );
or   ( new_n1874_, new_n1873_, new_n1857_ );
and  ( new_n1875_, new_n1873_, new_n1857_ );
or   ( new_n1876_, new_n755_, new_n419_ );
or   ( new_n1877_, new_n757_, new_n348_ );
and  ( new_n1878_, new_n1877_, new_n1876_ );
xor  ( new_n1879_, new_n1878_, new_n523_ );
or   ( new_n1880_, new_n524_, new_n509_ );
or   ( new_n1881_, new_n526_, new_n443_ );
and  ( new_n1882_, new_n1881_, new_n1880_ );
xor  ( new_n1883_, new_n1882_, new_n403_ );
nor  ( new_n1884_, new_n1883_, new_n1879_ );
and  ( new_n1885_, new_n1883_, new_n1879_ );
or   ( new_n1886_, new_n409_, new_n775_ );
or   ( new_n1887_, new_n411_, new_n515_ );
and  ( new_n1888_, new_n1887_, new_n1886_ );
xor  ( new_n1889_, new_n1888_, new_n328_ );
nor  ( new_n1890_, new_n1889_, new_n1885_ );
nor  ( new_n1891_, new_n1890_, new_n1884_ );
or   ( new_n1892_, new_n1891_, new_n1875_ );
and  ( new_n1893_, new_n1892_, new_n1874_ );
xnor ( new_n1894_, new_n1770_, new_n1769_ );
or   ( new_n1895_, new_n299_, new_n1523_ );
or   ( new_n1896_, new_n302_, new_n1525_ );
and  ( new_n1897_, new_n1896_, new_n1895_ );
xor  ( new_n1898_, new_n1897_, new_n293_ );
not  ( new_n1899_, RIbb2cc58_90 );
or   ( new_n1900_, new_n268_, new_n1899_ );
or   ( new_n1901_, new_n271_, new_n1754_ );
and  ( new_n1902_, new_n1901_, new_n1900_ );
xor  ( new_n1903_, new_n1902_, new_n263_ );
or   ( new_n1904_, new_n1903_, new_n1898_ );
and  ( new_n1905_, RIbb2cbe0_91, RIbb2f610_1 );
and  ( new_n1906_, new_n1903_, new_n1898_ );
or   ( new_n1907_, new_n1906_, new_n1905_ );
and  ( new_n1908_, new_n1907_, new_n1904_ );
or   ( new_n1909_, new_n1908_, new_n1894_ );
and  ( new_n1910_, new_n1908_, new_n1894_ );
or   ( new_n1911_, new_n337_, new_n886_ );
or   ( new_n1912_, new_n340_, new_n805_ );
and  ( new_n1913_, new_n1912_, new_n1911_ );
xor  ( new_n1914_, new_n1913_, new_n332_ );
or   ( new_n1915_, new_n317_, new_n1168_ );
or   ( new_n1916_, new_n320_, new_n986_ );
and  ( new_n1917_, new_n1916_, new_n1915_ );
xor  ( new_n1918_, new_n1917_, new_n312_ );
nor  ( new_n1919_, new_n1918_, new_n1914_ );
and  ( new_n1920_, new_n1918_, new_n1914_ );
or   ( new_n1921_, new_n283_, new_n1318_ );
or   ( new_n1922_, new_n286_, new_n1213_ );
and  ( new_n1923_, new_n1922_, new_n1921_ );
xor  ( new_n1924_, new_n1923_, new_n278_ );
nor  ( new_n1925_, new_n1924_, new_n1920_ );
nor  ( new_n1926_, new_n1925_, new_n1919_ );
or   ( new_n1927_, new_n1926_, new_n1910_ );
and  ( new_n1928_, new_n1927_, new_n1909_ );
and  ( new_n1929_, new_n1928_, new_n1893_ );
nor  ( new_n1930_, new_n1928_, new_n1893_ );
xnor ( new_n1931_, new_n1724_, new_n1720_ );
xor  ( new_n1932_, new_n1931_, new_n1730_ );
xnor ( new_n1933_, new_n1708_, new_n1704_ );
xor  ( new_n1934_, new_n1933_, new_n1714_ );
nor  ( new_n1935_, new_n1934_, new_n1932_ );
and  ( new_n1936_, new_n1934_, new_n1932_ );
xor  ( new_n1937_, new_n1779_, new_n1775_ );
xnor ( new_n1938_, new_n1937_, new_n1785_ );
nor  ( new_n1939_, new_n1938_, new_n1936_ );
nor  ( new_n1940_, new_n1939_, new_n1935_ );
nor  ( new_n1941_, new_n1940_, new_n1930_ );
nor  ( new_n1942_, new_n1941_, new_n1929_ );
nor  ( new_n1943_, new_n1942_, new_n1839_ );
nor  ( new_n1944_, new_n1943_, new_n1838_ );
or   ( new_n1945_, new_n1944_, new_n1824_ );
and  ( new_n1946_, new_n1945_, new_n1823_ );
or   ( new_n1947_, new_n1946_, new_n1819_ );
and  ( new_n1948_, new_n1947_, new_n1818_ );
nor  ( new_n1949_, new_n1948_, new_n1813_ );
xor  ( new_n1950_, new_n1817_, new_n1815_ );
xor  ( new_n1951_, new_n1950_, new_n1946_ );
xor  ( new_n1952_, new_n1732_, new_n1716_ );
xor  ( new_n1953_, new_n1952_, new_n1751_ );
xnor ( new_n1954_, new_n1928_, new_n1893_ );
xor  ( new_n1955_, new_n1954_, new_n1940_ );
and  ( new_n1956_, new_n1955_, new_n1953_ );
nor  ( new_n1957_, new_n1955_, new_n1953_ );
not  ( new_n1958_, new_n1957_ );
xor  ( new_n1959_, new_n1828_, new_n1826_ );
xor  ( new_n1960_, new_n1959_, new_n1833_ );
and  ( new_n1961_, new_n1960_, new_n1958_ );
nor  ( new_n1962_, new_n1961_, new_n1956_ );
xnor ( new_n1963_, new_n1763_, new_n1753_ );
xor  ( new_n1964_, new_n1963_, new_n1796_ );
xor  ( new_n1965_, new_n1964_, new_n1962_ );
xor  ( new_n1966_, new_n1787_, new_n1771_ );
xor  ( new_n1967_, new_n1966_, new_n1794_ );
xor  ( new_n1968_, new_n1743_, new_n1738_ );
xor  ( new_n1969_, new_n1968_, new_n1749_ );
xnor ( new_n1970_, new_n1934_, new_n1932_ );
xor  ( new_n1971_, new_n1970_, new_n1938_ );
nand ( new_n1972_, new_n1971_, new_n1969_ );
nor  ( new_n1973_, new_n1971_, new_n1969_ );
xor  ( new_n1974_, new_n1908_, new_n1894_ );
xnor ( new_n1975_, new_n1974_, new_n1926_ );
or   ( new_n1976_, new_n1975_, new_n1973_ );
and  ( new_n1977_, new_n1976_, new_n1972_ );
or   ( new_n1978_, new_n1977_, new_n1967_ );
and  ( new_n1979_, new_n1977_, new_n1967_ );
or   ( new_n1980_, new_n1364_, new_n301_ );
or   ( new_n1981_, new_n1366_, new_n279_ );
and  ( new_n1982_, new_n1981_, new_n1980_ );
xor  ( new_n1983_, new_n1982_, new_n1129_ );
or   ( new_n1984_, new_n1135_, new_n270_ );
or   ( new_n1985_, new_n1137_, new_n294_ );
and  ( new_n1986_, new_n1985_, new_n1984_ );
xor  ( new_n1987_, new_n1986_, new_n896_ );
or   ( new_n1988_, new_n1987_, new_n1983_ );
and  ( new_n1989_, new_n1987_, new_n1983_ );
or   ( new_n1990_, new_n897_, new_n348_ );
or   ( new_n1991_, new_n899_, new_n264_ );
and  ( new_n1992_, new_n1991_, new_n1990_ );
xor  ( new_n1993_, new_n1992_, new_n748_ );
or   ( new_n1994_, new_n1993_, new_n1989_ );
and  ( new_n1995_, new_n1994_, new_n1988_ );
or   ( new_n1996_, new_n1844_, new_n319_ );
or   ( new_n1997_, new_n1846_, new_n333_ );
and  ( new_n1998_, new_n1997_, new_n1996_ );
xor  ( new_n1999_, new_n1998_, new_n1585_ );
xor  ( new_n2000_, RIbb2e8f0_29, RIbb2e968_28 );
xor  ( new_n2001_, RIbb2e968_28, new_n1840_ );
nor  ( new_n2002_, new_n2001_, new_n2000_ );
and  ( new_n2003_, new_n2002_, RIbb2d810_65 );
xor  ( new_n2004_, new_n2003_, new_n1843_ );
nand ( new_n2005_, new_n2004_, new_n1999_ );
nor  ( new_n2006_, new_n2004_, new_n1999_ );
or   ( new_n2007_, new_n1593_, new_n285_ );
or   ( new_n2008_, new_n1595_, new_n313_ );
and  ( new_n2009_, new_n2008_, new_n2007_ );
xor  ( new_n2010_, new_n2009_, new_n1358_ );
or   ( new_n2011_, new_n2010_, new_n2006_ );
and  ( new_n2012_, new_n2011_, new_n2005_ );
or   ( new_n2013_, new_n2012_, new_n1995_ );
and  ( new_n2014_, new_n2012_, new_n1995_ );
or   ( new_n2015_, new_n755_, new_n443_ );
or   ( new_n2016_, new_n757_, new_n419_ );
and  ( new_n2017_, new_n2016_, new_n2015_ );
xor  ( new_n2018_, new_n2017_, new_n523_ );
or   ( new_n2019_, new_n524_, new_n515_ );
or   ( new_n2020_, new_n526_, new_n509_ );
and  ( new_n2021_, new_n2020_, new_n2019_ );
xor  ( new_n2022_, new_n2021_, new_n403_ );
nor  ( new_n2023_, new_n2022_, new_n2018_ );
and  ( new_n2024_, new_n2022_, new_n2018_ );
or   ( new_n2025_, new_n409_, new_n805_ );
or   ( new_n2026_, new_n411_, new_n775_ );
and  ( new_n2027_, new_n2026_, new_n2025_ );
xor  ( new_n2028_, new_n2027_, new_n328_ );
nor  ( new_n2029_, new_n2028_, new_n2024_ );
nor  ( new_n2030_, new_n2029_, new_n2023_ );
or   ( new_n2031_, new_n2030_, new_n2014_ );
and  ( new_n2032_, new_n2031_, new_n2013_ );
xor  ( new_n2033_, new_n1903_, new_n1898_ );
xor  ( new_n2034_, new_n2033_, new_n1905_ );
or   ( new_n2035_, new_n337_, new_n986_ );
or   ( new_n2036_, new_n340_, new_n886_ );
and  ( new_n2037_, new_n2036_, new_n2035_ );
xor  ( new_n2038_, new_n2037_, new_n332_ );
or   ( new_n2039_, new_n317_, new_n1213_ );
or   ( new_n2040_, new_n320_, new_n1168_ );
and  ( new_n2041_, new_n2040_, new_n2039_ );
xor  ( new_n2042_, new_n2041_, new_n312_ );
or   ( new_n2043_, new_n2042_, new_n2038_ );
and  ( new_n2044_, new_n2042_, new_n2038_ );
or   ( new_n2045_, new_n283_, new_n1525_ );
or   ( new_n2046_, new_n286_, new_n1318_ );
and  ( new_n2047_, new_n2046_, new_n2045_ );
xor  ( new_n2048_, new_n2047_, new_n278_ );
or   ( new_n2049_, new_n2048_, new_n2044_ );
and  ( new_n2050_, new_n2049_, new_n2043_ );
or   ( new_n2051_, new_n2050_, new_n2034_ );
and  ( new_n2052_, new_n2050_, new_n2034_ );
or   ( new_n2053_, new_n299_, new_n1754_ );
or   ( new_n2054_, new_n302_, new_n1523_ );
and  ( new_n2055_, new_n2054_, new_n2053_ );
xor  ( new_n2056_, new_n2055_, new_n293_ );
not  ( new_n2057_, RIbb2cbe0_91 );
or   ( new_n2058_, new_n268_, new_n2057_ );
or   ( new_n2059_, new_n271_, new_n1899_ );
and  ( new_n2060_, new_n2059_, new_n2058_ );
xor  ( new_n2061_, new_n2060_, new_n263_ );
nor  ( new_n2062_, new_n2061_, new_n2056_ );
and  ( new_n2063_, RIbb2cb68_92, RIbb2f610_1 );
and  ( new_n2064_, new_n2061_, new_n2056_ );
nor  ( new_n2065_, new_n2064_, new_n2063_ );
nor  ( new_n2066_, new_n2065_, new_n2062_ );
or   ( new_n2067_, new_n2066_, new_n2052_ );
and  ( new_n2068_, new_n2067_, new_n2051_ );
and  ( new_n2069_, new_n2068_, new_n2032_ );
nor  ( new_n2070_, new_n2068_, new_n2032_ );
xnor ( new_n2071_, new_n1865_, new_n1861_ );
xor  ( new_n2072_, new_n2071_, new_n1871_ );
xnor ( new_n2073_, new_n1918_, new_n1914_ );
xor  ( new_n2074_, new_n2073_, new_n1924_ );
nor  ( new_n2075_, new_n2074_, new_n2072_ );
and  ( new_n2076_, new_n2074_, new_n2072_ );
xor  ( new_n2077_, new_n1883_, new_n1879_ );
xnor ( new_n2078_, new_n2077_, new_n1889_ );
nor  ( new_n2079_, new_n2078_, new_n2076_ );
nor  ( new_n2080_, new_n2079_, new_n2075_ );
nor  ( new_n2081_, new_n2080_, new_n2070_ );
nor  ( new_n2082_, new_n2081_, new_n2069_ );
or   ( new_n2083_, new_n2082_, new_n1979_ );
and  ( new_n2084_, new_n2083_, new_n1978_ );
xor  ( new_n2085_, new_n2084_, new_n1965_ );
xnor ( new_n2086_, new_n1837_, new_n1835_ );
xor  ( new_n2087_, new_n2086_, new_n1942_ );
or   ( new_n2088_, new_n2087_, new_n2085_ );
and  ( new_n2089_, new_n2087_, new_n2085_ );
xor  ( new_n2090_, new_n1955_, new_n1953_ );
xor  ( new_n2091_, new_n2090_, new_n1960_ );
xor  ( new_n2092_, new_n2074_, new_n2072_ );
xor  ( new_n2093_, new_n2092_, new_n2078_ );
xnor ( new_n2094_, new_n2050_, new_n2034_ );
xor  ( new_n2095_, new_n2094_, new_n2066_ );
nor  ( new_n2096_, new_n2095_, new_n2093_ );
nand ( new_n2097_, new_n2095_, new_n2093_ );
xor  ( new_n2098_, new_n1849_, new_n1843_ );
xor  ( new_n2099_, new_n2098_, new_n1855_ );
and  ( new_n2100_, new_n2099_, new_n2097_ );
or   ( new_n2101_, new_n2100_, new_n2096_ );
or   ( new_n2102_, new_n1593_, new_n279_ );
or   ( new_n2103_, new_n1595_, new_n285_ );
and  ( new_n2104_, new_n2103_, new_n2102_ );
xor  ( new_n2105_, new_n2104_, new_n1358_ );
or   ( new_n2106_, new_n1364_, new_n294_ );
or   ( new_n2107_, new_n1366_, new_n301_ );
and  ( new_n2108_, new_n2107_, new_n2106_ );
xor  ( new_n2109_, new_n2108_, new_n1129_ );
nor  ( new_n2110_, new_n2109_, new_n2105_ );
and  ( new_n2111_, new_n2109_, new_n2105_ );
or   ( new_n2112_, new_n1135_, new_n264_ );
or   ( new_n2113_, new_n1137_, new_n270_ );
and  ( new_n2114_, new_n2113_, new_n2112_ );
xor  ( new_n2115_, new_n2114_, new_n896_ );
nor  ( new_n2116_, new_n2115_, new_n2111_ );
or   ( new_n2117_, new_n2116_, new_n2110_ );
not  ( new_n2118_, RIbb2e8f0_29 );
and  ( new_n2119_, RIbb2e800_31, RIbb2e878_30 );
nor  ( new_n2120_, new_n2119_, new_n2118_ );
not  ( new_n2121_, new_n2120_ );
not  ( new_n2122_, new_n2002_ );
or   ( new_n2123_, new_n2122_, new_n333_ );
not  ( new_n2124_, new_n2000_ );
or   ( new_n2125_, new_n2124_, new_n339_ );
and  ( new_n2126_, new_n2125_, new_n2123_ );
xor  ( new_n2127_, new_n2126_, new_n1843_ );
nand ( new_n2128_, new_n2127_, new_n2121_ );
or   ( new_n2129_, new_n2127_, new_n2121_ );
or   ( new_n2130_, new_n1844_, new_n313_ );
or   ( new_n2131_, new_n1846_, new_n319_ );
and  ( new_n2132_, new_n2131_, new_n2130_ );
xor  ( new_n2133_, new_n2132_, new_n1586_ );
nand ( new_n2134_, new_n2133_, new_n2129_ );
and  ( new_n2135_, new_n2134_, new_n2128_ );
and  ( new_n2136_, new_n2135_, new_n2117_ );
nor  ( new_n2137_, new_n2135_, new_n2117_ );
or   ( new_n2138_, new_n897_, new_n419_ );
or   ( new_n2139_, new_n899_, new_n348_ );
and  ( new_n2140_, new_n2139_, new_n2138_ );
xor  ( new_n2141_, new_n2140_, new_n748_ );
or   ( new_n2142_, new_n755_, new_n509_ );
or   ( new_n2143_, new_n757_, new_n443_ );
and  ( new_n2144_, new_n2143_, new_n2142_ );
xor  ( new_n2145_, new_n2144_, new_n523_ );
nor  ( new_n2146_, new_n2145_, new_n2141_ );
and  ( new_n2147_, new_n2145_, new_n2141_ );
or   ( new_n2148_, new_n524_, new_n775_ );
or   ( new_n2149_, new_n526_, new_n515_ );
and  ( new_n2150_, new_n2149_, new_n2148_ );
xor  ( new_n2151_, new_n2150_, new_n403_ );
nor  ( new_n2152_, new_n2151_, new_n2147_ );
nor  ( new_n2153_, new_n2152_, new_n2146_ );
nor  ( new_n2154_, new_n2153_, new_n2137_ );
or   ( new_n2155_, new_n2154_, new_n2136_ );
xnor ( new_n2156_, new_n2042_, new_n2038_ );
xor  ( new_n2157_, new_n2156_, new_n2048_ );
xnor ( new_n2158_, new_n2061_, new_n2056_ );
xor  ( new_n2159_, new_n2158_, new_n2063_ );
or   ( new_n2160_, new_n2159_, new_n2157_ );
and  ( new_n2161_, new_n2159_, new_n2157_ );
xor  ( new_n2162_, new_n2022_, new_n2018_ );
xnor ( new_n2163_, new_n2162_, new_n2028_ );
or   ( new_n2164_, new_n2163_, new_n2161_ );
and  ( new_n2165_, new_n2164_, new_n2160_ );
nand ( new_n2166_, new_n2165_, new_n2155_ );
or   ( new_n2167_, new_n2165_, new_n2155_ );
or   ( new_n2168_, new_n283_, new_n1523_ );
or   ( new_n2169_, new_n286_, new_n1525_ );
and  ( new_n2170_, new_n2169_, new_n2168_ );
xor  ( new_n2171_, new_n2170_, new_n278_ );
or   ( new_n2172_, new_n299_, new_n1899_ );
or   ( new_n2173_, new_n302_, new_n1754_ );
and  ( new_n2174_, new_n2173_, new_n2172_ );
xor  ( new_n2175_, new_n2174_, new_n293_ );
nor  ( new_n2176_, new_n2175_, new_n2171_ );
and  ( new_n2177_, new_n2175_, new_n2171_ );
not  ( new_n2178_, RIbb2cb68_92 );
or   ( new_n2179_, new_n268_, new_n2178_ );
or   ( new_n2180_, new_n271_, new_n2057_ );
and  ( new_n2181_, new_n2180_, new_n2179_ );
xor  ( new_n2182_, new_n2181_, new_n263_ );
nor  ( new_n2183_, new_n2182_, new_n2177_ );
nor  ( new_n2184_, new_n2183_, new_n2176_ );
or   ( new_n2185_, new_n409_, new_n886_ );
or   ( new_n2186_, new_n411_, new_n805_ );
and  ( new_n2187_, new_n2186_, new_n2185_ );
xor  ( new_n2188_, new_n2187_, new_n328_ );
or   ( new_n2189_, new_n337_, new_n1168_ );
or   ( new_n2190_, new_n340_, new_n986_ );
and  ( new_n2191_, new_n2190_, new_n2189_ );
xor  ( new_n2192_, new_n2191_, new_n332_ );
or   ( new_n2193_, new_n2192_, new_n2188_ );
and  ( new_n2194_, new_n2192_, new_n2188_ );
or   ( new_n2195_, new_n317_, new_n1318_ );
or   ( new_n2196_, new_n320_, new_n1213_ );
and  ( new_n2197_, new_n2196_, new_n2195_ );
xor  ( new_n2198_, new_n2197_, new_n312_ );
or   ( new_n2199_, new_n2198_, new_n2194_ );
and  ( new_n2200_, new_n2199_, new_n2193_ );
nor  ( new_n2201_, new_n2200_, new_n2184_ );
nand ( new_n2202_, new_n2201_, new_n2167_ );
and  ( new_n2203_, new_n2202_, new_n2166_ );
or   ( new_n2204_, new_n2203_, new_n2101_ );
nand ( new_n2205_, new_n2203_, new_n2101_ );
xor  ( new_n2206_, new_n1873_, new_n1857_ );
xnor ( new_n2207_, new_n2206_, new_n1891_ );
nand ( new_n2208_, new_n2207_, new_n2205_ );
and  ( new_n2209_, new_n2208_, new_n2204_ );
nor  ( new_n2210_, new_n2209_, new_n2091_ );
and  ( new_n2211_, new_n2209_, new_n2091_ );
xor  ( new_n2212_, new_n1977_, new_n1967_ );
xnor ( new_n2213_, new_n2212_, new_n2082_ );
nor  ( new_n2214_, new_n2213_, new_n2211_ );
nor  ( new_n2215_, new_n2214_, new_n2210_ );
or   ( new_n2216_, new_n2215_, new_n2089_ );
and  ( new_n2217_, new_n2216_, new_n2088_ );
xnor ( new_n2218_, new_n1822_, new_n1820_ );
xor  ( new_n2219_, new_n2218_, new_n1944_ );
nand ( new_n2220_, new_n2219_, new_n2217_ );
nor  ( new_n2221_, new_n2219_, new_n2217_ );
not  ( new_n2222_, new_n1962_ );
nand ( new_n2223_, new_n1964_, new_n2222_ );
nor  ( new_n2224_, new_n1964_, new_n2222_ );
or   ( new_n2225_, new_n2084_, new_n2224_ );
and  ( new_n2226_, new_n2225_, new_n2223_ );
or   ( new_n2227_, new_n2226_, new_n2221_ );
and  ( new_n2228_, new_n2227_, new_n2220_ );
nor  ( new_n2229_, new_n2228_, new_n1951_ );
xor  ( new_n2230_, new_n2203_, new_n2101_ );
xor  ( new_n2231_, new_n2230_, new_n2207_ );
not  ( new_n2232_, new_n2231_ );
xnor ( new_n2233_, new_n2068_, new_n2032_ );
xor  ( new_n2234_, new_n2233_, new_n2080_ );
and  ( new_n2235_, new_n2234_, new_n2232_ );
xnor ( new_n2236_, new_n1971_, new_n1969_ );
xor  ( new_n2237_, new_n2236_, new_n1975_ );
or   ( new_n2238_, new_n2122_, new_n319_ );
or   ( new_n2239_, new_n2124_, new_n333_ );
and  ( new_n2240_, new_n2239_, new_n2238_ );
xor  ( new_n2241_, new_n2240_, new_n1842_ );
xor  ( new_n2242_, RIbb2e800_31, RIbb2e878_30 );
xor  ( new_n2243_, RIbb2e878_30, new_n2118_ );
nor  ( new_n2244_, new_n2243_, new_n2242_ );
and  ( new_n2245_, new_n2244_, RIbb2d810_65 );
xor  ( new_n2246_, new_n2245_, new_n2121_ );
nand ( new_n2247_, new_n2246_, new_n2241_ );
nor  ( new_n2248_, new_n2246_, new_n2241_ );
or   ( new_n2249_, new_n1844_, new_n285_ );
or   ( new_n2250_, new_n1846_, new_n313_ );
and  ( new_n2251_, new_n2250_, new_n2249_ );
xor  ( new_n2252_, new_n2251_, new_n1586_ );
or   ( new_n2253_, new_n2252_, new_n2248_ );
and  ( new_n2254_, new_n2253_, new_n2247_ );
or   ( new_n2255_, new_n1593_, new_n301_ );
or   ( new_n2256_, new_n1595_, new_n279_ );
and  ( new_n2257_, new_n2256_, new_n2255_ );
xor  ( new_n2258_, new_n2257_, new_n1358_ );
or   ( new_n2259_, new_n1364_, new_n270_ );
or   ( new_n2260_, new_n1366_, new_n294_ );
and  ( new_n2261_, new_n2260_, new_n2259_ );
xor  ( new_n2262_, new_n2261_, new_n1129_ );
or   ( new_n2263_, new_n2262_, new_n2258_ );
and  ( new_n2264_, new_n2262_, new_n2258_ );
or   ( new_n2265_, new_n1135_, new_n348_ );
or   ( new_n2266_, new_n1137_, new_n264_ );
and  ( new_n2267_, new_n2266_, new_n2265_ );
xor  ( new_n2268_, new_n2267_, new_n896_ );
or   ( new_n2269_, new_n2268_, new_n2264_ );
and  ( new_n2270_, new_n2269_, new_n2263_ );
or   ( new_n2271_, new_n2270_, new_n2254_ );
and  ( new_n2272_, new_n2270_, new_n2254_ );
or   ( new_n2273_, new_n897_, new_n443_ );
or   ( new_n2274_, new_n899_, new_n419_ );
and  ( new_n2275_, new_n2274_, new_n2273_ );
xor  ( new_n2276_, new_n2275_, new_n748_ );
or   ( new_n2277_, new_n755_, new_n515_ );
or   ( new_n2278_, new_n757_, new_n509_ );
and  ( new_n2279_, new_n2278_, new_n2277_ );
xor  ( new_n2280_, new_n2279_, new_n523_ );
nor  ( new_n2281_, new_n2280_, new_n2276_ );
and  ( new_n2282_, new_n2280_, new_n2276_ );
or   ( new_n2283_, new_n524_, new_n805_ );
or   ( new_n2284_, new_n526_, new_n775_ );
and  ( new_n2285_, new_n2284_, new_n2283_ );
xor  ( new_n2286_, new_n2285_, new_n403_ );
nor  ( new_n2287_, new_n2286_, new_n2282_ );
nor  ( new_n2288_, new_n2287_, new_n2281_ );
or   ( new_n2289_, new_n2288_, new_n2272_ );
and  ( new_n2290_, new_n2289_, new_n2271_ );
not  ( new_n2291_, RIbb2caf0_93 );
or   ( new_n2292_, new_n2291_, new_n260_ );
xnor ( new_n2293_, new_n2175_, new_n2171_ );
xor  ( new_n2294_, new_n2293_, new_n2182_ );
nand ( new_n2295_, new_n2294_, new_n2292_ );
or   ( new_n2296_, new_n2294_, new_n2292_ );
xor  ( new_n2297_, new_n2192_, new_n2188_ );
xnor ( new_n2298_, new_n2297_, new_n2198_ );
nand ( new_n2299_, new_n2298_, new_n2296_ );
and  ( new_n2300_, new_n2299_, new_n2295_ );
nor  ( new_n2301_, new_n2300_, new_n2290_ );
nand ( new_n2302_, new_n2300_, new_n2290_ );
or   ( new_n2303_, new_n283_, new_n1754_ );
or   ( new_n2304_, new_n286_, new_n1523_ );
and  ( new_n2305_, new_n2304_, new_n2303_ );
xor  ( new_n2306_, new_n2305_, new_n278_ );
or   ( new_n2307_, new_n299_, new_n2057_ );
or   ( new_n2308_, new_n302_, new_n1899_ );
and  ( new_n2309_, new_n2308_, new_n2307_ );
xor  ( new_n2310_, new_n2309_, new_n293_ );
nor  ( new_n2311_, new_n2310_, new_n2306_ );
nand ( new_n2312_, new_n2310_, new_n2306_ );
or   ( new_n2313_, new_n268_, new_n2291_ );
or   ( new_n2314_, new_n271_, new_n2178_ );
and  ( new_n2315_, new_n2314_, new_n2313_ );
xor  ( new_n2316_, new_n2315_, new_n262_ );
and  ( new_n2317_, new_n2316_, new_n2312_ );
or   ( new_n2318_, new_n2317_, new_n2311_ );
and  ( new_n2319_, RIbb2ca78_94, RIbb2f610_1 );
not  ( new_n2320_, new_n2319_ );
or   ( new_n2321_, new_n409_, new_n986_ );
or   ( new_n2322_, new_n411_, new_n886_ );
and  ( new_n2323_, new_n2322_, new_n2321_ );
xor  ( new_n2324_, new_n2323_, new_n328_ );
or   ( new_n2325_, new_n337_, new_n1213_ );
or   ( new_n2326_, new_n340_, new_n1168_ );
and  ( new_n2327_, new_n2326_, new_n2325_ );
xor  ( new_n2328_, new_n2327_, new_n332_ );
nor  ( new_n2329_, new_n2328_, new_n2324_ );
and  ( new_n2330_, new_n2328_, new_n2324_ );
or   ( new_n2331_, new_n317_, new_n1525_ );
or   ( new_n2332_, new_n320_, new_n1318_ );
and  ( new_n2333_, new_n2332_, new_n2331_ );
xor  ( new_n2334_, new_n2333_, new_n312_ );
nor  ( new_n2335_, new_n2334_, new_n2330_ );
nor  ( new_n2336_, new_n2335_, new_n2329_ );
not  ( new_n2337_, new_n2336_ );
or   ( new_n2338_, new_n2337_, new_n2320_ );
and  ( new_n2339_, new_n2338_, new_n2318_ );
and  ( new_n2340_, new_n2337_, new_n2320_ );
or   ( new_n2341_, new_n2340_, new_n2339_ );
and  ( new_n2342_, new_n2341_, new_n2302_ );
or   ( new_n2343_, new_n2342_, new_n2301_ );
xnor ( new_n2344_, new_n2004_, new_n1999_ );
xor  ( new_n2345_, new_n2344_, new_n2010_ );
xor  ( new_n2346_, new_n2109_, new_n2105_ );
xor  ( new_n2347_, new_n2346_, new_n2115_ );
xor  ( new_n2348_, new_n2127_, new_n2121_ );
xor  ( new_n2349_, new_n2348_, new_n2133_ );
nand ( new_n2350_, new_n2349_, new_n2347_ );
nor  ( new_n2351_, new_n2349_, new_n2347_ );
xnor ( new_n2352_, new_n2145_, new_n2141_ );
xor  ( new_n2353_, new_n2352_, new_n2151_ );
or   ( new_n2354_, new_n2353_, new_n2351_ );
and  ( new_n2355_, new_n2354_, new_n2350_ );
or   ( new_n2356_, new_n2355_, new_n2345_ );
and  ( new_n2357_, new_n2355_, new_n2345_ );
xnor ( new_n2358_, new_n1987_, new_n1983_ );
xor  ( new_n2359_, new_n2358_, new_n1993_ );
or   ( new_n2360_, new_n2359_, new_n2357_ );
and  ( new_n2361_, new_n2360_, new_n2356_ );
nand ( new_n2362_, new_n2361_, new_n2343_ );
or   ( new_n2363_, new_n2361_, new_n2343_ );
xor  ( new_n2364_, new_n2135_, new_n2117_ );
xor  ( new_n2365_, new_n2364_, new_n2153_ );
xnor ( new_n2366_, new_n2159_, new_n2157_ );
xor  ( new_n2367_, new_n2366_, new_n2163_ );
and  ( new_n2368_, new_n2367_, new_n2365_ );
nor  ( new_n2369_, new_n2367_, new_n2365_ );
xor  ( new_n2370_, new_n2200_, new_n2184_ );
nor  ( new_n2371_, new_n2370_, new_n2369_ );
nor  ( new_n2372_, new_n2371_, new_n2368_ );
nand ( new_n2373_, new_n2372_, new_n2363_ );
and  ( new_n2374_, new_n2373_, new_n2362_ );
or   ( new_n2375_, new_n2374_, new_n2237_ );
and  ( new_n2376_, new_n2374_, new_n2237_ );
xnor ( new_n2377_, new_n2012_, new_n1995_ );
xor  ( new_n2378_, new_n2377_, new_n2030_ );
xor  ( new_n2379_, new_n2165_, new_n2155_ );
xor  ( new_n2380_, new_n2379_, new_n2201_ );
nor  ( new_n2381_, new_n2380_, new_n2378_ );
nand ( new_n2382_, new_n2380_, new_n2378_ );
xor  ( new_n2383_, new_n2095_, new_n2093_ );
xor  ( new_n2384_, new_n2383_, new_n2099_ );
and  ( new_n2385_, new_n2384_, new_n2382_ );
or   ( new_n2386_, new_n2385_, new_n2381_ );
or   ( new_n2387_, new_n2386_, new_n2376_ );
and  ( new_n2388_, new_n2387_, new_n2375_ );
nand ( new_n2389_, new_n2388_, new_n2235_ );
nor  ( new_n2390_, new_n2388_, new_n2235_ );
xor  ( new_n2391_, new_n2209_, new_n2091_ );
xnor ( new_n2392_, new_n2391_, new_n2213_ );
or   ( new_n2393_, new_n2392_, new_n2390_ );
and  ( new_n2394_, new_n2393_, new_n2389_ );
xnor ( new_n2395_, new_n2087_, new_n2085_ );
xor  ( new_n2396_, new_n2395_, new_n2215_ );
or   ( new_n2397_, new_n2396_, new_n2394_ );
xor  ( new_n2398_, new_n2219_, new_n2217_ );
xor  ( new_n2399_, new_n2398_, new_n2226_ );
nor  ( new_n2400_, new_n2399_, new_n2397_ );
xnor ( new_n2401_, new_n2388_, new_n2235_ );
xor  ( new_n2402_, new_n2401_, new_n2392_ );
xor  ( new_n2403_, new_n2374_, new_n2237_ );
xor  ( new_n2404_, new_n2403_, new_n2386_ );
or   ( new_n2405_, new_n1135_, new_n419_ );
or   ( new_n2406_, new_n1137_, new_n348_ );
and  ( new_n2407_, new_n2406_, new_n2405_ );
xor  ( new_n2408_, new_n2407_, new_n896_ );
or   ( new_n2409_, new_n897_, new_n509_ );
or   ( new_n2410_, new_n899_, new_n443_ );
and  ( new_n2411_, new_n2410_, new_n2409_ );
xor  ( new_n2412_, new_n2411_, new_n748_ );
nor  ( new_n2413_, new_n2412_, new_n2408_ );
and  ( new_n2414_, new_n2412_, new_n2408_ );
or   ( new_n2415_, new_n755_, new_n775_ );
or   ( new_n2416_, new_n757_, new_n515_ );
and  ( new_n2417_, new_n2416_, new_n2415_ );
xor  ( new_n2418_, new_n2417_, new_n523_ );
nor  ( new_n2419_, new_n2418_, new_n2414_ );
or   ( new_n2420_, new_n2419_, new_n2413_ );
not  ( new_n2421_, RIbb2e800_31 );
and  ( new_n2422_, RIbb2e710_33, RIbb2e788_32 );
nor  ( new_n2423_, new_n2422_, new_n2421_ );
not  ( new_n2424_, new_n2423_ );
not  ( new_n2425_, new_n2244_ );
or   ( new_n2426_, new_n2425_, new_n333_ );
not  ( new_n2427_, new_n2242_ );
or   ( new_n2428_, new_n2427_, new_n339_ );
and  ( new_n2429_, new_n2428_, new_n2426_ );
xor  ( new_n2430_, new_n2429_, new_n2121_ );
nand ( new_n2431_, new_n2430_, new_n2424_ );
or   ( new_n2432_, new_n2430_, new_n2424_ );
or   ( new_n2433_, new_n2122_, new_n313_ );
or   ( new_n2434_, new_n2124_, new_n319_ );
and  ( new_n2435_, new_n2434_, new_n2433_ );
xor  ( new_n2436_, new_n2435_, new_n1843_ );
nand ( new_n2437_, new_n2436_, new_n2432_ );
and  ( new_n2438_, new_n2437_, new_n2431_ );
nand ( new_n2439_, new_n2438_, new_n2420_ );
nor  ( new_n2440_, new_n2438_, new_n2420_ );
or   ( new_n2441_, new_n1844_, new_n279_ );
or   ( new_n2442_, new_n1846_, new_n285_ );
and  ( new_n2443_, new_n2442_, new_n2441_ );
xor  ( new_n2444_, new_n2443_, new_n1586_ );
or   ( new_n2445_, new_n1593_, new_n294_ );
or   ( new_n2446_, new_n1595_, new_n301_ );
and  ( new_n2447_, new_n2446_, new_n2445_ );
xor  ( new_n2448_, new_n2447_, new_n1358_ );
nor  ( new_n2449_, new_n2448_, new_n2444_ );
and  ( new_n2450_, new_n2448_, new_n2444_ );
or   ( new_n2451_, new_n1364_, new_n264_ );
or   ( new_n2452_, new_n1366_, new_n270_ );
and  ( new_n2453_, new_n2452_, new_n2451_ );
xor  ( new_n2454_, new_n2453_, new_n1129_ );
nor  ( new_n2455_, new_n2454_, new_n2450_ );
nor  ( new_n2456_, new_n2455_, new_n2449_ );
or   ( new_n2457_, new_n2456_, new_n2440_ );
and  ( new_n2458_, new_n2457_, new_n2439_ );
or   ( new_n2459_, new_n317_, new_n1523_ );
or   ( new_n2460_, new_n320_, new_n1525_ );
and  ( new_n2461_, new_n2460_, new_n2459_ );
xor  ( new_n2462_, new_n2461_, new_n312_ );
or   ( new_n2463_, new_n283_, new_n1899_ );
or   ( new_n2464_, new_n286_, new_n1754_ );
and  ( new_n2465_, new_n2464_, new_n2463_ );
xor  ( new_n2466_, new_n2465_, new_n278_ );
nor  ( new_n2467_, new_n2466_, new_n2462_ );
and  ( new_n2468_, new_n2466_, new_n2462_ );
or   ( new_n2469_, new_n299_, new_n2178_ );
or   ( new_n2470_, new_n302_, new_n2057_ );
and  ( new_n2471_, new_n2470_, new_n2469_ );
xor  ( new_n2472_, new_n2471_, new_n293_ );
nor  ( new_n2473_, new_n2472_, new_n2468_ );
nor  ( new_n2474_, new_n2473_, new_n2467_ );
not  ( new_n2475_, RIbb2ca78_94 );
or   ( new_n2476_, new_n268_, new_n2475_ );
or   ( new_n2477_, new_n271_, new_n2291_ );
and  ( new_n2478_, new_n2477_, new_n2476_ );
xor  ( new_n2479_, new_n2478_, new_n263_ );
and  ( new_n2480_, RIbb2ca00_95, RIbb2f610_1 );
and  ( new_n2481_, new_n2480_, new_n2479_ );
or   ( new_n2482_, new_n524_, new_n886_ );
or   ( new_n2483_, new_n526_, new_n805_ );
and  ( new_n2484_, new_n2483_, new_n2482_ );
xor  ( new_n2485_, new_n2484_, new_n403_ );
or   ( new_n2486_, new_n409_, new_n1168_ );
or   ( new_n2487_, new_n411_, new_n986_ );
and  ( new_n2488_, new_n2487_, new_n2486_ );
xor  ( new_n2489_, new_n2488_, new_n328_ );
or   ( new_n2490_, new_n2489_, new_n2485_ );
and  ( new_n2491_, new_n2489_, new_n2485_ );
or   ( new_n2492_, new_n337_, new_n1318_ );
or   ( new_n2493_, new_n340_, new_n1213_ );
and  ( new_n2494_, new_n2493_, new_n2492_ );
xor  ( new_n2495_, new_n2494_, new_n332_ );
or   ( new_n2496_, new_n2495_, new_n2491_ );
and  ( new_n2497_, new_n2496_, new_n2490_ );
and  ( new_n2498_, new_n2497_, new_n2481_ );
or   ( new_n2499_, new_n2498_, new_n2474_ );
or   ( new_n2500_, new_n2497_, new_n2481_ );
and  ( new_n2501_, new_n2500_, new_n2499_ );
nor  ( new_n2502_, new_n2501_, new_n2458_ );
nand ( new_n2503_, new_n2501_, new_n2458_ );
xor  ( new_n2504_, new_n2310_, new_n2306_ );
xor  ( new_n2505_, new_n2504_, new_n2316_ );
xnor ( new_n2506_, new_n2328_, new_n2324_ );
xor  ( new_n2507_, new_n2506_, new_n2334_ );
nor  ( new_n2508_, new_n2507_, new_n2505_ );
and  ( new_n2509_, new_n2507_, new_n2505_ );
nor  ( new_n2510_, new_n2509_, new_n2319_ );
nor  ( new_n2511_, new_n2510_, new_n2508_ );
and  ( new_n2512_, new_n2511_, new_n2503_ );
or   ( new_n2513_, new_n2512_, new_n2502_ );
xor  ( new_n2514_, new_n2349_, new_n2347_ );
xor  ( new_n2515_, new_n2514_, new_n2353_ );
xnor ( new_n2516_, new_n2262_, new_n2258_ );
xor  ( new_n2517_, new_n2516_, new_n2268_ );
xnor ( new_n2518_, new_n2246_, new_n2241_ );
xor  ( new_n2519_, new_n2518_, new_n2252_ );
or   ( new_n2520_, new_n2519_, new_n2517_ );
and  ( new_n2521_, new_n2519_, new_n2517_ );
xnor ( new_n2522_, new_n2280_, new_n2276_ );
xor  ( new_n2523_, new_n2522_, new_n2286_ );
or   ( new_n2524_, new_n2523_, new_n2521_ );
and  ( new_n2525_, new_n2524_, new_n2520_ );
or   ( new_n2526_, new_n2525_, new_n2515_ );
and  ( new_n2527_, new_n2525_, new_n2515_ );
xor  ( new_n2528_, new_n2294_, new_n2292_ );
xor  ( new_n2529_, new_n2528_, new_n2298_ );
or   ( new_n2530_, new_n2529_, new_n2527_ );
and  ( new_n2531_, new_n2530_, new_n2526_ );
and  ( new_n2532_, new_n2531_, new_n2513_ );
or   ( new_n2533_, new_n2531_, new_n2513_ );
xor  ( new_n2534_, new_n2270_, new_n2254_ );
xnor ( new_n2535_, new_n2534_, new_n2288_ );
not  ( new_n2536_, new_n2535_ );
xor  ( new_n2537_, new_n2336_, new_n2320_ );
xor  ( new_n2538_, new_n2537_, new_n2318_ );
and  ( new_n2539_, new_n2538_, new_n2536_ );
not  ( new_n2540_, new_n2539_ );
and  ( new_n2541_, new_n2540_, new_n2533_ );
or   ( new_n2542_, new_n2541_, new_n2532_ );
xor  ( new_n2543_, new_n2355_, new_n2345_ );
xor  ( new_n2544_, new_n2543_, new_n2359_ );
xor  ( new_n2545_, new_n2300_, new_n2290_ );
xor  ( new_n2546_, new_n2545_, new_n2341_ );
or   ( new_n2547_, new_n2546_, new_n2544_ );
and  ( new_n2548_, new_n2546_, new_n2544_ );
xor  ( new_n2549_, new_n2367_, new_n2365_ );
xor  ( new_n2550_, new_n2549_, new_n2370_ );
or   ( new_n2551_, new_n2550_, new_n2548_ );
and  ( new_n2552_, new_n2551_, new_n2547_ );
nand ( new_n2553_, new_n2552_, new_n2542_ );
or   ( new_n2554_, new_n2552_, new_n2542_ );
xor  ( new_n2555_, new_n2380_, new_n2378_ );
xnor ( new_n2556_, new_n2555_, new_n2384_ );
nand ( new_n2557_, new_n2556_, new_n2554_ );
and  ( new_n2558_, new_n2557_, new_n2553_ );
or   ( new_n2559_, new_n2558_, new_n2404_ );
and  ( new_n2560_, new_n2558_, new_n2404_ );
xor  ( new_n2561_, new_n2234_, new_n2232_ );
or   ( new_n2562_, new_n2561_, new_n2560_ );
and  ( new_n2563_, new_n2562_, new_n2559_ );
and  ( new_n2564_, new_n2563_, new_n2402_ );
xor  ( new_n2565_, new_n2396_, new_n2394_ );
and  ( new_n2566_, new_n2565_, new_n2564_ );
xor  ( new_n2567_, new_n2552_, new_n2542_ );
xor  ( new_n2568_, new_n2567_, new_n2556_ );
xor  ( new_n2569_, new_n2361_, new_n2343_ );
xor  ( new_n2570_, new_n2569_, new_n2372_ );
or   ( new_n2571_, new_n2570_, new_n2568_ );
and  ( new_n2572_, new_n2570_, new_n2568_ );
xnor ( new_n2573_, new_n2501_, new_n2458_ );
xor  ( new_n2574_, new_n2573_, new_n2511_ );
xnor ( new_n2575_, new_n2525_, new_n2515_ );
xor  ( new_n2576_, new_n2575_, new_n2529_ );
nor  ( new_n2577_, new_n2576_, new_n2574_ );
nand ( new_n2578_, new_n2576_, new_n2574_ );
xor  ( new_n2579_, new_n2538_, new_n2536_ );
not  ( new_n2580_, new_n2579_ );
and  ( new_n2581_, new_n2580_, new_n2578_ );
or   ( new_n2582_, new_n2581_, new_n2577_ );
xor  ( new_n2583_, new_n2546_, new_n2544_ );
xor  ( new_n2584_, new_n2583_, new_n2550_ );
nor  ( new_n2585_, new_n2584_, new_n2582_ );
and  ( new_n2586_, new_n2584_, new_n2582_ );
xor  ( new_n2587_, new_n2438_, new_n2420_ );
xnor ( new_n2588_, new_n2587_, new_n2456_ );
not  ( new_n2589_, new_n2588_ );
xor  ( new_n2590_, new_n2497_, new_n2481_ );
xor  ( new_n2591_, new_n2590_, new_n2474_ );
nand ( new_n2592_, new_n2591_, new_n2589_ );
or   ( new_n2593_, new_n1135_, new_n443_ );
or   ( new_n2594_, new_n1137_, new_n419_ );
and  ( new_n2595_, new_n2594_, new_n2593_ );
xor  ( new_n2596_, new_n2595_, new_n896_ );
or   ( new_n2597_, new_n897_, new_n515_ );
or   ( new_n2598_, new_n899_, new_n509_ );
and  ( new_n2599_, new_n2598_, new_n2597_ );
xor  ( new_n2600_, new_n2599_, new_n748_ );
or   ( new_n2601_, new_n2600_, new_n2596_ );
and  ( new_n2602_, new_n2600_, new_n2596_ );
or   ( new_n2603_, new_n755_, new_n805_ );
or   ( new_n2604_, new_n757_, new_n775_ );
and  ( new_n2605_, new_n2604_, new_n2603_ );
xor  ( new_n2606_, new_n2605_, new_n523_ );
or   ( new_n2607_, new_n2606_, new_n2602_ );
and  ( new_n2608_, new_n2607_, new_n2601_ );
or   ( new_n2609_, new_n2425_, new_n319_ );
or   ( new_n2610_, new_n2427_, new_n333_ );
and  ( new_n2611_, new_n2610_, new_n2609_ );
xor  ( new_n2612_, new_n2611_, new_n2120_ );
xor  ( new_n2613_, RIbb2e710_33, RIbb2e788_32 );
xor  ( new_n2614_, RIbb2e788_32, new_n2421_ );
nor  ( new_n2615_, new_n2614_, new_n2613_ );
and  ( new_n2616_, new_n2615_, RIbb2d810_65 );
xor  ( new_n2617_, new_n2616_, new_n2424_ );
nand ( new_n2618_, new_n2617_, new_n2612_ );
nor  ( new_n2619_, new_n2617_, new_n2612_ );
or   ( new_n2620_, new_n2122_, new_n285_ );
or   ( new_n2621_, new_n2124_, new_n313_ );
and  ( new_n2622_, new_n2621_, new_n2620_ );
xor  ( new_n2623_, new_n2622_, new_n1843_ );
or   ( new_n2624_, new_n2623_, new_n2619_ );
and  ( new_n2625_, new_n2624_, new_n2618_ );
or   ( new_n2626_, new_n2625_, new_n2608_ );
and  ( new_n2627_, new_n2625_, new_n2608_ );
or   ( new_n2628_, new_n1844_, new_n301_ );
or   ( new_n2629_, new_n1846_, new_n279_ );
and  ( new_n2630_, new_n2629_, new_n2628_ );
xor  ( new_n2631_, new_n2630_, new_n1586_ );
or   ( new_n2632_, new_n1593_, new_n270_ );
or   ( new_n2633_, new_n1595_, new_n294_ );
and  ( new_n2634_, new_n2633_, new_n2632_ );
xor  ( new_n2635_, new_n2634_, new_n1358_ );
nor  ( new_n2636_, new_n2635_, new_n2631_ );
and  ( new_n2637_, new_n2635_, new_n2631_ );
or   ( new_n2638_, new_n1364_, new_n348_ );
or   ( new_n2639_, new_n1366_, new_n264_ );
and  ( new_n2640_, new_n2639_, new_n2638_ );
xor  ( new_n2641_, new_n2640_, new_n1129_ );
nor  ( new_n2642_, new_n2641_, new_n2637_ );
nor  ( new_n2643_, new_n2642_, new_n2636_ );
or   ( new_n2644_, new_n2643_, new_n2627_ );
and  ( new_n2645_, new_n2644_, new_n2626_ );
not  ( new_n2646_, RIbb2ca00_95 );
or   ( new_n2647_, new_n268_, new_n2646_ );
or   ( new_n2648_, new_n271_, new_n2475_ );
and  ( new_n2649_, new_n2648_, new_n2647_ );
xor  ( new_n2650_, new_n2649_, new_n263_ );
and  ( new_n2651_, RIbb2c988_96, RIbb2f610_1 );
or   ( new_n2652_, new_n2651_, new_n2650_ );
or   ( new_n2653_, new_n317_, new_n1754_ );
or   ( new_n2654_, new_n320_, new_n1523_ );
and  ( new_n2655_, new_n2654_, new_n2653_ );
xor  ( new_n2656_, new_n2655_, new_n312_ );
or   ( new_n2657_, new_n283_, new_n2057_ );
or   ( new_n2658_, new_n286_, new_n1899_ );
and  ( new_n2659_, new_n2658_, new_n2657_ );
xor  ( new_n2660_, new_n2659_, new_n278_ );
or   ( new_n2661_, new_n2660_, new_n2656_ );
and  ( new_n2662_, new_n2660_, new_n2656_ );
or   ( new_n2663_, new_n299_, new_n2291_ );
or   ( new_n2664_, new_n302_, new_n2178_ );
and  ( new_n2665_, new_n2664_, new_n2663_ );
xor  ( new_n2666_, new_n2665_, new_n293_ );
or   ( new_n2667_, new_n2666_, new_n2662_ );
and  ( new_n2668_, new_n2667_, new_n2661_ );
or   ( new_n2669_, new_n2668_, new_n2652_ );
and  ( new_n2670_, new_n2668_, new_n2652_ );
or   ( new_n2671_, new_n524_, new_n986_ );
or   ( new_n2672_, new_n526_, new_n886_ );
and  ( new_n2673_, new_n2672_, new_n2671_ );
xor  ( new_n2674_, new_n2673_, new_n403_ );
or   ( new_n2675_, new_n409_, new_n1213_ );
or   ( new_n2676_, new_n411_, new_n1168_ );
and  ( new_n2677_, new_n2676_, new_n2675_ );
xor  ( new_n2678_, new_n2677_, new_n328_ );
nor  ( new_n2679_, new_n2678_, new_n2674_ );
and  ( new_n2680_, new_n2678_, new_n2674_ );
or   ( new_n2681_, new_n337_, new_n1525_ );
or   ( new_n2682_, new_n340_, new_n1318_ );
and  ( new_n2683_, new_n2682_, new_n2681_ );
xor  ( new_n2684_, new_n2683_, new_n332_ );
nor  ( new_n2685_, new_n2684_, new_n2680_ );
nor  ( new_n2686_, new_n2685_, new_n2679_ );
or   ( new_n2687_, new_n2686_, new_n2670_ );
and  ( new_n2688_, new_n2687_, new_n2669_ );
nand ( new_n2689_, new_n2688_, new_n2645_ );
nor  ( new_n2690_, new_n2688_, new_n2645_ );
xnor ( new_n2691_, new_n2466_, new_n2462_ );
xor  ( new_n2692_, new_n2691_, new_n2472_ );
xnor ( new_n2693_, new_n2489_, new_n2485_ );
xor  ( new_n2694_, new_n2693_, new_n2495_ );
nor  ( new_n2695_, new_n2694_, new_n2692_ );
and  ( new_n2696_, new_n2694_, new_n2692_ );
xor  ( new_n2697_, new_n2480_, new_n2479_ );
not  ( new_n2698_, new_n2697_ );
nor  ( new_n2699_, new_n2698_, new_n2696_ );
nor  ( new_n2700_, new_n2699_, new_n2695_ );
or   ( new_n2701_, new_n2700_, new_n2690_ );
and  ( new_n2702_, new_n2701_, new_n2689_ );
nor  ( new_n2703_, new_n2702_, new_n2592_ );
and  ( new_n2704_, new_n2702_, new_n2592_ );
xor  ( new_n2705_, new_n2519_, new_n2517_ );
xor  ( new_n2706_, new_n2705_, new_n2523_ );
xor  ( new_n2707_, new_n2412_, new_n2408_ );
xor  ( new_n2708_, new_n2707_, new_n2418_ );
xor  ( new_n2709_, new_n2430_, new_n2424_ );
xor  ( new_n2710_, new_n2709_, new_n2436_ );
nand ( new_n2711_, new_n2710_, new_n2708_ );
nor  ( new_n2712_, new_n2710_, new_n2708_ );
xnor ( new_n2713_, new_n2448_, new_n2444_ );
xor  ( new_n2714_, new_n2713_, new_n2454_ );
or   ( new_n2715_, new_n2714_, new_n2712_ );
and  ( new_n2716_, new_n2715_, new_n2711_ );
nor  ( new_n2717_, new_n2716_, new_n2706_ );
and  ( new_n2718_, new_n2716_, new_n2706_ );
xor  ( new_n2719_, new_n2507_, new_n2505_ );
xnor ( new_n2720_, new_n2719_, new_n2320_ );
nor  ( new_n2721_, new_n2720_, new_n2718_ );
nor  ( new_n2722_, new_n2721_, new_n2717_ );
nor  ( new_n2723_, new_n2722_, new_n2704_ );
nor  ( new_n2724_, new_n2723_, new_n2703_ );
nor  ( new_n2725_, new_n2724_, new_n2586_ );
nor  ( new_n2726_, new_n2725_, new_n2585_ );
or   ( new_n2727_, new_n2726_, new_n2572_ );
and  ( new_n2728_, new_n2727_, new_n2571_ );
xnor ( new_n2729_, new_n2558_, new_n2404_ );
xor  ( new_n2730_, new_n2729_, new_n2561_ );
nor  ( new_n2731_, new_n2730_, new_n2728_ );
xor  ( new_n2732_, new_n2563_, new_n2402_ );
and  ( new_n2733_, new_n2732_, new_n2731_ );
xnor ( new_n2734_, new_n2570_, new_n2568_ );
xor  ( new_n2735_, new_n2734_, new_n2726_ );
xnor ( new_n2736_, new_n2584_, new_n2582_ );
xor  ( new_n2737_, new_n2736_, new_n2724_ );
xnor ( new_n2738_, new_n2716_, new_n2706_ );
xor  ( new_n2739_, new_n2738_, new_n2720_ );
xnor ( new_n2740_, new_n2688_, new_n2645_ );
xor  ( new_n2741_, new_n2740_, new_n2700_ );
or   ( new_n2742_, new_n2741_, new_n2739_ );
and  ( new_n2743_, new_n2741_, new_n2739_ );
xor  ( new_n2744_, new_n2591_, new_n2589_ );
or   ( new_n2745_, new_n2744_, new_n2743_ );
and  ( new_n2746_, new_n2745_, new_n2742_ );
or   ( new_n2747_, new_n299_, new_n2475_ );
or   ( new_n2748_, new_n302_, new_n2291_ );
and  ( new_n2749_, new_n2748_, new_n2747_ );
xor  ( new_n2750_, new_n2749_, new_n293_ );
not  ( new_n2751_, RIbb2c988_96 );
or   ( new_n2752_, new_n268_, new_n2751_ );
or   ( new_n2753_, new_n271_, new_n2646_ );
and  ( new_n2754_, new_n2753_, new_n2752_ );
xor  ( new_n2755_, new_n2754_, new_n263_ );
or   ( new_n2756_, new_n2755_, new_n2750_ );
and  ( new_n2757_, RIbb2c910_97, RIbb2f610_1 );
and  ( new_n2758_, new_n2755_, new_n2750_ );
or   ( new_n2759_, new_n2758_, new_n2757_ );
and  ( new_n2760_, new_n2759_, new_n2756_ );
or   ( new_n2761_, new_n337_, new_n1523_ );
or   ( new_n2762_, new_n340_, new_n1525_ );
and  ( new_n2763_, new_n2762_, new_n2761_ );
xor  ( new_n2764_, new_n2763_, new_n332_ );
or   ( new_n2765_, new_n317_, new_n1899_ );
or   ( new_n2766_, new_n320_, new_n1754_ );
and  ( new_n2767_, new_n2766_, new_n2765_ );
xor  ( new_n2768_, new_n2767_, new_n312_ );
or   ( new_n2769_, new_n2768_, new_n2764_ );
and  ( new_n2770_, new_n2768_, new_n2764_ );
or   ( new_n2771_, new_n283_, new_n2178_ );
or   ( new_n2772_, new_n286_, new_n2057_ );
and  ( new_n2773_, new_n2772_, new_n2771_ );
xor  ( new_n2774_, new_n2773_, new_n278_ );
or   ( new_n2775_, new_n2774_, new_n2770_ );
and  ( new_n2776_, new_n2775_, new_n2769_ );
or   ( new_n2777_, new_n2776_, new_n2760_ );
and  ( new_n2778_, new_n2776_, new_n2760_ );
or   ( new_n2779_, new_n755_, new_n886_ );
or   ( new_n2780_, new_n757_, new_n805_ );
and  ( new_n2781_, new_n2780_, new_n2779_ );
xor  ( new_n2782_, new_n2781_, new_n523_ );
or   ( new_n2783_, new_n524_, new_n1168_ );
or   ( new_n2784_, new_n526_, new_n986_ );
and  ( new_n2785_, new_n2784_, new_n2783_ );
xor  ( new_n2786_, new_n2785_, new_n403_ );
nor  ( new_n2787_, new_n2786_, new_n2782_ );
and  ( new_n2788_, new_n2786_, new_n2782_ );
or   ( new_n2789_, new_n409_, new_n1318_ );
or   ( new_n2790_, new_n411_, new_n1213_ );
and  ( new_n2791_, new_n2790_, new_n2789_ );
xor  ( new_n2792_, new_n2791_, new_n328_ );
nor  ( new_n2793_, new_n2792_, new_n2788_ );
nor  ( new_n2794_, new_n2793_, new_n2787_ );
or   ( new_n2795_, new_n2794_, new_n2778_ );
and  ( new_n2796_, new_n2795_, new_n2777_ );
not  ( new_n2797_, RIbb2e710_33 );
and  ( new_n2798_, RIbb2e620_35, RIbb2e698_34 );
nor  ( new_n2799_, new_n2798_, new_n2797_ );
not  ( new_n2800_, new_n2799_ );
or   ( new_n2801_, new_n2425_, new_n313_ );
or   ( new_n2802_, new_n2427_, new_n319_ );
and  ( new_n2803_, new_n2802_, new_n2801_ );
xor  ( new_n2804_, new_n2803_, new_n2121_ );
and  ( new_n2805_, new_n2804_, new_n2800_ );
or   ( new_n2806_, new_n2804_, new_n2800_ );
not  ( new_n2807_, new_n2615_ );
or   ( new_n2808_, new_n2807_, new_n333_ );
not  ( new_n2809_, new_n2613_ );
or   ( new_n2810_, new_n2809_, new_n339_ );
and  ( new_n2811_, new_n2810_, new_n2808_ );
xor  ( new_n2812_, new_n2811_, new_n2424_ );
and  ( new_n2813_, new_n2812_, new_n2806_ );
or   ( new_n2814_, new_n2813_, new_n2805_ );
or   ( new_n2815_, new_n2122_, new_n279_ );
or   ( new_n2816_, new_n2124_, new_n285_ );
and  ( new_n2817_, new_n2816_, new_n2815_ );
xor  ( new_n2818_, new_n2817_, new_n1843_ );
or   ( new_n2819_, new_n1844_, new_n294_ );
or   ( new_n2820_, new_n1846_, new_n301_ );
and  ( new_n2821_, new_n2820_, new_n2819_ );
xor  ( new_n2822_, new_n2821_, new_n1586_ );
or   ( new_n2823_, new_n2822_, new_n2818_ );
and  ( new_n2824_, new_n2822_, new_n2818_ );
or   ( new_n2825_, new_n1593_, new_n264_ );
or   ( new_n2826_, new_n1595_, new_n270_ );
and  ( new_n2827_, new_n2826_, new_n2825_ );
xor  ( new_n2828_, new_n2827_, new_n1358_ );
or   ( new_n2829_, new_n2828_, new_n2824_ );
and  ( new_n2830_, new_n2829_, new_n2823_ );
or   ( new_n2831_, new_n2830_, new_n2814_ );
and  ( new_n2832_, new_n2830_, new_n2814_ );
or   ( new_n2833_, new_n1364_, new_n419_ );
or   ( new_n2834_, new_n1366_, new_n348_ );
and  ( new_n2835_, new_n2834_, new_n2833_ );
xor  ( new_n2836_, new_n2835_, new_n1129_ );
or   ( new_n2837_, new_n1135_, new_n509_ );
or   ( new_n2838_, new_n1137_, new_n443_ );
and  ( new_n2839_, new_n2838_, new_n2837_ );
xor  ( new_n2840_, new_n2839_, new_n896_ );
nor  ( new_n2841_, new_n2840_, new_n2836_ );
and  ( new_n2842_, new_n2840_, new_n2836_ );
or   ( new_n2843_, new_n897_, new_n775_ );
or   ( new_n2844_, new_n899_, new_n515_ );
and  ( new_n2845_, new_n2844_, new_n2843_ );
xor  ( new_n2846_, new_n2845_, new_n748_ );
nor  ( new_n2847_, new_n2846_, new_n2842_ );
nor  ( new_n2848_, new_n2847_, new_n2841_ );
or   ( new_n2849_, new_n2848_, new_n2832_ );
and  ( new_n2850_, new_n2849_, new_n2831_ );
nor  ( new_n2851_, new_n2850_, new_n2796_ );
nand ( new_n2852_, new_n2850_, new_n2796_ );
xnor ( new_n2853_, new_n2660_, new_n2656_ );
xor  ( new_n2854_, new_n2853_, new_n2666_ );
xnor ( new_n2855_, new_n2678_, new_n2674_ );
xor  ( new_n2856_, new_n2855_, new_n2684_ );
or   ( new_n2857_, new_n2856_, new_n2854_ );
and  ( new_n2858_, new_n2856_, new_n2854_ );
xor  ( new_n2859_, new_n2651_, new_n2650_ );
or   ( new_n2860_, new_n2859_, new_n2858_ );
and  ( new_n2861_, new_n2860_, new_n2857_ );
and  ( new_n2862_, new_n2861_, new_n2852_ );
or   ( new_n2863_, new_n2862_, new_n2851_ );
xor  ( new_n2864_, new_n2710_, new_n2708_ );
xor  ( new_n2865_, new_n2864_, new_n2714_ );
xnor ( new_n2866_, new_n2617_, new_n2612_ );
xor  ( new_n2867_, new_n2866_, new_n2623_ );
xnor ( new_n2868_, new_n2600_, new_n2596_ );
xor  ( new_n2869_, new_n2868_, new_n2606_ );
or   ( new_n2870_, new_n2869_, new_n2867_ );
and  ( new_n2871_, new_n2869_, new_n2867_ );
xnor ( new_n2872_, new_n2635_, new_n2631_ );
xor  ( new_n2873_, new_n2872_, new_n2641_ );
or   ( new_n2874_, new_n2873_, new_n2871_ );
and  ( new_n2875_, new_n2874_, new_n2870_ );
or   ( new_n2876_, new_n2875_, new_n2865_ );
and  ( new_n2877_, new_n2875_, new_n2865_ );
xor  ( new_n2878_, new_n2694_, new_n2692_ );
xor  ( new_n2879_, new_n2878_, new_n2698_ );
or   ( new_n2880_, new_n2879_, new_n2877_ );
and  ( new_n2881_, new_n2880_, new_n2876_ );
nand ( new_n2882_, new_n2881_, new_n2863_ );
nor  ( new_n2883_, new_n2881_, new_n2863_ );
xor  ( new_n2884_, new_n2625_, new_n2608_ );
xnor ( new_n2885_, new_n2884_, new_n2643_ );
xnor ( new_n2886_, new_n2668_, new_n2652_ );
xor  ( new_n2887_, new_n2886_, new_n2686_ );
nor  ( new_n2888_, new_n2887_, new_n2885_ );
or   ( new_n2889_, new_n2888_, new_n2883_ );
and  ( new_n2890_, new_n2889_, new_n2882_ );
or   ( new_n2891_, new_n2890_, new_n2746_ );
nand ( new_n2892_, new_n2890_, new_n2746_ );
xor  ( new_n2893_, new_n2576_, new_n2574_ );
xor  ( new_n2894_, new_n2893_, new_n2580_ );
nand ( new_n2895_, new_n2894_, new_n2892_ );
and  ( new_n2896_, new_n2895_, new_n2891_ );
or   ( new_n2897_, new_n2896_, new_n2737_ );
nand ( new_n2898_, new_n2896_, new_n2737_ );
xor  ( new_n2899_, new_n2531_, new_n2513_ );
xor  ( new_n2900_, new_n2899_, new_n2540_ );
nand ( new_n2901_, new_n2900_, new_n2898_ );
and  ( new_n2902_, new_n2901_, new_n2897_ );
and  ( new_n2903_, new_n2902_, new_n2735_ );
xor  ( new_n2904_, new_n2730_, new_n2728_ );
and  ( new_n2905_, new_n2904_, new_n2903_ );
xnor ( new_n2906_, new_n2741_, new_n2739_ );
xor  ( new_n2907_, new_n2906_, new_n2744_ );
xor  ( new_n2908_, new_n2850_, new_n2796_ );
xor  ( new_n2909_, new_n2908_, new_n2861_ );
xor  ( new_n2910_, new_n2875_, new_n2865_ );
xor  ( new_n2911_, new_n2910_, new_n2879_ );
or   ( new_n2912_, new_n2911_, new_n2909_ );
nand ( new_n2913_, new_n2911_, new_n2909_ );
xor  ( new_n2914_, new_n2887_, new_n2885_ );
nand ( new_n2915_, new_n2914_, new_n2913_ );
and  ( new_n2916_, new_n2915_, new_n2912_ );
nor  ( new_n2917_, new_n2916_, new_n2907_ );
nand ( new_n2918_, new_n2916_, new_n2907_ );
xnor ( new_n2919_, new_n2776_, new_n2760_ );
xor  ( new_n2920_, new_n2919_, new_n2794_ );
xnor ( new_n2921_, new_n2830_, new_n2814_ );
xor  ( new_n2922_, new_n2921_, new_n2848_ );
or   ( new_n2923_, new_n2922_, new_n2920_ );
or   ( new_n2924_, new_n2807_, new_n319_ );
or   ( new_n2925_, new_n2809_, new_n333_ );
and  ( new_n2926_, new_n2925_, new_n2924_ );
xor  ( new_n2927_, new_n2926_, new_n2423_ );
xor  ( new_n2928_, RIbb2e620_35, RIbb2e698_34 );
xor  ( new_n2929_, RIbb2e698_34, new_n2797_ );
nor  ( new_n2930_, new_n2929_, new_n2928_ );
and  ( new_n2931_, new_n2930_, RIbb2d810_65 );
xor  ( new_n2932_, new_n2931_, new_n2800_ );
nand ( new_n2933_, new_n2932_, new_n2927_ );
nor  ( new_n2934_, new_n2932_, new_n2927_ );
or   ( new_n2935_, new_n2425_, new_n285_ );
or   ( new_n2936_, new_n2427_, new_n313_ );
and  ( new_n2937_, new_n2936_, new_n2935_ );
xor  ( new_n2938_, new_n2937_, new_n2121_ );
or   ( new_n2939_, new_n2938_, new_n2934_ );
and  ( new_n2940_, new_n2939_, new_n2933_ );
or   ( new_n2941_, new_n2122_, new_n301_ );
or   ( new_n2942_, new_n2124_, new_n279_ );
and  ( new_n2943_, new_n2942_, new_n2941_ );
xor  ( new_n2944_, new_n2943_, new_n1843_ );
or   ( new_n2945_, new_n1844_, new_n270_ );
or   ( new_n2946_, new_n1846_, new_n294_ );
and  ( new_n2947_, new_n2946_, new_n2945_ );
xor  ( new_n2948_, new_n2947_, new_n1586_ );
or   ( new_n2949_, new_n2948_, new_n2944_ );
and  ( new_n2950_, new_n2948_, new_n2944_ );
or   ( new_n2951_, new_n1593_, new_n348_ );
or   ( new_n2952_, new_n1595_, new_n264_ );
and  ( new_n2953_, new_n2952_, new_n2951_ );
xor  ( new_n2954_, new_n2953_, new_n1358_ );
or   ( new_n2955_, new_n2954_, new_n2950_ );
and  ( new_n2956_, new_n2955_, new_n2949_ );
nor  ( new_n2957_, new_n2956_, new_n2940_ );
nand ( new_n2958_, new_n2956_, new_n2940_ );
or   ( new_n2959_, new_n1364_, new_n443_ );
or   ( new_n2960_, new_n1366_, new_n419_ );
and  ( new_n2961_, new_n2960_, new_n2959_ );
xor  ( new_n2962_, new_n2961_, new_n1129_ );
or   ( new_n2963_, new_n1135_, new_n515_ );
or   ( new_n2964_, new_n1137_, new_n509_ );
and  ( new_n2965_, new_n2964_, new_n2963_ );
xor  ( new_n2966_, new_n2965_, new_n896_ );
nor  ( new_n2967_, new_n2966_, new_n2962_ );
nand ( new_n2968_, new_n2966_, new_n2962_ );
or   ( new_n2969_, new_n897_, new_n805_ );
or   ( new_n2970_, new_n899_, new_n775_ );
and  ( new_n2971_, new_n2970_, new_n2969_ );
xor  ( new_n2972_, new_n2971_, new_n747_ );
and  ( new_n2973_, new_n2972_, new_n2968_ );
or   ( new_n2974_, new_n2973_, new_n2967_ );
and  ( new_n2975_, new_n2974_, new_n2958_ );
or   ( new_n2976_, new_n2975_, new_n2957_ );
or   ( new_n2977_, new_n299_, new_n2646_ );
or   ( new_n2978_, new_n302_, new_n2475_ );
and  ( new_n2979_, new_n2978_, new_n2977_ );
xor  ( new_n2980_, new_n2979_, new_n293_ );
not  ( new_n2981_, RIbb2c910_97 );
or   ( new_n2982_, new_n268_, new_n2981_ );
or   ( new_n2983_, new_n271_, new_n2751_ );
and  ( new_n2984_, new_n2983_, new_n2982_ );
xor  ( new_n2985_, new_n2984_, new_n263_ );
or   ( new_n2986_, new_n2985_, new_n2980_ );
and  ( new_n2987_, RIbb2c898_98, RIbb2f610_1 );
and  ( new_n2988_, new_n2985_, new_n2980_ );
or   ( new_n2989_, new_n2988_, new_n2987_ );
and  ( new_n2990_, new_n2989_, new_n2986_ );
or   ( new_n2991_, new_n337_, new_n1754_ );
or   ( new_n2992_, new_n340_, new_n1523_ );
and  ( new_n2993_, new_n2992_, new_n2991_ );
xor  ( new_n2994_, new_n2993_, new_n332_ );
or   ( new_n2995_, new_n317_, new_n2057_ );
or   ( new_n2996_, new_n320_, new_n1899_ );
and  ( new_n2997_, new_n2996_, new_n2995_ );
xor  ( new_n2998_, new_n2997_, new_n312_ );
or   ( new_n2999_, new_n2998_, new_n2994_ );
and  ( new_n3000_, new_n2998_, new_n2994_ );
or   ( new_n3001_, new_n283_, new_n2291_ );
or   ( new_n3002_, new_n286_, new_n2178_ );
and  ( new_n3003_, new_n3002_, new_n3001_ );
xor  ( new_n3004_, new_n3003_, new_n278_ );
or   ( new_n3005_, new_n3004_, new_n3000_ );
and  ( new_n3006_, new_n3005_, new_n2999_ );
nor  ( new_n3007_, new_n3006_, new_n2990_ );
and  ( new_n3008_, new_n3006_, new_n2990_ );
or   ( new_n3009_, new_n755_, new_n986_ );
or   ( new_n3010_, new_n757_, new_n886_ );
and  ( new_n3011_, new_n3010_, new_n3009_ );
xor  ( new_n3012_, new_n3011_, new_n523_ );
or   ( new_n3013_, new_n524_, new_n1213_ );
or   ( new_n3014_, new_n526_, new_n1168_ );
and  ( new_n3015_, new_n3014_, new_n3013_ );
xor  ( new_n3016_, new_n3015_, new_n403_ );
nor  ( new_n3017_, new_n3016_, new_n3012_ );
and  ( new_n3018_, new_n3016_, new_n3012_ );
or   ( new_n3019_, new_n409_, new_n1525_ );
or   ( new_n3020_, new_n411_, new_n1318_ );
and  ( new_n3021_, new_n3020_, new_n3019_ );
xor  ( new_n3022_, new_n3021_, new_n328_ );
nor  ( new_n3023_, new_n3022_, new_n3018_ );
nor  ( new_n3024_, new_n3023_, new_n3017_ );
nor  ( new_n3025_, new_n3024_, new_n3008_ );
nor  ( new_n3026_, new_n3025_, new_n3007_ );
not  ( new_n3027_, new_n3026_ );
or   ( new_n3028_, new_n3027_, new_n2976_ );
and  ( new_n3029_, new_n3027_, new_n2976_ );
xnor ( new_n3030_, new_n2755_, new_n2750_ );
xor  ( new_n3031_, new_n3030_, new_n2757_ );
xnor ( new_n3032_, new_n2768_, new_n2764_ );
xor  ( new_n3033_, new_n3032_, new_n2774_ );
or   ( new_n3034_, new_n3033_, new_n3031_ );
and  ( new_n3035_, new_n3033_, new_n3031_ );
xnor ( new_n3036_, new_n2786_, new_n2782_ );
xor  ( new_n3037_, new_n3036_, new_n2792_ );
or   ( new_n3038_, new_n3037_, new_n3035_ );
and  ( new_n3039_, new_n3038_, new_n3034_ );
or   ( new_n3040_, new_n3039_, new_n3029_ );
and  ( new_n3041_, new_n3040_, new_n3028_ );
nor  ( new_n3042_, new_n3041_, new_n2923_ );
nand ( new_n3043_, new_n3041_, new_n2923_ );
xor  ( new_n3044_, new_n2869_, new_n2867_ );
xor  ( new_n3045_, new_n3044_, new_n2873_ );
xnor ( new_n3046_, new_n2822_, new_n2818_ );
xor  ( new_n3047_, new_n3046_, new_n2828_ );
xnor ( new_n3048_, new_n2840_, new_n2836_ );
xor  ( new_n3049_, new_n3048_, new_n2846_ );
or   ( new_n3050_, new_n3049_, new_n3047_ );
and  ( new_n3051_, new_n3049_, new_n3047_ );
xor  ( new_n3052_, new_n2804_, new_n2799_ );
xor  ( new_n3053_, new_n3052_, new_n2812_ );
or   ( new_n3054_, new_n3053_, new_n3051_ );
and  ( new_n3055_, new_n3054_, new_n3050_ );
nor  ( new_n3056_, new_n3055_, new_n3045_ );
nand ( new_n3057_, new_n3055_, new_n3045_ );
xnor ( new_n3058_, new_n2856_, new_n2854_ );
xor  ( new_n3059_, new_n3058_, new_n2859_ );
and  ( new_n3060_, new_n3059_, new_n3057_ );
or   ( new_n3061_, new_n3060_, new_n3056_ );
and  ( new_n3062_, new_n3061_, new_n3043_ );
or   ( new_n3063_, new_n3062_, new_n3042_ );
and  ( new_n3064_, new_n3063_, new_n2918_ );
or   ( new_n3065_, new_n3064_, new_n2917_ );
xnor ( new_n3066_, new_n2702_, new_n2592_ );
xor  ( new_n3067_, new_n3066_, new_n2722_ );
nand ( new_n3068_, new_n3067_, new_n3065_ );
nor  ( new_n3069_, new_n3067_, new_n3065_ );
xor  ( new_n3070_, new_n2890_, new_n2746_ );
xor  ( new_n3071_, new_n3070_, new_n2894_ );
or   ( new_n3072_, new_n3071_, new_n3069_ );
and  ( new_n3073_, new_n3072_, new_n3068_ );
xor  ( new_n3074_, new_n2896_, new_n2737_ );
xor  ( new_n3075_, new_n3074_, new_n2900_ );
nor  ( new_n3076_, new_n3075_, new_n3073_ );
xor  ( new_n3077_, new_n2902_, new_n2735_ );
and  ( new_n3078_, new_n3077_, new_n3076_ );
xnor ( new_n3079_, new_n3067_, new_n3065_ );
xor  ( new_n3080_, new_n3079_, new_n3071_ );
xor  ( new_n3081_, new_n2916_, new_n2907_ );
xor  ( new_n3082_, new_n3081_, new_n3063_ );
xor  ( new_n3083_, new_n3026_, new_n2976_ );
xor  ( new_n3084_, new_n3083_, new_n3039_ );
xor  ( new_n3085_, new_n3055_, new_n3045_ );
xor  ( new_n3086_, new_n3085_, new_n3059_ );
or   ( new_n3087_, new_n3086_, new_n3084_ );
and  ( new_n3088_, new_n3086_, new_n3084_ );
xor  ( new_n3089_, new_n2922_, new_n2920_ );
or   ( new_n3090_, new_n3089_, new_n3088_ );
and  ( new_n3091_, new_n3090_, new_n3087_ );
xor  ( new_n3092_, new_n2985_, new_n2980_ );
xnor ( new_n3093_, new_n3092_, new_n2987_ );
xnor ( new_n3094_, new_n2998_, new_n2994_ );
xor  ( new_n3095_, new_n3094_, new_n3004_ );
nand ( new_n3096_, new_n3095_, new_n3093_ );
or   ( new_n3097_, new_n1593_, new_n419_ );
or   ( new_n3098_, new_n1595_, new_n348_ );
and  ( new_n3099_, new_n3098_, new_n3097_ );
xor  ( new_n3100_, new_n3099_, new_n1358_ );
or   ( new_n3101_, new_n1364_, new_n509_ );
or   ( new_n3102_, new_n1366_, new_n443_ );
and  ( new_n3103_, new_n3102_, new_n3101_ );
xor  ( new_n3104_, new_n3103_, new_n1129_ );
nor  ( new_n3105_, new_n3104_, new_n3100_ );
or   ( new_n3106_, new_n1135_, new_n775_ );
or   ( new_n3107_, new_n1137_, new_n515_ );
and  ( new_n3108_, new_n3107_, new_n3106_ );
xor  ( new_n3109_, new_n3108_, new_n895_ );
nand ( new_n3110_, new_n3104_, new_n3100_ );
and  ( new_n3111_, new_n3110_, new_n3109_ );
or   ( new_n3112_, new_n3111_, new_n3105_ );
not  ( new_n3113_, RIbb2e620_35 );
and  ( new_n3114_, RIbb2e530_37, RIbb2e5a8_36 );
nor  ( new_n3115_, new_n3114_, new_n3113_ );
not  ( new_n3116_, new_n3115_ );
not  ( new_n3117_, new_n2930_ );
or   ( new_n3118_, new_n3117_, new_n333_ );
not  ( new_n3119_, new_n2928_ );
or   ( new_n3120_, new_n3119_, new_n339_ );
and  ( new_n3121_, new_n3120_, new_n3118_ );
xor  ( new_n3122_, new_n3121_, new_n2800_ );
nand ( new_n3123_, new_n3122_, new_n3116_ );
or   ( new_n3124_, new_n2807_, new_n313_ );
or   ( new_n3125_, new_n2809_, new_n319_ );
and  ( new_n3126_, new_n3125_, new_n3124_ );
xor  ( new_n3127_, new_n3126_, new_n2423_ );
nor  ( new_n3128_, new_n3122_, new_n3116_ );
or   ( new_n3129_, new_n3128_, new_n3127_ );
and  ( new_n3130_, new_n3129_, new_n3123_ );
nand ( new_n3131_, new_n3130_, new_n3112_ );
nor  ( new_n3132_, new_n3130_, new_n3112_ );
or   ( new_n3133_, new_n2425_, new_n279_ );
or   ( new_n3134_, new_n2427_, new_n285_ );
and  ( new_n3135_, new_n3134_, new_n3133_ );
xor  ( new_n3136_, new_n3135_, new_n2121_ );
or   ( new_n3137_, new_n2122_, new_n294_ );
or   ( new_n3138_, new_n2124_, new_n301_ );
and  ( new_n3139_, new_n3138_, new_n3137_ );
xor  ( new_n3140_, new_n3139_, new_n1843_ );
nor  ( new_n3141_, new_n3140_, new_n3136_ );
or   ( new_n3142_, new_n1844_, new_n264_ );
or   ( new_n3143_, new_n1846_, new_n270_ );
and  ( new_n3144_, new_n3143_, new_n3142_ );
xor  ( new_n3145_, new_n3144_, new_n1586_ );
and  ( new_n3146_, new_n3140_, new_n3136_ );
nor  ( new_n3147_, new_n3146_, new_n3145_ );
nor  ( new_n3148_, new_n3147_, new_n3141_ );
or   ( new_n3149_, new_n3148_, new_n3132_ );
and  ( new_n3150_, new_n3149_, new_n3131_ );
nor  ( new_n3151_, new_n3150_, new_n3096_ );
nand ( new_n3152_, new_n3150_, new_n3096_ );
or   ( new_n3153_, new_n897_, new_n886_ );
or   ( new_n3154_, new_n899_, new_n805_ );
and  ( new_n3155_, new_n3154_, new_n3153_ );
xor  ( new_n3156_, new_n3155_, new_n748_ );
or   ( new_n3157_, new_n755_, new_n1168_ );
or   ( new_n3158_, new_n757_, new_n986_ );
and  ( new_n3159_, new_n3158_, new_n3157_ );
xor  ( new_n3160_, new_n3159_, new_n523_ );
or   ( new_n3161_, new_n3160_, new_n3156_ );
or   ( new_n3162_, new_n524_, new_n1318_ );
or   ( new_n3163_, new_n526_, new_n1213_ );
and  ( new_n3164_, new_n3163_, new_n3162_ );
xor  ( new_n3165_, new_n3164_, new_n403_ );
and  ( new_n3166_, new_n3160_, new_n3156_ );
or   ( new_n3167_, new_n3166_, new_n3165_ );
and  ( new_n3168_, new_n3167_, new_n3161_ );
or   ( new_n3169_, new_n283_, new_n2475_ );
or   ( new_n3170_, new_n286_, new_n2291_ );
and  ( new_n3171_, new_n3170_, new_n3169_ );
xor  ( new_n3172_, new_n3171_, new_n278_ );
or   ( new_n3173_, new_n299_, new_n2751_ );
or   ( new_n3174_, new_n302_, new_n2646_ );
and  ( new_n3175_, new_n3174_, new_n3173_ );
xor  ( new_n3176_, new_n3175_, new_n293_ );
or   ( new_n3177_, new_n3176_, new_n3172_ );
not  ( new_n3178_, RIbb2c898_98 );
or   ( new_n3179_, new_n268_, new_n3178_ );
or   ( new_n3180_, new_n271_, new_n2981_ );
and  ( new_n3181_, new_n3180_, new_n3179_ );
xor  ( new_n3182_, new_n3181_, new_n263_ );
and  ( new_n3183_, new_n3176_, new_n3172_ );
or   ( new_n3184_, new_n3183_, new_n3182_ );
and  ( new_n3185_, new_n3184_, new_n3177_ );
nor  ( new_n3186_, new_n3185_, new_n3168_ );
nand ( new_n3187_, new_n3185_, new_n3168_ );
or   ( new_n3188_, new_n409_, new_n1523_ );
or   ( new_n3189_, new_n411_, new_n1525_ );
and  ( new_n3190_, new_n3189_, new_n3188_ );
xor  ( new_n3191_, new_n3190_, new_n328_ );
or   ( new_n3192_, new_n337_, new_n1899_ );
or   ( new_n3193_, new_n340_, new_n1754_ );
and  ( new_n3194_, new_n3193_, new_n3192_ );
xor  ( new_n3195_, new_n3194_, new_n332_ );
nor  ( new_n3196_, new_n3195_, new_n3191_ );
or   ( new_n3197_, new_n317_, new_n2178_ );
or   ( new_n3198_, new_n320_, new_n2057_ );
and  ( new_n3199_, new_n3198_, new_n3197_ );
xor  ( new_n3200_, new_n3199_, new_n312_ );
not  ( new_n3201_, new_n3200_ );
nand ( new_n3202_, new_n3195_, new_n3191_ );
and  ( new_n3203_, new_n3202_, new_n3201_ );
or   ( new_n3204_, new_n3203_, new_n3196_ );
and  ( new_n3205_, new_n3204_, new_n3187_ );
or   ( new_n3206_, new_n3205_, new_n3186_ );
and  ( new_n3207_, new_n3206_, new_n3152_ );
or   ( new_n3208_, new_n3207_, new_n3151_ );
xor  ( new_n3209_, new_n3033_, new_n3031_ );
xor  ( new_n3210_, new_n3209_, new_n3037_ );
xnor ( new_n3211_, new_n2948_, new_n2944_ );
xor  ( new_n3212_, new_n3211_, new_n2954_ );
xor  ( new_n3213_, new_n2966_, new_n2962_ );
xor  ( new_n3214_, new_n3213_, new_n2972_ );
or   ( new_n3215_, new_n3214_, new_n3212_ );
and  ( new_n3216_, new_n3214_, new_n3212_ );
xnor ( new_n3217_, new_n3016_, new_n3012_ );
xor  ( new_n3218_, new_n3217_, new_n3022_ );
or   ( new_n3219_, new_n3218_, new_n3216_ );
and  ( new_n3220_, new_n3219_, new_n3215_ );
or   ( new_n3221_, new_n3220_, new_n3210_ );
and  ( new_n3222_, new_n3220_, new_n3210_ );
xor  ( new_n3223_, new_n3049_, new_n3047_ );
xor  ( new_n3224_, new_n3223_, new_n3053_ );
or   ( new_n3225_, new_n3224_, new_n3222_ );
and  ( new_n3226_, new_n3225_, new_n3221_ );
nand ( new_n3227_, new_n3226_, new_n3208_ );
nor  ( new_n3228_, new_n3226_, new_n3208_ );
xor  ( new_n3229_, new_n3006_, new_n2990_ );
xnor ( new_n3230_, new_n3229_, new_n3024_ );
xor  ( new_n3231_, new_n2956_, new_n2940_ );
xor  ( new_n3232_, new_n3231_, new_n2974_ );
nor  ( new_n3233_, new_n3232_, new_n3230_ );
or   ( new_n3234_, new_n3233_, new_n3228_ );
and  ( new_n3235_, new_n3234_, new_n3227_ );
or   ( new_n3236_, new_n3235_, new_n3091_ );
and  ( new_n3237_, new_n3235_, new_n3091_ );
xor  ( new_n3238_, new_n2911_, new_n2909_ );
xor  ( new_n3239_, new_n3238_, new_n2914_ );
or   ( new_n3240_, new_n3239_, new_n3237_ );
and  ( new_n3241_, new_n3240_, new_n3236_ );
or   ( new_n3242_, new_n3241_, new_n3082_ );
nand ( new_n3243_, new_n3241_, new_n3082_ );
xor  ( new_n3244_, new_n2881_, new_n2863_ );
xnor ( new_n3245_, new_n3244_, new_n2888_ );
nand ( new_n3246_, new_n3245_, new_n3243_ );
and  ( new_n3247_, new_n3246_, new_n3242_ );
and  ( new_n3248_, new_n3247_, new_n3080_ );
xor  ( new_n3249_, new_n3075_, new_n3073_ );
and  ( new_n3250_, new_n3249_, new_n3248_ );
xor  ( new_n3251_, new_n3086_, new_n3084_ );
xor  ( new_n3252_, new_n3251_, new_n3089_ );
or   ( new_n3253_, new_n2425_, new_n301_ );
or   ( new_n3254_, new_n2427_, new_n279_ );
and  ( new_n3255_, new_n3254_, new_n3253_ );
xor  ( new_n3256_, new_n3255_, new_n2121_ );
or   ( new_n3257_, new_n2122_, new_n270_ );
or   ( new_n3258_, new_n2124_, new_n294_ );
and  ( new_n3259_, new_n3258_, new_n3257_ );
xor  ( new_n3260_, new_n3259_, new_n1843_ );
or   ( new_n3261_, new_n3260_, new_n3256_ );
or   ( new_n3262_, new_n1844_, new_n348_ );
or   ( new_n3263_, new_n1846_, new_n264_ );
and  ( new_n3264_, new_n3263_, new_n3262_ );
xor  ( new_n3265_, new_n3264_, new_n1586_ );
and  ( new_n3266_, new_n3260_, new_n3256_ );
or   ( new_n3267_, new_n3266_, new_n3265_ );
and  ( new_n3268_, new_n3267_, new_n3261_ );
or   ( new_n3269_, new_n1593_, new_n443_ );
or   ( new_n3270_, new_n1595_, new_n419_ );
and  ( new_n3271_, new_n3270_, new_n3269_ );
xor  ( new_n3272_, new_n3271_, new_n1358_ );
or   ( new_n3273_, new_n1364_, new_n515_ );
or   ( new_n3274_, new_n1366_, new_n509_ );
and  ( new_n3275_, new_n3274_, new_n3273_ );
xor  ( new_n3276_, new_n3275_, new_n1129_ );
or   ( new_n3277_, new_n3276_, new_n3272_ );
or   ( new_n3278_, new_n1135_, new_n805_ );
or   ( new_n3279_, new_n1137_, new_n775_ );
and  ( new_n3280_, new_n3279_, new_n3278_ );
xor  ( new_n3281_, new_n3280_, new_n896_ );
and  ( new_n3282_, new_n3276_, new_n3272_ );
or   ( new_n3283_, new_n3282_, new_n3281_ );
and  ( new_n3284_, new_n3283_, new_n3277_ );
or   ( new_n3285_, new_n3284_, new_n3268_ );
and  ( new_n3286_, new_n3284_, new_n3268_ );
or   ( new_n3287_, new_n3117_, new_n319_ );
or   ( new_n3288_, new_n3119_, new_n333_ );
and  ( new_n3289_, new_n3288_, new_n3287_ );
xor  ( new_n3290_, new_n3289_, new_n2799_ );
xor  ( new_n3291_, RIbb2e530_37, RIbb2e5a8_36 );
xor  ( new_n3292_, RIbb2e5a8_36, new_n3113_ );
nor  ( new_n3293_, new_n3292_, new_n3291_ );
and  ( new_n3294_, new_n3293_, RIbb2d810_65 );
xor  ( new_n3295_, new_n3294_, new_n3116_ );
and  ( new_n3296_, new_n3295_, new_n3290_ );
or   ( new_n3297_, new_n2807_, new_n285_ );
or   ( new_n3298_, new_n2809_, new_n313_ );
and  ( new_n3299_, new_n3298_, new_n3297_ );
xor  ( new_n3300_, new_n3299_, new_n2424_ );
nor  ( new_n3301_, new_n3295_, new_n3290_ );
nor  ( new_n3302_, new_n3301_, new_n3300_ );
nor  ( new_n3303_, new_n3302_, new_n3296_ );
or   ( new_n3304_, new_n3303_, new_n3286_ );
and  ( new_n3305_, new_n3304_, new_n3285_ );
not  ( new_n3306_, RIbb2c820_99 );
or   ( new_n3307_, new_n3306_, new_n260_ );
xnor ( new_n3308_, new_n3176_, new_n3172_ );
xor  ( new_n3309_, new_n3308_, new_n3182_ );
nand ( new_n3310_, new_n3309_, new_n3307_ );
or   ( new_n3311_, new_n3309_, new_n3307_ );
xor  ( new_n3312_, new_n3195_, new_n3191_ );
xor  ( new_n3313_, new_n3312_, new_n3201_ );
nand ( new_n3314_, new_n3313_, new_n3311_ );
and  ( new_n3315_, new_n3314_, new_n3310_ );
nor  ( new_n3316_, new_n3315_, new_n3305_ );
nand ( new_n3317_, new_n3315_, new_n3305_ );
or   ( new_n3318_, new_n283_, new_n2646_ );
or   ( new_n3319_, new_n286_, new_n2475_ );
and  ( new_n3320_, new_n3319_, new_n3318_ );
xor  ( new_n3321_, new_n3320_, new_n278_ );
or   ( new_n3322_, new_n299_, new_n2981_ );
or   ( new_n3323_, new_n302_, new_n2751_ );
and  ( new_n3324_, new_n3323_, new_n3322_ );
xor  ( new_n3325_, new_n3324_, new_n293_ );
or   ( new_n3326_, new_n3325_, new_n3321_ );
or   ( new_n3327_, new_n268_, new_n3306_ );
or   ( new_n3328_, new_n271_, new_n3178_ );
and  ( new_n3329_, new_n3328_, new_n3327_ );
xor  ( new_n3330_, new_n3329_, new_n263_ );
and  ( new_n3331_, new_n3325_, new_n3321_ );
or   ( new_n3332_, new_n3331_, new_n3330_ );
and  ( new_n3333_, new_n3332_, new_n3326_ );
or   ( new_n3334_, new_n897_, new_n986_ );
or   ( new_n3335_, new_n899_, new_n886_ );
and  ( new_n3336_, new_n3335_, new_n3334_ );
xor  ( new_n3337_, new_n3336_, new_n748_ );
or   ( new_n3338_, new_n755_, new_n1213_ );
or   ( new_n3339_, new_n757_, new_n1168_ );
and  ( new_n3340_, new_n3339_, new_n3338_ );
xor  ( new_n3341_, new_n3340_, new_n523_ );
or   ( new_n3342_, new_n3341_, new_n3337_ );
or   ( new_n3343_, new_n524_, new_n1525_ );
or   ( new_n3344_, new_n526_, new_n1318_ );
and  ( new_n3345_, new_n3344_, new_n3343_ );
xor  ( new_n3346_, new_n3345_, new_n403_ );
and  ( new_n3347_, new_n3341_, new_n3337_ );
or   ( new_n3348_, new_n3347_, new_n3346_ );
and  ( new_n3349_, new_n3348_, new_n3342_ );
nor  ( new_n3350_, new_n3349_, new_n3333_ );
nand ( new_n3351_, new_n3349_, new_n3333_ );
or   ( new_n3352_, new_n409_, new_n1754_ );
or   ( new_n3353_, new_n411_, new_n1523_ );
and  ( new_n3354_, new_n3353_, new_n3352_ );
xor  ( new_n3355_, new_n3354_, new_n328_ );
or   ( new_n3356_, new_n337_, new_n2057_ );
or   ( new_n3357_, new_n340_, new_n1899_ );
and  ( new_n3358_, new_n3357_, new_n3356_ );
xor  ( new_n3359_, new_n3358_, new_n332_ );
nor  ( new_n3360_, new_n3359_, new_n3355_ );
or   ( new_n3361_, new_n317_, new_n2291_ );
or   ( new_n3362_, new_n320_, new_n2178_ );
and  ( new_n3363_, new_n3362_, new_n3361_ );
xor  ( new_n3364_, new_n3363_, new_n312_ );
not  ( new_n3365_, new_n3364_ );
nand ( new_n3366_, new_n3359_, new_n3355_ );
and  ( new_n3367_, new_n3366_, new_n3365_ );
or   ( new_n3368_, new_n3367_, new_n3360_ );
and  ( new_n3369_, new_n3368_, new_n3351_ );
or   ( new_n3370_, new_n3369_, new_n3350_ );
and  ( new_n3371_, new_n3370_, new_n3317_ );
or   ( new_n3372_, new_n3371_, new_n3316_ );
xnor ( new_n3373_, new_n2932_, new_n2927_ );
xor  ( new_n3374_, new_n3373_, new_n2938_ );
xor  ( new_n3375_, new_n3104_, new_n3100_ );
xor  ( new_n3376_, new_n3375_, new_n3109_ );
xnor ( new_n3377_, new_n3160_, new_n3156_ );
xor  ( new_n3378_, new_n3377_, new_n3165_ );
or   ( new_n3379_, new_n3378_, new_n3376_ );
and  ( new_n3380_, new_n3378_, new_n3376_ );
xor  ( new_n3381_, new_n3140_, new_n3136_ );
xnor ( new_n3382_, new_n3381_, new_n3145_ );
or   ( new_n3383_, new_n3382_, new_n3380_ );
and  ( new_n3384_, new_n3383_, new_n3379_ );
or   ( new_n3385_, new_n3384_, new_n3374_ );
and  ( new_n3386_, new_n3384_, new_n3374_ );
xor  ( new_n3387_, new_n3214_, new_n3212_ );
xor  ( new_n3388_, new_n3387_, new_n3218_ );
or   ( new_n3389_, new_n3388_, new_n3386_ );
and  ( new_n3390_, new_n3389_, new_n3385_ );
nand ( new_n3391_, new_n3390_, new_n3372_ );
or   ( new_n3392_, new_n3390_, new_n3372_ );
xnor ( new_n3393_, new_n3130_, new_n3112_ );
xor  ( new_n3394_, new_n3393_, new_n3148_ );
xor  ( new_n3395_, new_n3185_, new_n3168_ );
xor  ( new_n3396_, new_n3395_, new_n3204_ );
nor  ( new_n3397_, new_n3396_, new_n3394_ );
and  ( new_n3398_, new_n3396_, new_n3394_ );
xor  ( new_n3399_, new_n3095_, new_n3093_ );
nor  ( new_n3400_, new_n3399_, new_n3398_ );
nor  ( new_n3401_, new_n3400_, new_n3397_ );
nand ( new_n3402_, new_n3401_, new_n3392_ );
and  ( new_n3403_, new_n3402_, new_n3391_ );
or   ( new_n3404_, new_n3403_, new_n3252_ );
nand ( new_n3405_, new_n3403_, new_n3252_ );
xor  ( new_n3406_, new_n3220_, new_n3210_ );
xor  ( new_n3407_, new_n3406_, new_n3224_ );
xor  ( new_n3408_, new_n3150_, new_n3096_ );
xor  ( new_n3409_, new_n3408_, new_n3206_ );
nor  ( new_n3410_, new_n3409_, new_n3407_ );
and  ( new_n3411_, new_n3409_, new_n3407_ );
not  ( new_n3412_, new_n3411_ );
xor  ( new_n3413_, new_n3232_, new_n3230_ );
and  ( new_n3414_, new_n3413_, new_n3412_ );
nor  ( new_n3415_, new_n3414_, new_n3410_ );
nand ( new_n3416_, new_n3415_, new_n3405_ );
and  ( new_n3417_, new_n3416_, new_n3404_ );
xor  ( new_n3418_, new_n3041_, new_n2923_ );
xor  ( new_n3419_, new_n3418_, new_n3061_ );
nand ( new_n3420_, new_n3419_, new_n3417_ );
nor  ( new_n3421_, new_n3419_, new_n3417_ );
xnor ( new_n3422_, new_n3235_, new_n3091_ );
xor  ( new_n3423_, new_n3422_, new_n3239_ );
or   ( new_n3424_, new_n3423_, new_n3421_ );
and  ( new_n3425_, new_n3424_, new_n3420_ );
xor  ( new_n3426_, new_n3241_, new_n3082_ );
xor  ( new_n3427_, new_n3426_, new_n3245_ );
nor  ( new_n3428_, new_n3427_, new_n3425_ );
xor  ( new_n3429_, new_n3247_, new_n3080_ );
and  ( new_n3430_, new_n3429_, new_n3428_ );
xor  ( new_n3431_, new_n3419_, new_n3417_ );
xor  ( new_n3432_, new_n3431_, new_n3423_ );
xor  ( new_n3433_, new_n3122_, new_n3116_ );
xor  ( new_n3434_, new_n3433_, new_n3127_ );
xnor ( new_n3435_, new_n3276_, new_n3272_ );
xor  ( new_n3436_, new_n3435_, new_n3281_ );
xnor ( new_n3437_, new_n3341_, new_n3337_ );
xor  ( new_n3438_, new_n3437_, new_n3346_ );
or   ( new_n3439_, new_n3438_, new_n3436_ );
and  ( new_n3440_, new_n3438_, new_n3436_ );
xor  ( new_n3441_, new_n3359_, new_n3355_ );
xor  ( new_n3442_, new_n3441_, new_n3365_ );
or   ( new_n3443_, new_n3442_, new_n3440_ );
and  ( new_n3444_, new_n3443_, new_n3439_ );
nor  ( new_n3445_, new_n3444_, new_n3434_ );
and  ( new_n3446_, new_n3444_, new_n3434_ );
xor  ( new_n3447_, new_n3378_, new_n3376_ );
xnor ( new_n3448_, new_n3447_, new_n3382_ );
not  ( new_n3449_, new_n3448_ );
nor  ( new_n3450_, new_n3449_, new_n3446_ );
nor  ( new_n3451_, new_n3450_, new_n3445_ );
and  ( new_n3452_, RIbb2c7a8_100, RIbb2f610_1 );
not  ( new_n3453_, new_n3452_ );
xnor ( new_n3454_, new_n3325_, new_n3321_ );
xor  ( new_n3455_, new_n3454_, new_n3330_ );
nand ( new_n3456_, new_n3455_, new_n3453_ );
not  ( new_n3457_, RIbb2e530_37 );
and  ( new_n3458_, RIbb2e440_39, RIbb2e4b8_38 );
nor  ( new_n3459_, new_n3458_, new_n3457_ );
not  ( new_n3460_, new_n3459_ );
not  ( new_n3461_, new_n3293_ );
or   ( new_n3462_, new_n3461_, new_n333_ );
not  ( new_n3463_, new_n3291_ );
or   ( new_n3464_, new_n3463_, new_n339_ );
and  ( new_n3465_, new_n3464_, new_n3462_ );
xor  ( new_n3466_, new_n3465_, new_n3116_ );
and  ( new_n3467_, new_n3466_, new_n3460_ );
or   ( new_n3468_, new_n3117_, new_n313_ );
or   ( new_n3469_, new_n3119_, new_n319_ );
and  ( new_n3470_, new_n3469_, new_n3468_ );
xor  ( new_n3471_, new_n3470_, new_n2800_ );
or   ( new_n3472_, new_n3466_, new_n3460_ );
and  ( new_n3473_, new_n3472_, new_n3471_ );
or   ( new_n3474_, new_n3473_, new_n3467_ );
or   ( new_n3475_, new_n2807_, new_n279_ );
or   ( new_n3476_, new_n2809_, new_n285_ );
and  ( new_n3477_, new_n3476_, new_n3475_ );
xor  ( new_n3478_, new_n3477_, new_n2424_ );
or   ( new_n3479_, new_n2425_, new_n294_ );
or   ( new_n3480_, new_n2427_, new_n301_ );
and  ( new_n3481_, new_n3480_, new_n3479_ );
xor  ( new_n3482_, new_n3481_, new_n2121_ );
or   ( new_n3483_, new_n3482_, new_n3478_ );
or   ( new_n3484_, new_n2122_, new_n264_ );
or   ( new_n3485_, new_n2124_, new_n270_ );
and  ( new_n3486_, new_n3485_, new_n3484_ );
xor  ( new_n3487_, new_n3486_, new_n1843_ );
and  ( new_n3488_, new_n3482_, new_n3478_ );
or   ( new_n3489_, new_n3488_, new_n3487_ );
and  ( new_n3490_, new_n3489_, new_n3483_ );
or   ( new_n3491_, new_n3490_, new_n3474_ );
and  ( new_n3492_, new_n3490_, new_n3474_ );
or   ( new_n3493_, new_n1844_, new_n419_ );
or   ( new_n3494_, new_n1846_, new_n348_ );
and  ( new_n3495_, new_n3494_, new_n3493_ );
xor  ( new_n3496_, new_n3495_, new_n1586_ );
or   ( new_n3497_, new_n1593_, new_n509_ );
or   ( new_n3498_, new_n1595_, new_n443_ );
and  ( new_n3499_, new_n3498_, new_n3497_ );
xor  ( new_n3500_, new_n3499_, new_n1358_ );
nor  ( new_n3501_, new_n3500_, new_n3496_ );
or   ( new_n3502_, new_n1364_, new_n775_ );
or   ( new_n3503_, new_n1366_, new_n515_ );
and  ( new_n3504_, new_n3503_, new_n3502_ );
xor  ( new_n3505_, new_n3504_, new_n1129_ );
and  ( new_n3506_, new_n3500_, new_n3496_ );
nor  ( new_n3507_, new_n3506_, new_n3505_ );
nor  ( new_n3508_, new_n3507_, new_n3501_ );
or   ( new_n3509_, new_n3508_, new_n3492_ );
and  ( new_n3510_, new_n3509_, new_n3491_ );
and  ( new_n3511_, new_n3510_, new_n3456_ );
or   ( new_n3512_, new_n1135_, new_n886_ );
or   ( new_n3513_, new_n1137_, new_n805_ );
and  ( new_n3514_, new_n3513_, new_n3512_ );
xor  ( new_n3515_, new_n3514_, new_n896_ );
or   ( new_n3516_, new_n897_, new_n1168_ );
or   ( new_n3517_, new_n899_, new_n986_ );
and  ( new_n3518_, new_n3517_, new_n3516_ );
xor  ( new_n3519_, new_n3518_, new_n748_ );
or   ( new_n3520_, new_n3519_, new_n3515_ );
or   ( new_n3521_, new_n755_, new_n1318_ );
or   ( new_n3522_, new_n757_, new_n1213_ );
and  ( new_n3523_, new_n3522_, new_n3521_ );
xor  ( new_n3524_, new_n3523_, new_n523_ );
and  ( new_n3525_, new_n3519_, new_n3515_ );
or   ( new_n3526_, new_n3525_, new_n3524_ );
and  ( new_n3527_, new_n3526_, new_n3520_ );
or   ( new_n3528_, new_n524_, new_n1523_ );
or   ( new_n3529_, new_n526_, new_n1525_ );
and  ( new_n3530_, new_n3529_, new_n3528_ );
xor  ( new_n3531_, new_n3530_, new_n403_ );
or   ( new_n3532_, new_n409_, new_n1899_ );
or   ( new_n3533_, new_n411_, new_n1754_ );
and  ( new_n3534_, new_n3533_, new_n3532_ );
xor  ( new_n3535_, new_n3534_, new_n328_ );
or   ( new_n3536_, new_n3535_, new_n3531_ );
or   ( new_n3537_, new_n337_, new_n2178_ );
or   ( new_n3538_, new_n340_, new_n2057_ );
and  ( new_n3539_, new_n3538_, new_n3537_ );
xor  ( new_n3540_, new_n3539_, new_n332_ );
and  ( new_n3541_, new_n3535_, new_n3531_ );
or   ( new_n3542_, new_n3541_, new_n3540_ );
and  ( new_n3543_, new_n3542_, new_n3536_ );
nor  ( new_n3544_, new_n3543_, new_n3527_ );
and  ( new_n3545_, new_n3543_, new_n3527_ );
or   ( new_n3546_, new_n317_, new_n2475_ );
or   ( new_n3547_, new_n320_, new_n2291_ );
and  ( new_n3548_, new_n3547_, new_n3546_ );
xor  ( new_n3549_, new_n3548_, new_n312_ );
or   ( new_n3550_, new_n283_, new_n2751_ );
or   ( new_n3551_, new_n286_, new_n2646_ );
and  ( new_n3552_, new_n3551_, new_n3550_ );
xor  ( new_n3553_, new_n3552_, new_n278_ );
nor  ( new_n3554_, new_n3553_, new_n3549_ );
or   ( new_n3555_, new_n299_, new_n3178_ );
or   ( new_n3556_, new_n302_, new_n2981_ );
and  ( new_n3557_, new_n3556_, new_n3555_ );
xor  ( new_n3558_, new_n3557_, new_n293_ );
and  ( new_n3559_, new_n3553_, new_n3549_ );
nor  ( new_n3560_, new_n3559_, new_n3558_ );
nor  ( new_n3561_, new_n3560_, new_n3554_ );
nor  ( new_n3562_, new_n3561_, new_n3545_ );
nor  ( new_n3563_, new_n3562_, new_n3544_ );
not  ( new_n3564_, new_n3563_ );
nor  ( new_n3565_, new_n3510_, new_n3456_ );
nor  ( new_n3566_, new_n3565_, new_n3564_ );
nor  ( new_n3567_, new_n3566_, new_n3511_ );
and  ( new_n3568_, new_n3567_, new_n3451_ );
not  ( new_n3569_, new_n3568_ );
xnor ( new_n3570_, new_n3284_, new_n3268_ );
xor  ( new_n3571_, new_n3570_, new_n3303_ );
xor  ( new_n3572_, new_n3349_, new_n3333_ );
xor  ( new_n3573_, new_n3572_, new_n3368_ );
nor  ( new_n3574_, new_n3573_, new_n3571_ );
and  ( new_n3575_, new_n3573_, new_n3571_ );
xor  ( new_n3576_, new_n3309_, new_n3307_ );
xor  ( new_n3577_, new_n3576_, new_n3313_ );
nor  ( new_n3578_, new_n3577_, new_n3575_ );
nor  ( new_n3579_, new_n3578_, new_n3574_ );
not  ( new_n3580_, new_n3579_ );
and  ( new_n3581_, new_n3580_, new_n3569_ );
nor  ( new_n3582_, new_n3567_, new_n3451_ );
or   ( new_n3583_, new_n3582_, new_n3581_ );
xor  ( new_n3584_, new_n3409_, new_n3407_ );
xor  ( new_n3585_, new_n3584_, new_n3413_ );
nor  ( new_n3586_, new_n3585_, new_n3583_ );
nand ( new_n3587_, new_n3585_, new_n3583_ );
xor  ( new_n3588_, new_n3384_, new_n3374_ );
xor  ( new_n3589_, new_n3588_, new_n3388_ );
xor  ( new_n3590_, new_n3315_, new_n3305_ );
xor  ( new_n3591_, new_n3590_, new_n3370_ );
nor  ( new_n3592_, new_n3591_, new_n3589_ );
and  ( new_n3593_, new_n3591_, new_n3589_ );
xor  ( new_n3594_, new_n3396_, new_n3394_ );
xor  ( new_n3595_, new_n3594_, new_n3399_ );
nor  ( new_n3596_, new_n3595_, new_n3593_ );
nor  ( new_n3597_, new_n3596_, new_n3592_ );
and  ( new_n3598_, new_n3597_, new_n3587_ );
or   ( new_n3599_, new_n3598_, new_n3586_ );
xnor ( new_n3600_, new_n3226_, new_n3208_ );
xor  ( new_n3601_, new_n3600_, new_n3233_ );
or   ( new_n3602_, new_n3601_, new_n3599_ );
and  ( new_n3603_, new_n3601_, new_n3599_ );
xor  ( new_n3604_, new_n3403_, new_n3252_ );
xor  ( new_n3605_, new_n3604_, new_n3415_ );
or   ( new_n3606_, new_n3605_, new_n3603_ );
and  ( new_n3607_, new_n3606_, new_n3602_ );
nor  ( new_n3608_, new_n3607_, new_n3432_ );
xor  ( new_n3609_, new_n3427_, new_n3425_ );
and  ( new_n3610_, new_n3609_, new_n3608_ );
xnor ( new_n3611_, new_n3585_, new_n3583_ );
xor  ( new_n3612_, new_n3611_, new_n3597_ );
xnor ( new_n3613_, new_n3591_, new_n3589_ );
xor  ( new_n3614_, new_n3613_, new_n3595_ );
xnor ( new_n3615_, new_n3260_, new_n3256_ );
xor  ( new_n3616_, new_n3615_, new_n3265_ );
xor  ( new_n3617_, new_n3466_, new_n3459_ );
xor  ( new_n3618_, new_n3617_, new_n3471_ );
xnor ( new_n3619_, new_n3482_, new_n3478_ );
xor  ( new_n3620_, new_n3619_, new_n3487_ );
or   ( new_n3621_, new_n3620_, new_n3618_ );
and  ( new_n3622_, new_n3620_, new_n3618_ );
xnor ( new_n3623_, new_n3500_, new_n3496_ );
xor  ( new_n3624_, new_n3623_, new_n3505_ );
or   ( new_n3625_, new_n3624_, new_n3622_ );
and  ( new_n3626_, new_n3625_, new_n3621_ );
nor  ( new_n3627_, new_n3626_, new_n3616_ );
nand ( new_n3628_, new_n3626_, new_n3616_ );
xnor ( new_n3629_, new_n3535_, new_n3531_ );
xor  ( new_n3630_, new_n3629_, new_n3540_ );
xnor ( new_n3631_, new_n3519_, new_n3515_ );
xor  ( new_n3632_, new_n3631_, new_n3524_ );
nor  ( new_n3633_, new_n3632_, new_n3630_ );
and  ( new_n3634_, new_n3632_, new_n3630_ );
xor  ( new_n3635_, new_n3553_, new_n3549_ );
xnor ( new_n3636_, new_n3635_, new_n3558_ );
nor  ( new_n3637_, new_n3636_, new_n3634_ );
nor  ( new_n3638_, new_n3637_, new_n3633_ );
not  ( new_n3639_, new_n3638_ );
and  ( new_n3640_, new_n3639_, new_n3628_ );
or   ( new_n3641_, new_n3640_, new_n3627_ );
or   ( new_n3642_, new_n524_, new_n1754_ );
or   ( new_n3643_, new_n526_, new_n1523_ );
and  ( new_n3644_, new_n3643_, new_n3642_ );
xor  ( new_n3645_, new_n3644_, new_n403_ );
or   ( new_n3646_, new_n409_, new_n2057_ );
or   ( new_n3647_, new_n411_, new_n1899_ );
and  ( new_n3648_, new_n3647_, new_n3646_ );
xor  ( new_n3649_, new_n3648_, new_n328_ );
or   ( new_n3650_, new_n3649_, new_n3645_ );
or   ( new_n3651_, new_n337_, new_n2291_ );
or   ( new_n3652_, new_n340_, new_n2178_ );
and  ( new_n3653_, new_n3652_, new_n3651_ );
xor  ( new_n3654_, new_n3653_, new_n332_ );
and  ( new_n3655_, new_n3649_, new_n3645_ );
or   ( new_n3656_, new_n3655_, new_n3654_ );
and  ( new_n3657_, new_n3656_, new_n3650_ );
or   ( new_n3658_, new_n1135_, new_n986_ );
or   ( new_n3659_, new_n1137_, new_n886_ );
and  ( new_n3660_, new_n3659_, new_n3658_ );
xor  ( new_n3661_, new_n3660_, new_n896_ );
or   ( new_n3662_, new_n897_, new_n1213_ );
or   ( new_n3663_, new_n899_, new_n1168_ );
and  ( new_n3664_, new_n3663_, new_n3662_ );
xor  ( new_n3665_, new_n3664_, new_n748_ );
or   ( new_n3666_, new_n3665_, new_n3661_ );
or   ( new_n3667_, new_n755_, new_n1525_ );
or   ( new_n3668_, new_n757_, new_n1318_ );
and  ( new_n3669_, new_n3668_, new_n3667_ );
xor  ( new_n3670_, new_n3669_, new_n523_ );
and  ( new_n3671_, new_n3665_, new_n3661_ );
or   ( new_n3672_, new_n3671_, new_n3670_ );
and  ( new_n3673_, new_n3672_, new_n3666_ );
nor  ( new_n3674_, new_n3673_, new_n3657_ );
and  ( new_n3675_, new_n3673_, new_n3657_ );
or   ( new_n3676_, new_n317_, new_n2646_ );
or   ( new_n3677_, new_n320_, new_n2475_ );
and  ( new_n3678_, new_n3677_, new_n3676_ );
xor  ( new_n3679_, new_n3678_, new_n312_ );
or   ( new_n3680_, new_n283_, new_n2981_ );
or   ( new_n3681_, new_n286_, new_n2751_ );
and  ( new_n3682_, new_n3681_, new_n3680_ );
xor  ( new_n3683_, new_n3682_, new_n278_ );
nor  ( new_n3684_, new_n3683_, new_n3679_ );
or   ( new_n3685_, new_n299_, new_n3306_ );
or   ( new_n3686_, new_n302_, new_n3178_ );
and  ( new_n3687_, new_n3686_, new_n3685_ );
xor  ( new_n3688_, new_n3687_, new_n293_ );
and  ( new_n3689_, new_n3683_, new_n3679_ );
nor  ( new_n3690_, new_n3689_, new_n3688_ );
nor  ( new_n3691_, new_n3690_, new_n3684_ );
nor  ( new_n3692_, new_n3691_, new_n3675_ );
nor  ( new_n3693_, new_n3692_, new_n3674_ );
not  ( new_n3694_, RIbb2c730_101 );
or   ( new_n3695_, new_n268_, new_n3694_ );
not  ( new_n3696_, RIbb2c7a8_100 );
or   ( new_n3697_, new_n271_, new_n3696_ );
and  ( new_n3698_, new_n3697_, new_n3695_ );
xor  ( new_n3699_, new_n3698_, new_n263_ );
and  ( new_n3700_, RIbb2c6b8_102, RIbb2f610_1 );
or   ( new_n3701_, new_n3700_, new_n3699_ );
or   ( new_n3702_, new_n268_, new_n3696_ );
or   ( new_n3703_, new_n271_, new_n3306_ );
and  ( new_n3704_, new_n3703_, new_n3702_ );
xor  ( new_n3705_, new_n3704_, new_n263_ );
or   ( new_n3706_, new_n3705_, new_n3701_ );
and  ( new_n3707_, RIbb2c730_101, RIbb2f610_1 );
and  ( new_n3708_, new_n3705_, new_n3701_ );
or   ( new_n3709_, new_n3708_, new_n3707_ );
and  ( new_n3710_, new_n3709_, new_n3706_ );
or   ( new_n3711_, new_n2807_, new_n301_ );
or   ( new_n3712_, new_n2809_, new_n279_ );
and  ( new_n3713_, new_n3712_, new_n3711_ );
xor  ( new_n3714_, new_n3713_, new_n2424_ );
or   ( new_n3715_, new_n2425_, new_n270_ );
or   ( new_n3716_, new_n2427_, new_n294_ );
and  ( new_n3717_, new_n3716_, new_n3715_ );
xor  ( new_n3718_, new_n3717_, new_n2121_ );
or   ( new_n3719_, new_n3718_, new_n3714_ );
or   ( new_n3720_, new_n2122_, new_n348_ );
or   ( new_n3721_, new_n2124_, new_n264_ );
and  ( new_n3722_, new_n3721_, new_n3720_ );
xor  ( new_n3723_, new_n3722_, new_n1843_ );
and  ( new_n3724_, new_n3718_, new_n3714_ );
or   ( new_n3725_, new_n3724_, new_n3723_ );
and  ( new_n3726_, new_n3725_, new_n3719_ );
or   ( new_n3727_, new_n3461_, new_n319_ );
or   ( new_n3728_, new_n3463_, new_n333_ );
and  ( new_n3729_, new_n3728_, new_n3727_ );
xor  ( new_n3730_, new_n3729_, new_n3115_ );
xor  ( new_n3731_, RIbb2e440_39, RIbb2e4b8_38 );
xor  ( new_n3732_, RIbb2e4b8_38, new_n3457_ );
nor  ( new_n3733_, new_n3732_, new_n3731_ );
and  ( new_n3734_, new_n3733_, RIbb2d810_65 );
xor  ( new_n3735_, new_n3734_, new_n3460_ );
nand ( new_n3736_, new_n3735_, new_n3730_ );
or   ( new_n3737_, new_n3117_, new_n285_ );
or   ( new_n3738_, new_n3119_, new_n313_ );
and  ( new_n3739_, new_n3738_, new_n3737_ );
xor  ( new_n3740_, new_n3739_, new_n2800_ );
nor  ( new_n3741_, new_n3735_, new_n3730_ );
or   ( new_n3742_, new_n3741_, new_n3740_ );
and  ( new_n3743_, new_n3742_, new_n3736_ );
or   ( new_n3744_, new_n3743_, new_n3726_ );
and  ( new_n3745_, new_n3743_, new_n3726_ );
or   ( new_n3746_, new_n1844_, new_n443_ );
or   ( new_n3747_, new_n1846_, new_n419_ );
and  ( new_n3748_, new_n3747_, new_n3746_ );
xor  ( new_n3749_, new_n3748_, new_n1586_ );
or   ( new_n3750_, new_n1593_, new_n515_ );
or   ( new_n3751_, new_n1595_, new_n509_ );
and  ( new_n3752_, new_n3751_, new_n3750_ );
xor  ( new_n3753_, new_n3752_, new_n1358_ );
nor  ( new_n3754_, new_n3753_, new_n3749_ );
or   ( new_n3755_, new_n1364_, new_n805_ );
or   ( new_n3756_, new_n1366_, new_n775_ );
and  ( new_n3757_, new_n3756_, new_n3755_ );
xor  ( new_n3758_, new_n3757_, new_n1129_ );
and  ( new_n3759_, new_n3753_, new_n3749_ );
nor  ( new_n3760_, new_n3759_, new_n3758_ );
nor  ( new_n3761_, new_n3760_, new_n3754_ );
or   ( new_n3762_, new_n3761_, new_n3745_ );
and  ( new_n3763_, new_n3762_, new_n3744_ );
and  ( new_n3764_, new_n3763_, new_n3710_ );
or   ( new_n3765_, new_n3764_, new_n3693_ );
or   ( new_n3766_, new_n3763_, new_n3710_ );
and  ( new_n3767_, new_n3766_, new_n3765_ );
or   ( new_n3768_, new_n3767_, new_n3641_ );
nand ( new_n3769_, new_n3767_, new_n3641_ );
xor  ( new_n3770_, new_n3295_, new_n3290_ );
xor  ( new_n3771_, new_n3770_, new_n3300_ );
xnor ( new_n3772_, new_n3438_, new_n3436_ );
xor  ( new_n3773_, new_n3772_, new_n3442_ );
and  ( new_n3774_, new_n3773_, new_n3771_ );
xor  ( new_n3775_, new_n3455_, new_n3453_ );
nor  ( new_n3776_, new_n3773_, new_n3771_ );
nor  ( new_n3777_, new_n3776_, new_n3775_ );
nor  ( new_n3778_, new_n3777_, new_n3774_ );
nand ( new_n3779_, new_n3778_, new_n3769_ );
and  ( new_n3780_, new_n3779_, new_n3768_ );
or   ( new_n3781_, new_n3780_, new_n3614_ );
nand ( new_n3782_, new_n3780_, new_n3614_ );
xor  ( new_n3783_, new_n3510_, new_n3456_ );
xor  ( new_n3784_, new_n3783_, new_n3564_ );
xor  ( new_n3785_, new_n3444_, new_n3434_ );
xor  ( new_n3786_, new_n3785_, new_n3449_ );
nor  ( new_n3787_, new_n3786_, new_n3784_ );
and  ( new_n3788_, new_n3786_, new_n3784_ );
not  ( new_n3789_, new_n3788_ );
xor  ( new_n3790_, new_n3573_, new_n3571_ );
xnor ( new_n3791_, new_n3790_, new_n3577_ );
and  ( new_n3792_, new_n3791_, new_n3789_ );
nor  ( new_n3793_, new_n3792_, new_n3787_ );
nand ( new_n3794_, new_n3793_, new_n3782_ );
and  ( new_n3795_, new_n3794_, new_n3781_ );
or   ( new_n3796_, new_n3795_, new_n3612_ );
nand ( new_n3797_, new_n3795_, new_n3612_ );
xor  ( new_n3798_, new_n3390_, new_n3372_ );
xor  ( new_n3799_, new_n3798_, new_n3401_ );
nand ( new_n3800_, new_n3799_, new_n3797_ );
and  ( new_n3801_, new_n3800_, new_n3796_ );
xnor ( new_n3802_, new_n3601_, new_n3599_ );
xor  ( new_n3803_, new_n3802_, new_n3605_ );
and  ( new_n3804_, new_n3803_, new_n3801_ );
xor  ( new_n3805_, new_n3607_, new_n3432_ );
and  ( new_n3806_, new_n3805_, new_n3804_ );
xor  ( new_n3807_, new_n3795_, new_n3612_ );
xor  ( new_n3808_, new_n3807_, new_n3799_ );
xor  ( new_n3809_, new_n3567_, new_n3451_ );
or   ( new_n3810_, new_n3809_, new_n3580_ );
not  ( new_n3811_, new_n3581_ );
or   ( new_n3812_, new_n3582_, new_n3811_ );
and  ( new_n3813_, new_n3812_, new_n3810_ );
xor  ( new_n3814_, new_n3786_, new_n3784_ );
xor  ( new_n3815_, new_n3814_, new_n3791_ );
or   ( new_n3816_, new_n299_, new_n3696_ );
or   ( new_n3817_, new_n302_, new_n3306_ );
and  ( new_n3818_, new_n3817_, new_n3816_ );
xor  ( new_n3819_, new_n3818_, new_n293_ );
not  ( new_n3820_, RIbb2c6b8_102 );
or   ( new_n3821_, new_n268_, new_n3820_ );
or   ( new_n3822_, new_n271_, new_n3694_ );
and  ( new_n3823_, new_n3822_, new_n3821_ );
xor  ( new_n3824_, new_n3823_, new_n263_ );
nor  ( new_n3825_, new_n3824_, new_n3819_ );
and  ( new_n3826_, RIbb2c640_103, RIbb2f610_1 );
not  ( new_n3827_, new_n3826_ );
nand ( new_n3828_, new_n3824_, new_n3819_ );
and  ( new_n3829_, new_n3828_, new_n3827_ );
or   ( new_n3830_, new_n3829_, new_n3825_ );
xnor ( new_n3831_, new_n3683_, new_n3679_ );
xor  ( new_n3832_, new_n3831_, new_n3688_ );
nor  ( new_n3833_, new_n3832_, new_n3830_ );
xor  ( new_n3834_, new_n3700_, new_n3699_ );
and  ( new_n3835_, new_n3832_, new_n3830_ );
nor  ( new_n3836_, new_n3835_, new_n3834_ );
or   ( new_n3837_, new_n3836_, new_n3833_ );
or   ( new_n3838_, new_n1364_, new_n886_ );
or   ( new_n3839_, new_n1366_, new_n805_ );
and  ( new_n3840_, new_n3839_, new_n3838_ );
xor  ( new_n3841_, new_n3840_, new_n1129_ );
or   ( new_n3842_, new_n1135_, new_n1168_ );
or   ( new_n3843_, new_n1137_, new_n986_ );
and  ( new_n3844_, new_n3843_, new_n3842_ );
xor  ( new_n3845_, new_n3844_, new_n896_ );
or   ( new_n3846_, new_n3845_, new_n3841_ );
and  ( new_n3847_, new_n3845_, new_n3841_ );
or   ( new_n3848_, new_n897_, new_n1318_ );
or   ( new_n3849_, new_n899_, new_n1213_ );
and  ( new_n3850_, new_n3849_, new_n3848_ );
xor  ( new_n3851_, new_n3850_, new_n748_ );
or   ( new_n3852_, new_n3851_, new_n3847_ );
and  ( new_n3853_, new_n3852_, new_n3846_ );
or   ( new_n3854_, new_n755_, new_n1523_ );
or   ( new_n3855_, new_n757_, new_n1525_ );
and  ( new_n3856_, new_n3855_, new_n3854_ );
xor  ( new_n3857_, new_n3856_, new_n523_ );
or   ( new_n3858_, new_n524_, new_n1899_ );
or   ( new_n3859_, new_n526_, new_n1754_ );
and  ( new_n3860_, new_n3859_, new_n3858_ );
xor  ( new_n3861_, new_n3860_, new_n403_ );
or   ( new_n3862_, new_n3861_, new_n3857_ );
and  ( new_n3863_, new_n3861_, new_n3857_ );
or   ( new_n3864_, new_n409_, new_n2178_ );
or   ( new_n3865_, new_n411_, new_n2057_ );
and  ( new_n3866_, new_n3865_, new_n3864_ );
xor  ( new_n3867_, new_n3866_, new_n328_ );
or   ( new_n3868_, new_n3867_, new_n3863_ );
and  ( new_n3869_, new_n3868_, new_n3862_ );
or   ( new_n3870_, new_n3869_, new_n3853_ );
and  ( new_n3871_, new_n3869_, new_n3853_ );
or   ( new_n3872_, new_n337_, new_n2475_ );
or   ( new_n3873_, new_n340_, new_n2291_ );
and  ( new_n3874_, new_n3873_, new_n3872_ );
xor  ( new_n3875_, new_n3874_, new_n332_ );
or   ( new_n3876_, new_n317_, new_n2751_ );
or   ( new_n3877_, new_n320_, new_n2646_ );
and  ( new_n3878_, new_n3877_, new_n3876_ );
xor  ( new_n3879_, new_n3878_, new_n312_ );
nor  ( new_n3880_, new_n3879_, new_n3875_ );
or   ( new_n3881_, new_n283_, new_n3178_ );
or   ( new_n3882_, new_n286_, new_n2981_ );
and  ( new_n3883_, new_n3882_, new_n3881_ );
xor  ( new_n3884_, new_n3883_, new_n278_ );
and  ( new_n3885_, new_n3879_, new_n3875_ );
nor  ( new_n3886_, new_n3885_, new_n3884_ );
nor  ( new_n3887_, new_n3886_, new_n3880_ );
or   ( new_n3888_, new_n3887_, new_n3871_ );
and  ( new_n3889_, new_n3888_, new_n3870_ );
nor  ( new_n3890_, new_n3889_, new_n3837_ );
nand ( new_n3891_, new_n3889_, new_n3837_ );
not  ( new_n3892_, RIbb2e440_39 );
and  ( new_n3893_, RIbb2e350_41, RIbb2e3c8_40 );
nor  ( new_n3894_, new_n3893_, new_n3892_ );
not  ( new_n3895_, new_n3894_ );
not  ( new_n3896_, new_n3733_ );
or   ( new_n3897_, new_n3896_, new_n333_ );
not  ( new_n3898_, new_n3731_ );
or   ( new_n3899_, new_n3898_, new_n339_ );
and  ( new_n3900_, new_n3899_, new_n3897_ );
xor  ( new_n3901_, new_n3900_, new_n3460_ );
and  ( new_n3902_, new_n3901_, new_n3895_ );
or   ( new_n3903_, new_n3901_, new_n3895_ );
or   ( new_n3904_, new_n3461_, new_n313_ );
or   ( new_n3905_, new_n3463_, new_n319_ );
and  ( new_n3906_, new_n3905_, new_n3904_ );
xor  ( new_n3907_, new_n3906_, new_n3116_ );
and  ( new_n3908_, new_n3907_, new_n3903_ );
or   ( new_n3909_, new_n3908_, new_n3902_ );
or   ( new_n3910_, new_n3117_, new_n279_ );
or   ( new_n3911_, new_n3119_, new_n285_ );
and  ( new_n3912_, new_n3911_, new_n3910_ );
xor  ( new_n3913_, new_n3912_, new_n2800_ );
or   ( new_n3914_, new_n2807_, new_n294_ );
or   ( new_n3915_, new_n2809_, new_n301_ );
and  ( new_n3916_, new_n3915_, new_n3914_ );
xor  ( new_n3917_, new_n3916_, new_n2424_ );
or   ( new_n3918_, new_n3917_, new_n3913_ );
and  ( new_n3919_, new_n3917_, new_n3913_ );
or   ( new_n3920_, new_n2425_, new_n264_ );
or   ( new_n3921_, new_n2427_, new_n270_ );
and  ( new_n3922_, new_n3921_, new_n3920_ );
xor  ( new_n3923_, new_n3922_, new_n2121_ );
or   ( new_n3924_, new_n3923_, new_n3919_ );
and  ( new_n3925_, new_n3924_, new_n3918_ );
nor  ( new_n3926_, new_n3925_, new_n3909_ );
and  ( new_n3927_, new_n3925_, new_n3909_ );
or   ( new_n3928_, new_n2122_, new_n419_ );
or   ( new_n3929_, new_n2124_, new_n348_ );
and  ( new_n3930_, new_n3929_, new_n3928_ );
xor  ( new_n3931_, new_n3930_, new_n1843_ );
or   ( new_n3932_, new_n1844_, new_n509_ );
or   ( new_n3933_, new_n1846_, new_n443_ );
and  ( new_n3934_, new_n3933_, new_n3932_ );
xor  ( new_n3935_, new_n3934_, new_n1586_ );
nor  ( new_n3936_, new_n3935_, new_n3931_ );
and  ( new_n3937_, new_n3935_, new_n3931_ );
or   ( new_n3938_, new_n1593_, new_n775_ );
or   ( new_n3939_, new_n1595_, new_n515_ );
and  ( new_n3940_, new_n3939_, new_n3938_ );
xor  ( new_n3941_, new_n3940_, new_n1358_ );
nor  ( new_n3942_, new_n3941_, new_n3937_ );
nor  ( new_n3943_, new_n3942_, new_n3936_ );
nor  ( new_n3944_, new_n3943_, new_n3927_ );
nor  ( new_n3945_, new_n3944_, new_n3926_ );
not  ( new_n3946_, new_n3945_ );
and  ( new_n3947_, new_n3946_, new_n3891_ );
or   ( new_n3948_, new_n3947_, new_n3890_ );
xor  ( new_n3949_, new_n3735_, new_n3730_ );
xnor ( new_n3950_, new_n3949_, new_n3740_ );
xnor ( new_n3951_, new_n3718_, new_n3714_ );
xor  ( new_n3952_, new_n3951_, new_n3723_ );
or   ( new_n3953_, new_n3952_, new_n3950_ );
xnor ( new_n3954_, new_n3665_, new_n3661_ );
xor  ( new_n3955_, new_n3954_, new_n3670_ );
xnor ( new_n3956_, new_n3649_, new_n3645_ );
xor  ( new_n3957_, new_n3956_, new_n3654_ );
or   ( new_n3958_, new_n3957_, new_n3955_ );
and  ( new_n3959_, new_n3957_, new_n3955_ );
xnor ( new_n3960_, new_n3753_, new_n3749_ );
xor  ( new_n3961_, new_n3960_, new_n3758_ );
or   ( new_n3962_, new_n3961_, new_n3959_ );
and  ( new_n3963_, new_n3962_, new_n3958_ );
or   ( new_n3964_, new_n3963_, new_n3953_ );
and  ( new_n3965_, new_n3963_, new_n3953_ );
xor  ( new_n3966_, new_n3620_, new_n3618_ );
xor  ( new_n3967_, new_n3966_, new_n3624_ );
or   ( new_n3968_, new_n3967_, new_n3965_ );
and  ( new_n3969_, new_n3968_, new_n3964_ );
nand ( new_n3970_, new_n3969_, new_n3948_ );
or   ( new_n3971_, new_n3969_, new_n3948_ );
xnor ( new_n3972_, new_n3673_, new_n3657_ );
xor  ( new_n3973_, new_n3972_, new_n3691_ );
xnor ( new_n3974_, new_n3705_, new_n3701_ );
xor  ( new_n3975_, new_n3974_, new_n3707_ );
nor  ( new_n3976_, new_n3975_, new_n3973_ );
and  ( new_n3977_, new_n3975_, new_n3973_ );
xor  ( new_n3978_, new_n3632_, new_n3630_ );
xnor ( new_n3979_, new_n3978_, new_n3636_ );
not  ( new_n3980_, new_n3979_ );
nor  ( new_n3981_, new_n3980_, new_n3977_ );
nor  ( new_n3982_, new_n3981_, new_n3976_ );
nand ( new_n3983_, new_n3982_, new_n3971_ );
and  ( new_n3984_, new_n3983_, new_n3970_ );
or   ( new_n3985_, new_n3984_, new_n3815_ );
nand ( new_n3986_, new_n3984_, new_n3815_ );
xnor ( new_n3987_, new_n3490_, new_n3474_ );
xor  ( new_n3988_, new_n3987_, new_n3508_ );
xnor ( new_n3989_, new_n3543_, new_n3527_ );
xor  ( new_n3990_, new_n3989_, new_n3561_ );
nor  ( new_n3991_, new_n3990_, new_n3988_ );
and  ( new_n3992_, new_n3990_, new_n3988_ );
xor  ( new_n3993_, new_n3773_, new_n3771_ );
xnor ( new_n3994_, new_n3993_, new_n3775_ );
not  ( new_n3995_, new_n3994_ );
nor  ( new_n3996_, new_n3995_, new_n3992_ );
nor  ( new_n3997_, new_n3996_, new_n3991_ );
nand ( new_n3998_, new_n3997_, new_n3986_ );
and  ( new_n3999_, new_n3998_, new_n3985_ );
nand ( new_n4000_, new_n3999_, new_n3813_ );
nor  ( new_n4001_, new_n3999_, new_n3813_ );
xor  ( new_n4002_, new_n3780_, new_n3614_ );
xor  ( new_n4003_, new_n4002_, new_n3793_ );
or   ( new_n4004_, new_n4003_, new_n4001_ );
and  ( new_n4005_, new_n4004_, new_n4000_ );
nor  ( new_n4006_, new_n4005_, new_n3808_ );
xor  ( new_n4007_, new_n3803_, new_n3801_ );
and  ( new_n4008_, new_n4007_, new_n4006_ );
xor  ( new_n4009_, new_n3767_, new_n3641_ );
xor  ( new_n4010_, new_n4009_, new_n3778_ );
not  ( new_n4011_, new_n4010_ );
or   ( new_n4012_, new_n3117_, new_n301_ );
or   ( new_n4013_, new_n3119_, new_n279_ );
and  ( new_n4014_, new_n4013_, new_n4012_ );
xor  ( new_n4015_, new_n4014_, new_n2800_ );
or   ( new_n4016_, new_n2807_, new_n270_ );
or   ( new_n4017_, new_n2809_, new_n294_ );
and  ( new_n4018_, new_n4017_, new_n4016_ );
xor  ( new_n4019_, new_n4018_, new_n2424_ );
or   ( new_n4020_, new_n4019_, new_n4015_ );
and  ( new_n4021_, new_n4019_, new_n4015_ );
or   ( new_n4022_, new_n2425_, new_n348_ );
or   ( new_n4023_, new_n2427_, new_n264_ );
and  ( new_n4024_, new_n4023_, new_n4022_ );
xor  ( new_n4025_, new_n4024_, new_n2121_ );
or   ( new_n4026_, new_n4025_, new_n4021_ );
and  ( new_n4027_, new_n4026_, new_n4020_ );
or   ( new_n4028_, new_n3896_, new_n319_ );
or   ( new_n4029_, new_n3898_, new_n333_ );
and  ( new_n4030_, new_n4029_, new_n4028_ );
xor  ( new_n4031_, new_n4030_, new_n3459_ );
xor  ( new_n4032_, RIbb2e350_41, RIbb2e3c8_40 );
xor  ( new_n4033_, RIbb2e3c8_40, new_n3892_ );
nor  ( new_n4034_, new_n4033_, new_n4032_ );
and  ( new_n4035_, new_n4034_, RIbb2d810_65 );
xor  ( new_n4036_, new_n4035_, new_n3895_ );
nand ( new_n4037_, new_n4036_, new_n4031_ );
nor  ( new_n4038_, new_n4036_, new_n4031_ );
or   ( new_n4039_, new_n3461_, new_n285_ );
or   ( new_n4040_, new_n3463_, new_n313_ );
and  ( new_n4041_, new_n4040_, new_n4039_ );
xor  ( new_n4042_, new_n4041_, new_n3116_ );
or   ( new_n4043_, new_n4042_, new_n4038_ );
and  ( new_n4044_, new_n4043_, new_n4037_ );
or   ( new_n4045_, new_n4044_, new_n4027_ );
and  ( new_n4046_, new_n4044_, new_n4027_ );
or   ( new_n4047_, new_n2122_, new_n443_ );
or   ( new_n4048_, new_n2124_, new_n419_ );
and  ( new_n4049_, new_n4048_, new_n4047_ );
xor  ( new_n4050_, new_n4049_, new_n1843_ );
or   ( new_n4051_, new_n1844_, new_n515_ );
or   ( new_n4052_, new_n1846_, new_n509_ );
and  ( new_n4053_, new_n4052_, new_n4051_ );
xor  ( new_n4054_, new_n4053_, new_n1586_ );
nor  ( new_n4055_, new_n4054_, new_n4050_ );
and  ( new_n4056_, new_n4054_, new_n4050_ );
or   ( new_n4057_, new_n1593_, new_n805_ );
or   ( new_n4058_, new_n1595_, new_n775_ );
and  ( new_n4059_, new_n4058_, new_n4057_ );
xor  ( new_n4060_, new_n4059_, new_n1358_ );
nor  ( new_n4061_, new_n4060_, new_n4056_ );
nor  ( new_n4062_, new_n4061_, new_n4055_ );
or   ( new_n4063_, new_n4062_, new_n4046_ );
and  ( new_n4064_, new_n4063_, new_n4045_ );
or   ( new_n4065_, new_n299_, new_n3694_ );
or   ( new_n4066_, new_n302_, new_n3696_ );
and  ( new_n4067_, new_n4066_, new_n4065_ );
xor  ( new_n4068_, new_n4067_, new_n293_ );
not  ( new_n4069_, RIbb2c640_103 );
or   ( new_n4070_, new_n268_, new_n4069_ );
or   ( new_n4071_, new_n271_, new_n3820_ );
and  ( new_n4072_, new_n4071_, new_n4070_ );
xor  ( new_n4073_, new_n4072_, new_n263_ );
nor  ( new_n4074_, new_n4073_, new_n4068_ );
and  ( new_n4075_, RIbb2c5c8_104, RIbb2f610_1 );
not  ( new_n4076_, new_n4075_ );
nand ( new_n4077_, new_n4073_, new_n4068_ );
and  ( new_n4078_, new_n4077_, new_n4076_ );
or   ( new_n4079_, new_n4078_, new_n4074_ );
xnor ( new_n4080_, new_n3879_, new_n3875_ );
xor  ( new_n4081_, new_n4080_, new_n3884_ );
nand ( new_n4082_, new_n4081_, new_n4079_ );
or   ( new_n4083_, new_n4081_, new_n4079_ );
xor  ( new_n4084_, new_n3824_, new_n3819_ );
xor  ( new_n4085_, new_n4084_, new_n3827_ );
nand ( new_n4086_, new_n4085_, new_n4083_ );
and  ( new_n4087_, new_n4086_, new_n4082_ );
nor  ( new_n4088_, new_n4087_, new_n4064_ );
nand ( new_n4089_, new_n4087_, new_n4064_ );
or   ( new_n4090_, new_n1364_, new_n986_ );
or   ( new_n4091_, new_n1366_, new_n886_ );
and  ( new_n4092_, new_n4091_, new_n4090_ );
xor  ( new_n4093_, new_n4092_, new_n1129_ );
or   ( new_n4094_, new_n1135_, new_n1213_ );
or   ( new_n4095_, new_n1137_, new_n1168_ );
and  ( new_n4096_, new_n4095_, new_n4094_ );
xor  ( new_n4097_, new_n4096_, new_n896_ );
or   ( new_n4098_, new_n4097_, new_n4093_ );
and  ( new_n4099_, new_n4097_, new_n4093_ );
or   ( new_n4100_, new_n897_, new_n1525_ );
or   ( new_n4101_, new_n899_, new_n1318_ );
and  ( new_n4102_, new_n4101_, new_n4100_ );
xor  ( new_n4103_, new_n4102_, new_n748_ );
or   ( new_n4104_, new_n4103_, new_n4099_ );
and  ( new_n4105_, new_n4104_, new_n4098_ );
or   ( new_n4106_, new_n337_, new_n2646_ );
or   ( new_n4107_, new_n340_, new_n2475_ );
and  ( new_n4108_, new_n4107_, new_n4106_ );
xor  ( new_n4109_, new_n4108_, new_n332_ );
or   ( new_n4110_, new_n317_, new_n2981_ );
or   ( new_n4111_, new_n320_, new_n2751_ );
and  ( new_n4112_, new_n4111_, new_n4110_ );
xor  ( new_n4113_, new_n4112_, new_n312_ );
or   ( new_n4114_, new_n4113_, new_n4109_ );
and  ( new_n4115_, new_n4113_, new_n4109_ );
or   ( new_n4116_, new_n283_, new_n3306_ );
or   ( new_n4117_, new_n286_, new_n3178_ );
and  ( new_n4118_, new_n4117_, new_n4116_ );
xor  ( new_n4119_, new_n4118_, new_n278_ );
or   ( new_n4120_, new_n4119_, new_n4115_ );
and  ( new_n4121_, new_n4120_, new_n4114_ );
nor  ( new_n4122_, new_n4121_, new_n4105_ );
nand ( new_n4123_, new_n4121_, new_n4105_ );
or   ( new_n4124_, new_n755_, new_n1754_ );
or   ( new_n4125_, new_n757_, new_n1523_ );
and  ( new_n4126_, new_n4125_, new_n4124_ );
xor  ( new_n4127_, new_n4126_, new_n523_ );
or   ( new_n4128_, new_n524_, new_n2057_ );
or   ( new_n4129_, new_n526_, new_n1899_ );
and  ( new_n4130_, new_n4129_, new_n4128_ );
xor  ( new_n4131_, new_n4130_, new_n403_ );
nor  ( new_n4132_, new_n4131_, new_n4127_ );
nand ( new_n4133_, new_n4131_, new_n4127_ );
or   ( new_n4134_, new_n409_, new_n2291_ );
or   ( new_n4135_, new_n411_, new_n2178_ );
and  ( new_n4136_, new_n4135_, new_n4134_ );
xor  ( new_n4137_, new_n4136_, new_n328_ );
not  ( new_n4138_, new_n4137_ );
and  ( new_n4139_, new_n4138_, new_n4133_ );
or   ( new_n4140_, new_n4139_, new_n4132_ );
and  ( new_n4141_, new_n4140_, new_n4123_ );
or   ( new_n4142_, new_n4141_, new_n4122_ );
and  ( new_n4143_, new_n4142_, new_n4089_ );
or   ( new_n4144_, new_n4143_, new_n4088_ );
xnor ( new_n4145_, new_n3869_, new_n3853_ );
xor  ( new_n4146_, new_n4145_, new_n3887_ );
xnor ( new_n4147_, new_n3925_, new_n3909_ );
xor  ( new_n4148_, new_n4147_, new_n3943_ );
or   ( new_n4149_, new_n4148_, new_n4146_ );
and  ( new_n4150_, new_n4148_, new_n4146_ );
xor  ( new_n4151_, new_n3832_, new_n3830_ );
xor  ( new_n4152_, new_n4151_, new_n3834_ );
or   ( new_n4153_, new_n4152_, new_n4150_ );
and  ( new_n4154_, new_n4153_, new_n4149_ );
and  ( new_n4155_, new_n4154_, new_n4144_ );
nor  ( new_n4156_, new_n4154_, new_n4144_ );
xor  ( new_n4157_, new_n3957_, new_n3955_ );
xor  ( new_n4158_, new_n4157_, new_n3961_ );
xnor ( new_n4159_, new_n3861_, new_n3857_ );
xor  ( new_n4160_, new_n4159_, new_n3867_ );
xnor ( new_n4161_, new_n3845_, new_n3841_ );
xor  ( new_n4162_, new_n4161_, new_n3851_ );
or   ( new_n4163_, new_n4162_, new_n4160_ );
and  ( new_n4164_, new_n4162_, new_n4160_ );
xor  ( new_n4165_, new_n3935_, new_n3931_ );
xnor ( new_n4166_, new_n4165_, new_n3941_ );
or   ( new_n4167_, new_n4166_, new_n4164_ );
and  ( new_n4168_, new_n4167_, new_n4163_ );
nor  ( new_n4169_, new_n4168_, new_n4158_ );
and  ( new_n4170_, new_n4168_, new_n4158_ );
xor  ( new_n4171_, new_n3952_, new_n3950_ );
not  ( new_n4172_, new_n4171_ );
nor  ( new_n4173_, new_n4172_, new_n4170_ );
nor  ( new_n4174_, new_n4173_, new_n4169_ );
not  ( new_n4175_, new_n4174_ );
nor  ( new_n4176_, new_n4175_, new_n4156_ );
nor  ( new_n4177_, new_n4176_, new_n4155_ );
xor  ( new_n4178_, new_n3626_, new_n3616_ );
xor  ( new_n4179_, new_n4178_, new_n3639_ );
and  ( new_n4180_, new_n4179_, new_n4177_ );
xnor ( new_n4181_, new_n3743_, new_n3726_ );
xor  ( new_n4182_, new_n4181_, new_n3761_ );
xor  ( new_n4183_, new_n3963_, new_n3953_ );
xor  ( new_n4184_, new_n4183_, new_n3967_ );
nor  ( new_n4185_, new_n4184_, new_n4182_ );
and  ( new_n4186_, new_n4184_, new_n4182_ );
xor  ( new_n4187_, new_n3975_, new_n3973_ );
xor  ( new_n4188_, new_n4187_, new_n3980_ );
nor  ( new_n4189_, new_n4188_, new_n4186_ );
nor  ( new_n4190_, new_n4189_, new_n4185_ );
not  ( new_n4191_, new_n4177_ );
not  ( new_n4192_, new_n4179_ );
and  ( new_n4193_, new_n4192_, new_n4191_ );
nor  ( new_n4194_, new_n4193_, new_n4190_ );
nor  ( new_n4195_, new_n4194_, new_n4180_ );
not  ( new_n4196_, new_n4195_ );
and  ( new_n4197_, new_n4196_, new_n4011_ );
not  ( new_n4198_, new_n4197_ );
and  ( new_n4199_, new_n4195_, new_n4010_ );
xnor ( new_n4200_, new_n3763_, new_n3693_ );
xor  ( new_n4201_, new_n4200_, new_n3710_ );
xor  ( new_n4202_, new_n3969_, new_n3948_ );
xor  ( new_n4203_, new_n4202_, new_n3982_ );
nor  ( new_n4204_, new_n4203_, new_n4201_ );
and  ( new_n4205_, new_n4203_, new_n4201_ );
xor  ( new_n4206_, new_n3990_, new_n3988_ );
xor  ( new_n4207_, new_n4206_, new_n3995_ );
nor  ( new_n4208_, new_n4207_, new_n4205_ );
nor  ( new_n4209_, new_n4208_, new_n4204_ );
nor  ( new_n4210_, new_n4209_, new_n4199_ );
not  ( new_n4211_, new_n4210_ );
and  ( new_n4212_, new_n4211_, new_n4198_ );
xnor ( new_n4213_, new_n3999_, new_n3813_ );
xnor ( new_n4214_, new_n4213_, new_n4003_ );
nor  ( new_n4215_, new_n4214_, new_n4212_ );
xor  ( new_n4216_, new_n4005_, new_n3808_ );
and  ( new_n4217_, new_n4216_, new_n4215_ );
xnor ( new_n4218_, new_n4214_, new_n4212_ );
xor  ( new_n4219_, new_n4154_, new_n4144_ );
xor  ( new_n4220_, new_n4219_, new_n4174_ );
not  ( new_n4221_, new_n4220_ );
xnor ( new_n4222_, new_n4184_, new_n4182_ );
xor  ( new_n4223_, new_n4222_, new_n4188_ );
and  ( new_n4224_, new_n4223_, new_n4221_ );
xnor ( new_n4225_, new_n4203_, new_n4201_ );
xor  ( new_n4226_, new_n4225_, new_n4207_ );
or   ( new_n4227_, new_n4226_, new_n4224_ );
and  ( new_n4228_, new_n4226_, new_n4224_ );
xnor ( new_n4229_, new_n3917_, new_n3913_ );
xor  ( new_n4230_, new_n4229_, new_n3923_ );
xnor ( new_n4231_, new_n4036_, new_n4031_ );
xor  ( new_n4232_, new_n4231_, new_n4042_ );
xnor ( new_n4233_, new_n4019_, new_n4015_ );
xor  ( new_n4234_, new_n4233_, new_n4025_ );
or   ( new_n4235_, new_n4234_, new_n4232_ );
and  ( new_n4236_, new_n4234_, new_n4232_ );
xnor ( new_n4237_, new_n4054_, new_n4050_ );
xor  ( new_n4238_, new_n4237_, new_n4060_ );
or   ( new_n4239_, new_n4238_, new_n4236_ );
and  ( new_n4240_, new_n4239_, new_n4235_ );
nor  ( new_n4241_, new_n4240_, new_n4230_ );
and  ( new_n4242_, new_n4240_, new_n4230_ );
xnor ( new_n4243_, new_n4113_, new_n4109_ );
xor  ( new_n4244_, new_n4243_, new_n4119_ );
xnor ( new_n4245_, new_n4097_, new_n4093_ );
xor  ( new_n4246_, new_n4245_, new_n4103_ );
nor  ( new_n4247_, new_n4246_, new_n4244_ );
and  ( new_n4248_, new_n4246_, new_n4244_ );
xor  ( new_n4249_, new_n4131_, new_n4127_ );
xor  ( new_n4250_, new_n4249_, new_n4138_ );
nor  ( new_n4251_, new_n4250_, new_n4248_ );
nor  ( new_n4252_, new_n4251_, new_n4247_ );
nor  ( new_n4253_, new_n4252_, new_n4242_ );
or   ( new_n4254_, new_n4253_, new_n4241_ );
xor  ( new_n4255_, new_n4073_, new_n4068_ );
xor  ( new_n4256_, new_n4255_, new_n4076_ );
not  ( new_n4257_, new_n4256_ );
or   ( new_n4258_, new_n283_, new_n3696_ );
or   ( new_n4259_, new_n286_, new_n3306_ );
and  ( new_n4260_, new_n4259_, new_n4258_ );
xor  ( new_n4261_, new_n4260_, new_n278_ );
or   ( new_n4262_, new_n299_, new_n3820_ );
or   ( new_n4263_, new_n302_, new_n3694_ );
and  ( new_n4264_, new_n4263_, new_n4262_ );
xor  ( new_n4265_, new_n4264_, new_n293_ );
or   ( new_n4266_, new_n4265_, new_n4261_ );
not  ( new_n4267_, RIbb2c5c8_104 );
or   ( new_n4268_, new_n268_, new_n4267_ );
or   ( new_n4269_, new_n271_, new_n4069_ );
and  ( new_n4270_, new_n4269_, new_n4268_ );
xor  ( new_n4271_, new_n4270_, new_n263_ );
and  ( new_n4272_, new_n4265_, new_n4261_ );
or   ( new_n4273_, new_n4272_, new_n4271_ );
and  ( new_n4274_, new_n4273_, new_n4266_ );
or   ( new_n4275_, new_n4274_, new_n4257_ );
or   ( new_n4276_, new_n2425_, new_n419_ );
or   ( new_n4277_, new_n2427_, new_n348_ );
and  ( new_n4278_, new_n4277_, new_n4276_ );
xor  ( new_n4279_, new_n4278_, new_n2121_ );
or   ( new_n4280_, new_n2122_, new_n509_ );
or   ( new_n4281_, new_n2124_, new_n443_ );
and  ( new_n4282_, new_n4281_, new_n4280_ );
xor  ( new_n4283_, new_n4282_, new_n1843_ );
nor  ( new_n4284_, new_n4283_, new_n4279_ );
or   ( new_n4285_, new_n1844_, new_n775_ );
or   ( new_n4286_, new_n1846_, new_n515_ );
and  ( new_n4287_, new_n4286_, new_n4285_ );
xor  ( new_n4288_, new_n4287_, new_n1585_ );
nand ( new_n4289_, new_n4283_, new_n4279_ );
and  ( new_n4290_, new_n4289_, new_n4288_ );
or   ( new_n4291_, new_n4290_, new_n4284_ );
not  ( new_n4292_, RIbb2e350_41 );
and  ( new_n4293_, RIbb2e260_43, RIbb2e2d8_42 );
nor  ( new_n4294_, new_n4293_, new_n4292_ );
not  ( new_n4295_, new_n4294_ );
or   ( new_n4296_, new_n3896_, new_n313_ );
or   ( new_n4297_, new_n3898_, new_n319_ );
and  ( new_n4298_, new_n4297_, new_n4296_ );
xor  ( new_n4299_, new_n4298_, new_n3460_ );
nand ( new_n4300_, new_n4299_, new_n4295_ );
nor  ( new_n4301_, new_n4299_, new_n4295_ );
not  ( new_n4302_, new_n4034_ );
or   ( new_n4303_, new_n4302_, new_n333_ );
not  ( new_n4304_, new_n4032_ );
or   ( new_n4305_, new_n4304_, new_n339_ );
and  ( new_n4306_, new_n4305_, new_n4303_ );
xor  ( new_n4307_, new_n4306_, new_n3894_ );
or   ( new_n4308_, new_n4307_, new_n4301_ );
and  ( new_n4309_, new_n4308_, new_n4300_ );
nand ( new_n4310_, new_n4309_, new_n4291_ );
nor  ( new_n4311_, new_n4309_, new_n4291_ );
or   ( new_n4312_, new_n3461_, new_n279_ );
or   ( new_n4313_, new_n3463_, new_n285_ );
and  ( new_n4314_, new_n4313_, new_n4312_ );
xor  ( new_n4315_, new_n4314_, new_n3116_ );
or   ( new_n4316_, new_n3117_, new_n294_ );
or   ( new_n4317_, new_n3119_, new_n301_ );
and  ( new_n4318_, new_n4317_, new_n4316_ );
xor  ( new_n4319_, new_n4318_, new_n2800_ );
or   ( new_n4320_, new_n4319_, new_n4315_ );
or   ( new_n4321_, new_n2807_, new_n264_ );
or   ( new_n4322_, new_n2809_, new_n270_ );
and  ( new_n4323_, new_n4322_, new_n4321_ );
xor  ( new_n4324_, new_n4323_, new_n2424_ );
and  ( new_n4325_, new_n4319_, new_n4315_ );
or   ( new_n4326_, new_n4325_, new_n4324_ );
and  ( new_n4327_, new_n4326_, new_n4320_ );
or   ( new_n4328_, new_n4327_, new_n4311_ );
and  ( new_n4329_, new_n4328_, new_n4310_ );
or   ( new_n4330_, new_n4329_, new_n4275_ );
and  ( new_n4331_, new_n4329_, new_n4275_ );
or   ( new_n4332_, new_n1593_, new_n886_ );
or   ( new_n4333_, new_n1595_, new_n805_ );
and  ( new_n4334_, new_n4333_, new_n4332_ );
xor  ( new_n4335_, new_n4334_, new_n1358_ );
or   ( new_n4336_, new_n1364_, new_n1168_ );
or   ( new_n4337_, new_n1366_, new_n986_ );
and  ( new_n4338_, new_n4337_, new_n4336_ );
xor  ( new_n4339_, new_n4338_, new_n1129_ );
or   ( new_n4340_, new_n4339_, new_n4335_ );
or   ( new_n4341_, new_n1135_, new_n1318_ );
or   ( new_n4342_, new_n1137_, new_n1213_ );
and  ( new_n4343_, new_n4342_, new_n4341_ );
xor  ( new_n4344_, new_n4343_, new_n896_ );
and  ( new_n4345_, new_n4339_, new_n4335_ );
or   ( new_n4346_, new_n4345_, new_n4344_ );
and  ( new_n4347_, new_n4346_, new_n4340_ );
or   ( new_n4348_, new_n409_, new_n2475_ );
or   ( new_n4349_, new_n411_, new_n2291_ );
and  ( new_n4350_, new_n4349_, new_n4348_ );
xor  ( new_n4351_, new_n4350_, new_n328_ );
or   ( new_n4352_, new_n337_, new_n2751_ );
or   ( new_n4353_, new_n340_, new_n2646_ );
and  ( new_n4354_, new_n4353_, new_n4352_ );
xor  ( new_n4355_, new_n4354_, new_n332_ );
or   ( new_n4356_, new_n4355_, new_n4351_ );
or   ( new_n4357_, new_n317_, new_n3178_ );
or   ( new_n4358_, new_n320_, new_n2981_ );
and  ( new_n4359_, new_n4358_, new_n4357_ );
xor  ( new_n4360_, new_n4359_, new_n312_ );
and  ( new_n4361_, new_n4355_, new_n4351_ );
or   ( new_n4362_, new_n4361_, new_n4360_ );
and  ( new_n4363_, new_n4362_, new_n4356_ );
nor  ( new_n4364_, new_n4363_, new_n4347_ );
and  ( new_n4365_, new_n4363_, new_n4347_ );
or   ( new_n4366_, new_n897_, new_n1523_ );
or   ( new_n4367_, new_n899_, new_n1525_ );
and  ( new_n4368_, new_n4367_, new_n4366_ );
xor  ( new_n4369_, new_n4368_, new_n748_ );
or   ( new_n4370_, new_n755_, new_n1899_ );
or   ( new_n4371_, new_n757_, new_n1754_ );
and  ( new_n4372_, new_n4371_, new_n4370_ );
xor  ( new_n4373_, new_n4372_, new_n523_ );
nor  ( new_n4374_, new_n4373_, new_n4369_ );
or   ( new_n4375_, new_n524_, new_n2178_ );
or   ( new_n4376_, new_n526_, new_n2057_ );
and  ( new_n4377_, new_n4376_, new_n4375_ );
xor  ( new_n4378_, new_n4377_, new_n403_ );
and  ( new_n4379_, new_n4373_, new_n4369_ );
nor  ( new_n4380_, new_n4379_, new_n4378_ );
nor  ( new_n4381_, new_n4380_, new_n4374_ );
nor  ( new_n4382_, new_n4381_, new_n4365_ );
nor  ( new_n4383_, new_n4382_, new_n4364_ );
or   ( new_n4384_, new_n4383_, new_n4331_ );
and  ( new_n4385_, new_n4384_, new_n4330_ );
nor  ( new_n4386_, new_n4385_, new_n4254_ );
nand ( new_n4387_, new_n4385_, new_n4254_ );
xor  ( new_n4388_, new_n3901_, new_n3895_ );
xor  ( new_n4389_, new_n4388_, new_n3907_ );
xnor ( new_n4390_, new_n4162_, new_n4160_ );
xor  ( new_n4391_, new_n4390_, new_n4166_ );
nor  ( new_n4392_, new_n4391_, new_n4389_ );
nand ( new_n4393_, new_n4391_, new_n4389_ );
xor  ( new_n4394_, new_n4081_, new_n4079_ );
xor  ( new_n4395_, new_n4394_, new_n4085_ );
and  ( new_n4396_, new_n4395_, new_n4393_ );
or   ( new_n4397_, new_n4396_, new_n4392_ );
and  ( new_n4398_, new_n4397_, new_n4387_ );
or   ( new_n4399_, new_n4398_, new_n4386_ );
xor  ( new_n4400_, new_n4148_, new_n4146_ );
xor  ( new_n4401_, new_n4400_, new_n4152_ );
xor  ( new_n4402_, new_n4087_, new_n4064_ );
xor  ( new_n4403_, new_n4402_, new_n4142_ );
or   ( new_n4404_, new_n4403_, new_n4401_ );
and  ( new_n4405_, new_n4403_, new_n4401_ );
xor  ( new_n4406_, new_n4168_, new_n4158_ );
xor  ( new_n4407_, new_n4406_, new_n4172_ );
or   ( new_n4408_, new_n4407_, new_n4405_ );
and  ( new_n4409_, new_n4408_, new_n4404_ );
and  ( new_n4410_, new_n4409_, new_n4399_ );
nor  ( new_n4411_, new_n4409_, new_n4399_ );
not  ( new_n4412_, new_n4411_ );
xor  ( new_n4413_, new_n3889_, new_n3837_ );
xor  ( new_n4414_, new_n4413_, new_n3946_ );
and  ( new_n4415_, new_n4414_, new_n4412_ );
nor  ( new_n4416_, new_n4415_, new_n4410_ );
or   ( new_n4417_, new_n4416_, new_n4228_ );
and  ( new_n4418_, new_n4417_, new_n4227_ );
xor  ( new_n4419_, new_n4195_, new_n4011_ );
nand ( new_n4420_, new_n4419_, new_n4209_ );
or   ( new_n4421_, new_n4211_, new_n4197_ );
and  ( new_n4422_, new_n4421_, new_n4420_ );
nand ( new_n4423_, new_n4422_, new_n4418_ );
nor  ( new_n4424_, new_n4422_, new_n4418_ );
xor  ( new_n4425_, new_n3984_, new_n3815_ );
xor  ( new_n4426_, new_n4425_, new_n3997_ );
or   ( new_n4427_, new_n4426_, new_n4424_ );
and  ( new_n4428_, new_n4427_, new_n4423_ );
nor  ( new_n4429_, new_n4428_, new_n4218_ );
xor  ( new_n4430_, new_n4422_, new_n4418_ );
xor  ( new_n4431_, new_n4430_, new_n4426_ );
xor  ( new_n4432_, new_n4190_, new_n4192_ );
xor  ( new_n4433_, new_n4432_, new_n4191_ );
xor  ( new_n4434_, new_n4403_, new_n4401_ );
xor  ( new_n4435_, new_n4434_, new_n4407_ );
xnor ( new_n4436_, new_n4044_, new_n4027_ );
xor  ( new_n4437_, new_n4436_, new_n4062_ );
xor  ( new_n4438_, new_n4121_, new_n4105_ );
xor  ( new_n4439_, new_n4438_, new_n4140_ );
or   ( new_n4440_, new_n4439_, new_n4437_ );
and  ( new_n4441_, new_n4439_, new_n4437_ );
xor  ( new_n4442_, new_n4391_, new_n4389_ );
xor  ( new_n4443_, new_n4442_, new_n4395_ );
or   ( new_n4444_, new_n4443_, new_n4441_ );
and  ( new_n4445_, new_n4444_, new_n4440_ );
or   ( new_n4446_, new_n4445_, new_n4435_ );
and  ( new_n4447_, new_n4445_, new_n4435_ );
xor  ( new_n4448_, new_n4234_, new_n4232_ );
xor  ( new_n4449_, new_n4448_, new_n4238_ );
xor  ( new_n4450_, new_n4283_, new_n4279_ );
xor  ( new_n4451_, new_n4450_, new_n4288_ );
xnor ( new_n4452_, new_n4339_, new_n4335_ );
xor  ( new_n4453_, new_n4452_, new_n4344_ );
or   ( new_n4454_, new_n4453_, new_n4451_ );
and  ( new_n4455_, new_n4453_, new_n4451_ );
xor  ( new_n4456_, new_n4319_, new_n4315_ );
xnor ( new_n4457_, new_n4456_, new_n4324_ );
or   ( new_n4458_, new_n4457_, new_n4455_ );
and  ( new_n4459_, new_n4458_, new_n4454_ );
or   ( new_n4460_, new_n4459_, new_n4449_ );
and  ( new_n4461_, new_n4459_, new_n4449_ );
xnor ( new_n4462_, new_n4355_, new_n4351_ );
xor  ( new_n4463_, new_n4462_, new_n4360_ );
xnor ( new_n4464_, new_n4373_, new_n4369_ );
xor  ( new_n4465_, new_n4464_, new_n4378_ );
nor  ( new_n4466_, new_n4465_, new_n4463_ );
and  ( new_n4467_, new_n4465_, new_n4463_ );
xor  ( new_n4468_, new_n4265_, new_n4261_ );
xnor ( new_n4469_, new_n4468_, new_n4271_ );
nor  ( new_n4470_, new_n4469_, new_n4467_ );
nor  ( new_n4471_, new_n4470_, new_n4466_ );
or   ( new_n4472_, new_n4471_, new_n4461_ );
and  ( new_n4473_, new_n4472_, new_n4460_ );
xor  ( new_n4474_, new_n4363_, new_n4347_ );
xor  ( new_n4475_, new_n4474_, new_n4381_ );
xnor ( new_n4476_, new_n4246_, new_n4244_ );
xor  ( new_n4477_, new_n4476_, new_n4250_ );
nand ( new_n4478_, new_n4477_, new_n4475_ );
nor  ( new_n4479_, new_n4477_, new_n4475_ );
xor  ( new_n4480_, new_n4274_, new_n4257_ );
or   ( new_n4481_, new_n4480_, new_n4479_ );
and  ( new_n4482_, new_n4481_, new_n4478_ );
and  ( new_n4483_, new_n4482_, new_n4473_ );
or   ( new_n4484_, new_n4482_, new_n4473_ );
or   ( new_n4485_, new_n897_, new_n1754_ );
or   ( new_n4486_, new_n899_, new_n1523_ );
and  ( new_n4487_, new_n4486_, new_n4485_ );
xor  ( new_n4488_, new_n4487_, new_n748_ );
or   ( new_n4489_, new_n755_, new_n2057_ );
or   ( new_n4490_, new_n757_, new_n1899_ );
and  ( new_n4491_, new_n4490_, new_n4489_ );
xor  ( new_n4492_, new_n4491_, new_n523_ );
or   ( new_n4493_, new_n4492_, new_n4488_ );
and  ( new_n4494_, new_n4492_, new_n4488_ );
or   ( new_n4495_, new_n524_, new_n2291_ );
or   ( new_n4496_, new_n526_, new_n2178_ );
and  ( new_n4497_, new_n4496_, new_n4495_ );
xor  ( new_n4498_, new_n4497_, new_n403_ );
or   ( new_n4499_, new_n4498_, new_n4494_ );
and  ( new_n4500_, new_n4499_, new_n4493_ );
or   ( new_n4501_, new_n409_, new_n2646_ );
or   ( new_n4502_, new_n411_, new_n2475_ );
and  ( new_n4503_, new_n4502_, new_n4501_ );
xor  ( new_n4504_, new_n4503_, new_n328_ );
or   ( new_n4505_, new_n337_, new_n2981_ );
or   ( new_n4506_, new_n340_, new_n2751_ );
and  ( new_n4507_, new_n4506_, new_n4505_ );
xor  ( new_n4508_, new_n4507_, new_n332_ );
or   ( new_n4509_, new_n4508_, new_n4504_ );
and  ( new_n4510_, new_n4508_, new_n4504_ );
or   ( new_n4511_, new_n317_, new_n3306_ );
or   ( new_n4512_, new_n320_, new_n3178_ );
and  ( new_n4513_, new_n4512_, new_n4511_ );
xor  ( new_n4514_, new_n4513_, new_n312_ );
or   ( new_n4515_, new_n4514_, new_n4510_ );
and  ( new_n4516_, new_n4515_, new_n4509_ );
or   ( new_n4517_, new_n4516_, new_n4500_ );
and  ( new_n4518_, new_n4516_, new_n4500_ );
or   ( new_n4519_, new_n1593_, new_n986_ );
or   ( new_n4520_, new_n1595_, new_n886_ );
and  ( new_n4521_, new_n4520_, new_n4519_ );
xor  ( new_n4522_, new_n4521_, new_n1358_ );
or   ( new_n4523_, new_n1364_, new_n1213_ );
or   ( new_n4524_, new_n1366_, new_n1168_ );
and  ( new_n4525_, new_n4524_, new_n4523_ );
xor  ( new_n4526_, new_n4525_, new_n1129_ );
nor  ( new_n4527_, new_n4526_, new_n4522_ );
and  ( new_n4528_, new_n4526_, new_n4522_ );
or   ( new_n4529_, new_n1135_, new_n1525_ );
or   ( new_n4530_, new_n1137_, new_n1318_ );
and  ( new_n4531_, new_n4530_, new_n4529_ );
xor  ( new_n4532_, new_n4531_, new_n896_ );
nor  ( new_n4533_, new_n4532_, new_n4528_ );
nor  ( new_n4534_, new_n4533_, new_n4527_ );
or   ( new_n4535_, new_n4534_, new_n4518_ );
and  ( new_n4536_, new_n4535_, new_n4517_ );
or   ( new_n4537_, new_n4302_, new_n319_ );
or   ( new_n4538_, new_n4304_, new_n333_ );
and  ( new_n4539_, new_n4538_, new_n4537_ );
xor  ( new_n4540_, new_n4539_, new_n3894_ );
xor  ( new_n4541_, RIbb2e260_43, RIbb2e2d8_42 );
xor  ( new_n4542_, RIbb2e2d8_42, new_n4292_ );
nor  ( new_n4543_, new_n4542_, new_n4541_ );
and  ( new_n4544_, new_n4543_, RIbb2d810_65 );
xor  ( new_n4545_, new_n4544_, new_n4295_ );
nand ( new_n4546_, new_n4545_, new_n4540_ );
nor  ( new_n4547_, new_n4545_, new_n4540_ );
or   ( new_n4548_, new_n3896_, new_n285_ );
or   ( new_n4549_, new_n3898_, new_n313_ );
and  ( new_n4550_, new_n4549_, new_n4548_ );
xor  ( new_n4551_, new_n4550_, new_n3460_ );
or   ( new_n4552_, new_n4551_, new_n4547_ );
and  ( new_n4553_, new_n4552_, new_n4546_ );
or   ( new_n4554_, new_n2425_, new_n443_ );
or   ( new_n4555_, new_n2427_, new_n419_ );
and  ( new_n4556_, new_n4555_, new_n4554_ );
xor  ( new_n4557_, new_n4556_, new_n2121_ );
or   ( new_n4558_, new_n2122_, new_n515_ );
or   ( new_n4559_, new_n2124_, new_n509_ );
and  ( new_n4560_, new_n4559_, new_n4558_ );
xor  ( new_n4561_, new_n4560_, new_n1843_ );
or   ( new_n4562_, new_n4561_, new_n4557_ );
and  ( new_n4563_, new_n4561_, new_n4557_ );
or   ( new_n4564_, new_n1844_, new_n805_ );
or   ( new_n4565_, new_n1846_, new_n775_ );
and  ( new_n4566_, new_n4565_, new_n4564_ );
xor  ( new_n4567_, new_n4566_, new_n1586_ );
or   ( new_n4568_, new_n4567_, new_n4563_ );
and  ( new_n4569_, new_n4568_, new_n4562_ );
or   ( new_n4570_, new_n4569_, new_n4553_ );
and  ( new_n4571_, new_n4569_, new_n4553_ );
or   ( new_n4572_, new_n3461_, new_n301_ );
or   ( new_n4573_, new_n3463_, new_n279_ );
and  ( new_n4574_, new_n4573_, new_n4572_ );
xor  ( new_n4575_, new_n4574_, new_n3116_ );
or   ( new_n4576_, new_n3117_, new_n270_ );
or   ( new_n4577_, new_n3119_, new_n294_ );
and  ( new_n4578_, new_n4577_, new_n4576_ );
xor  ( new_n4579_, new_n4578_, new_n2800_ );
nor  ( new_n4580_, new_n4579_, new_n4575_ );
and  ( new_n4581_, new_n4579_, new_n4575_ );
or   ( new_n4582_, new_n2807_, new_n348_ );
or   ( new_n4583_, new_n2809_, new_n264_ );
and  ( new_n4584_, new_n4583_, new_n4582_ );
xor  ( new_n4585_, new_n4584_, new_n2424_ );
nor  ( new_n4586_, new_n4585_, new_n4581_ );
nor  ( new_n4587_, new_n4586_, new_n4580_ );
or   ( new_n4588_, new_n4587_, new_n4571_ );
and  ( new_n4589_, new_n4588_, new_n4570_ );
nor  ( new_n4590_, new_n4589_, new_n4536_ );
nand ( new_n4591_, new_n4589_, new_n4536_ );
and  ( new_n4592_, RIbb2c4d8_106, RIbb2f610_1 );
or   ( new_n4593_, new_n283_, new_n3694_ );
or   ( new_n4594_, new_n286_, new_n3696_ );
and  ( new_n4595_, new_n4594_, new_n4593_ );
xor  ( new_n4596_, new_n4595_, new_n278_ );
or   ( new_n4597_, new_n299_, new_n4069_ );
or   ( new_n4598_, new_n302_, new_n3820_ );
and  ( new_n4599_, new_n4598_, new_n4597_ );
xor  ( new_n4600_, new_n4599_, new_n293_ );
or   ( new_n4601_, new_n4600_, new_n4596_ );
and  ( new_n4602_, new_n4600_, new_n4596_ );
not  ( new_n4603_, RIbb2c550_105 );
or   ( new_n4604_, new_n268_, new_n4603_ );
or   ( new_n4605_, new_n271_, new_n4267_ );
and  ( new_n4606_, new_n4605_, new_n4604_ );
xor  ( new_n4607_, new_n4606_, new_n263_ );
or   ( new_n4608_, new_n4607_, new_n4602_ );
and  ( new_n4609_, new_n4608_, new_n4601_ );
nor  ( new_n4610_, new_n4609_, new_n4592_ );
and  ( new_n4611_, new_n4609_, new_n4592_ );
and  ( new_n4612_, RIbb2c550_105, RIbb2f610_1 );
nor  ( new_n4613_, new_n4612_, new_n4611_ );
or   ( new_n4614_, new_n4613_, new_n4610_ );
and  ( new_n4615_, new_n4614_, new_n4591_ );
or   ( new_n4616_, new_n4615_, new_n4590_ );
and  ( new_n4617_, new_n4616_, new_n4484_ );
or   ( new_n4618_, new_n4617_, new_n4483_ );
or   ( new_n4619_, new_n4618_, new_n4447_ );
and  ( new_n4620_, new_n4619_, new_n4446_ );
xor  ( new_n4621_, new_n4409_, new_n4399_ );
xor  ( new_n4622_, new_n4621_, new_n4414_ );
or   ( new_n4623_, new_n4622_, new_n4620_ );
nand ( new_n4624_, new_n4622_, new_n4620_ );
xor  ( new_n4625_, new_n4223_, new_n4221_ );
nand ( new_n4626_, new_n4625_, new_n4624_ );
and  ( new_n4627_, new_n4626_, new_n4623_ );
or   ( new_n4628_, new_n4627_, new_n4433_ );
and  ( new_n4629_, new_n4627_, new_n4433_ );
xor  ( new_n4630_, new_n4226_, new_n4224_ );
xnor ( new_n4631_, new_n4630_, new_n4416_ );
or   ( new_n4632_, new_n4631_, new_n4629_ );
and  ( new_n4633_, new_n4632_, new_n4628_ );
nor  ( new_n4634_, new_n4633_, new_n4431_ );
xnor ( new_n4635_, new_n4627_, new_n4433_ );
xor  ( new_n4636_, new_n4635_, new_n4631_ );
or   ( new_n4637_, new_n524_, new_n2475_ );
or   ( new_n4638_, new_n526_, new_n2291_ );
and  ( new_n4639_, new_n4638_, new_n4637_ );
xor  ( new_n4640_, new_n4639_, new_n403_ );
or   ( new_n4641_, new_n409_, new_n2751_ );
or   ( new_n4642_, new_n411_, new_n2646_ );
and  ( new_n4643_, new_n4642_, new_n4641_ );
xor  ( new_n4644_, new_n4643_, new_n328_ );
or   ( new_n4645_, new_n4644_, new_n4640_ );
and  ( new_n4646_, new_n4644_, new_n4640_ );
or   ( new_n4647_, new_n337_, new_n3178_ );
or   ( new_n4648_, new_n340_, new_n2981_ );
and  ( new_n4649_, new_n4648_, new_n4647_ );
xor  ( new_n4650_, new_n4649_, new_n332_ );
or   ( new_n4651_, new_n4650_, new_n4646_ );
and  ( new_n4652_, new_n4651_, new_n4645_ );
or   ( new_n4653_, new_n1844_, new_n886_ );
or   ( new_n4654_, new_n1846_, new_n805_ );
and  ( new_n4655_, new_n4654_, new_n4653_ );
xor  ( new_n4656_, new_n4655_, new_n1586_ );
or   ( new_n4657_, new_n1593_, new_n1168_ );
or   ( new_n4658_, new_n1595_, new_n986_ );
and  ( new_n4659_, new_n4658_, new_n4657_ );
xor  ( new_n4660_, new_n4659_, new_n1358_ );
or   ( new_n4661_, new_n4660_, new_n4656_ );
and  ( new_n4662_, new_n4660_, new_n4656_ );
or   ( new_n4663_, new_n1364_, new_n1318_ );
or   ( new_n4664_, new_n1366_, new_n1213_ );
and  ( new_n4665_, new_n4664_, new_n4663_ );
xor  ( new_n4666_, new_n4665_, new_n1129_ );
or   ( new_n4667_, new_n4666_, new_n4662_ );
and  ( new_n4668_, new_n4667_, new_n4661_ );
or   ( new_n4669_, new_n4668_, new_n4652_ );
and  ( new_n4670_, new_n4668_, new_n4652_ );
or   ( new_n4671_, new_n1135_, new_n1523_ );
or   ( new_n4672_, new_n1137_, new_n1525_ );
and  ( new_n4673_, new_n4672_, new_n4671_ );
xor  ( new_n4674_, new_n4673_, new_n896_ );
or   ( new_n4675_, new_n897_, new_n1899_ );
or   ( new_n4676_, new_n899_, new_n1754_ );
and  ( new_n4677_, new_n4676_, new_n4675_ );
xor  ( new_n4678_, new_n4677_, new_n748_ );
or   ( new_n4679_, new_n4678_, new_n4674_ );
and  ( new_n4680_, new_n4678_, new_n4674_ );
or   ( new_n4681_, new_n755_, new_n2178_ );
or   ( new_n4682_, new_n757_, new_n2057_ );
and  ( new_n4683_, new_n4682_, new_n4681_ );
xor  ( new_n4684_, new_n4683_, new_n523_ );
or   ( new_n4685_, new_n4684_, new_n4680_ );
and  ( new_n4686_, new_n4685_, new_n4679_ );
or   ( new_n4687_, new_n4686_, new_n4670_ );
and  ( new_n4688_, new_n4687_, new_n4669_ );
or   ( new_n4689_, new_n2807_, new_n419_ );
or   ( new_n4690_, new_n2809_, new_n348_ );
and  ( new_n4691_, new_n4690_, new_n4689_ );
xor  ( new_n4692_, new_n4691_, new_n2424_ );
or   ( new_n4693_, new_n2425_, new_n509_ );
or   ( new_n4694_, new_n2427_, new_n443_ );
and  ( new_n4695_, new_n4694_, new_n4693_ );
xor  ( new_n4696_, new_n4695_, new_n2121_ );
nor  ( new_n4697_, new_n4696_, new_n4692_ );
nand ( new_n4698_, new_n4696_, new_n4692_ );
or   ( new_n4699_, new_n2122_, new_n775_ );
or   ( new_n4700_, new_n2124_, new_n515_ );
and  ( new_n4701_, new_n4700_, new_n4699_ );
xor  ( new_n4702_, new_n4701_, new_n1842_ );
and  ( new_n4703_, new_n4702_, new_n4698_ );
or   ( new_n4704_, new_n4703_, new_n4697_ );
not  ( new_n4705_, RIbb2e260_43 );
and  ( new_n4706_, RIbb2e170_45, RIbb2e1e8_44 );
nor  ( new_n4707_, new_n4706_, new_n4705_ );
not  ( new_n4708_, new_n4707_ );
not  ( new_n4709_, new_n4543_ );
or   ( new_n4710_, new_n4709_, new_n333_ );
not  ( new_n4711_, new_n4541_ );
or   ( new_n4712_, new_n4711_, new_n339_ );
and  ( new_n4713_, new_n4712_, new_n4710_ );
xor  ( new_n4714_, new_n4713_, new_n4295_ );
nand ( new_n4715_, new_n4714_, new_n4708_ );
nor  ( new_n4716_, new_n4714_, new_n4708_ );
or   ( new_n4717_, new_n4302_, new_n313_ );
or   ( new_n4718_, new_n4304_, new_n319_ );
and  ( new_n4719_, new_n4718_, new_n4717_ );
xor  ( new_n4720_, new_n4719_, new_n3894_ );
or   ( new_n4721_, new_n4720_, new_n4716_ );
and  ( new_n4722_, new_n4721_, new_n4715_ );
nand ( new_n4723_, new_n4722_, new_n4704_ );
nor  ( new_n4724_, new_n4722_, new_n4704_ );
or   ( new_n4725_, new_n3896_, new_n279_ );
or   ( new_n4726_, new_n3898_, new_n285_ );
and  ( new_n4727_, new_n4726_, new_n4725_ );
xor  ( new_n4728_, new_n4727_, new_n3460_ );
or   ( new_n4729_, new_n3461_, new_n294_ );
or   ( new_n4730_, new_n3463_, new_n301_ );
and  ( new_n4731_, new_n4730_, new_n4729_ );
xor  ( new_n4732_, new_n4731_, new_n3116_ );
nor  ( new_n4733_, new_n4732_, new_n4728_ );
and  ( new_n4734_, new_n4732_, new_n4728_ );
or   ( new_n4735_, new_n3117_, new_n264_ );
or   ( new_n4736_, new_n3119_, new_n270_ );
and  ( new_n4737_, new_n4736_, new_n4735_ );
xor  ( new_n4738_, new_n4737_, new_n2800_ );
nor  ( new_n4739_, new_n4738_, new_n4734_ );
nor  ( new_n4740_, new_n4739_, new_n4733_ );
or   ( new_n4741_, new_n4740_, new_n4724_ );
and  ( new_n4742_, new_n4741_, new_n4723_ );
nor  ( new_n4743_, new_n4742_, new_n4688_ );
nand ( new_n4744_, new_n4742_, new_n4688_ );
not  ( new_n4745_, new_n4592_ );
or   ( new_n4746_, new_n317_, new_n3696_ );
or   ( new_n4747_, new_n320_, new_n3306_ );
and  ( new_n4748_, new_n4747_, new_n4746_ );
xor  ( new_n4749_, new_n4748_, new_n312_ );
or   ( new_n4750_, new_n283_, new_n3820_ );
or   ( new_n4751_, new_n286_, new_n3694_ );
and  ( new_n4752_, new_n4751_, new_n4750_ );
xor  ( new_n4753_, new_n4752_, new_n278_ );
or   ( new_n4754_, new_n4753_, new_n4749_ );
and  ( new_n4755_, new_n4753_, new_n4749_ );
or   ( new_n4756_, new_n299_, new_n4267_ );
or   ( new_n4757_, new_n302_, new_n4069_ );
and  ( new_n4758_, new_n4757_, new_n4756_ );
xor  ( new_n4759_, new_n4758_, new_n293_ );
or   ( new_n4760_, new_n4759_, new_n4755_ );
and  ( new_n4761_, new_n4760_, new_n4754_ );
nor  ( new_n4762_, new_n4761_, new_n4745_ );
nand ( new_n4763_, new_n4761_, new_n4745_ );
xor  ( new_n4764_, new_n4600_, new_n4596_ );
xnor ( new_n4765_, new_n4764_, new_n4607_ );
and  ( new_n4766_, new_n4765_, new_n4763_ );
or   ( new_n4767_, new_n4766_, new_n4762_ );
and  ( new_n4768_, new_n4767_, new_n4744_ );
or   ( new_n4769_, new_n4768_, new_n4743_ );
xor  ( new_n4770_, new_n4299_, new_n4295_ );
xor  ( new_n4771_, new_n4770_, new_n4307_ );
xnor ( new_n4772_, new_n4508_, new_n4504_ );
xor  ( new_n4773_, new_n4772_, new_n4514_ );
xnor ( new_n4774_, new_n4492_, new_n4488_ );
xor  ( new_n4775_, new_n4774_, new_n4498_ );
or   ( new_n4776_, new_n4775_, new_n4773_ );
and  ( new_n4777_, new_n4775_, new_n4773_ );
xor  ( new_n4778_, new_n4526_, new_n4522_ );
xnor ( new_n4779_, new_n4778_, new_n4532_ );
or   ( new_n4780_, new_n4779_, new_n4777_ );
and  ( new_n4781_, new_n4780_, new_n4776_ );
or   ( new_n4782_, new_n4781_, new_n4771_ );
and  ( new_n4783_, new_n4781_, new_n4771_ );
xnor ( new_n4784_, new_n4561_, new_n4557_ );
xor  ( new_n4785_, new_n4784_, new_n4567_ );
xnor ( new_n4786_, new_n4545_, new_n4540_ );
xor  ( new_n4787_, new_n4786_, new_n4551_ );
nor  ( new_n4788_, new_n4787_, new_n4785_ );
and  ( new_n4789_, new_n4787_, new_n4785_ );
xor  ( new_n4790_, new_n4579_, new_n4575_ );
xnor ( new_n4791_, new_n4790_, new_n4585_ );
nor  ( new_n4792_, new_n4791_, new_n4789_ );
nor  ( new_n4793_, new_n4792_, new_n4788_ );
or   ( new_n4794_, new_n4793_, new_n4783_ );
and  ( new_n4795_, new_n4794_, new_n4782_ );
or   ( new_n4796_, new_n4795_, new_n4769_ );
and  ( new_n4797_, new_n4795_, new_n4769_ );
xor  ( new_n4798_, new_n4609_, new_n4592_ );
xor  ( new_n4799_, new_n4798_, new_n4612_ );
xnor ( new_n4800_, new_n4465_, new_n4463_ );
xor  ( new_n4801_, new_n4800_, new_n4469_ );
and  ( new_n4802_, new_n4801_, new_n4799_ );
nor  ( new_n4803_, new_n4801_, new_n4799_ );
xor  ( new_n4804_, new_n4453_, new_n4451_ );
xnor ( new_n4805_, new_n4804_, new_n4457_ );
not  ( new_n4806_, new_n4805_ );
nor  ( new_n4807_, new_n4806_, new_n4803_ );
nor  ( new_n4808_, new_n4807_, new_n4802_ );
or   ( new_n4809_, new_n4808_, new_n4797_ );
and  ( new_n4810_, new_n4809_, new_n4796_ );
xor  ( new_n4811_, new_n4309_, new_n4291_ );
xor  ( new_n4812_, new_n4811_, new_n4327_ );
xnor ( new_n4813_, new_n4459_, new_n4449_ );
xor  ( new_n4814_, new_n4813_, new_n4471_ );
nand ( new_n4815_, new_n4814_, new_n4812_ );
or   ( new_n4816_, new_n4814_, new_n4812_ );
xor  ( new_n4817_, new_n4477_, new_n4475_ );
xnor ( new_n4818_, new_n4817_, new_n4480_ );
nand ( new_n4819_, new_n4818_, new_n4816_ );
and  ( new_n4820_, new_n4819_, new_n4815_ );
and  ( new_n4821_, new_n4820_, new_n4810_ );
or   ( new_n4822_, new_n4820_, new_n4810_ );
xor  ( new_n4823_, new_n4240_, new_n4230_ );
xor  ( new_n4824_, new_n4823_, new_n4252_ );
and  ( new_n4825_, new_n4824_, new_n4822_ );
or   ( new_n4826_, new_n4825_, new_n4821_ );
xor  ( new_n4827_, new_n4482_, new_n4473_ );
xor  ( new_n4828_, new_n4827_, new_n4616_ );
xnor ( new_n4829_, new_n4329_, new_n4275_ );
xor  ( new_n4830_, new_n4829_, new_n4383_ );
or   ( new_n4831_, new_n4830_, new_n4828_ );
and  ( new_n4832_, new_n4830_, new_n4828_ );
xor  ( new_n4833_, new_n4439_, new_n4437_ );
xor  ( new_n4834_, new_n4833_, new_n4443_ );
or   ( new_n4835_, new_n4834_, new_n4832_ );
and  ( new_n4836_, new_n4835_, new_n4831_ );
or   ( new_n4837_, new_n4836_, new_n4826_ );
and  ( new_n4838_, new_n4836_, new_n4826_ );
xor  ( new_n4839_, new_n4385_, new_n4254_ );
xor  ( new_n4840_, new_n4839_, new_n4397_ );
or   ( new_n4841_, new_n4840_, new_n4838_ );
and  ( new_n4842_, new_n4841_, new_n4837_ );
xor  ( new_n4843_, new_n4836_, new_n4826_ );
xor  ( new_n4844_, new_n4843_, new_n4840_ );
xor  ( new_n4845_, new_n4589_, new_n4536_ );
xor  ( new_n4846_, new_n4845_, new_n4614_ );
xnor ( new_n4847_, new_n4569_, new_n4553_ );
xor  ( new_n4848_, new_n4847_, new_n4587_ );
xnor ( new_n4849_, new_n4516_, new_n4500_ );
xor  ( new_n4850_, new_n4849_, new_n4534_ );
or   ( new_n4851_, new_n4850_, new_n4848_ );
and  ( new_n4852_, new_n4850_, new_n4848_ );
xor  ( new_n4853_, new_n4801_, new_n4799_ );
xor  ( new_n4854_, new_n4853_, new_n4806_ );
or   ( new_n4855_, new_n4854_, new_n4852_ );
and  ( new_n4856_, new_n4855_, new_n4851_ );
or   ( new_n4857_, new_n4856_, new_n4846_ );
and  ( new_n4858_, new_n4856_, new_n4846_ );
not  ( new_n4859_, RIbb2c460_107 );
or   ( new_n4860_, new_n4859_, new_n260_ );
xnor ( new_n4861_, new_n4753_, new_n4749_ );
xor  ( new_n4862_, new_n4861_, new_n4759_ );
and  ( new_n4863_, new_n4862_, new_n4860_ );
or   ( new_n4864_, new_n4862_, new_n4860_ );
xnor ( new_n4865_, new_n4644_, new_n4640_ );
xor  ( new_n4866_, new_n4865_, new_n4650_ );
and  ( new_n4867_, new_n4866_, new_n4864_ );
or   ( new_n4868_, new_n4867_, new_n4863_ );
xnor ( new_n4869_, new_n4660_, new_n4656_ );
xor  ( new_n4870_, new_n4869_, new_n4666_ );
xor  ( new_n4871_, new_n4696_, new_n4692_ );
xor  ( new_n4872_, new_n4871_, new_n4702_ );
or   ( new_n4873_, new_n4872_, new_n4870_ );
and  ( new_n4874_, new_n4872_, new_n4870_ );
xor  ( new_n4875_, new_n4678_, new_n4674_ );
xnor ( new_n4876_, new_n4875_, new_n4684_ );
or   ( new_n4877_, new_n4876_, new_n4874_ );
and  ( new_n4878_, new_n4877_, new_n4873_ );
and  ( new_n4879_, new_n4878_, new_n4868_ );
nor  ( new_n4880_, new_n4878_, new_n4868_ );
xor  ( new_n4881_, new_n4787_, new_n4785_ );
xnor ( new_n4882_, new_n4881_, new_n4791_ );
nor  ( new_n4883_, new_n4882_, new_n4880_ );
or   ( new_n4884_, new_n4883_, new_n4879_ );
or   ( new_n4885_, new_n1135_, new_n1754_ );
or   ( new_n4886_, new_n1137_, new_n1523_ );
and  ( new_n4887_, new_n4886_, new_n4885_ );
xor  ( new_n4888_, new_n4887_, new_n896_ );
or   ( new_n4889_, new_n897_, new_n2057_ );
or   ( new_n4890_, new_n899_, new_n1899_ );
and  ( new_n4891_, new_n4890_, new_n4889_ );
xor  ( new_n4892_, new_n4891_, new_n748_ );
or   ( new_n4893_, new_n4892_, new_n4888_ );
and  ( new_n4894_, new_n4892_, new_n4888_ );
or   ( new_n4895_, new_n755_, new_n2291_ );
or   ( new_n4896_, new_n757_, new_n2178_ );
and  ( new_n4897_, new_n4896_, new_n4895_ );
xor  ( new_n4898_, new_n4897_, new_n523_ );
or   ( new_n4899_, new_n4898_, new_n4894_ );
and  ( new_n4900_, new_n4899_, new_n4893_ );
or   ( new_n4901_, new_n1844_, new_n986_ );
or   ( new_n4902_, new_n1846_, new_n886_ );
and  ( new_n4903_, new_n4902_, new_n4901_ );
xor  ( new_n4904_, new_n4903_, new_n1586_ );
or   ( new_n4905_, new_n1593_, new_n1213_ );
or   ( new_n4906_, new_n1595_, new_n1168_ );
and  ( new_n4907_, new_n4906_, new_n4905_ );
xor  ( new_n4908_, new_n4907_, new_n1358_ );
or   ( new_n4909_, new_n4908_, new_n4904_ );
and  ( new_n4910_, new_n4908_, new_n4904_ );
or   ( new_n4911_, new_n1364_, new_n1525_ );
or   ( new_n4912_, new_n1366_, new_n1318_ );
and  ( new_n4913_, new_n4912_, new_n4911_ );
xor  ( new_n4914_, new_n4913_, new_n1129_ );
or   ( new_n4915_, new_n4914_, new_n4910_ );
and  ( new_n4916_, new_n4915_, new_n4909_ );
nor  ( new_n4917_, new_n4916_, new_n4900_ );
nand ( new_n4918_, new_n4916_, new_n4900_ );
or   ( new_n4919_, new_n524_, new_n2646_ );
or   ( new_n4920_, new_n526_, new_n2475_ );
and  ( new_n4921_, new_n4920_, new_n4919_ );
xor  ( new_n4922_, new_n4921_, new_n403_ );
or   ( new_n4923_, new_n409_, new_n2981_ );
or   ( new_n4924_, new_n411_, new_n2751_ );
and  ( new_n4925_, new_n4924_, new_n4923_ );
xor  ( new_n4926_, new_n4925_, new_n328_ );
nor  ( new_n4927_, new_n4926_, new_n4922_ );
and  ( new_n4928_, new_n4926_, new_n4922_ );
or   ( new_n4929_, new_n337_, new_n3306_ );
or   ( new_n4930_, new_n340_, new_n3178_ );
and  ( new_n4931_, new_n4930_, new_n4929_ );
xor  ( new_n4932_, new_n4931_, new_n332_ );
nor  ( new_n4933_, new_n4932_, new_n4928_ );
nor  ( new_n4934_, new_n4933_, new_n4927_ );
not  ( new_n4935_, new_n4934_ );
and  ( new_n4936_, new_n4935_, new_n4918_ );
or   ( new_n4937_, new_n4936_, new_n4917_ );
or   ( new_n4938_, new_n2807_, new_n443_ );
or   ( new_n4939_, new_n2809_, new_n419_ );
and  ( new_n4940_, new_n4939_, new_n4938_ );
xor  ( new_n4941_, new_n4940_, new_n2424_ );
or   ( new_n4942_, new_n2425_, new_n515_ );
or   ( new_n4943_, new_n2427_, new_n509_ );
and  ( new_n4944_, new_n4943_, new_n4942_ );
xor  ( new_n4945_, new_n4944_, new_n2121_ );
or   ( new_n4946_, new_n4945_, new_n4941_ );
and  ( new_n4947_, new_n4945_, new_n4941_ );
or   ( new_n4948_, new_n2122_, new_n805_ );
or   ( new_n4949_, new_n2124_, new_n775_ );
and  ( new_n4950_, new_n4949_, new_n4948_ );
xor  ( new_n4951_, new_n4950_, new_n1843_ );
or   ( new_n4952_, new_n4951_, new_n4947_ );
and  ( new_n4953_, new_n4952_, new_n4946_ );
or   ( new_n4954_, new_n4709_, new_n319_ );
or   ( new_n4955_, new_n4711_, new_n333_ );
and  ( new_n4956_, new_n4955_, new_n4954_ );
xor  ( new_n4957_, new_n4956_, new_n4294_ );
xor  ( new_n4958_, RIbb2e170_45, RIbb2e1e8_44 );
xor  ( new_n4959_, RIbb2e1e8_44, new_n4705_ );
nor  ( new_n4960_, new_n4959_, new_n4958_ );
and  ( new_n4961_, new_n4960_, RIbb2d810_65 );
xor  ( new_n4962_, new_n4961_, new_n4708_ );
nand ( new_n4963_, new_n4962_, new_n4957_ );
nor  ( new_n4964_, new_n4962_, new_n4957_ );
or   ( new_n4965_, new_n4302_, new_n285_ );
or   ( new_n4966_, new_n4304_, new_n313_ );
and  ( new_n4967_, new_n4966_, new_n4965_ );
xor  ( new_n4968_, new_n4967_, new_n3895_ );
or   ( new_n4969_, new_n4968_, new_n4964_ );
and  ( new_n4970_, new_n4969_, new_n4963_ );
nor  ( new_n4971_, new_n4970_, new_n4953_ );
and  ( new_n4972_, new_n4970_, new_n4953_ );
or   ( new_n4973_, new_n3896_, new_n301_ );
or   ( new_n4974_, new_n3898_, new_n279_ );
and  ( new_n4975_, new_n4974_, new_n4973_ );
xor  ( new_n4976_, new_n4975_, new_n3460_ );
or   ( new_n4977_, new_n3461_, new_n270_ );
or   ( new_n4978_, new_n3463_, new_n294_ );
and  ( new_n4979_, new_n4978_, new_n4977_ );
xor  ( new_n4980_, new_n4979_, new_n3116_ );
nor  ( new_n4981_, new_n4980_, new_n4976_ );
and  ( new_n4982_, new_n4980_, new_n4976_ );
or   ( new_n4983_, new_n3117_, new_n348_ );
or   ( new_n4984_, new_n3119_, new_n264_ );
and  ( new_n4985_, new_n4984_, new_n4983_ );
xor  ( new_n4986_, new_n4985_, new_n2800_ );
nor  ( new_n4987_, new_n4986_, new_n4982_ );
nor  ( new_n4988_, new_n4987_, new_n4981_ );
nor  ( new_n4989_, new_n4988_, new_n4972_ );
nor  ( new_n4990_, new_n4989_, new_n4971_ );
not  ( new_n4991_, new_n4990_ );
or   ( new_n4992_, new_n4991_, new_n4937_ );
and  ( new_n4993_, new_n4991_, new_n4937_ );
or   ( new_n4994_, new_n268_, new_n4859_ );
not  ( new_n4995_, RIbb2c4d8_106 );
or   ( new_n4996_, new_n271_, new_n4995_ );
and  ( new_n4997_, new_n4996_, new_n4994_ );
xor  ( new_n4998_, new_n4997_, new_n263_ );
and  ( new_n4999_, RIbb2c3e8_108, RIbb2f610_1 );
or   ( new_n5000_, new_n4999_, new_n4998_ );
or   ( new_n5001_, new_n317_, new_n3694_ );
or   ( new_n5002_, new_n320_, new_n3696_ );
and  ( new_n5003_, new_n5002_, new_n5001_ );
xor  ( new_n5004_, new_n5003_, new_n312_ );
or   ( new_n5005_, new_n283_, new_n4069_ );
or   ( new_n5006_, new_n286_, new_n3820_ );
and  ( new_n5007_, new_n5006_, new_n5005_ );
xor  ( new_n5008_, new_n5007_, new_n278_ );
or   ( new_n5009_, new_n5008_, new_n5004_ );
and  ( new_n5010_, new_n5008_, new_n5004_ );
or   ( new_n5011_, new_n299_, new_n4603_ );
or   ( new_n5012_, new_n302_, new_n4267_ );
and  ( new_n5013_, new_n5012_, new_n5011_ );
xor  ( new_n5014_, new_n5013_, new_n293_ );
or   ( new_n5015_, new_n5014_, new_n5010_ );
and  ( new_n5016_, new_n5015_, new_n5009_ );
and  ( new_n5017_, new_n5016_, new_n5000_ );
nor  ( new_n5018_, new_n5016_, new_n5000_ );
not  ( new_n5019_, new_n5018_ );
or   ( new_n5020_, new_n268_, new_n4995_ );
or   ( new_n5021_, new_n271_, new_n4603_ );
and  ( new_n5022_, new_n5021_, new_n5020_ );
xor  ( new_n5023_, new_n5022_, new_n263_ );
and  ( new_n5024_, new_n5023_, new_n5019_ );
nor  ( new_n5025_, new_n5024_, new_n5017_ );
or   ( new_n5026_, new_n5025_, new_n4993_ );
and  ( new_n5027_, new_n5026_, new_n4992_ );
nor  ( new_n5028_, new_n5027_, new_n4884_ );
and  ( new_n5029_, new_n5027_, new_n4884_ );
xor  ( new_n5030_, new_n4668_, new_n4652_ );
xor  ( new_n5031_, new_n5030_, new_n4686_ );
xnor ( new_n5032_, new_n4775_, new_n4773_ );
xor  ( new_n5033_, new_n5032_, new_n4779_ );
and  ( new_n5034_, new_n5033_, new_n5031_ );
nor  ( new_n5035_, new_n5033_, new_n5031_ );
xor  ( new_n5036_, new_n4761_, new_n4745_ );
xor  ( new_n5037_, new_n5036_, new_n4765_ );
nor  ( new_n5038_, new_n5037_, new_n5035_ );
nor  ( new_n5039_, new_n5038_, new_n5034_ );
nor  ( new_n5040_, new_n5039_, new_n5029_ );
nor  ( new_n5041_, new_n5040_, new_n5028_ );
or   ( new_n5042_, new_n5041_, new_n4858_ );
and  ( new_n5043_, new_n5042_, new_n4857_ );
xor  ( new_n5044_, new_n4820_, new_n4810_ );
xor  ( new_n5045_, new_n5044_, new_n4824_ );
or   ( new_n5046_, new_n5045_, new_n5043_ );
and  ( new_n5047_, new_n5045_, new_n5043_ );
xor  ( new_n5048_, new_n4830_, new_n4828_ );
xor  ( new_n5049_, new_n5048_, new_n4834_ );
or   ( new_n5050_, new_n5049_, new_n5047_ );
and  ( new_n5051_, new_n5050_, new_n5046_ );
or   ( new_n5052_, new_n5051_, new_n4844_ );
and  ( new_n5053_, new_n5051_, new_n4844_ );
xor  ( new_n5054_, new_n4445_, new_n4435_ );
xor  ( new_n5055_, new_n5054_, new_n4618_ );
or   ( new_n5056_, new_n5055_, new_n5053_ );
and  ( new_n5057_, new_n5056_, new_n5052_ );
nand ( new_n5058_, new_n5057_, new_n4842_ );
nor  ( new_n5059_, new_n5057_, new_n4842_ );
xor  ( new_n5060_, new_n4622_, new_n4620_ );
xor  ( new_n5061_, new_n5060_, new_n4625_ );
or   ( new_n5062_, new_n5061_, new_n5059_ );
and  ( new_n5063_, new_n5062_, new_n5058_ );
and  ( new_n5064_, new_n5063_, new_n4636_ );
xor  ( new_n5065_, new_n5051_, new_n4844_ );
xor  ( new_n5066_, new_n5065_, new_n5055_ );
xor  ( new_n5067_, new_n4795_, new_n4769_ );
xnor ( new_n5068_, new_n5067_, new_n4808_ );
xnor ( new_n5069_, new_n4856_, new_n4846_ );
xor  ( new_n5070_, new_n5069_, new_n5041_ );
and  ( new_n5071_, new_n5070_, new_n5068_ );
xor  ( new_n5072_, new_n4814_, new_n4812_ );
xor  ( new_n5073_, new_n5072_, new_n4818_ );
xor  ( new_n5074_, new_n4850_, new_n4848_ );
xor  ( new_n5075_, new_n5074_, new_n4854_ );
xor  ( new_n5076_, new_n4742_, new_n4688_ );
xor  ( new_n5077_, new_n5076_, new_n4767_ );
nand ( new_n5078_, new_n5077_, new_n5075_ );
nor  ( new_n5079_, new_n5077_, new_n5075_ );
xor  ( new_n5080_, new_n5027_, new_n4884_ );
xnor ( new_n5081_, new_n5080_, new_n5039_ );
or   ( new_n5082_, new_n5081_, new_n5079_ );
and  ( new_n5083_, new_n5082_, new_n5078_ );
or   ( new_n5084_, new_n5083_, new_n5073_ );
and  ( new_n5085_, new_n5083_, new_n5073_ );
xnor ( new_n5086_, new_n4781_, new_n4771_ );
xor  ( new_n5087_, new_n5086_, new_n4793_ );
xnor ( new_n5088_, new_n4732_, new_n4728_ );
xor  ( new_n5089_, new_n5088_, new_n4738_ );
xnor ( new_n5090_, new_n4908_, new_n4904_ );
xor  ( new_n5091_, new_n5090_, new_n4914_ );
xnor ( new_n5092_, new_n4945_, new_n4941_ );
xor  ( new_n5093_, new_n5092_, new_n4951_ );
or   ( new_n5094_, new_n5093_, new_n5091_ );
and  ( new_n5095_, new_n5093_, new_n5091_ );
xor  ( new_n5096_, new_n4980_, new_n4976_ );
xnor ( new_n5097_, new_n5096_, new_n4986_ );
or   ( new_n5098_, new_n5097_, new_n5095_ );
and  ( new_n5099_, new_n5098_, new_n5094_ );
nor  ( new_n5100_, new_n5099_, new_n5089_ );
nand ( new_n5101_, new_n5099_, new_n5089_ );
xnor ( new_n5102_, new_n5008_, new_n5004_ );
xor  ( new_n5103_, new_n5102_, new_n5014_ );
xnor ( new_n5104_, new_n4892_, new_n4888_ );
xor  ( new_n5105_, new_n5104_, new_n4898_ );
nor  ( new_n5106_, new_n5105_, new_n5103_ );
nand ( new_n5107_, new_n5105_, new_n5103_ );
xor  ( new_n5108_, new_n4926_, new_n4922_ );
xor  ( new_n5109_, new_n5108_, new_n4932_ );
and  ( new_n5110_, new_n5109_, new_n5107_ );
or   ( new_n5111_, new_n5110_, new_n5106_ );
and  ( new_n5112_, new_n5111_, new_n5101_ );
or   ( new_n5113_, new_n5112_, new_n5100_ );
or   ( new_n5114_, new_n1364_, new_n1523_ );
or   ( new_n5115_, new_n1366_, new_n1525_ );
and  ( new_n5116_, new_n5115_, new_n5114_ );
xor  ( new_n5117_, new_n5116_, new_n1129_ );
or   ( new_n5118_, new_n1135_, new_n1899_ );
or   ( new_n5119_, new_n1137_, new_n1754_ );
and  ( new_n5120_, new_n5119_, new_n5118_ );
xor  ( new_n5121_, new_n5120_, new_n896_ );
or   ( new_n5122_, new_n5121_, new_n5117_ );
and  ( new_n5123_, new_n5121_, new_n5117_ );
or   ( new_n5124_, new_n897_, new_n2178_ );
or   ( new_n5125_, new_n899_, new_n2057_ );
and  ( new_n5126_, new_n5125_, new_n5124_ );
xor  ( new_n5127_, new_n5126_, new_n748_ );
or   ( new_n5128_, new_n5127_, new_n5123_ );
and  ( new_n5129_, new_n5128_, new_n5122_ );
or   ( new_n5130_, new_n2122_, new_n886_ );
or   ( new_n5131_, new_n2124_, new_n805_ );
and  ( new_n5132_, new_n5131_, new_n5130_ );
xor  ( new_n5133_, new_n5132_, new_n1843_ );
or   ( new_n5134_, new_n1844_, new_n1168_ );
or   ( new_n5135_, new_n1846_, new_n986_ );
and  ( new_n5136_, new_n5135_, new_n5134_ );
xor  ( new_n5137_, new_n5136_, new_n1586_ );
or   ( new_n5138_, new_n5137_, new_n5133_ );
and  ( new_n5139_, new_n5137_, new_n5133_ );
or   ( new_n5140_, new_n1593_, new_n1318_ );
or   ( new_n5141_, new_n1595_, new_n1213_ );
and  ( new_n5142_, new_n5141_, new_n5140_ );
xor  ( new_n5143_, new_n5142_, new_n1358_ );
or   ( new_n5144_, new_n5143_, new_n5139_ );
and  ( new_n5145_, new_n5144_, new_n5138_ );
or   ( new_n5146_, new_n5145_, new_n5129_ );
and  ( new_n5147_, new_n5145_, new_n5129_ );
or   ( new_n5148_, new_n755_, new_n2475_ );
or   ( new_n5149_, new_n757_, new_n2291_ );
and  ( new_n5150_, new_n5149_, new_n5148_ );
xor  ( new_n5151_, new_n5150_, new_n523_ );
or   ( new_n5152_, new_n524_, new_n2751_ );
or   ( new_n5153_, new_n526_, new_n2646_ );
and  ( new_n5154_, new_n5153_, new_n5152_ );
xor  ( new_n5155_, new_n5154_, new_n403_ );
nor  ( new_n5156_, new_n5155_, new_n5151_ );
and  ( new_n5157_, new_n5155_, new_n5151_ );
or   ( new_n5158_, new_n409_, new_n3178_ );
or   ( new_n5159_, new_n411_, new_n2981_ );
and  ( new_n5160_, new_n5159_, new_n5158_ );
xor  ( new_n5161_, new_n5160_, new_n328_ );
nor  ( new_n5162_, new_n5161_, new_n5157_ );
nor  ( new_n5163_, new_n5162_, new_n5156_ );
or   ( new_n5164_, new_n5163_, new_n5147_ );
and  ( new_n5165_, new_n5164_, new_n5146_ );
xnor ( new_n5166_, new_n4999_, new_n4998_ );
or   ( new_n5167_, new_n299_, new_n4995_ );
or   ( new_n5168_, new_n302_, new_n4603_ );
and  ( new_n5169_, new_n5168_, new_n5167_ );
xor  ( new_n5170_, new_n5169_, new_n293_ );
not  ( new_n5171_, RIbb2c3e8_108 );
or   ( new_n5172_, new_n268_, new_n5171_ );
or   ( new_n5173_, new_n271_, new_n4859_ );
and  ( new_n5174_, new_n5173_, new_n5172_ );
xor  ( new_n5175_, new_n5174_, new_n263_ );
or   ( new_n5176_, new_n5175_, new_n5170_ );
and  ( new_n5177_, RIbb2c370_109, RIbb2f610_1 );
and  ( new_n5178_, new_n5175_, new_n5170_ );
or   ( new_n5179_, new_n5178_, new_n5177_ );
and  ( new_n5180_, new_n5179_, new_n5176_ );
or   ( new_n5181_, new_n5180_, new_n5166_ );
and  ( new_n5182_, new_n5180_, new_n5166_ );
or   ( new_n5183_, new_n337_, new_n3696_ );
or   ( new_n5184_, new_n340_, new_n3306_ );
and  ( new_n5185_, new_n5184_, new_n5183_ );
xor  ( new_n5186_, new_n5185_, new_n332_ );
or   ( new_n5187_, new_n317_, new_n3820_ );
or   ( new_n5188_, new_n320_, new_n3694_ );
and  ( new_n5189_, new_n5188_, new_n5187_ );
xor  ( new_n5190_, new_n5189_, new_n312_ );
nor  ( new_n5191_, new_n5190_, new_n5186_ );
and  ( new_n5192_, new_n5190_, new_n5186_ );
or   ( new_n5193_, new_n283_, new_n4267_ );
or   ( new_n5194_, new_n286_, new_n4069_ );
and  ( new_n5195_, new_n5194_, new_n5193_ );
xor  ( new_n5196_, new_n5195_, new_n278_ );
nor  ( new_n5197_, new_n5196_, new_n5192_ );
nor  ( new_n5198_, new_n5197_, new_n5191_ );
or   ( new_n5199_, new_n5198_, new_n5182_ );
and  ( new_n5200_, new_n5199_, new_n5181_ );
or   ( new_n5201_, new_n5200_, new_n5165_ );
and  ( new_n5202_, new_n5200_, new_n5165_ );
not  ( new_n5203_, RIbb2e170_45 );
and  ( new_n5204_, RIbb2e080_47, RIbb2e0f8_46 );
nor  ( new_n5205_, new_n5204_, new_n5203_ );
not  ( new_n5206_, new_n5205_ );
not  ( new_n5207_, new_n4960_ );
or   ( new_n5208_, new_n5207_, new_n333_ );
not  ( new_n5209_, new_n4958_ );
or   ( new_n5210_, new_n5209_, new_n339_ );
and  ( new_n5211_, new_n5210_, new_n5208_ );
xor  ( new_n5212_, new_n5211_, new_n4708_ );
and  ( new_n5213_, new_n5212_, new_n5206_ );
or   ( new_n5214_, new_n5212_, new_n5206_ );
or   ( new_n5215_, new_n4709_, new_n313_ );
or   ( new_n5216_, new_n4711_, new_n319_ );
and  ( new_n5217_, new_n5216_, new_n5215_ );
xor  ( new_n5218_, new_n5217_, new_n4295_ );
and  ( new_n5219_, new_n5218_, new_n5214_ );
or   ( new_n5220_, new_n5219_, new_n5213_ );
or   ( new_n5221_, new_n4302_, new_n279_ );
or   ( new_n5222_, new_n4304_, new_n285_ );
and  ( new_n5223_, new_n5222_, new_n5221_ );
xor  ( new_n5224_, new_n5223_, new_n3895_ );
or   ( new_n5225_, new_n3896_, new_n294_ );
or   ( new_n5226_, new_n3898_, new_n301_ );
and  ( new_n5227_, new_n5226_, new_n5225_ );
xor  ( new_n5228_, new_n5227_, new_n3460_ );
or   ( new_n5229_, new_n5228_, new_n5224_ );
and  ( new_n5230_, new_n5228_, new_n5224_ );
or   ( new_n5231_, new_n3461_, new_n264_ );
or   ( new_n5232_, new_n3463_, new_n270_ );
and  ( new_n5233_, new_n5232_, new_n5231_ );
xor  ( new_n5234_, new_n5233_, new_n3116_ );
or   ( new_n5235_, new_n5234_, new_n5230_ );
and  ( new_n5236_, new_n5235_, new_n5229_ );
nor  ( new_n5237_, new_n5236_, new_n5220_ );
and  ( new_n5238_, new_n5236_, new_n5220_ );
or   ( new_n5239_, new_n3117_, new_n419_ );
or   ( new_n5240_, new_n3119_, new_n348_ );
and  ( new_n5241_, new_n5240_, new_n5239_ );
xor  ( new_n5242_, new_n5241_, new_n2800_ );
or   ( new_n5243_, new_n2807_, new_n509_ );
or   ( new_n5244_, new_n2809_, new_n443_ );
and  ( new_n5245_, new_n5244_, new_n5243_ );
xor  ( new_n5246_, new_n5245_, new_n2424_ );
nor  ( new_n5247_, new_n5246_, new_n5242_ );
and  ( new_n5248_, new_n5246_, new_n5242_ );
or   ( new_n5249_, new_n2425_, new_n775_ );
or   ( new_n5250_, new_n2427_, new_n515_ );
and  ( new_n5251_, new_n5250_, new_n5249_ );
xor  ( new_n5252_, new_n5251_, new_n2121_ );
nor  ( new_n5253_, new_n5252_, new_n5248_ );
nor  ( new_n5254_, new_n5253_, new_n5247_ );
nor  ( new_n5255_, new_n5254_, new_n5238_ );
nor  ( new_n5256_, new_n5255_, new_n5237_ );
or   ( new_n5257_, new_n5256_, new_n5202_ );
and  ( new_n5258_, new_n5257_, new_n5201_ );
or   ( new_n5259_, new_n5258_, new_n5113_ );
nand ( new_n5260_, new_n5258_, new_n5113_ );
xor  ( new_n5261_, new_n4714_, new_n4708_ );
xor  ( new_n5262_, new_n5261_, new_n4720_ );
xor  ( new_n5263_, new_n4862_, new_n4860_ );
xor  ( new_n5264_, new_n5263_, new_n4866_ );
nor  ( new_n5265_, new_n5264_, new_n5262_ );
and  ( new_n5266_, new_n5264_, new_n5262_ );
xor  ( new_n5267_, new_n4872_, new_n4870_ );
xnor ( new_n5268_, new_n5267_, new_n4876_ );
not  ( new_n5269_, new_n5268_ );
nor  ( new_n5270_, new_n5269_, new_n5266_ );
nor  ( new_n5271_, new_n5270_, new_n5265_ );
nand ( new_n5272_, new_n5271_, new_n5260_ );
and  ( new_n5273_, new_n5272_, new_n5259_ );
nor  ( new_n5274_, new_n5273_, new_n5087_ );
and  ( new_n5275_, new_n5273_, new_n5087_ );
xnor ( new_n5276_, new_n4722_, new_n4704_ );
xor  ( new_n5277_, new_n5276_, new_n4740_ );
xor  ( new_n5278_, new_n4970_, new_n4953_ );
xor  ( new_n5279_, new_n5278_, new_n4988_ );
xor  ( new_n5280_, new_n5016_, new_n5000_ );
xor  ( new_n5281_, new_n5280_, new_n5023_ );
nand ( new_n5282_, new_n5281_, new_n5279_ );
nor  ( new_n5283_, new_n5281_, new_n5279_ );
xor  ( new_n5284_, new_n4916_, new_n4900_ );
xor  ( new_n5285_, new_n5284_, new_n4935_ );
or   ( new_n5286_, new_n5285_, new_n5283_ );
and  ( new_n5287_, new_n5286_, new_n5282_ );
nor  ( new_n5288_, new_n5287_, new_n5277_ );
and  ( new_n5289_, new_n5287_, new_n5277_ );
xor  ( new_n5290_, new_n5033_, new_n5031_ );
xnor ( new_n5291_, new_n5290_, new_n5037_ );
not  ( new_n5292_, new_n5291_ );
nor  ( new_n5293_, new_n5292_, new_n5289_ );
nor  ( new_n5294_, new_n5293_, new_n5288_ );
not  ( new_n5295_, new_n5294_ );
nor  ( new_n5296_, new_n5295_, new_n5275_ );
nor  ( new_n5297_, new_n5296_, new_n5274_ );
or   ( new_n5298_, new_n5297_, new_n5085_ );
and  ( new_n5299_, new_n5298_, new_n5084_ );
nand ( new_n5300_, new_n5299_, new_n5071_ );
nor  ( new_n5301_, new_n5299_, new_n5071_ );
xor  ( new_n5302_, new_n5045_, new_n5043_ );
xor  ( new_n5303_, new_n5302_, new_n5049_ );
or   ( new_n5304_, new_n5303_, new_n5301_ );
and  ( new_n5305_, new_n5304_, new_n5300_ );
or   ( new_n5306_, new_n5305_, new_n5066_ );
xnor ( new_n5307_, new_n5057_, new_n4842_ );
xor  ( new_n5308_, new_n5307_, new_n5061_ );
nor  ( new_n5309_, new_n5308_, new_n5306_ );
xor  ( new_n5310_, new_n5299_, new_n5071_ );
xor  ( new_n5311_, new_n5310_, new_n5303_ );
xor  ( new_n5312_, new_n4991_, new_n4937_ );
xor  ( new_n5313_, new_n5312_, new_n5025_ );
xor  ( new_n5314_, new_n5258_, new_n5113_ );
xor  ( new_n5315_, new_n5314_, new_n5271_ );
nor  ( new_n5316_, new_n5315_, new_n5313_ );
nand ( new_n5317_, new_n5315_, new_n5313_ );
xor  ( new_n5318_, new_n5287_, new_n5277_ );
xor  ( new_n5319_, new_n5318_, new_n5292_ );
not  ( new_n5320_, new_n5319_ );
and  ( new_n5321_, new_n5320_, new_n5317_ );
or   ( new_n5322_, new_n5321_, new_n5316_ );
xor  ( new_n5323_, new_n4878_, new_n4868_ );
xor  ( new_n5324_, new_n5323_, new_n4882_ );
xnor ( new_n5325_, new_n4962_, new_n4957_ );
xor  ( new_n5326_, new_n5325_, new_n4968_ );
xnor ( new_n5327_, new_n5121_, new_n5117_ );
xor  ( new_n5328_, new_n5327_, new_n5127_ );
xnor ( new_n5329_, new_n5155_, new_n5151_ );
xor  ( new_n5330_, new_n5329_, new_n5161_ );
or   ( new_n5331_, new_n5330_, new_n5328_ );
and  ( new_n5332_, new_n5330_, new_n5328_ );
xor  ( new_n5333_, new_n5190_, new_n5186_ );
xnor ( new_n5334_, new_n5333_, new_n5196_ );
or   ( new_n5335_, new_n5334_, new_n5332_ );
and  ( new_n5336_, new_n5335_, new_n5331_ );
nor  ( new_n5337_, new_n5336_, new_n5326_ );
and  ( new_n5338_, new_n5336_, new_n5326_ );
xnor ( new_n5339_, new_n5137_, new_n5133_ );
xor  ( new_n5340_, new_n5339_, new_n5143_ );
xnor ( new_n5341_, new_n5228_, new_n5224_ );
xor  ( new_n5342_, new_n5341_, new_n5234_ );
nor  ( new_n5343_, new_n5342_, new_n5340_ );
and  ( new_n5344_, new_n5342_, new_n5340_ );
xor  ( new_n5345_, new_n5246_, new_n5242_ );
xnor ( new_n5346_, new_n5345_, new_n5252_ );
nor  ( new_n5347_, new_n5346_, new_n5344_ );
nor  ( new_n5348_, new_n5347_, new_n5343_ );
nor  ( new_n5349_, new_n5348_, new_n5338_ );
or   ( new_n5350_, new_n5349_, new_n5337_ );
or   ( new_n5351_, new_n4302_, new_n301_ );
or   ( new_n5352_, new_n4304_, new_n279_ );
and  ( new_n5353_, new_n5352_, new_n5351_ );
xor  ( new_n5354_, new_n5353_, new_n3895_ );
or   ( new_n5355_, new_n3896_, new_n270_ );
or   ( new_n5356_, new_n3898_, new_n294_ );
and  ( new_n5357_, new_n5356_, new_n5355_ );
xor  ( new_n5358_, new_n5357_, new_n3460_ );
or   ( new_n5359_, new_n5358_, new_n5354_ );
and  ( new_n5360_, new_n5358_, new_n5354_ );
or   ( new_n5361_, new_n3461_, new_n348_ );
or   ( new_n5362_, new_n3463_, new_n264_ );
and  ( new_n5363_, new_n5362_, new_n5361_ );
xor  ( new_n5364_, new_n5363_, new_n3116_ );
or   ( new_n5365_, new_n5364_, new_n5360_ );
and  ( new_n5366_, new_n5365_, new_n5359_ );
or   ( new_n5367_, new_n5207_, new_n319_ );
or   ( new_n5368_, new_n5209_, new_n333_ );
and  ( new_n5369_, new_n5368_, new_n5367_ );
xor  ( new_n5370_, new_n5369_, new_n4707_ );
xor  ( new_n5371_, RIbb2e080_47, RIbb2e0f8_46 );
xor  ( new_n5372_, RIbb2e0f8_46, new_n5203_ );
nor  ( new_n5373_, new_n5372_, new_n5371_ );
and  ( new_n5374_, new_n5373_, RIbb2d810_65 );
xor  ( new_n5375_, new_n5374_, new_n5206_ );
nand ( new_n5376_, new_n5375_, new_n5370_ );
nor  ( new_n5377_, new_n5375_, new_n5370_ );
or   ( new_n5378_, new_n4709_, new_n285_ );
or   ( new_n5379_, new_n4711_, new_n313_ );
and  ( new_n5380_, new_n5379_, new_n5378_ );
xor  ( new_n5381_, new_n5380_, new_n4295_ );
or   ( new_n5382_, new_n5381_, new_n5377_ );
and  ( new_n5383_, new_n5382_, new_n5376_ );
or   ( new_n5384_, new_n5383_, new_n5366_ );
and  ( new_n5385_, new_n5383_, new_n5366_ );
or   ( new_n5386_, new_n3117_, new_n443_ );
or   ( new_n5387_, new_n3119_, new_n419_ );
and  ( new_n5388_, new_n5387_, new_n5386_ );
xor  ( new_n5389_, new_n5388_, new_n2800_ );
or   ( new_n5390_, new_n2807_, new_n515_ );
or   ( new_n5391_, new_n2809_, new_n509_ );
and  ( new_n5392_, new_n5391_, new_n5390_ );
xor  ( new_n5393_, new_n5392_, new_n2424_ );
nor  ( new_n5394_, new_n5393_, new_n5389_ );
and  ( new_n5395_, new_n5393_, new_n5389_ );
or   ( new_n5396_, new_n2425_, new_n805_ );
or   ( new_n5397_, new_n2427_, new_n775_ );
and  ( new_n5398_, new_n5397_, new_n5396_ );
xor  ( new_n5399_, new_n5398_, new_n2121_ );
nor  ( new_n5400_, new_n5399_, new_n5395_ );
nor  ( new_n5401_, new_n5400_, new_n5394_ );
or   ( new_n5402_, new_n5401_, new_n5385_ );
and  ( new_n5403_, new_n5402_, new_n5384_ );
xor  ( new_n5404_, new_n5175_, new_n5170_ );
xor  ( new_n5405_, new_n5404_, new_n5177_ );
or   ( new_n5406_, new_n337_, new_n3694_ );
or   ( new_n5407_, new_n340_, new_n3696_ );
and  ( new_n5408_, new_n5407_, new_n5406_ );
xor  ( new_n5409_, new_n5408_, new_n332_ );
or   ( new_n5410_, new_n317_, new_n4069_ );
or   ( new_n5411_, new_n320_, new_n3820_ );
and  ( new_n5412_, new_n5411_, new_n5410_ );
xor  ( new_n5413_, new_n5412_, new_n312_ );
or   ( new_n5414_, new_n5413_, new_n5409_ );
and  ( new_n5415_, new_n5413_, new_n5409_ );
or   ( new_n5416_, new_n283_, new_n4603_ );
or   ( new_n5417_, new_n286_, new_n4267_ );
and  ( new_n5418_, new_n5417_, new_n5416_ );
xor  ( new_n5419_, new_n5418_, new_n278_ );
or   ( new_n5420_, new_n5419_, new_n5415_ );
and  ( new_n5421_, new_n5420_, new_n5414_ );
or   ( new_n5422_, new_n5421_, new_n5405_ );
and  ( new_n5423_, new_n5421_, new_n5405_ );
or   ( new_n5424_, new_n299_, new_n4859_ );
or   ( new_n5425_, new_n302_, new_n4995_ );
and  ( new_n5426_, new_n5425_, new_n5424_ );
xor  ( new_n5427_, new_n5426_, new_n293_ );
not  ( new_n5428_, RIbb2c370_109 );
or   ( new_n5429_, new_n268_, new_n5428_ );
or   ( new_n5430_, new_n271_, new_n5171_ );
and  ( new_n5431_, new_n5430_, new_n5429_ );
xor  ( new_n5432_, new_n5431_, new_n263_ );
nor  ( new_n5433_, new_n5432_, new_n5427_ );
and  ( new_n5434_, RIbb2c2f8_110, RIbb2f610_1 );
and  ( new_n5435_, new_n5432_, new_n5427_ );
nor  ( new_n5436_, new_n5435_, new_n5434_ );
nor  ( new_n5437_, new_n5436_, new_n5433_ );
or   ( new_n5438_, new_n5437_, new_n5423_ );
and  ( new_n5439_, new_n5438_, new_n5422_ );
or   ( new_n5440_, new_n5439_, new_n5403_ );
and  ( new_n5441_, new_n5439_, new_n5403_ );
or   ( new_n5442_, new_n1364_, new_n1754_ );
or   ( new_n5443_, new_n1366_, new_n1523_ );
and  ( new_n5444_, new_n5443_, new_n5442_ );
xor  ( new_n5445_, new_n5444_, new_n1129_ );
or   ( new_n5446_, new_n1135_, new_n2057_ );
or   ( new_n5447_, new_n1137_, new_n1899_ );
and  ( new_n5448_, new_n5447_, new_n5446_ );
xor  ( new_n5449_, new_n5448_, new_n896_ );
or   ( new_n5450_, new_n5449_, new_n5445_ );
and  ( new_n5451_, new_n5449_, new_n5445_ );
or   ( new_n5452_, new_n897_, new_n2291_ );
or   ( new_n5453_, new_n899_, new_n2178_ );
and  ( new_n5454_, new_n5453_, new_n5452_ );
xor  ( new_n5455_, new_n5454_, new_n748_ );
or   ( new_n5456_, new_n5455_, new_n5451_ );
and  ( new_n5457_, new_n5456_, new_n5450_ );
or   ( new_n5458_, new_n2122_, new_n986_ );
or   ( new_n5459_, new_n2124_, new_n886_ );
and  ( new_n5460_, new_n5459_, new_n5458_ );
xor  ( new_n5461_, new_n5460_, new_n1843_ );
or   ( new_n5462_, new_n1844_, new_n1213_ );
or   ( new_n5463_, new_n1846_, new_n1168_ );
and  ( new_n5464_, new_n5463_, new_n5462_ );
xor  ( new_n5465_, new_n5464_, new_n1586_ );
or   ( new_n5466_, new_n5465_, new_n5461_ );
and  ( new_n5467_, new_n5465_, new_n5461_ );
or   ( new_n5468_, new_n1593_, new_n1525_ );
or   ( new_n5469_, new_n1595_, new_n1318_ );
and  ( new_n5470_, new_n5469_, new_n5468_ );
xor  ( new_n5471_, new_n5470_, new_n1358_ );
or   ( new_n5472_, new_n5471_, new_n5467_ );
and  ( new_n5473_, new_n5472_, new_n5466_ );
nor  ( new_n5474_, new_n5473_, new_n5457_ );
and  ( new_n5475_, new_n5473_, new_n5457_ );
or   ( new_n5476_, new_n755_, new_n2646_ );
or   ( new_n5477_, new_n757_, new_n2475_ );
and  ( new_n5478_, new_n5477_, new_n5476_ );
xor  ( new_n5479_, new_n5478_, new_n523_ );
or   ( new_n5480_, new_n524_, new_n2981_ );
or   ( new_n5481_, new_n526_, new_n2751_ );
and  ( new_n5482_, new_n5481_, new_n5480_ );
xor  ( new_n5483_, new_n5482_, new_n403_ );
nor  ( new_n5484_, new_n5483_, new_n5479_ );
and  ( new_n5485_, new_n5483_, new_n5479_ );
or   ( new_n5486_, new_n409_, new_n3306_ );
or   ( new_n5487_, new_n411_, new_n3178_ );
and  ( new_n5488_, new_n5487_, new_n5486_ );
xor  ( new_n5489_, new_n5488_, new_n328_ );
nor  ( new_n5490_, new_n5489_, new_n5485_ );
nor  ( new_n5491_, new_n5490_, new_n5484_ );
nor  ( new_n5492_, new_n5491_, new_n5475_ );
nor  ( new_n5493_, new_n5492_, new_n5474_ );
or   ( new_n5494_, new_n5493_, new_n5441_ );
and  ( new_n5495_, new_n5494_, new_n5440_ );
or   ( new_n5496_, new_n5495_, new_n5350_ );
nand ( new_n5497_, new_n5495_, new_n5350_ );
xor  ( new_n5498_, new_n5105_, new_n5103_ );
xor  ( new_n5499_, new_n5498_, new_n5109_ );
xnor ( new_n5500_, new_n5093_, new_n5091_ );
xor  ( new_n5501_, new_n5500_, new_n5097_ );
and  ( new_n5502_, new_n5501_, new_n5499_ );
nor  ( new_n5503_, new_n5501_, new_n5499_ );
xor  ( new_n5504_, new_n5180_, new_n5166_ );
xnor ( new_n5505_, new_n5504_, new_n5198_ );
nor  ( new_n5506_, new_n5505_, new_n5503_ );
nor  ( new_n5507_, new_n5506_, new_n5502_ );
nand ( new_n5508_, new_n5507_, new_n5497_ );
and  ( new_n5509_, new_n5508_, new_n5496_ );
or   ( new_n5510_, new_n5509_, new_n5324_ );
nand ( new_n5511_, new_n5509_, new_n5324_ );
xor  ( new_n5512_, new_n5099_, new_n5089_ );
xor  ( new_n5513_, new_n5512_, new_n5111_ );
xnor ( new_n5514_, new_n5281_, new_n5279_ );
xor  ( new_n5515_, new_n5514_, new_n5285_ );
and  ( new_n5516_, new_n5515_, new_n5513_ );
nor  ( new_n5517_, new_n5515_, new_n5513_ );
xor  ( new_n5518_, new_n5264_, new_n5262_ );
xor  ( new_n5519_, new_n5518_, new_n5269_ );
nor  ( new_n5520_, new_n5519_, new_n5517_ );
nor  ( new_n5521_, new_n5520_, new_n5516_ );
nand ( new_n5522_, new_n5521_, new_n5511_ );
and  ( new_n5523_, new_n5522_, new_n5510_ );
nor  ( new_n5524_, new_n5523_, new_n5322_ );
nand ( new_n5525_, new_n5523_, new_n5322_ );
xor  ( new_n5526_, new_n5077_, new_n5075_ );
xnor ( new_n5527_, new_n5526_, new_n5081_ );
and  ( new_n5528_, new_n5527_, new_n5525_ );
or   ( new_n5529_, new_n5528_, new_n5524_ );
xnor ( new_n5530_, new_n5083_, new_n5073_ );
xor  ( new_n5531_, new_n5530_, new_n5297_ );
or   ( new_n5532_, new_n5531_, new_n5529_ );
nand ( new_n5533_, new_n5531_, new_n5529_ );
xor  ( new_n5534_, new_n5070_, new_n5068_ );
nand ( new_n5535_, new_n5534_, new_n5533_ );
and  ( new_n5536_, new_n5535_, new_n5532_ );
nor  ( new_n5537_, new_n5536_, new_n5311_ );
xor  ( new_n5538_, new_n5305_, new_n5066_ );
and  ( new_n5539_, new_n5538_, new_n5537_ );
xor  ( new_n5540_, new_n5531_, new_n5529_ );
xor  ( new_n5541_, new_n5540_, new_n5534_ );
xnor ( new_n5542_, new_n5523_, new_n5322_ );
xor  ( new_n5543_, new_n5542_, new_n5527_ );
or   ( new_n5544_, new_n409_, new_n3696_ );
or   ( new_n5545_, new_n411_, new_n3306_ );
and  ( new_n5546_, new_n5545_, new_n5544_ );
xor  ( new_n5547_, new_n5546_, new_n328_ );
or   ( new_n5548_, new_n337_, new_n3820_ );
or   ( new_n5549_, new_n340_, new_n3694_ );
and  ( new_n5550_, new_n5549_, new_n5548_ );
xor  ( new_n5551_, new_n5550_, new_n332_ );
nor  ( new_n5552_, new_n5551_, new_n5547_ );
and  ( new_n5553_, new_n5551_, new_n5547_ );
or   ( new_n5554_, new_n317_, new_n4267_ );
or   ( new_n5555_, new_n320_, new_n4069_ );
and  ( new_n5556_, new_n5555_, new_n5554_ );
xor  ( new_n5557_, new_n5556_, new_n312_ );
nor  ( new_n5558_, new_n5557_, new_n5553_ );
nor  ( new_n5559_, new_n5558_, new_n5552_ );
or   ( new_n5560_, new_n283_, new_n4995_ );
or   ( new_n5561_, new_n286_, new_n4603_ );
and  ( new_n5562_, new_n5561_, new_n5560_ );
xor  ( new_n5563_, new_n5562_, new_n278_ );
or   ( new_n5564_, new_n299_, new_n5171_ );
or   ( new_n5565_, new_n302_, new_n4859_ );
and  ( new_n5566_, new_n5565_, new_n5564_ );
xor  ( new_n5567_, new_n5566_, new_n293_ );
or   ( new_n5568_, new_n5567_, new_n5563_ );
and  ( new_n5569_, new_n5567_, new_n5563_ );
not  ( new_n5570_, RIbb2c2f8_110 );
or   ( new_n5571_, new_n268_, new_n5570_ );
or   ( new_n5572_, new_n271_, new_n5428_ );
and  ( new_n5573_, new_n5572_, new_n5571_ );
xor  ( new_n5574_, new_n5573_, new_n263_ );
or   ( new_n5575_, new_n5574_, new_n5569_ );
and  ( new_n5576_, new_n5575_, new_n5568_ );
or   ( new_n5577_, new_n5576_, new_n5559_ );
or   ( new_n5578_, new_n4709_, new_n279_ );
or   ( new_n5579_, new_n4711_, new_n285_ );
and  ( new_n5580_, new_n5579_, new_n5578_ );
xor  ( new_n5581_, new_n5580_, new_n4295_ );
or   ( new_n5582_, new_n4302_, new_n294_ );
or   ( new_n5583_, new_n4304_, new_n301_ );
and  ( new_n5584_, new_n5583_, new_n5582_ );
xor  ( new_n5585_, new_n5584_, new_n3895_ );
nor  ( new_n5586_, new_n5585_, new_n5581_ );
and  ( new_n5587_, new_n5585_, new_n5581_ );
or   ( new_n5588_, new_n3896_, new_n264_ );
or   ( new_n5589_, new_n3898_, new_n270_ );
and  ( new_n5590_, new_n5589_, new_n5588_ );
xor  ( new_n5591_, new_n5590_, new_n3460_ );
nor  ( new_n5592_, new_n5591_, new_n5587_ );
or   ( new_n5593_, new_n5592_, new_n5586_ );
not  ( new_n5594_, RIbb2e080_47 );
and  ( new_n5595_, RIbb2df90_49, RIbb2e008_48 );
nor  ( new_n5596_, new_n5595_, new_n5594_ );
not  ( new_n5597_, new_n5596_ );
or   ( new_n5598_, new_n5207_, new_n313_ );
or   ( new_n5599_, new_n5209_, new_n319_ );
and  ( new_n5600_, new_n5599_, new_n5598_ );
xor  ( new_n5601_, new_n5600_, new_n4708_ );
nand ( new_n5602_, new_n5601_, new_n5597_ );
or   ( new_n5603_, new_n5601_, new_n5597_ );
not  ( new_n5604_, new_n5373_ );
or   ( new_n5605_, new_n5604_, new_n333_ );
not  ( new_n5606_, new_n5371_ );
or   ( new_n5607_, new_n5606_, new_n339_ );
and  ( new_n5608_, new_n5607_, new_n5605_ );
xor  ( new_n5609_, new_n5608_, new_n5206_ );
nand ( new_n5610_, new_n5609_, new_n5603_ );
and  ( new_n5611_, new_n5610_, new_n5602_ );
nand ( new_n5612_, new_n5611_, new_n5593_ );
nor  ( new_n5613_, new_n5611_, new_n5593_ );
or   ( new_n5614_, new_n3461_, new_n419_ );
or   ( new_n5615_, new_n3463_, new_n348_ );
and  ( new_n5616_, new_n5615_, new_n5614_ );
xor  ( new_n5617_, new_n5616_, new_n3116_ );
or   ( new_n5618_, new_n3117_, new_n509_ );
or   ( new_n5619_, new_n3119_, new_n443_ );
and  ( new_n5620_, new_n5619_, new_n5618_ );
xor  ( new_n5621_, new_n5620_, new_n2800_ );
nor  ( new_n5622_, new_n5621_, new_n5617_ );
and  ( new_n5623_, new_n5621_, new_n5617_ );
or   ( new_n5624_, new_n2807_, new_n775_ );
or   ( new_n5625_, new_n2809_, new_n515_ );
and  ( new_n5626_, new_n5625_, new_n5624_ );
xor  ( new_n5627_, new_n5626_, new_n2424_ );
nor  ( new_n5628_, new_n5627_, new_n5623_ );
nor  ( new_n5629_, new_n5628_, new_n5622_ );
or   ( new_n5630_, new_n5629_, new_n5613_ );
and  ( new_n5631_, new_n5630_, new_n5612_ );
nor  ( new_n5632_, new_n5631_, new_n5577_ );
nand ( new_n5633_, new_n5631_, new_n5577_ );
or   ( new_n5634_, new_n1593_, new_n1523_ );
or   ( new_n5635_, new_n1595_, new_n1525_ );
and  ( new_n5636_, new_n5635_, new_n5634_ );
xor  ( new_n5637_, new_n5636_, new_n1358_ );
or   ( new_n5638_, new_n1364_, new_n1899_ );
or   ( new_n5639_, new_n1366_, new_n1754_ );
and  ( new_n5640_, new_n5639_, new_n5638_ );
xor  ( new_n5641_, new_n5640_, new_n1129_ );
or   ( new_n5642_, new_n5641_, new_n5637_ );
and  ( new_n5643_, new_n5641_, new_n5637_ );
or   ( new_n5644_, new_n1135_, new_n2178_ );
or   ( new_n5645_, new_n1137_, new_n2057_ );
and  ( new_n5646_, new_n5645_, new_n5644_ );
xor  ( new_n5647_, new_n5646_, new_n896_ );
or   ( new_n5648_, new_n5647_, new_n5643_ );
and  ( new_n5649_, new_n5648_, new_n5642_ );
or   ( new_n5650_, new_n897_, new_n2475_ );
or   ( new_n5651_, new_n899_, new_n2291_ );
and  ( new_n5652_, new_n5651_, new_n5650_ );
xor  ( new_n5653_, new_n5652_, new_n748_ );
or   ( new_n5654_, new_n755_, new_n2751_ );
or   ( new_n5655_, new_n757_, new_n2646_ );
and  ( new_n5656_, new_n5655_, new_n5654_ );
xor  ( new_n5657_, new_n5656_, new_n523_ );
or   ( new_n5658_, new_n5657_, new_n5653_ );
and  ( new_n5659_, new_n5657_, new_n5653_ );
or   ( new_n5660_, new_n524_, new_n3178_ );
or   ( new_n5661_, new_n526_, new_n2981_ );
and  ( new_n5662_, new_n5661_, new_n5660_ );
xor  ( new_n5663_, new_n5662_, new_n403_ );
or   ( new_n5664_, new_n5663_, new_n5659_ );
and  ( new_n5665_, new_n5664_, new_n5658_ );
nor  ( new_n5666_, new_n5665_, new_n5649_ );
and  ( new_n5667_, new_n5665_, new_n5649_ );
or   ( new_n5668_, new_n2425_, new_n886_ );
or   ( new_n5669_, new_n2427_, new_n805_ );
and  ( new_n5670_, new_n5669_, new_n5668_ );
xor  ( new_n5671_, new_n5670_, new_n2121_ );
or   ( new_n5672_, new_n2122_, new_n1168_ );
or   ( new_n5673_, new_n2124_, new_n986_ );
and  ( new_n5674_, new_n5673_, new_n5672_ );
xor  ( new_n5675_, new_n5674_, new_n1843_ );
nor  ( new_n5676_, new_n5675_, new_n5671_ );
and  ( new_n5677_, new_n5675_, new_n5671_ );
or   ( new_n5678_, new_n1844_, new_n1318_ );
or   ( new_n5679_, new_n1846_, new_n1213_ );
and  ( new_n5680_, new_n5679_, new_n5678_ );
xor  ( new_n5681_, new_n5680_, new_n1586_ );
nor  ( new_n5682_, new_n5681_, new_n5677_ );
nor  ( new_n5683_, new_n5682_, new_n5676_ );
nor  ( new_n5684_, new_n5683_, new_n5667_ );
nor  ( new_n5685_, new_n5684_, new_n5666_ );
not  ( new_n5686_, new_n5685_ );
and  ( new_n5687_, new_n5686_, new_n5633_ );
or   ( new_n5688_, new_n5687_, new_n5632_ );
xor  ( new_n5689_, new_n5375_, new_n5370_ );
xnor ( new_n5690_, new_n5689_, new_n5381_ );
xnor ( new_n5691_, new_n5358_, new_n5354_ );
xor  ( new_n5692_, new_n5691_, new_n5364_ );
or   ( new_n5693_, new_n5692_, new_n5690_ );
xnor ( new_n5694_, new_n5465_, new_n5461_ );
xor  ( new_n5695_, new_n5694_, new_n5471_ );
xnor ( new_n5696_, new_n5449_, new_n5445_ );
xor  ( new_n5697_, new_n5696_, new_n5455_ );
or   ( new_n5698_, new_n5697_, new_n5695_ );
and  ( new_n5699_, new_n5697_, new_n5695_ );
xor  ( new_n5700_, new_n5393_, new_n5389_ );
xnor ( new_n5701_, new_n5700_, new_n5399_ );
or   ( new_n5702_, new_n5701_, new_n5699_ );
and  ( new_n5703_, new_n5702_, new_n5698_ );
or   ( new_n5704_, new_n5703_, new_n5693_ );
and  ( new_n5705_, new_n5703_, new_n5693_ );
xnor ( new_n5706_, new_n5483_, new_n5479_ );
xor  ( new_n5707_, new_n5706_, new_n5489_ );
xnor ( new_n5708_, new_n5413_, new_n5409_ );
xor  ( new_n5709_, new_n5708_, new_n5419_ );
nor  ( new_n5710_, new_n5709_, new_n5707_ );
and  ( new_n5711_, new_n5709_, new_n5707_ );
xor  ( new_n5712_, new_n5432_, new_n5427_ );
xnor ( new_n5713_, new_n5712_, new_n5434_ );
nor  ( new_n5714_, new_n5713_, new_n5711_ );
nor  ( new_n5715_, new_n5714_, new_n5710_ );
or   ( new_n5716_, new_n5715_, new_n5705_ );
and  ( new_n5717_, new_n5716_, new_n5704_ );
or   ( new_n5718_, new_n5717_, new_n5688_ );
nand ( new_n5719_, new_n5717_, new_n5688_ );
xor  ( new_n5720_, new_n5212_, new_n5206_ );
xor  ( new_n5721_, new_n5720_, new_n5218_ );
xnor ( new_n5722_, new_n5342_, new_n5340_ );
xor  ( new_n5723_, new_n5722_, new_n5346_ );
nor  ( new_n5724_, new_n5723_, new_n5721_ );
and  ( new_n5725_, new_n5723_, new_n5721_ );
xor  ( new_n5726_, new_n5330_, new_n5328_ );
xnor ( new_n5727_, new_n5726_, new_n5334_ );
nor  ( new_n5728_, new_n5727_, new_n5725_ );
nor  ( new_n5729_, new_n5728_, new_n5724_ );
nand ( new_n5730_, new_n5729_, new_n5719_ );
and  ( new_n5731_, new_n5730_, new_n5718_ );
xnor ( new_n5732_, new_n5236_, new_n5220_ );
xor  ( new_n5733_, new_n5732_, new_n5254_ );
xnor ( new_n5734_, new_n5383_, new_n5366_ );
xor  ( new_n5735_, new_n5734_, new_n5401_ );
xnor ( new_n5736_, new_n5473_, new_n5457_ );
xor  ( new_n5737_, new_n5736_, new_n5491_ );
or   ( new_n5738_, new_n5737_, new_n5735_ );
and  ( new_n5739_, new_n5737_, new_n5735_ );
xnor ( new_n5740_, new_n5421_, new_n5405_ );
xor  ( new_n5741_, new_n5740_, new_n5437_ );
or   ( new_n5742_, new_n5741_, new_n5739_ );
and  ( new_n5743_, new_n5742_, new_n5738_ );
or   ( new_n5744_, new_n5743_, new_n5733_ );
and  ( new_n5745_, new_n5743_, new_n5733_ );
xor  ( new_n5746_, new_n5145_, new_n5129_ );
xnor ( new_n5747_, new_n5746_, new_n5163_ );
or   ( new_n5748_, new_n5747_, new_n5745_ );
and  ( new_n5749_, new_n5748_, new_n5744_ );
or   ( new_n5750_, new_n5749_, new_n5731_ );
and  ( new_n5751_, new_n5749_, new_n5731_ );
xor  ( new_n5752_, new_n5336_, new_n5326_ );
xor  ( new_n5753_, new_n5752_, new_n5348_ );
xnor ( new_n5754_, new_n5439_, new_n5403_ );
xor  ( new_n5755_, new_n5754_, new_n5493_ );
nor  ( new_n5756_, new_n5755_, new_n5753_ );
and  ( new_n5757_, new_n5755_, new_n5753_ );
xor  ( new_n5758_, new_n5501_, new_n5499_ );
xnor ( new_n5759_, new_n5758_, new_n5505_ );
not  ( new_n5760_, new_n5759_ );
nor  ( new_n5761_, new_n5760_, new_n5757_ );
nor  ( new_n5762_, new_n5761_, new_n5756_ );
or   ( new_n5763_, new_n5762_, new_n5751_ );
and  ( new_n5764_, new_n5763_, new_n5750_ );
xor  ( new_n5765_, new_n5495_, new_n5350_ );
xor  ( new_n5766_, new_n5765_, new_n5507_ );
xnor ( new_n5767_, new_n5200_, new_n5165_ );
xor  ( new_n5768_, new_n5767_, new_n5256_ );
or   ( new_n5769_, new_n5768_, new_n5766_ );
and  ( new_n5770_, new_n5768_, new_n5766_ );
xor  ( new_n5771_, new_n5515_, new_n5513_ );
xor  ( new_n5772_, new_n5771_, new_n5519_ );
or   ( new_n5773_, new_n5772_, new_n5770_ );
and  ( new_n5774_, new_n5773_, new_n5769_ );
nand ( new_n5775_, new_n5774_, new_n5764_ );
nor  ( new_n5776_, new_n5774_, new_n5764_ );
xor  ( new_n5777_, new_n5315_, new_n5313_ );
xor  ( new_n5778_, new_n5777_, new_n5320_ );
or   ( new_n5779_, new_n5778_, new_n5776_ );
and  ( new_n5780_, new_n5779_, new_n5775_ );
or   ( new_n5781_, new_n5780_, new_n5543_ );
nand ( new_n5782_, new_n5780_, new_n5543_ );
xor  ( new_n5783_, new_n5273_, new_n5087_ );
xor  ( new_n5784_, new_n5783_, new_n5294_ );
nand ( new_n5785_, new_n5784_, new_n5782_ );
and  ( new_n5786_, new_n5785_, new_n5781_ );
and  ( new_n5787_, new_n5786_, new_n5541_ );
xor  ( new_n5788_, new_n5536_, new_n5311_ );
and  ( new_n5789_, new_n5788_, new_n5787_ );
xor  ( new_n5790_, new_n5768_, new_n5766_ );
xor  ( new_n5791_, new_n5790_, new_n5772_ );
xor  ( new_n5792_, new_n5717_, new_n5688_ );
xor  ( new_n5793_, new_n5792_, new_n5729_ );
xnor ( new_n5794_, new_n5743_, new_n5733_ );
xor  ( new_n5795_, new_n5794_, new_n5747_ );
nand ( new_n5796_, new_n5795_, new_n5793_ );
nor  ( new_n5797_, new_n5795_, new_n5793_ );
xor  ( new_n5798_, new_n5755_, new_n5753_ );
xor  ( new_n5799_, new_n5798_, new_n5760_ );
or   ( new_n5800_, new_n5799_, new_n5797_ );
and  ( new_n5801_, new_n5800_, new_n5796_ );
or   ( new_n5802_, new_n5801_, new_n5791_ );
and  ( new_n5803_, new_n5801_, new_n5791_ );
xor  ( new_n5804_, new_n5631_, new_n5577_ );
xor  ( new_n5805_, new_n5804_, new_n5686_ );
not  ( new_n5806_, new_n5805_ );
xnor ( new_n5807_, new_n5703_, new_n5693_ );
xor  ( new_n5808_, new_n5807_, new_n5715_ );
nand ( new_n5809_, new_n5808_, new_n5806_ );
xnor ( new_n5810_, new_n5697_, new_n5695_ );
xor  ( new_n5811_, new_n5810_, new_n5701_ );
xnor ( new_n5812_, new_n5709_, new_n5707_ );
xor  ( new_n5813_, new_n5812_, new_n5713_ );
nor  ( new_n5814_, new_n5813_, new_n5811_ );
nand ( new_n5815_, new_n5813_, new_n5811_ );
xor  ( new_n5816_, new_n5692_, new_n5690_ );
not  ( new_n5817_, new_n5816_ );
and  ( new_n5818_, new_n5817_, new_n5815_ );
or   ( new_n5819_, new_n5818_, new_n5814_ );
or   ( new_n5820_, new_n2425_, new_n986_ );
or   ( new_n5821_, new_n2427_, new_n886_ );
and  ( new_n5822_, new_n5821_, new_n5820_ );
xor  ( new_n5823_, new_n5822_, new_n2121_ );
or   ( new_n5824_, new_n2122_, new_n1213_ );
or   ( new_n5825_, new_n2124_, new_n1168_ );
and  ( new_n5826_, new_n5825_, new_n5824_ );
xor  ( new_n5827_, new_n5826_, new_n1843_ );
or   ( new_n5828_, new_n5827_, new_n5823_ );
and  ( new_n5829_, new_n5827_, new_n5823_ );
or   ( new_n5830_, new_n1844_, new_n1525_ );
or   ( new_n5831_, new_n1846_, new_n1318_ );
and  ( new_n5832_, new_n5831_, new_n5830_ );
xor  ( new_n5833_, new_n5832_, new_n1586_ );
or   ( new_n5834_, new_n5833_, new_n5829_ );
and  ( new_n5835_, new_n5834_, new_n5828_ );
or   ( new_n5836_, new_n1593_, new_n1754_ );
or   ( new_n5837_, new_n1595_, new_n1523_ );
and  ( new_n5838_, new_n5837_, new_n5836_ );
xor  ( new_n5839_, new_n5838_, new_n1358_ );
or   ( new_n5840_, new_n1364_, new_n2057_ );
or   ( new_n5841_, new_n1366_, new_n1899_ );
and  ( new_n5842_, new_n5841_, new_n5840_ );
xor  ( new_n5843_, new_n5842_, new_n1129_ );
or   ( new_n5844_, new_n5843_, new_n5839_ );
and  ( new_n5845_, new_n5843_, new_n5839_ );
or   ( new_n5846_, new_n1135_, new_n2291_ );
or   ( new_n5847_, new_n1137_, new_n2178_ );
and  ( new_n5848_, new_n5847_, new_n5846_ );
xor  ( new_n5849_, new_n5848_, new_n896_ );
or   ( new_n5850_, new_n5849_, new_n5845_ );
and  ( new_n5851_, new_n5850_, new_n5844_ );
or   ( new_n5852_, new_n5851_, new_n5835_ );
and  ( new_n5853_, new_n5851_, new_n5835_ );
or   ( new_n5854_, new_n897_, new_n2646_ );
or   ( new_n5855_, new_n899_, new_n2475_ );
and  ( new_n5856_, new_n5855_, new_n5854_ );
xor  ( new_n5857_, new_n5856_, new_n748_ );
or   ( new_n5858_, new_n755_, new_n2981_ );
or   ( new_n5859_, new_n757_, new_n2751_ );
and  ( new_n5860_, new_n5859_, new_n5858_ );
xor  ( new_n5861_, new_n5860_, new_n523_ );
nor  ( new_n5862_, new_n5861_, new_n5857_ );
and  ( new_n5863_, new_n5861_, new_n5857_ );
or   ( new_n5864_, new_n524_, new_n3306_ );
or   ( new_n5865_, new_n526_, new_n3178_ );
and  ( new_n5866_, new_n5865_, new_n5864_ );
xor  ( new_n5867_, new_n5866_, new_n403_ );
nor  ( new_n5868_, new_n5867_, new_n5863_ );
nor  ( new_n5869_, new_n5868_, new_n5862_ );
or   ( new_n5870_, new_n5869_, new_n5853_ );
and  ( new_n5871_, new_n5870_, new_n5852_ );
or   ( new_n5872_, new_n409_, new_n3694_ );
or   ( new_n5873_, new_n411_, new_n3696_ );
and  ( new_n5874_, new_n5873_, new_n5872_ );
xor  ( new_n5875_, new_n5874_, new_n328_ );
or   ( new_n5876_, new_n337_, new_n4069_ );
or   ( new_n5877_, new_n340_, new_n3820_ );
and  ( new_n5878_, new_n5877_, new_n5876_ );
xor  ( new_n5879_, new_n5878_, new_n332_ );
or   ( new_n5880_, new_n5879_, new_n5875_ );
and  ( new_n5881_, new_n5879_, new_n5875_ );
or   ( new_n5882_, new_n317_, new_n4603_ );
or   ( new_n5883_, new_n320_, new_n4267_ );
and  ( new_n5884_, new_n5883_, new_n5882_ );
xor  ( new_n5885_, new_n5884_, new_n312_ );
or   ( new_n5886_, new_n5885_, new_n5881_ );
and  ( new_n5887_, new_n5886_, new_n5880_ );
and  ( new_n5888_, RIbb2c208_112, RIbb2f610_1 );
or   ( new_n5889_, new_n283_, new_n4859_ );
or   ( new_n5890_, new_n286_, new_n4995_ );
and  ( new_n5891_, new_n5890_, new_n5889_ );
xor  ( new_n5892_, new_n5891_, new_n278_ );
or   ( new_n5893_, new_n299_, new_n5428_ );
or   ( new_n5894_, new_n302_, new_n5171_ );
and  ( new_n5895_, new_n5894_, new_n5893_ );
xor  ( new_n5896_, new_n5895_, new_n293_ );
or   ( new_n5897_, new_n5896_, new_n5892_ );
and  ( new_n5898_, new_n5896_, new_n5892_ );
not  ( new_n5899_, RIbb2c280_111 );
or   ( new_n5900_, new_n268_, new_n5899_ );
or   ( new_n5901_, new_n271_, new_n5570_ );
and  ( new_n5902_, new_n5901_, new_n5900_ );
xor  ( new_n5903_, new_n5902_, new_n263_ );
or   ( new_n5904_, new_n5903_, new_n5898_ );
and  ( new_n5905_, new_n5904_, new_n5897_ );
and  ( new_n5906_, new_n5905_, new_n5888_ );
or   ( new_n5907_, new_n5906_, new_n5887_ );
or   ( new_n5908_, new_n5905_, new_n5888_ );
and  ( new_n5909_, new_n5908_, new_n5907_ );
nor  ( new_n5910_, new_n5909_, new_n5871_ );
or   ( new_n5911_, new_n5604_, new_n319_ );
or   ( new_n5912_, new_n5606_, new_n333_ );
and  ( new_n5913_, new_n5912_, new_n5911_ );
xor  ( new_n5914_, new_n5913_, new_n5205_ );
xor  ( new_n5915_, RIbb2df90_49, RIbb2e008_48 );
xor  ( new_n5916_, RIbb2e008_48, new_n5594_ );
nor  ( new_n5917_, new_n5916_, new_n5915_ );
and  ( new_n5918_, new_n5917_, RIbb2d810_65 );
xor  ( new_n5919_, new_n5918_, new_n5597_ );
nand ( new_n5920_, new_n5919_, new_n5914_ );
nor  ( new_n5921_, new_n5919_, new_n5914_ );
or   ( new_n5922_, new_n5207_, new_n285_ );
or   ( new_n5923_, new_n5209_, new_n313_ );
and  ( new_n5924_, new_n5923_, new_n5922_ );
xor  ( new_n5925_, new_n5924_, new_n4708_ );
or   ( new_n5926_, new_n5925_, new_n5921_ );
and  ( new_n5927_, new_n5926_, new_n5920_ );
or   ( new_n5928_, new_n4709_, new_n301_ );
or   ( new_n5929_, new_n4711_, new_n279_ );
and  ( new_n5930_, new_n5929_, new_n5928_ );
xor  ( new_n5931_, new_n5930_, new_n4295_ );
or   ( new_n5932_, new_n4302_, new_n270_ );
or   ( new_n5933_, new_n4304_, new_n294_ );
and  ( new_n5934_, new_n5933_, new_n5932_ );
xor  ( new_n5935_, new_n5934_, new_n3895_ );
or   ( new_n5936_, new_n5935_, new_n5931_ );
and  ( new_n5937_, new_n5935_, new_n5931_ );
or   ( new_n5938_, new_n3896_, new_n348_ );
or   ( new_n5939_, new_n3898_, new_n264_ );
and  ( new_n5940_, new_n5939_, new_n5938_ );
xor  ( new_n5941_, new_n5940_, new_n3460_ );
or   ( new_n5942_, new_n5941_, new_n5937_ );
and  ( new_n5943_, new_n5942_, new_n5936_ );
nor  ( new_n5944_, new_n5943_, new_n5927_ );
and  ( new_n5945_, new_n5943_, new_n5927_ );
or   ( new_n5946_, new_n3461_, new_n443_ );
or   ( new_n5947_, new_n3463_, new_n419_ );
and  ( new_n5948_, new_n5947_, new_n5946_ );
xor  ( new_n5949_, new_n5948_, new_n3116_ );
or   ( new_n5950_, new_n3117_, new_n515_ );
or   ( new_n5951_, new_n3119_, new_n509_ );
and  ( new_n5952_, new_n5951_, new_n5950_ );
xor  ( new_n5953_, new_n5952_, new_n2800_ );
nor  ( new_n5954_, new_n5953_, new_n5949_ );
and  ( new_n5955_, new_n5953_, new_n5949_ );
or   ( new_n5956_, new_n2807_, new_n805_ );
or   ( new_n5957_, new_n2809_, new_n775_ );
and  ( new_n5958_, new_n5957_, new_n5956_ );
xor  ( new_n5959_, new_n5958_, new_n2424_ );
nor  ( new_n5960_, new_n5959_, new_n5955_ );
nor  ( new_n5961_, new_n5960_, new_n5954_ );
nor  ( new_n5962_, new_n5961_, new_n5945_ );
nor  ( new_n5963_, new_n5962_, new_n5944_ );
and  ( new_n5964_, new_n5909_, new_n5871_ );
nor  ( new_n5965_, new_n5964_, new_n5963_ );
nor  ( new_n5966_, new_n5965_, new_n5910_ );
not  ( new_n5967_, new_n5966_ );
or   ( new_n5968_, new_n5967_, new_n5819_ );
and  ( new_n5969_, new_n5967_, new_n5819_ );
xor  ( new_n5970_, new_n5621_, new_n5617_ );
xor  ( new_n5971_, new_n5970_, new_n5627_ );
xor  ( new_n5972_, new_n5601_, new_n5597_ );
xor  ( new_n5973_, new_n5972_, new_n5609_ );
and  ( new_n5974_, new_n5973_, new_n5971_ );
or   ( new_n5975_, new_n5973_, new_n5971_ );
xor  ( new_n5976_, new_n5585_, new_n5581_ );
xor  ( new_n5977_, new_n5976_, new_n5591_ );
and  ( new_n5978_, new_n5977_, new_n5975_ );
or   ( new_n5979_, new_n5978_, new_n5974_ );
or   ( new_n5980_, new_n5899_, new_n260_ );
xnor ( new_n5981_, new_n5551_, new_n5547_ );
xor  ( new_n5982_, new_n5981_, new_n5557_ );
nand ( new_n5983_, new_n5982_, new_n5980_ );
or   ( new_n5984_, new_n5982_, new_n5980_ );
xor  ( new_n5985_, new_n5567_, new_n5563_ );
xnor ( new_n5986_, new_n5985_, new_n5574_ );
nand ( new_n5987_, new_n5986_, new_n5984_ );
and  ( new_n5988_, new_n5987_, new_n5983_ );
nand ( new_n5989_, new_n5988_, new_n5979_ );
nor  ( new_n5990_, new_n5988_, new_n5979_ );
xnor ( new_n5991_, new_n5657_, new_n5653_ );
xor  ( new_n5992_, new_n5991_, new_n5663_ );
xnor ( new_n5993_, new_n5641_, new_n5637_ );
xor  ( new_n5994_, new_n5993_, new_n5647_ );
nor  ( new_n5995_, new_n5994_, new_n5992_ );
and  ( new_n5996_, new_n5994_, new_n5992_ );
xor  ( new_n5997_, new_n5675_, new_n5671_ );
xnor ( new_n5998_, new_n5997_, new_n5681_ );
nor  ( new_n5999_, new_n5998_, new_n5996_ );
nor  ( new_n6000_, new_n5999_, new_n5995_ );
or   ( new_n6001_, new_n6000_, new_n5990_ );
and  ( new_n6002_, new_n6001_, new_n5989_ );
or   ( new_n6003_, new_n6002_, new_n5969_ );
and  ( new_n6004_, new_n6003_, new_n5968_ );
or   ( new_n6005_, new_n6004_, new_n5809_ );
and  ( new_n6006_, new_n6004_, new_n5809_ );
xor  ( new_n6007_, new_n5737_, new_n5735_ );
xor  ( new_n6008_, new_n6007_, new_n5741_ );
xnor ( new_n6009_, new_n5723_, new_n5721_ );
xor  ( new_n6010_, new_n6009_, new_n5727_ );
nor  ( new_n6011_, new_n6010_, new_n6008_ );
and  ( new_n6012_, new_n6010_, new_n6008_ );
xnor ( new_n6013_, new_n5611_, new_n5593_ );
xor  ( new_n6014_, new_n6013_, new_n5629_ );
xnor ( new_n6015_, new_n5665_, new_n5649_ );
xor  ( new_n6016_, new_n6015_, new_n5683_ );
nor  ( new_n6017_, new_n6016_, new_n6014_ );
and  ( new_n6018_, new_n6016_, new_n6014_ );
xor  ( new_n6019_, new_n5576_, new_n5559_ );
nor  ( new_n6020_, new_n6019_, new_n6018_ );
nor  ( new_n6021_, new_n6020_, new_n6017_ );
nor  ( new_n6022_, new_n6021_, new_n6012_ );
nor  ( new_n6023_, new_n6022_, new_n6011_ );
or   ( new_n6024_, new_n6023_, new_n6006_ );
and  ( new_n6025_, new_n6024_, new_n6005_ );
or   ( new_n6026_, new_n6025_, new_n5803_ );
and  ( new_n6027_, new_n6026_, new_n5802_ );
xor  ( new_n6028_, new_n5509_, new_n5324_ );
xor  ( new_n6029_, new_n6028_, new_n5521_ );
or   ( new_n6030_, new_n6029_, new_n6027_ );
and  ( new_n6031_, new_n6029_, new_n6027_ );
xnor ( new_n6032_, new_n5774_, new_n5764_ );
xor  ( new_n6033_, new_n6032_, new_n5778_ );
or   ( new_n6034_, new_n6033_, new_n6031_ );
and  ( new_n6035_, new_n6034_, new_n6030_ );
xor  ( new_n6036_, new_n5780_, new_n5543_ );
xor  ( new_n6037_, new_n6036_, new_n5784_ );
nor  ( new_n6038_, new_n6037_, new_n6035_ );
xor  ( new_n6039_, new_n5786_, new_n5541_ );
and  ( new_n6040_, new_n6039_, new_n6038_ );
xor  ( new_n6041_, new_n6029_, new_n6027_ );
xor  ( new_n6042_, new_n6041_, new_n6033_ );
xor  ( new_n6043_, new_n5966_, new_n5819_ );
xor  ( new_n6044_, new_n6043_, new_n6002_ );
xnor ( new_n6045_, new_n6010_, new_n6008_ );
xor  ( new_n6046_, new_n6045_, new_n6021_ );
or   ( new_n6047_, new_n6046_, new_n6044_ );
and  ( new_n6048_, new_n6046_, new_n6044_ );
xor  ( new_n6049_, new_n5808_, new_n5806_ );
or   ( new_n6050_, new_n6049_, new_n6048_ );
and  ( new_n6051_, new_n6050_, new_n6047_ );
xnor ( new_n6052_, new_n5795_, new_n5793_ );
xor  ( new_n6053_, new_n6052_, new_n5799_ );
and  ( new_n6054_, new_n6053_, new_n6051_ );
or   ( new_n6055_, new_n6053_, new_n6051_ );
xor  ( new_n6056_, new_n5909_, new_n5871_ );
xnor ( new_n6057_, new_n6056_, new_n5963_ );
xnor ( new_n6058_, new_n5988_, new_n5979_ );
xnor ( new_n6059_, new_n6058_, new_n6000_ );
or   ( new_n6060_, new_n6059_, new_n6057_ );
xnor ( new_n6061_, new_n5935_, new_n5931_ );
xor  ( new_n6062_, new_n6061_, new_n5941_ );
xnor ( new_n6063_, new_n5919_, new_n5914_ );
xor  ( new_n6064_, new_n6063_, new_n5925_ );
or   ( new_n6065_, new_n6064_, new_n6062_ );
and  ( new_n6066_, new_n6064_, new_n6062_ );
xor  ( new_n6067_, new_n5953_, new_n5949_ );
xnor ( new_n6068_, new_n6067_, new_n5959_ );
or   ( new_n6069_, new_n6068_, new_n6066_ );
and  ( new_n6070_, new_n6069_, new_n6065_ );
xnor ( new_n6071_, new_n5879_, new_n5875_ );
xor  ( new_n6072_, new_n6071_, new_n5885_ );
xnor ( new_n6073_, new_n5896_, new_n5892_ );
xor  ( new_n6074_, new_n6073_, new_n5903_ );
or   ( new_n6075_, new_n6074_, new_n6072_ );
and  ( new_n6076_, new_n6074_, new_n6072_ );
or   ( new_n6077_, new_n6076_, new_n5888_ );
and  ( new_n6078_, new_n6077_, new_n6075_ );
nor  ( new_n6079_, new_n6078_, new_n6070_ );
nand ( new_n6080_, new_n6078_, new_n6070_ );
xnor ( new_n6081_, new_n5843_, new_n5839_ );
xor  ( new_n6082_, new_n6081_, new_n5849_ );
xnor ( new_n6083_, new_n5827_, new_n5823_ );
xor  ( new_n6084_, new_n6083_, new_n5833_ );
nor  ( new_n6085_, new_n6084_, new_n6082_ );
and  ( new_n6086_, new_n6084_, new_n6082_ );
xor  ( new_n6087_, new_n5861_, new_n5857_ );
xnor ( new_n6088_, new_n6087_, new_n5867_ );
nor  ( new_n6089_, new_n6088_, new_n6086_ );
nor  ( new_n6090_, new_n6089_, new_n6085_ );
not  ( new_n6091_, new_n6090_ );
and  ( new_n6092_, new_n6091_, new_n6080_ );
or   ( new_n6093_, new_n6092_, new_n6079_ );
or   ( new_n6094_, new_n1844_, new_n1523_ );
or   ( new_n6095_, new_n1846_, new_n1525_ );
and  ( new_n6096_, new_n6095_, new_n6094_ );
xor  ( new_n6097_, new_n6096_, new_n1586_ );
or   ( new_n6098_, new_n1593_, new_n1899_ );
or   ( new_n6099_, new_n1595_, new_n1754_ );
and  ( new_n6100_, new_n6099_, new_n6098_ );
xor  ( new_n6101_, new_n6100_, new_n1358_ );
or   ( new_n6102_, new_n6101_, new_n6097_ );
and  ( new_n6103_, new_n6101_, new_n6097_ );
or   ( new_n6104_, new_n1364_, new_n2178_ );
or   ( new_n6105_, new_n1366_, new_n2057_ );
and  ( new_n6106_, new_n6105_, new_n6104_ );
xor  ( new_n6107_, new_n6106_, new_n1129_ );
or   ( new_n6108_, new_n6107_, new_n6103_ );
and  ( new_n6109_, new_n6108_, new_n6102_ );
or   ( new_n6110_, new_n2807_, new_n886_ );
or   ( new_n6111_, new_n2809_, new_n805_ );
and  ( new_n6112_, new_n6111_, new_n6110_ );
xor  ( new_n6113_, new_n6112_, new_n2424_ );
or   ( new_n6114_, new_n2425_, new_n1168_ );
or   ( new_n6115_, new_n2427_, new_n986_ );
and  ( new_n6116_, new_n6115_, new_n6114_ );
xor  ( new_n6117_, new_n6116_, new_n2121_ );
or   ( new_n6118_, new_n6117_, new_n6113_ );
and  ( new_n6119_, new_n6117_, new_n6113_ );
or   ( new_n6120_, new_n2122_, new_n1318_ );
or   ( new_n6121_, new_n2124_, new_n1213_ );
and  ( new_n6122_, new_n6121_, new_n6120_ );
xor  ( new_n6123_, new_n6122_, new_n1843_ );
or   ( new_n6124_, new_n6123_, new_n6119_ );
and  ( new_n6125_, new_n6124_, new_n6118_ );
or   ( new_n6126_, new_n6125_, new_n6109_ );
and  ( new_n6127_, new_n6125_, new_n6109_ );
or   ( new_n6128_, new_n1135_, new_n2475_ );
or   ( new_n6129_, new_n1137_, new_n2291_ );
and  ( new_n6130_, new_n6129_, new_n6128_ );
xor  ( new_n6131_, new_n6130_, new_n896_ );
or   ( new_n6132_, new_n897_, new_n2751_ );
or   ( new_n6133_, new_n899_, new_n2646_ );
and  ( new_n6134_, new_n6133_, new_n6132_ );
xor  ( new_n6135_, new_n6134_, new_n748_ );
nor  ( new_n6136_, new_n6135_, new_n6131_ );
and  ( new_n6137_, new_n6135_, new_n6131_ );
or   ( new_n6138_, new_n755_, new_n3178_ );
or   ( new_n6139_, new_n757_, new_n2981_ );
and  ( new_n6140_, new_n6139_, new_n6138_ );
xor  ( new_n6141_, new_n6140_, new_n523_ );
nor  ( new_n6142_, new_n6141_, new_n6137_ );
nor  ( new_n6143_, new_n6142_, new_n6136_ );
or   ( new_n6144_, new_n6143_, new_n6127_ );
and  ( new_n6145_, new_n6144_, new_n6126_ );
or   ( new_n6146_, new_n5207_, new_n279_ );
or   ( new_n6147_, new_n5209_, new_n285_ );
and  ( new_n6148_, new_n6147_, new_n6146_ );
xor  ( new_n6149_, new_n6148_, new_n4708_ );
or   ( new_n6150_, new_n4709_, new_n294_ );
or   ( new_n6151_, new_n4711_, new_n301_ );
and  ( new_n6152_, new_n6151_, new_n6150_ );
xor  ( new_n6153_, new_n6152_, new_n4295_ );
nor  ( new_n6154_, new_n6153_, new_n6149_ );
nand ( new_n6155_, new_n6153_, new_n6149_ );
or   ( new_n6156_, new_n4302_, new_n264_ );
or   ( new_n6157_, new_n4304_, new_n270_ );
and  ( new_n6158_, new_n6157_, new_n6156_ );
xor  ( new_n6159_, new_n6158_, new_n3895_ );
not  ( new_n6160_, new_n6159_ );
and  ( new_n6161_, new_n6160_, new_n6155_ );
or   ( new_n6162_, new_n6161_, new_n6154_ );
not  ( new_n6163_, RIbb2df90_49 );
and  ( new_n6164_, RIbb2dea0_51, RIbb2df18_50 );
nor  ( new_n6165_, new_n6164_, new_n6163_ );
not  ( new_n6166_, new_n6165_ );
or   ( new_n6167_, new_n5604_, new_n313_ );
or   ( new_n6168_, new_n5606_, new_n319_ );
and  ( new_n6169_, new_n6168_, new_n6167_ );
xor  ( new_n6170_, new_n6169_, new_n5206_ );
nand ( new_n6171_, new_n6170_, new_n6166_ );
or   ( new_n6172_, new_n6170_, new_n6166_ );
not  ( new_n6173_, new_n5917_ );
or   ( new_n6174_, new_n6173_, new_n333_ );
not  ( new_n6175_, new_n5915_ );
or   ( new_n6176_, new_n6175_, new_n339_ );
and  ( new_n6177_, new_n6176_, new_n6174_ );
xor  ( new_n6178_, new_n6177_, new_n5597_ );
nand ( new_n6179_, new_n6178_, new_n6172_ );
and  ( new_n6180_, new_n6179_, new_n6171_ );
nand ( new_n6181_, new_n6180_, new_n6162_ );
nor  ( new_n6182_, new_n6180_, new_n6162_ );
or   ( new_n6183_, new_n3896_, new_n419_ );
or   ( new_n6184_, new_n3898_, new_n348_ );
and  ( new_n6185_, new_n6184_, new_n6183_ );
xor  ( new_n6186_, new_n6185_, new_n3460_ );
or   ( new_n6187_, new_n3461_, new_n509_ );
or   ( new_n6188_, new_n3463_, new_n443_ );
and  ( new_n6189_, new_n6188_, new_n6187_ );
xor  ( new_n6190_, new_n6189_, new_n3116_ );
or   ( new_n6191_, new_n6190_, new_n6186_ );
and  ( new_n6192_, new_n6190_, new_n6186_ );
or   ( new_n6193_, new_n3117_, new_n775_ );
or   ( new_n6194_, new_n3119_, new_n515_ );
and  ( new_n6195_, new_n6194_, new_n6193_ );
xor  ( new_n6196_, new_n6195_, new_n2800_ );
or   ( new_n6197_, new_n6196_, new_n6192_ );
and  ( new_n6198_, new_n6197_, new_n6191_ );
or   ( new_n6199_, new_n6198_, new_n6182_ );
and  ( new_n6200_, new_n6199_, new_n6181_ );
or   ( new_n6201_, new_n6200_, new_n6145_ );
and  ( new_n6202_, new_n6200_, new_n6145_ );
or   ( new_n6203_, new_n524_, new_n3696_ );
or   ( new_n6204_, new_n526_, new_n3306_ );
and  ( new_n6205_, new_n6204_, new_n6203_ );
xor  ( new_n6206_, new_n6205_, new_n403_ );
or   ( new_n6207_, new_n409_, new_n3820_ );
or   ( new_n6208_, new_n411_, new_n3694_ );
and  ( new_n6209_, new_n6208_, new_n6207_ );
xor  ( new_n6210_, new_n6209_, new_n328_ );
nor  ( new_n6211_, new_n6210_, new_n6206_ );
and  ( new_n6212_, new_n6210_, new_n6206_ );
or   ( new_n6213_, new_n337_, new_n4267_ );
or   ( new_n6214_, new_n340_, new_n4069_ );
and  ( new_n6215_, new_n6214_, new_n6213_ );
xor  ( new_n6216_, new_n6215_, new_n332_ );
nor  ( new_n6217_, new_n6216_, new_n6212_ );
nor  ( new_n6218_, new_n6217_, new_n6211_ );
not  ( new_n6219_, RIbb2c208_112 );
or   ( new_n6220_, new_n268_, new_n6219_ );
or   ( new_n6221_, new_n271_, new_n5899_ );
and  ( new_n6222_, new_n6221_, new_n6220_ );
xor  ( new_n6223_, new_n6222_, new_n263_ );
and  ( new_n6224_, RIbb2c190_113, RIbb2f610_1 );
and  ( new_n6225_, new_n6224_, new_n6223_ );
or   ( new_n6226_, new_n317_, new_n4995_ );
or   ( new_n6227_, new_n320_, new_n4603_ );
and  ( new_n6228_, new_n6227_, new_n6226_ );
xor  ( new_n6229_, new_n6228_, new_n312_ );
or   ( new_n6230_, new_n283_, new_n5171_ );
or   ( new_n6231_, new_n286_, new_n4859_ );
and  ( new_n6232_, new_n6231_, new_n6230_ );
xor  ( new_n6233_, new_n6232_, new_n278_ );
nor  ( new_n6234_, new_n6233_, new_n6229_ );
and  ( new_n6235_, new_n6233_, new_n6229_ );
or   ( new_n6236_, new_n299_, new_n5570_ );
or   ( new_n6237_, new_n302_, new_n5428_ );
and  ( new_n6238_, new_n6237_, new_n6236_ );
xor  ( new_n6239_, new_n6238_, new_n293_ );
nor  ( new_n6240_, new_n6239_, new_n6235_ );
nor  ( new_n6241_, new_n6240_, new_n6234_ );
and  ( new_n6242_, new_n6241_, new_n6225_ );
nor  ( new_n6243_, new_n6242_, new_n6218_ );
nor  ( new_n6244_, new_n6241_, new_n6225_ );
nor  ( new_n6245_, new_n6244_, new_n6243_ );
or   ( new_n6246_, new_n6245_, new_n6202_ );
and  ( new_n6247_, new_n6246_, new_n6201_ );
nand ( new_n6248_, new_n6247_, new_n6093_ );
nor  ( new_n6249_, new_n6247_, new_n6093_ );
xnor ( new_n6250_, new_n5994_, new_n5992_ );
xor  ( new_n6251_, new_n6250_, new_n5998_ );
xor  ( new_n6252_, new_n5973_, new_n5971_ );
xor  ( new_n6253_, new_n6252_, new_n5977_ );
and  ( new_n6254_, new_n6253_, new_n6251_ );
nor  ( new_n6255_, new_n6253_, new_n6251_ );
xor  ( new_n6256_, new_n5982_, new_n5980_ );
xor  ( new_n6257_, new_n6256_, new_n5986_ );
nor  ( new_n6258_, new_n6257_, new_n6255_ );
nor  ( new_n6259_, new_n6258_, new_n6254_ );
or   ( new_n6260_, new_n6259_, new_n6249_ );
and  ( new_n6261_, new_n6260_, new_n6248_ );
nor  ( new_n6262_, new_n6261_, new_n6060_ );
and  ( new_n6263_, new_n6261_, new_n6060_ );
xor  ( new_n6264_, new_n6016_, new_n6014_ );
xor  ( new_n6265_, new_n6264_, new_n6019_ );
not  ( new_n6266_, new_n5888_ );
xor  ( new_n6267_, new_n5905_, new_n6266_ );
xor  ( new_n6268_, new_n6267_, new_n5887_ );
xnor ( new_n6269_, new_n5851_, new_n5835_ );
xor  ( new_n6270_, new_n6269_, new_n5869_ );
or   ( new_n6271_, new_n6270_, new_n6268_ );
and  ( new_n6272_, new_n6270_, new_n6268_ );
xor  ( new_n6273_, new_n5943_, new_n5927_ );
xnor ( new_n6274_, new_n6273_, new_n5961_ );
or   ( new_n6275_, new_n6274_, new_n6272_ );
and  ( new_n6276_, new_n6275_, new_n6271_ );
nor  ( new_n6277_, new_n6276_, new_n6265_ );
and  ( new_n6278_, new_n6276_, new_n6265_ );
xor  ( new_n6279_, new_n5813_, new_n5811_ );
xor  ( new_n6280_, new_n6279_, new_n5817_ );
nor  ( new_n6281_, new_n6280_, new_n6278_ );
nor  ( new_n6282_, new_n6281_, new_n6277_ );
nor  ( new_n6283_, new_n6282_, new_n6263_ );
nor  ( new_n6284_, new_n6283_, new_n6262_ );
not  ( new_n6285_, new_n6284_ );
and  ( new_n6286_, new_n6285_, new_n6055_ );
or   ( new_n6287_, new_n6286_, new_n6054_ );
xnor ( new_n6288_, new_n5749_, new_n5731_ );
xor  ( new_n6289_, new_n6288_, new_n5762_ );
nand ( new_n6290_, new_n6289_, new_n6287_ );
nor  ( new_n6291_, new_n6289_, new_n6287_ );
xor  ( new_n6292_, new_n5801_, new_n5791_ );
xor  ( new_n6293_, new_n6292_, new_n6025_ );
or   ( new_n6294_, new_n6293_, new_n6291_ );
and  ( new_n6295_, new_n6294_, new_n6290_ );
nor  ( new_n6296_, new_n6295_, new_n6042_ );
xor  ( new_n6297_, new_n6037_, new_n6035_ );
and  ( new_n6298_, new_n6297_, new_n6296_ );
xor  ( new_n6299_, new_n6289_, new_n6287_ );
xor  ( new_n6300_, new_n6299_, new_n6293_ );
xnor ( new_n6301_, new_n6276_, new_n6265_ );
xor  ( new_n6302_, new_n6301_, new_n6280_ );
xnor ( new_n6303_, new_n6247_, new_n6093_ );
xor  ( new_n6304_, new_n6303_, new_n6259_ );
nor  ( new_n6305_, new_n6304_, new_n6302_ );
nand ( new_n6306_, new_n6304_, new_n6302_ );
xnor ( new_n6307_, new_n6059_, new_n6057_ );
and  ( new_n6308_, new_n6307_, new_n6306_ );
or   ( new_n6309_, new_n6308_, new_n6305_ );
xnor ( new_n6310_, new_n6046_, new_n6044_ );
xor  ( new_n6311_, new_n6310_, new_n6049_ );
nor  ( new_n6312_, new_n6311_, new_n6309_ );
nand ( new_n6313_, new_n6311_, new_n6309_ );
xor  ( new_n6314_, new_n6078_, new_n6070_ );
xor  ( new_n6315_, new_n6314_, new_n6091_ );
xnor ( new_n6316_, new_n6200_, new_n6145_ );
xnor ( new_n6317_, new_n6316_, new_n6245_ );
nand ( new_n6318_, new_n6317_, new_n6315_ );
xnor ( new_n6319_, new_n6253_, new_n6251_ );
xor  ( new_n6320_, new_n6319_, new_n6257_ );
xnor ( new_n6321_, new_n6270_, new_n6268_ );
xor  ( new_n6322_, new_n6321_, new_n6274_ );
nand ( new_n6323_, new_n6322_, new_n6320_ );
nor  ( new_n6324_, new_n6322_, new_n6320_ );
xor  ( new_n6325_, new_n6180_, new_n6162_ );
xor  ( new_n6326_, new_n6325_, new_n6198_ );
xor  ( new_n6327_, new_n6241_, new_n6225_ );
xor  ( new_n6328_, new_n6327_, new_n6218_ );
and  ( new_n6329_, new_n6328_, new_n6326_ );
nor  ( new_n6330_, new_n6328_, new_n6326_ );
xor  ( new_n6331_, new_n6125_, new_n6109_ );
xnor ( new_n6332_, new_n6331_, new_n6143_ );
nor  ( new_n6333_, new_n6332_, new_n6330_ );
nor  ( new_n6334_, new_n6333_, new_n6329_ );
or   ( new_n6335_, new_n6334_, new_n6324_ );
and  ( new_n6336_, new_n6335_, new_n6323_ );
nor  ( new_n6337_, new_n6336_, new_n6318_ );
and  ( new_n6338_, new_n6336_, new_n6318_ );
xor  ( new_n6339_, new_n6190_, new_n6186_ );
xor  ( new_n6340_, new_n6339_, new_n6196_ );
xor  ( new_n6341_, new_n6170_, new_n6166_ );
xor  ( new_n6342_, new_n6341_, new_n6178_ );
nand ( new_n6343_, new_n6342_, new_n6340_ );
nor  ( new_n6344_, new_n6342_, new_n6340_ );
xor  ( new_n6345_, new_n6153_, new_n6149_ );
xor  ( new_n6346_, new_n6345_, new_n6160_ );
or   ( new_n6347_, new_n6346_, new_n6344_ );
and  ( new_n6348_, new_n6347_, new_n6343_ );
xnor ( new_n6349_, new_n6210_, new_n6206_ );
xor  ( new_n6350_, new_n6349_, new_n6216_ );
xnor ( new_n6351_, new_n6233_, new_n6229_ );
xor  ( new_n6352_, new_n6351_, new_n6239_ );
or   ( new_n6353_, new_n6352_, new_n6350_ );
nand ( new_n6354_, new_n6352_, new_n6350_ );
xor  ( new_n6355_, new_n6224_, new_n6223_ );
nand ( new_n6356_, new_n6355_, new_n6354_ );
and  ( new_n6357_, new_n6356_, new_n6353_ );
nor  ( new_n6358_, new_n6357_, new_n6348_ );
nand ( new_n6359_, new_n6357_, new_n6348_ );
xnor ( new_n6360_, new_n6117_, new_n6113_ );
xor  ( new_n6361_, new_n6360_, new_n6123_ );
xnor ( new_n6362_, new_n6101_, new_n6097_ );
xor  ( new_n6363_, new_n6362_, new_n6107_ );
nor  ( new_n6364_, new_n6363_, new_n6361_ );
and  ( new_n6365_, new_n6363_, new_n6361_ );
xor  ( new_n6366_, new_n6135_, new_n6131_ );
xnor ( new_n6367_, new_n6366_, new_n6141_ );
nor  ( new_n6368_, new_n6367_, new_n6365_ );
nor  ( new_n6369_, new_n6368_, new_n6364_ );
not  ( new_n6370_, new_n6369_ );
and  ( new_n6371_, new_n6370_, new_n6359_ );
or   ( new_n6372_, new_n6371_, new_n6358_ );
or   ( new_n6373_, new_n1135_, new_n2646_ );
or   ( new_n6374_, new_n1137_, new_n2475_ );
and  ( new_n6375_, new_n6374_, new_n6373_ );
xor  ( new_n6376_, new_n6375_, new_n896_ );
or   ( new_n6377_, new_n897_, new_n2981_ );
or   ( new_n6378_, new_n899_, new_n2751_ );
and  ( new_n6379_, new_n6378_, new_n6377_ );
xor  ( new_n6380_, new_n6379_, new_n748_ );
or   ( new_n6381_, new_n6380_, new_n6376_ );
and  ( new_n6382_, new_n6380_, new_n6376_ );
or   ( new_n6383_, new_n755_, new_n3306_ );
or   ( new_n6384_, new_n757_, new_n3178_ );
and  ( new_n6385_, new_n6384_, new_n6383_ );
xor  ( new_n6386_, new_n6385_, new_n523_ );
or   ( new_n6387_, new_n6386_, new_n6382_ );
and  ( new_n6388_, new_n6387_, new_n6381_ );
or   ( new_n6389_, new_n1844_, new_n1754_ );
or   ( new_n6390_, new_n1846_, new_n1523_ );
and  ( new_n6391_, new_n6390_, new_n6389_ );
xor  ( new_n6392_, new_n6391_, new_n1586_ );
or   ( new_n6393_, new_n1593_, new_n2057_ );
or   ( new_n6394_, new_n1595_, new_n1899_ );
and  ( new_n6395_, new_n6394_, new_n6393_ );
xor  ( new_n6396_, new_n6395_, new_n1358_ );
or   ( new_n6397_, new_n6396_, new_n6392_ );
and  ( new_n6398_, new_n6396_, new_n6392_ );
or   ( new_n6399_, new_n1364_, new_n2291_ );
or   ( new_n6400_, new_n1366_, new_n2178_ );
and  ( new_n6401_, new_n6400_, new_n6399_ );
xor  ( new_n6402_, new_n6401_, new_n1129_ );
or   ( new_n6403_, new_n6402_, new_n6398_ );
and  ( new_n6404_, new_n6403_, new_n6397_ );
or   ( new_n6405_, new_n6404_, new_n6388_ );
and  ( new_n6406_, new_n6404_, new_n6388_ );
or   ( new_n6407_, new_n2807_, new_n986_ );
or   ( new_n6408_, new_n2809_, new_n886_ );
and  ( new_n6409_, new_n6408_, new_n6407_ );
xor  ( new_n6410_, new_n6409_, new_n2424_ );
or   ( new_n6411_, new_n2425_, new_n1213_ );
or   ( new_n6412_, new_n2427_, new_n1168_ );
and  ( new_n6413_, new_n6412_, new_n6411_ );
xor  ( new_n6414_, new_n6413_, new_n2121_ );
nor  ( new_n6415_, new_n6414_, new_n6410_ );
and  ( new_n6416_, new_n6414_, new_n6410_ );
or   ( new_n6417_, new_n2122_, new_n1525_ );
or   ( new_n6418_, new_n2124_, new_n1318_ );
and  ( new_n6419_, new_n6418_, new_n6417_ );
xor  ( new_n6420_, new_n6419_, new_n1843_ );
nor  ( new_n6421_, new_n6420_, new_n6416_ );
nor  ( new_n6422_, new_n6421_, new_n6415_ );
or   ( new_n6423_, new_n6422_, new_n6406_ );
and  ( new_n6424_, new_n6423_, new_n6405_ );
not  ( new_n6425_, RIbb2c190_113 );
or   ( new_n6426_, new_n268_, new_n6425_ );
or   ( new_n6427_, new_n271_, new_n6219_ );
and  ( new_n6428_, new_n6427_, new_n6426_ );
xor  ( new_n6429_, new_n6428_, new_n263_ );
and  ( new_n6430_, RIbb2c118_114, RIbb2f610_1 );
or   ( new_n6431_, new_n6430_, new_n6429_ );
or   ( new_n6432_, new_n524_, new_n3694_ );
or   ( new_n6433_, new_n526_, new_n3696_ );
and  ( new_n6434_, new_n6433_, new_n6432_ );
xor  ( new_n6435_, new_n6434_, new_n403_ );
or   ( new_n6436_, new_n409_, new_n4069_ );
or   ( new_n6437_, new_n411_, new_n3820_ );
and  ( new_n6438_, new_n6437_, new_n6436_ );
xor  ( new_n6439_, new_n6438_, new_n328_ );
or   ( new_n6440_, new_n6439_, new_n6435_ );
and  ( new_n6441_, new_n6439_, new_n6435_ );
or   ( new_n6442_, new_n337_, new_n4603_ );
or   ( new_n6443_, new_n340_, new_n4267_ );
and  ( new_n6444_, new_n6443_, new_n6442_ );
xor  ( new_n6445_, new_n6444_, new_n332_ );
or   ( new_n6446_, new_n6445_, new_n6441_ );
and  ( new_n6447_, new_n6446_, new_n6440_ );
or   ( new_n6448_, new_n6447_, new_n6431_ );
and  ( new_n6449_, new_n6447_, new_n6431_ );
or   ( new_n6450_, new_n317_, new_n4859_ );
or   ( new_n6451_, new_n320_, new_n4995_ );
and  ( new_n6452_, new_n6451_, new_n6450_ );
xor  ( new_n6453_, new_n6452_, new_n312_ );
or   ( new_n6454_, new_n283_, new_n5428_ );
or   ( new_n6455_, new_n286_, new_n5171_ );
and  ( new_n6456_, new_n6455_, new_n6454_ );
xor  ( new_n6457_, new_n6456_, new_n278_ );
nor  ( new_n6458_, new_n6457_, new_n6453_ );
and  ( new_n6459_, new_n6457_, new_n6453_ );
or   ( new_n6460_, new_n299_, new_n5899_ );
or   ( new_n6461_, new_n302_, new_n5570_ );
and  ( new_n6462_, new_n6461_, new_n6460_ );
xor  ( new_n6463_, new_n6462_, new_n293_ );
nor  ( new_n6464_, new_n6463_, new_n6459_ );
nor  ( new_n6465_, new_n6464_, new_n6458_ );
or   ( new_n6466_, new_n6465_, new_n6449_ );
and  ( new_n6467_, new_n6466_, new_n6448_ );
or   ( new_n6468_, new_n6467_, new_n6424_ );
and  ( new_n6469_, new_n6467_, new_n6424_ );
or   ( new_n6470_, new_n5207_, new_n301_ );
or   ( new_n6471_, new_n5209_, new_n279_ );
and  ( new_n6472_, new_n6471_, new_n6470_ );
xor  ( new_n6473_, new_n6472_, new_n4708_ );
or   ( new_n6474_, new_n4709_, new_n270_ );
or   ( new_n6475_, new_n4711_, new_n294_ );
and  ( new_n6476_, new_n6475_, new_n6474_ );
xor  ( new_n6477_, new_n6476_, new_n4295_ );
or   ( new_n6478_, new_n6477_, new_n6473_ );
and  ( new_n6479_, new_n6477_, new_n6473_ );
or   ( new_n6480_, new_n4302_, new_n348_ );
or   ( new_n6481_, new_n4304_, new_n264_ );
and  ( new_n6482_, new_n6481_, new_n6480_ );
xor  ( new_n6483_, new_n6482_, new_n3895_ );
or   ( new_n6484_, new_n6483_, new_n6479_ );
and  ( new_n6485_, new_n6484_, new_n6478_ );
or   ( new_n6486_, new_n3896_, new_n443_ );
or   ( new_n6487_, new_n3898_, new_n419_ );
and  ( new_n6488_, new_n6487_, new_n6486_ );
xor  ( new_n6489_, new_n6488_, new_n3460_ );
or   ( new_n6490_, new_n3461_, new_n515_ );
or   ( new_n6491_, new_n3463_, new_n509_ );
and  ( new_n6492_, new_n6491_, new_n6490_ );
xor  ( new_n6493_, new_n6492_, new_n3116_ );
or   ( new_n6494_, new_n6493_, new_n6489_ );
and  ( new_n6495_, new_n6493_, new_n6489_ );
or   ( new_n6496_, new_n3117_, new_n805_ );
or   ( new_n6497_, new_n3119_, new_n775_ );
and  ( new_n6498_, new_n6497_, new_n6496_ );
xor  ( new_n6499_, new_n6498_, new_n2800_ );
or   ( new_n6500_, new_n6499_, new_n6495_ );
and  ( new_n6501_, new_n6500_, new_n6494_ );
nor  ( new_n6502_, new_n6501_, new_n6485_ );
and  ( new_n6503_, new_n6501_, new_n6485_ );
or   ( new_n6504_, new_n6173_, new_n319_ );
or   ( new_n6505_, new_n6175_, new_n333_ );
and  ( new_n6506_, new_n6505_, new_n6504_ );
xor  ( new_n6507_, new_n6506_, new_n5596_ );
xor  ( new_n6508_, RIbb2dea0_51, RIbb2df18_50 );
xor  ( new_n6509_, RIbb2df18_50, new_n6163_ );
nor  ( new_n6510_, new_n6509_, new_n6508_ );
and  ( new_n6511_, new_n6510_, RIbb2d810_65 );
xor  ( new_n6512_, new_n6511_, new_n6166_ );
and  ( new_n6513_, new_n6512_, new_n6507_ );
nor  ( new_n6514_, new_n6512_, new_n6507_ );
or   ( new_n6515_, new_n5604_, new_n285_ );
or   ( new_n6516_, new_n5606_, new_n313_ );
and  ( new_n6517_, new_n6516_, new_n6515_ );
xor  ( new_n6518_, new_n6517_, new_n5206_ );
nor  ( new_n6519_, new_n6518_, new_n6514_ );
nor  ( new_n6520_, new_n6519_, new_n6513_ );
nor  ( new_n6521_, new_n6520_, new_n6503_ );
nor  ( new_n6522_, new_n6521_, new_n6502_ );
or   ( new_n6523_, new_n6522_, new_n6469_ );
and  ( new_n6524_, new_n6523_, new_n6468_ );
and  ( new_n6525_, new_n6524_, new_n6372_ );
nor  ( new_n6526_, new_n6524_, new_n6372_ );
xnor ( new_n6527_, new_n6084_, new_n6082_ );
xor  ( new_n6528_, new_n6527_, new_n6088_ );
xnor ( new_n6529_, new_n6064_, new_n6062_ );
xor  ( new_n6530_, new_n6529_, new_n6068_ );
and  ( new_n6531_, new_n6530_, new_n6528_ );
nor  ( new_n6532_, new_n6530_, new_n6528_ );
xor  ( new_n6533_, new_n6074_, new_n6072_ );
xnor ( new_n6534_, new_n6533_, new_n6266_ );
nor  ( new_n6535_, new_n6534_, new_n6532_ );
nor  ( new_n6536_, new_n6535_, new_n6531_ );
nor  ( new_n6537_, new_n6536_, new_n6526_ );
nor  ( new_n6538_, new_n6537_, new_n6525_ );
nor  ( new_n6539_, new_n6538_, new_n6338_ );
nor  ( new_n6540_, new_n6539_, new_n6337_ );
not  ( new_n6541_, new_n6540_ );
and  ( new_n6542_, new_n6541_, new_n6313_ );
or   ( new_n6543_, new_n6542_, new_n6312_ );
xnor ( new_n6544_, new_n6004_, new_n5809_ );
xor  ( new_n6545_, new_n6544_, new_n6023_ );
nand ( new_n6546_, new_n6545_, new_n6543_ );
or   ( new_n6547_, new_n6545_, new_n6543_ );
xor  ( new_n6548_, new_n6053_, new_n6051_ );
xor  ( new_n6549_, new_n6548_, new_n6285_ );
nand ( new_n6550_, new_n6549_, new_n6547_ );
and  ( new_n6551_, new_n6550_, new_n6546_ );
nor  ( new_n6552_, new_n6551_, new_n6300_ );
xor  ( new_n6553_, new_n6295_, new_n6042_ );
and  ( new_n6554_, new_n6553_, new_n6552_ );
xnor ( new_n6555_, new_n6261_, new_n6060_ );
xor  ( new_n6556_, new_n6555_, new_n6282_ );
xnor ( new_n6557_, new_n6524_, new_n6372_ );
xor  ( new_n6558_, new_n6557_, new_n6536_ );
xnor ( new_n6559_, new_n6322_, new_n6320_ );
xor  ( new_n6560_, new_n6559_, new_n6334_ );
nor  ( new_n6561_, new_n6560_, new_n6558_ );
nand ( new_n6562_, new_n6560_, new_n6558_ );
xnor ( new_n6563_, new_n6317_, new_n6315_ );
and  ( new_n6564_, new_n6563_, new_n6562_ );
or   ( new_n6565_, new_n6564_, new_n6561_ );
xor  ( new_n6566_, new_n6304_, new_n6302_ );
xor  ( new_n6567_, new_n6566_, new_n6307_ );
nand ( new_n6568_, new_n6567_, new_n6565_ );
nor  ( new_n6569_, new_n6567_, new_n6565_ );
xor  ( new_n6570_, new_n6357_, new_n6348_ );
xor  ( new_n6571_, new_n6570_, new_n6370_ );
xnor ( new_n6572_, new_n6467_, new_n6424_ );
xnor ( new_n6573_, new_n6572_, new_n6522_ );
and  ( new_n6574_, new_n6573_, new_n6571_ );
xnor ( new_n6575_, new_n6363_, new_n6361_ );
xor  ( new_n6576_, new_n6575_, new_n6367_ );
xnor ( new_n6577_, new_n6342_, new_n6340_ );
xor  ( new_n6578_, new_n6577_, new_n6346_ );
or   ( new_n6579_, new_n6578_, new_n6576_ );
and  ( new_n6580_, new_n6578_, new_n6576_ );
xor  ( new_n6581_, new_n6352_, new_n6350_ );
xor  ( new_n6582_, new_n6581_, new_n6355_ );
or   ( new_n6583_, new_n6582_, new_n6580_ );
and  ( new_n6584_, new_n6583_, new_n6579_ );
or   ( new_n6585_, new_n299_, new_n6219_ );
or   ( new_n6586_, new_n302_, new_n5899_ );
and  ( new_n6587_, new_n6586_, new_n6585_ );
xor  ( new_n6588_, new_n6587_, new_n293_ );
not  ( new_n6589_, RIbb2c118_114 );
or   ( new_n6590_, new_n268_, new_n6589_ );
or   ( new_n6591_, new_n271_, new_n6425_ );
and  ( new_n6592_, new_n6591_, new_n6590_ );
xor  ( new_n6593_, new_n6592_, new_n263_ );
or   ( new_n6594_, new_n6593_, new_n6588_ );
and  ( new_n6595_, RIbb2c0a0_115, RIbb2f610_1 );
and  ( new_n6596_, new_n6593_, new_n6588_ );
or   ( new_n6597_, new_n6596_, new_n6595_ );
and  ( new_n6598_, new_n6597_, new_n6594_ );
or   ( new_n6599_, new_n755_, new_n3696_ );
or   ( new_n6600_, new_n757_, new_n3306_ );
and  ( new_n6601_, new_n6600_, new_n6599_ );
xor  ( new_n6602_, new_n6601_, new_n523_ );
or   ( new_n6603_, new_n524_, new_n3820_ );
or   ( new_n6604_, new_n526_, new_n3694_ );
and  ( new_n6605_, new_n6604_, new_n6603_ );
xor  ( new_n6606_, new_n6605_, new_n403_ );
or   ( new_n6607_, new_n6606_, new_n6602_ );
and  ( new_n6608_, new_n6606_, new_n6602_ );
or   ( new_n6609_, new_n409_, new_n4267_ );
or   ( new_n6610_, new_n411_, new_n4069_ );
and  ( new_n6611_, new_n6610_, new_n6609_ );
xor  ( new_n6612_, new_n6611_, new_n328_ );
or   ( new_n6613_, new_n6612_, new_n6608_ );
and  ( new_n6614_, new_n6613_, new_n6607_ );
or   ( new_n6615_, new_n6614_, new_n6598_ );
and  ( new_n6616_, new_n6614_, new_n6598_ );
or   ( new_n6617_, new_n337_, new_n4995_ );
or   ( new_n6618_, new_n340_, new_n4603_ );
and  ( new_n6619_, new_n6618_, new_n6617_ );
xor  ( new_n6620_, new_n6619_, new_n332_ );
or   ( new_n6621_, new_n317_, new_n5171_ );
or   ( new_n6622_, new_n320_, new_n4859_ );
and  ( new_n6623_, new_n6622_, new_n6621_ );
xor  ( new_n6624_, new_n6623_, new_n312_ );
nor  ( new_n6625_, new_n6624_, new_n6620_ );
and  ( new_n6626_, new_n6624_, new_n6620_ );
or   ( new_n6627_, new_n283_, new_n5570_ );
or   ( new_n6628_, new_n286_, new_n5428_ );
and  ( new_n6629_, new_n6628_, new_n6627_ );
xor  ( new_n6630_, new_n6629_, new_n278_ );
nor  ( new_n6631_, new_n6630_, new_n6626_ );
nor  ( new_n6632_, new_n6631_, new_n6625_ );
or   ( new_n6633_, new_n6632_, new_n6616_ );
and  ( new_n6634_, new_n6633_, new_n6615_ );
not  ( new_n6635_, RIbb2dea0_51 );
and  ( new_n6636_, RIbb2ddb0_53, RIbb2de28_52 );
nor  ( new_n6637_, new_n6636_, new_n6635_ );
not  ( new_n6638_, new_n6637_ );
or   ( new_n6639_, new_n6173_, new_n313_ );
or   ( new_n6640_, new_n6175_, new_n319_ );
and  ( new_n6641_, new_n6640_, new_n6639_ );
xor  ( new_n6642_, new_n6641_, new_n5597_ );
and  ( new_n6643_, new_n6642_, new_n6638_ );
or   ( new_n6644_, new_n6642_, new_n6638_ );
not  ( new_n6645_, new_n6510_ );
or   ( new_n6646_, new_n6645_, new_n333_ );
not  ( new_n6647_, new_n6508_ );
or   ( new_n6648_, new_n6647_, new_n339_ );
and  ( new_n6649_, new_n6648_, new_n6646_ );
xor  ( new_n6650_, new_n6649_, new_n6166_ );
and  ( new_n6651_, new_n6650_, new_n6644_ );
or   ( new_n6652_, new_n6651_, new_n6643_ );
or   ( new_n6653_, new_n5604_, new_n279_ );
or   ( new_n6654_, new_n5606_, new_n285_ );
and  ( new_n6655_, new_n6654_, new_n6653_ );
xor  ( new_n6656_, new_n6655_, new_n5206_ );
or   ( new_n6657_, new_n5207_, new_n294_ );
or   ( new_n6658_, new_n5209_, new_n301_ );
and  ( new_n6659_, new_n6658_, new_n6657_ );
xor  ( new_n6660_, new_n6659_, new_n4708_ );
or   ( new_n6661_, new_n6660_, new_n6656_ );
and  ( new_n6662_, new_n6660_, new_n6656_ );
or   ( new_n6663_, new_n4709_, new_n264_ );
or   ( new_n6664_, new_n4711_, new_n270_ );
and  ( new_n6665_, new_n6664_, new_n6663_ );
xor  ( new_n6666_, new_n6665_, new_n4295_ );
or   ( new_n6667_, new_n6666_, new_n6662_ );
and  ( new_n6668_, new_n6667_, new_n6661_ );
or   ( new_n6669_, new_n6668_, new_n6652_ );
and  ( new_n6670_, new_n6668_, new_n6652_ );
or   ( new_n6671_, new_n4302_, new_n419_ );
or   ( new_n6672_, new_n4304_, new_n348_ );
and  ( new_n6673_, new_n6672_, new_n6671_ );
xor  ( new_n6674_, new_n6673_, new_n3895_ );
or   ( new_n6675_, new_n3896_, new_n509_ );
or   ( new_n6676_, new_n3898_, new_n443_ );
and  ( new_n6677_, new_n6676_, new_n6675_ );
xor  ( new_n6678_, new_n6677_, new_n3460_ );
nor  ( new_n6679_, new_n6678_, new_n6674_ );
and  ( new_n6680_, new_n6678_, new_n6674_ );
or   ( new_n6681_, new_n3461_, new_n775_ );
or   ( new_n6682_, new_n3463_, new_n515_ );
and  ( new_n6683_, new_n6682_, new_n6681_ );
xor  ( new_n6684_, new_n6683_, new_n3116_ );
nor  ( new_n6685_, new_n6684_, new_n6680_ );
nor  ( new_n6686_, new_n6685_, new_n6679_ );
or   ( new_n6687_, new_n6686_, new_n6670_ );
and  ( new_n6688_, new_n6687_, new_n6669_ );
or   ( new_n6689_, new_n6688_, new_n6634_ );
and  ( new_n6690_, new_n6688_, new_n6634_ );
or   ( new_n6691_, new_n2122_, new_n1523_ );
or   ( new_n6692_, new_n2124_, new_n1525_ );
and  ( new_n6693_, new_n6692_, new_n6691_ );
xor  ( new_n6694_, new_n6693_, new_n1843_ );
or   ( new_n6695_, new_n1844_, new_n1899_ );
or   ( new_n6696_, new_n1846_, new_n1754_ );
and  ( new_n6697_, new_n6696_, new_n6695_ );
xor  ( new_n6698_, new_n6697_, new_n1586_ );
or   ( new_n6699_, new_n6698_, new_n6694_ );
and  ( new_n6700_, new_n6698_, new_n6694_ );
or   ( new_n6701_, new_n1593_, new_n2178_ );
or   ( new_n6702_, new_n1595_, new_n2057_ );
and  ( new_n6703_, new_n6702_, new_n6701_ );
xor  ( new_n6704_, new_n6703_, new_n1358_ );
or   ( new_n6705_, new_n6704_, new_n6700_ );
and  ( new_n6706_, new_n6705_, new_n6699_ );
or   ( new_n6707_, new_n3117_, new_n886_ );
or   ( new_n6708_, new_n3119_, new_n805_ );
and  ( new_n6709_, new_n6708_, new_n6707_ );
xor  ( new_n6710_, new_n6709_, new_n2800_ );
or   ( new_n6711_, new_n2807_, new_n1168_ );
or   ( new_n6712_, new_n2809_, new_n986_ );
and  ( new_n6713_, new_n6712_, new_n6711_ );
xor  ( new_n6714_, new_n6713_, new_n2424_ );
or   ( new_n6715_, new_n6714_, new_n6710_ );
and  ( new_n6716_, new_n6714_, new_n6710_ );
or   ( new_n6717_, new_n2425_, new_n1318_ );
or   ( new_n6718_, new_n2427_, new_n1213_ );
and  ( new_n6719_, new_n6718_, new_n6717_ );
xor  ( new_n6720_, new_n6719_, new_n2121_ );
or   ( new_n6721_, new_n6720_, new_n6716_ );
and  ( new_n6722_, new_n6721_, new_n6715_ );
nor  ( new_n6723_, new_n6722_, new_n6706_ );
and  ( new_n6724_, new_n6722_, new_n6706_ );
or   ( new_n6725_, new_n1364_, new_n2475_ );
or   ( new_n6726_, new_n1366_, new_n2291_ );
and  ( new_n6727_, new_n6726_, new_n6725_ );
xor  ( new_n6728_, new_n6727_, new_n1129_ );
or   ( new_n6729_, new_n1135_, new_n2751_ );
or   ( new_n6730_, new_n1137_, new_n2646_ );
and  ( new_n6731_, new_n6730_, new_n6729_ );
xor  ( new_n6732_, new_n6731_, new_n896_ );
nor  ( new_n6733_, new_n6732_, new_n6728_ );
and  ( new_n6734_, new_n6732_, new_n6728_ );
or   ( new_n6735_, new_n897_, new_n3178_ );
or   ( new_n6736_, new_n899_, new_n2981_ );
and  ( new_n6737_, new_n6736_, new_n6735_ );
xor  ( new_n6738_, new_n6737_, new_n748_ );
nor  ( new_n6739_, new_n6738_, new_n6734_ );
nor  ( new_n6740_, new_n6739_, new_n6733_ );
nor  ( new_n6741_, new_n6740_, new_n6724_ );
nor  ( new_n6742_, new_n6741_, new_n6723_ );
or   ( new_n6743_, new_n6742_, new_n6690_ );
and  ( new_n6744_, new_n6743_, new_n6689_ );
or   ( new_n6745_, new_n6744_, new_n6584_ );
nand ( new_n6746_, new_n6744_, new_n6584_ );
xnor ( new_n6747_, new_n6493_, new_n6489_ );
xor  ( new_n6748_, new_n6747_, new_n6499_ );
xnor ( new_n6749_, new_n6477_, new_n6473_ );
xor  ( new_n6750_, new_n6749_, new_n6483_ );
or   ( new_n6751_, new_n6750_, new_n6748_ );
and  ( new_n6752_, new_n6750_, new_n6748_ );
xor  ( new_n6753_, new_n6512_, new_n6507_ );
xnor ( new_n6754_, new_n6753_, new_n6518_ );
or   ( new_n6755_, new_n6754_, new_n6752_ );
and  ( new_n6756_, new_n6755_, new_n6751_ );
xnor ( new_n6757_, new_n6439_, new_n6435_ );
xor  ( new_n6758_, new_n6757_, new_n6445_ );
xnor ( new_n6759_, new_n6457_, new_n6453_ );
xor  ( new_n6760_, new_n6759_, new_n6463_ );
or   ( new_n6761_, new_n6760_, new_n6758_ );
and  ( new_n6762_, new_n6760_, new_n6758_ );
xor  ( new_n6763_, new_n6430_, new_n6429_ );
or   ( new_n6764_, new_n6763_, new_n6762_ );
and  ( new_n6765_, new_n6764_, new_n6761_ );
nor  ( new_n6766_, new_n6765_, new_n6756_ );
and  ( new_n6767_, new_n6765_, new_n6756_ );
xnor ( new_n6768_, new_n6396_, new_n6392_ );
xor  ( new_n6769_, new_n6768_, new_n6402_ );
xnor ( new_n6770_, new_n6380_, new_n6376_ );
xor  ( new_n6771_, new_n6770_, new_n6386_ );
nor  ( new_n6772_, new_n6771_, new_n6769_ );
and  ( new_n6773_, new_n6771_, new_n6769_ );
xor  ( new_n6774_, new_n6414_, new_n6410_ );
xnor ( new_n6775_, new_n6774_, new_n6420_ );
nor  ( new_n6776_, new_n6775_, new_n6773_ );
nor  ( new_n6777_, new_n6776_, new_n6772_ );
nor  ( new_n6778_, new_n6777_, new_n6767_ );
nor  ( new_n6779_, new_n6778_, new_n6766_ );
nand ( new_n6780_, new_n6779_, new_n6746_ );
and  ( new_n6781_, new_n6780_, new_n6745_ );
nor  ( new_n6782_, new_n6781_, new_n6574_ );
and  ( new_n6783_, new_n6781_, new_n6574_ );
xnor ( new_n6784_, new_n6404_, new_n6388_ );
xor  ( new_n6785_, new_n6784_, new_n6422_ );
xnor ( new_n6786_, new_n6447_, new_n6431_ );
xor  ( new_n6787_, new_n6786_, new_n6465_ );
nor  ( new_n6788_, new_n6787_, new_n6785_ );
nand ( new_n6789_, new_n6787_, new_n6785_ );
xor  ( new_n6790_, new_n6501_, new_n6485_ );
xor  ( new_n6791_, new_n6790_, new_n6520_ );
and  ( new_n6792_, new_n6791_, new_n6789_ );
or   ( new_n6793_, new_n6792_, new_n6788_ );
xnor ( new_n6794_, new_n6530_, new_n6528_ );
xor  ( new_n6795_, new_n6794_, new_n6534_ );
nor  ( new_n6796_, new_n6795_, new_n6793_ );
and  ( new_n6797_, new_n6795_, new_n6793_ );
xor  ( new_n6798_, new_n6328_, new_n6326_ );
xnor ( new_n6799_, new_n6798_, new_n6332_ );
nor  ( new_n6800_, new_n6799_, new_n6797_ );
nor  ( new_n6801_, new_n6800_, new_n6796_ );
nor  ( new_n6802_, new_n6801_, new_n6783_ );
nor  ( new_n6803_, new_n6802_, new_n6782_ );
or   ( new_n6804_, new_n6803_, new_n6569_ );
and  ( new_n6805_, new_n6804_, new_n6568_ );
or   ( new_n6806_, new_n6805_, new_n6556_ );
and  ( new_n6807_, new_n6805_, new_n6556_ );
xor  ( new_n6808_, new_n6311_, new_n6309_ );
xor  ( new_n6809_, new_n6808_, new_n6541_ );
or   ( new_n6810_, new_n6809_, new_n6807_ );
and  ( new_n6811_, new_n6810_, new_n6806_ );
xor  ( new_n6812_, new_n6545_, new_n6543_ );
xor  ( new_n6813_, new_n6812_, new_n6549_ );
and  ( new_n6814_, new_n6813_, new_n6811_ );
xor  ( new_n6815_, new_n6551_, new_n6300_ );
and  ( new_n6816_, new_n6815_, new_n6814_ );
xor  ( new_n6817_, new_n6560_, new_n6558_ );
xor  ( new_n6818_, new_n6817_, new_n6563_ );
xor  ( new_n6819_, new_n6744_, new_n6584_ );
xor  ( new_n6820_, new_n6819_, new_n6779_ );
xnor ( new_n6821_, new_n6795_, new_n6793_ );
xor  ( new_n6822_, new_n6821_, new_n6799_ );
or   ( new_n6823_, new_n6822_, new_n6820_ );
and  ( new_n6824_, new_n6822_, new_n6820_ );
xnor ( new_n6825_, new_n6573_, new_n6571_ );
or   ( new_n6826_, new_n6825_, new_n6824_ );
and  ( new_n6827_, new_n6826_, new_n6823_ );
nor  ( new_n6828_, new_n6827_, new_n6818_ );
and  ( new_n6829_, new_n6827_, new_n6818_ );
xor  ( new_n6830_, new_n6765_, new_n6756_ );
xnor ( new_n6831_, new_n6830_, new_n6777_ );
xnor ( new_n6832_, new_n6688_, new_n6634_ );
xnor ( new_n6833_, new_n6832_, new_n6742_ );
and  ( new_n6834_, new_n6833_, new_n6831_ );
xnor ( new_n6835_, new_n6714_, new_n6710_ );
xor  ( new_n6836_, new_n6835_, new_n6720_ );
xnor ( new_n6837_, new_n6698_, new_n6694_ );
xor  ( new_n6838_, new_n6837_, new_n6704_ );
or   ( new_n6839_, new_n6838_, new_n6836_ );
and  ( new_n6840_, new_n6838_, new_n6836_ );
xor  ( new_n6841_, new_n6732_, new_n6728_ );
xnor ( new_n6842_, new_n6841_, new_n6738_ );
or   ( new_n6843_, new_n6842_, new_n6840_ );
and  ( new_n6844_, new_n6843_, new_n6839_ );
xnor ( new_n6845_, new_n6660_, new_n6656_ );
xor  ( new_n6846_, new_n6845_, new_n6666_ );
xnor ( new_n6847_, new_n6678_, new_n6674_ );
xor  ( new_n6848_, new_n6847_, new_n6684_ );
or   ( new_n6849_, new_n6848_, new_n6846_ );
and  ( new_n6850_, new_n6848_, new_n6846_ );
xor  ( new_n6851_, new_n6642_, new_n6638_ );
xor  ( new_n6852_, new_n6851_, new_n6650_ );
not  ( new_n6853_, new_n6852_ );
or   ( new_n6854_, new_n6853_, new_n6850_ );
and  ( new_n6855_, new_n6854_, new_n6849_ );
nor  ( new_n6856_, new_n6855_, new_n6844_ );
nand ( new_n6857_, new_n6855_, new_n6844_ );
xnor ( new_n6858_, new_n6593_, new_n6588_ );
xor  ( new_n6859_, new_n6858_, new_n6595_ );
xnor ( new_n6860_, new_n6606_, new_n6602_ );
xor  ( new_n6861_, new_n6860_, new_n6612_ );
nor  ( new_n6862_, new_n6861_, new_n6859_ );
nand ( new_n6863_, new_n6861_, new_n6859_ );
xor  ( new_n6864_, new_n6624_, new_n6620_ );
xor  ( new_n6865_, new_n6864_, new_n6630_ );
and  ( new_n6866_, new_n6865_, new_n6863_ );
or   ( new_n6867_, new_n6866_, new_n6862_ );
and  ( new_n6868_, new_n6867_, new_n6857_ );
or   ( new_n6869_, new_n6868_, new_n6856_ );
or   ( new_n6870_, new_n4302_, new_n443_ );
or   ( new_n6871_, new_n4304_, new_n419_ );
and  ( new_n6872_, new_n6871_, new_n6870_ );
xor  ( new_n6873_, new_n6872_, new_n3895_ );
or   ( new_n6874_, new_n3896_, new_n515_ );
or   ( new_n6875_, new_n3898_, new_n509_ );
and  ( new_n6876_, new_n6875_, new_n6874_ );
xor  ( new_n6877_, new_n6876_, new_n3460_ );
or   ( new_n6878_, new_n6877_, new_n6873_ );
and  ( new_n6879_, new_n6877_, new_n6873_ );
or   ( new_n6880_, new_n3461_, new_n805_ );
or   ( new_n6881_, new_n3463_, new_n775_ );
and  ( new_n6882_, new_n6881_, new_n6880_ );
xor  ( new_n6883_, new_n6882_, new_n3116_ );
or   ( new_n6884_, new_n6883_, new_n6879_ );
and  ( new_n6885_, new_n6884_, new_n6878_ );
or   ( new_n6886_, new_n5604_, new_n301_ );
or   ( new_n6887_, new_n5606_, new_n279_ );
and  ( new_n6888_, new_n6887_, new_n6886_ );
xor  ( new_n6889_, new_n6888_, new_n5206_ );
or   ( new_n6890_, new_n5207_, new_n270_ );
or   ( new_n6891_, new_n5209_, new_n294_ );
and  ( new_n6892_, new_n6891_, new_n6890_ );
xor  ( new_n6893_, new_n6892_, new_n4708_ );
or   ( new_n6894_, new_n6893_, new_n6889_ );
and  ( new_n6895_, new_n6893_, new_n6889_ );
or   ( new_n6896_, new_n4709_, new_n348_ );
or   ( new_n6897_, new_n4711_, new_n264_ );
and  ( new_n6898_, new_n6897_, new_n6896_ );
xor  ( new_n6899_, new_n6898_, new_n4295_ );
or   ( new_n6900_, new_n6899_, new_n6895_ );
and  ( new_n6901_, new_n6900_, new_n6894_ );
or   ( new_n6902_, new_n6901_, new_n6885_ );
and  ( new_n6903_, new_n6901_, new_n6885_ );
or   ( new_n6904_, new_n6645_, new_n319_ );
or   ( new_n6905_, new_n6647_, new_n333_ );
and  ( new_n6906_, new_n6905_, new_n6904_ );
xor  ( new_n6907_, new_n6906_, new_n6165_ );
xor  ( new_n6908_, RIbb2ddb0_53, RIbb2de28_52 );
xor  ( new_n6909_, RIbb2de28_52, new_n6635_ );
nor  ( new_n6910_, new_n6909_, new_n6908_ );
and  ( new_n6911_, new_n6910_, RIbb2d810_65 );
xor  ( new_n6912_, new_n6911_, new_n6638_ );
and  ( new_n6913_, new_n6912_, new_n6907_ );
nor  ( new_n6914_, new_n6912_, new_n6907_ );
or   ( new_n6915_, new_n6173_, new_n285_ );
or   ( new_n6916_, new_n6175_, new_n313_ );
and  ( new_n6917_, new_n6916_, new_n6915_ );
xor  ( new_n6918_, new_n6917_, new_n5597_ );
nor  ( new_n6919_, new_n6918_, new_n6914_ );
nor  ( new_n6920_, new_n6919_, new_n6913_ );
or   ( new_n6921_, new_n6920_, new_n6903_ );
and  ( new_n6922_, new_n6921_, new_n6902_ );
or   ( new_n6923_, new_n755_, new_n3694_ );
or   ( new_n6924_, new_n757_, new_n3696_ );
and  ( new_n6925_, new_n6924_, new_n6923_ );
xor  ( new_n6926_, new_n6925_, new_n523_ );
or   ( new_n6927_, new_n524_, new_n4069_ );
or   ( new_n6928_, new_n526_, new_n3820_ );
and  ( new_n6929_, new_n6928_, new_n6927_ );
xor  ( new_n6930_, new_n6929_, new_n403_ );
or   ( new_n6931_, new_n6930_, new_n6926_ );
and  ( new_n6932_, new_n6930_, new_n6926_ );
or   ( new_n6933_, new_n409_, new_n4603_ );
or   ( new_n6934_, new_n411_, new_n4267_ );
and  ( new_n6935_, new_n6934_, new_n6933_ );
xor  ( new_n6936_, new_n6935_, new_n328_ );
or   ( new_n6937_, new_n6936_, new_n6932_ );
and  ( new_n6938_, new_n6937_, new_n6931_ );
or   ( new_n6939_, new_n299_, new_n6425_ );
or   ( new_n6940_, new_n302_, new_n6219_ );
and  ( new_n6941_, new_n6940_, new_n6939_ );
xor  ( new_n6942_, new_n6941_, new_n293_ );
not  ( new_n6943_, RIbb2c0a0_115 );
or   ( new_n6944_, new_n268_, new_n6943_ );
or   ( new_n6945_, new_n271_, new_n6589_ );
and  ( new_n6946_, new_n6945_, new_n6944_ );
xor  ( new_n6947_, new_n6946_, new_n263_ );
nor  ( new_n6948_, new_n6947_, new_n6942_ );
and  ( new_n6949_, RIbb2c028_116, RIbb2f610_1 );
and  ( new_n6950_, new_n6947_, new_n6942_ );
nor  ( new_n6951_, new_n6950_, new_n6949_ );
nor  ( new_n6952_, new_n6951_, new_n6948_ );
or   ( new_n6953_, new_n337_, new_n4859_ );
or   ( new_n6954_, new_n340_, new_n4995_ );
and  ( new_n6955_, new_n6954_, new_n6953_ );
xor  ( new_n6956_, new_n6955_, new_n332_ );
or   ( new_n6957_, new_n317_, new_n5428_ );
or   ( new_n6958_, new_n320_, new_n5171_ );
and  ( new_n6959_, new_n6958_, new_n6957_ );
xor  ( new_n6960_, new_n6959_, new_n312_ );
or   ( new_n6961_, new_n6960_, new_n6956_ );
and  ( new_n6962_, new_n6960_, new_n6956_ );
or   ( new_n6963_, new_n283_, new_n5899_ );
or   ( new_n6964_, new_n286_, new_n5570_ );
and  ( new_n6965_, new_n6964_, new_n6963_ );
xor  ( new_n6966_, new_n6965_, new_n278_ );
or   ( new_n6967_, new_n6966_, new_n6962_ );
and  ( new_n6968_, new_n6967_, new_n6961_ );
and  ( new_n6969_, new_n6968_, new_n6952_ );
or   ( new_n6970_, new_n6969_, new_n6938_ );
or   ( new_n6971_, new_n6968_, new_n6952_ );
and  ( new_n6972_, new_n6971_, new_n6970_ );
or   ( new_n6973_, new_n6972_, new_n6922_ );
or   ( new_n6974_, new_n2122_, new_n1754_ );
or   ( new_n6975_, new_n2124_, new_n1523_ );
and  ( new_n6976_, new_n6975_, new_n6974_ );
xor  ( new_n6977_, new_n6976_, new_n1843_ );
or   ( new_n6978_, new_n1844_, new_n2057_ );
or   ( new_n6979_, new_n1846_, new_n1899_ );
and  ( new_n6980_, new_n6979_, new_n6978_ );
xor  ( new_n6981_, new_n6980_, new_n1586_ );
or   ( new_n6982_, new_n6981_, new_n6977_ );
and  ( new_n6983_, new_n6981_, new_n6977_ );
or   ( new_n6984_, new_n1593_, new_n2291_ );
or   ( new_n6985_, new_n1595_, new_n2178_ );
and  ( new_n6986_, new_n6985_, new_n6984_ );
xor  ( new_n6987_, new_n6986_, new_n1358_ );
or   ( new_n6988_, new_n6987_, new_n6983_ );
and  ( new_n6989_, new_n6988_, new_n6982_ );
or   ( new_n6990_, new_n3117_, new_n986_ );
or   ( new_n6991_, new_n3119_, new_n886_ );
and  ( new_n6992_, new_n6991_, new_n6990_ );
xor  ( new_n6993_, new_n6992_, new_n2800_ );
or   ( new_n6994_, new_n2807_, new_n1213_ );
or   ( new_n6995_, new_n2809_, new_n1168_ );
and  ( new_n6996_, new_n6995_, new_n6994_ );
xor  ( new_n6997_, new_n6996_, new_n2424_ );
or   ( new_n6998_, new_n6997_, new_n6993_ );
and  ( new_n6999_, new_n6997_, new_n6993_ );
or   ( new_n7000_, new_n2425_, new_n1525_ );
or   ( new_n7001_, new_n2427_, new_n1318_ );
and  ( new_n7002_, new_n7001_, new_n7000_ );
xor  ( new_n7003_, new_n7002_, new_n2121_ );
or   ( new_n7004_, new_n7003_, new_n6999_ );
and  ( new_n7005_, new_n7004_, new_n6998_ );
nor  ( new_n7006_, new_n7005_, new_n6989_ );
and  ( new_n7007_, new_n7005_, new_n6989_ );
or   ( new_n7008_, new_n1364_, new_n2646_ );
or   ( new_n7009_, new_n1366_, new_n2475_ );
and  ( new_n7010_, new_n7009_, new_n7008_ );
xor  ( new_n7011_, new_n7010_, new_n1129_ );
or   ( new_n7012_, new_n1135_, new_n2981_ );
or   ( new_n7013_, new_n1137_, new_n2751_ );
and  ( new_n7014_, new_n7013_, new_n7012_ );
xor  ( new_n7015_, new_n7014_, new_n896_ );
nor  ( new_n7016_, new_n7015_, new_n7011_ );
and  ( new_n7017_, new_n7015_, new_n7011_ );
or   ( new_n7018_, new_n897_, new_n3306_ );
or   ( new_n7019_, new_n899_, new_n3178_ );
and  ( new_n7020_, new_n7019_, new_n7018_ );
xor  ( new_n7021_, new_n7020_, new_n748_ );
nor  ( new_n7022_, new_n7021_, new_n7017_ );
nor  ( new_n7023_, new_n7022_, new_n7016_ );
nor  ( new_n7024_, new_n7023_, new_n7007_ );
nor  ( new_n7025_, new_n7024_, new_n7006_ );
and  ( new_n7026_, new_n6972_, new_n6922_ );
or   ( new_n7027_, new_n7026_, new_n7025_ );
and  ( new_n7028_, new_n7027_, new_n6973_ );
or   ( new_n7029_, new_n7028_, new_n6869_ );
and  ( new_n7030_, new_n7028_, new_n6869_ );
xnor ( new_n7031_, new_n6771_, new_n6769_ );
xor  ( new_n7032_, new_n7031_, new_n6775_ );
xnor ( new_n7033_, new_n6750_, new_n6748_ );
xor  ( new_n7034_, new_n7033_, new_n6754_ );
and  ( new_n7035_, new_n7034_, new_n7032_ );
or   ( new_n7036_, new_n7034_, new_n7032_ );
xor  ( new_n7037_, new_n6760_, new_n6758_ );
xor  ( new_n7038_, new_n7037_, new_n6763_ );
not  ( new_n7039_, new_n7038_ );
and  ( new_n7040_, new_n7039_, new_n7036_ );
or   ( new_n7041_, new_n7040_, new_n7035_ );
or   ( new_n7042_, new_n7041_, new_n7030_ );
and  ( new_n7043_, new_n7042_, new_n7029_ );
and  ( new_n7044_, new_n7043_, new_n6834_ );
nor  ( new_n7045_, new_n7043_, new_n6834_ );
xnor ( new_n7046_, new_n6614_, new_n6598_ );
xor  ( new_n7047_, new_n7046_, new_n6632_ );
xnor ( new_n7048_, new_n6668_, new_n6652_ );
xor  ( new_n7049_, new_n7048_, new_n6686_ );
nor  ( new_n7050_, new_n7049_, new_n7047_ );
nand ( new_n7051_, new_n7049_, new_n7047_ );
xor  ( new_n7052_, new_n6722_, new_n6706_ );
xor  ( new_n7053_, new_n7052_, new_n6740_ );
and  ( new_n7054_, new_n7053_, new_n7051_ );
or   ( new_n7055_, new_n7054_, new_n7050_ );
xor  ( new_n7056_, new_n6787_, new_n6785_ );
xor  ( new_n7057_, new_n7056_, new_n6791_ );
and  ( new_n7058_, new_n7057_, new_n7055_ );
nor  ( new_n7059_, new_n7057_, new_n7055_ );
xor  ( new_n7060_, new_n6578_, new_n6576_ );
xnor ( new_n7061_, new_n7060_, new_n6582_ );
nor  ( new_n7062_, new_n7061_, new_n7059_ );
nor  ( new_n7063_, new_n7062_, new_n7058_ );
nor  ( new_n7064_, new_n7063_, new_n7045_ );
nor  ( new_n7065_, new_n7064_, new_n7044_ );
nor  ( new_n7066_, new_n7065_, new_n6829_ );
or   ( new_n7067_, new_n7066_, new_n6828_ );
xnor ( new_n7068_, new_n6336_, new_n6318_ );
xor  ( new_n7069_, new_n7068_, new_n6538_ );
nor  ( new_n7070_, new_n7069_, new_n7067_ );
nand ( new_n7071_, new_n7069_, new_n7067_ );
xnor ( new_n7072_, new_n6567_, new_n6565_ );
xor  ( new_n7073_, new_n7072_, new_n6803_ );
and  ( new_n7074_, new_n7073_, new_n7071_ );
or   ( new_n7075_, new_n7074_, new_n7070_ );
xnor ( new_n7076_, new_n6805_, new_n6556_ );
xor  ( new_n7077_, new_n7076_, new_n6809_ );
nor  ( new_n7078_, new_n7077_, new_n7075_ );
xor  ( new_n7079_, new_n6813_, new_n6811_ );
and  ( new_n7080_, new_n7079_, new_n7078_ );
xor  ( new_n7081_, new_n6827_, new_n6818_ );
xor  ( new_n7082_, new_n7081_, new_n7065_ );
xnor ( new_n7083_, new_n6781_, new_n6574_ );
xor  ( new_n7084_, new_n7083_, new_n6801_ );
or   ( new_n7085_, new_n7084_, new_n7082_ );
and  ( new_n7086_, new_n7084_, new_n7082_ );
xor  ( new_n7087_, new_n6822_, new_n6820_ );
xor  ( new_n7088_, new_n7087_, new_n6825_ );
xor  ( new_n7089_, new_n7028_, new_n6869_ );
xor  ( new_n7090_, new_n7089_, new_n7041_ );
xnor ( new_n7091_, new_n7057_, new_n7055_ );
xor  ( new_n7092_, new_n7091_, new_n7061_ );
nand ( new_n7093_, new_n7092_, new_n7090_ );
nor  ( new_n7094_, new_n7092_, new_n7090_ );
xnor ( new_n7095_, new_n6833_, new_n6831_ );
or   ( new_n7096_, new_n7095_, new_n7094_ );
and  ( new_n7097_, new_n7096_, new_n7093_ );
nor  ( new_n7098_, new_n7097_, new_n7088_ );
and  ( new_n7099_, new_n7097_, new_n7088_ );
xor  ( new_n7100_, new_n6972_, new_n6922_ );
xnor ( new_n7101_, new_n7100_, new_n7025_ );
xor  ( new_n7102_, new_n6855_, new_n6844_ );
xnor ( new_n7103_, new_n7102_, new_n6867_ );
or   ( new_n7104_, new_n7103_, new_n7101_ );
or   ( new_n7105_, new_n409_, new_n4995_ );
or   ( new_n7106_, new_n411_, new_n4603_ );
and  ( new_n7107_, new_n7106_, new_n7105_ );
xor  ( new_n7108_, new_n7107_, new_n328_ );
or   ( new_n7109_, new_n337_, new_n5171_ );
or   ( new_n7110_, new_n340_, new_n4859_ );
and  ( new_n7111_, new_n7110_, new_n7109_ );
xor  ( new_n7112_, new_n7111_, new_n332_ );
or   ( new_n7113_, new_n7112_, new_n7108_ );
and  ( new_n7114_, new_n7112_, new_n7108_ );
or   ( new_n7115_, new_n317_, new_n5570_ );
or   ( new_n7116_, new_n320_, new_n5428_ );
and  ( new_n7117_, new_n7116_, new_n7115_ );
xor  ( new_n7118_, new_n7117_, new_n312_ );
or   ( new_n7119_, new_n7118_, new_n7114_ );
and  ( new_n7120_, new_n7119_, new_n7113_ );
or   ( new_n7121_, new_n897_, new_n3696_ );
or   ( new_n7122_, new_n899_, new_n3306_ );
and  ( new_n7123_, new_n7122_, new_n7121_ );
xor  ( new_n7124_, new_n7123_, new_n748_ );
or   ( new_n7125_, new_n755_, new_n3820_ );
or   ( new_n7126_, new_n757_, new_n3694_ );
and  ( new_n7127_, new_n7126_, new_n7125_ );
xor  ( new_n7128_, new_n7127_, new_n523_ );
or   ( new_n7129_, new_n7128_, new_n7124_ );
and  ( new_n7130_, new_n7128_, new_n7124_ );
or   ( new_n7131_, new_n524_, new_n4267_ );
or   ( new_n7132_, new_n526_, new_n4069_ );
and  ( new_n7133_, new_n7132_, new_n7131_ );
xor  ( new_n7134_, new_n7133_, new_n403_ );
or   ( new_n7135_, new_n7134_, new_n7130_ );
and  ( new_n7136_, new_n7135_, new_n7129_ );
or   ( new_n7137_, new_n7136_, new_n7120_ );
and  ( new_n7138_, new_n7136_, new_n7120_ );
or   ( new_n7139_, new_n283_, new_n6219_ );
or   ( new_n7140_, new_n286_, new_n5899_ );
and  ( new_n7141_, new_n7140_, new_n7139_ );
xor  ( new_n7142_, new_n7141_, new_n278_ );
or   ( new_n7143_, new_n299_, new_n6589_ );
or   ( new_n7144_, new_n302_, new_n6425_ );
and  ( new_n7145_, new_n7144_, new_n7143_ );
xor  ( new_n7146_, new_n7145_, new_n293_ );
nor  ( new_n7147_, new_n7146_, new_n7142_ );
and  ( new_n7148_, new_n7146_, new_n7142_ );
not  ( new_n7149_, RIbb2c028_116 );
or   ( new_n7150_, new_n268_, new_n7149_ );
or   ( new_n7151_, new_n271_, new_n6943_ );
and  ( new_n7152_, new_n7151_, new_n7150_ );
xor  ( new_n7153_, new_n7152_, new_n263_ );
nor  ( new_n7154_, new_n7153_, new_n7148_ );
nor  ( new_n7155_, new_n7154_, new_n7147_ );
or   ( new_n7156_, new_n7155_, new_n7138_ );
and  ( new_n7157_, new_n7156_, new_n7137_ );
or   ( new_n7158_, new_n6173_, new_n279_ );
or   ( new_n7159_, new_n6175_, new_n285_ );
and  ( new_n7160_, new_n7159_, new_n7158_ );
xor  ( new_n7161_, new_n7160_, new_n5597_ );
or   ( new_n7162_, new_n5604_, new_n294_ );
or   ( new_n7163_, new_n5606_, new_n301_ );
and  ( new_n7164_, new_n7163_, new_n7162_ );
xor  ( new_n7165_, new_n7164_, new_n5206_ );
nor  ( new_n7166_, new_n7165_, new_n7161_ );
nand ( new_n7167_, new_n7165_, new_n7161_ );
or   ( new_n7168_, new_n5207_, new_n264_ );
or   ( new_n7169_, new_n5209_, new_n270_ );
and  ( new_n7170_, new_n7169_, new_n7168_ );
xor  ( new_n7171_, new_n7170_, new_n4707_ );
and  ( new_n7172_, new_n7171_, new_n7167_ );
or   ( new_n7173_, new_n7172_, new_n7166_ );
not  ( new_n7174_, RIbb2ddb0_53 );
and  ( new_n7175_, RIbb2dcc0_55, RIbb2dd38_54 );
nor  ( new_n7176_, new_n7175_, new_n7174_ );
not  ( new_n7177_, new_n7176_ );
or   ( new_n7178_, new_n6645_, new_n313_ );
or   ( new_n7179_, new_n6647_, new_n319_ );
and  ( new_n7180_, new_n7179_, new_n7178_ );
xor  ( new_n7181_, new_n7180_, new_n6166_ );
nand ( new_n7182_, new_n7181_, new_n7177_ );
or   ( new_n7183_, new_n7181_, new_n7177_ );
not  ( new_n7184_, new_n6910_ );
or   ( new_n7185_, new_n7184_, new_n333_ );
not  ( new_n7186_, new_n6908_ );
or   ( new_n7187_, new_n7186_, new_n339_ );
and  ( new_n7188_, new_n7187_, new_n7185_ );
xor  ( new_n7189_, new_n7188_, new_n6638_ );
nand ( new_n7190_, new_n7189_, new_n7183_ );
and  ( new_n7191_, new_n7190_, new_n7182_ );
nand ( new_n7192_, new_n7191_, new_n7173_ );
nor  ( new_n7193_, new_n7191_, new_n7173_ );
or   ( new_n7194_, new_n4709_, new_n419_ );
or   ( new_n7195_, new_n4711_, new_n348_ );
and  ( new_n7196_, new_n7195_, new_n7194_ );
xor  ( new_n7197_, new_n7196_, new_n4295_ );
or   ( new_n7198_, new_n4302_, new_n509_ );
or   ( new_n7199_, new_n4304_, new_n443_ );
and  ( new_n7200_, new_n7199_, new_n7198_ );
xor  ( new_n7201_, new_n7200_, new_n3895_ );
nor  ( new_n7202_, new_n7201_, new_n7197_ );
and  ( new_n7203_, new_n7201_, new_n7197_ );
or   ( new_n7204_, new_n3896_, new_n775_ );
or   ( new_n7205_, new_n3898_, new_n515_ );
and  ( new_n7206_, new_n7205_, new_n7204_ );
xor  ( new_n7207_, new_n7206_, new_n3460_ );
nor  ( new_n7208_, new_n7207_, new_n7203_ );
nor  ( new_n7209_, new_n7208_, new_n7202_ );
or   ( new_n7210_, new_n7209_, new_n7193_ );
and  ( new_n7211_, new_n7210_, new_n7192_ );
nor  ( new_n7212_, new_n7211_, new_n7157_ );
nand ( new_n7213_, new_n7211_, new_n7157_ );
or   ( new_n7214_, new_n3461_, new_n886_ );
or   ( new_n7215_, new_n3463_, new_n805_ );
and  ( new_n7216_, new_n7215_, new_n7214_ );
xor  ( new_n7217_, new_n7216_, new_n3116_ );
or   ( new_n7218_, new_n3117_, new_n1168_ );
or   ( new_n7219_, new_n3119_, new_n986_ );
and  ( new_n7220_, new_n7219_, new_n7218_ );
xor  ( new_n7221_, new_n7220_, new_n2800_ );
or   ( new_n7222_, new_n7221_, new_n7217_ );
and  ( new_n7223_, new_n7221_, new_n7217_ );
or   ( new_n7224_, new_n2807_, new_n1318_ );
or   ( new_n7225_, new_n2809_, new_n1213_ );
and  ( new_n7226_, new_n7225_, new_n7224_ );
xor  ( new_n7227_, new_n7226_, new_n2424_ );
or   ( new_n7228_, new_n7227_, new_n7223_ );
and  ( new_n7229_, new_n7228_, new_n7222_ );
or   ( new_n7230_, new_n2425_, new_n1523_ );
or   ( new_n7231_, new_n2427_, new_n1525_ );
and  ( new_n7232_, new_n7231_, new_n7230_ );
xor  ( new_n7233_, new_n7232_, new_n2121_ );
or   ( new_n7234_, new_n2122_, new_n1899_ );
or   ( new_n7235_, new_n2124_, new_n1754_ );
and  ( new_n7236_, new_n7235_, new_n7234_ );
xor  ( new_n7237_, new_n7236_, new_n1843_ );
or   ( new_n7238_, new_n7237_, new_n7233_ );
and  ( new_n7239_, new_n7237_, new_n7233_ );
or   ( new_n7240_, new_n1844_, new_n2178_ );
or   ( new_n7241_, new_n1846_, new_n2057_ );
and  ( new_n7242_, new_n7241_, new_n7240_ );
xor  ( new_n7243_, new_n7242_, new_n1586_ );
or   ( new_n7244_, new_n7243_, new_n7239_ );
and  ( new_n7245_, new_n7244_, new_n7238_ );
nor  ( new_n7246_, new_n7245_, new_n7229_ );
nand ( new_n7247_, new_n7245_, new_n7229_ );
or   ( new_n7248_, new_n1593_, new_n2475_ );
or   ( new_n7249_, new_n1595_, new_n2291_ );
and  ( new_n7250_, new_n7249_, new_n7248_ );
xor  ( new_n7251_, new_n7250_, new_n1358_ );
or   ( new_n7252_, new_n1364_, new_n2751_ );
or   ( new_n7253_, new_n1366_, new_n2646_ );
and  ( new_n7254_, new_n7253_, new_n7252_ );
xor  ( new_n7255_, new_n7254_, new_n1129_ );
nor  ( new_n7256_, new_n7255_, new_n7251_ );
and  ( new_n7257_, new_n7255_, new_n7251_ );
or   ( new_n7258_, new_n1135_, new_n3178_ );
or   ( new_n7259_, new_n1137_, new_n2981_ );
and  ( new_n7260_, new_n7259_, new_n7258_ );
xor  ( new_n7261_, new_n7260_, new_n896_ );
nor  ( new_n7262_, new_n7261_, new_n7257_ );
or   ( new_n7263_, new_n7262_, new_n7256_ );
and  ( new_n7264_, new_n7263_, new_n7247_ );
or   ( new_n7265_, new_n7264_, new_n7246_ );
and  ( new_n7266_, new_n7265_, new_n7213_ );
or   ( new_n7267_, new_n7266_, new_n7212_ );
xor  ( new_n7268_, new_n6861_, new_n6859_ );
xor  ( new_n7269_, new_n7268_, new_n6865_ );
xnor ( new_n7270_, new_n6838_, new_n6836_ );
xor  ( new_n7271_, new_n7270_, new_n6842_ );
nand ( new_n7272_, new_n7271_, new_n7269_ );
nor  ( new_n7273_, new_n7271_, new_n7269_ );
xor  ( new_n7274_, new_n6848_, new_n6846_ );
xor  ( new_n7275_, new_n7274_, new_n6853_ );
or   ( new_n7276_, new_n7275_, new_n7273_ );
and  ( new_n7277_, new_n7276_, new_n7272_ );
or   ( new_n7278_, new_n7277_, new_n7267_ );
and  ( new_n7279_, new_n7277_, new_n7267_ );
xor  ( new_n7280_, new_n6947_, new_n6942_ );
xnor ( new_n7281_, new_n7280_, new_n6949_ );
xnor ( new_n7282_, new_n6960_, new_n6956_ );
xor  ( new_n7283_, new_n7282_, new_n6966_ );
and  ( new_n7284_, new_n7283_, new_n7281_ );
xnor ( new_n7285_, new_n6981_, new_n6977_ );
xor  ( new_n7286_, new_n7285_, new_n6987_ );
xnor ( new_n7287_, new_n6930_, new_n6926_ );
xor  ( new_n7288_, new_n7287_, new_n6936_ );
or   ( new_n7289_, new_n7288_, new_n7286_ );
and  ( new_n7290_, new_n7288_, new_n7286_ );
xor  ( new_n7291_, new_n7015_, new_n7011_ );
xnor ( new_n7292_, new_n7291_, new_n7021_ );
or   ( new_n7293_, new_n7292_, new_n7290_ );
and  ( new_n7294_, new_n7293_, new_n7289_ );
or   ( new_n7295_, new_n7294_, new_n7284_ );
and  ( new_n7296_, new_n7294_, new_n7284_ );
xnor ( new_n7297_, new_n6893_, new_n6889_ );
xor  ( new_n7298_, new_n7297_, new_n6899_ );
xnor ( new_n7299_, new_n6997_, new_n6993_ );
xor  ( new_n7300_, new_n7299_, new_n7003_ );
nor  ( new_n7301_, new_n7300_, new_n7298_ );
and  ( new_n7302_, new_n7300_, new_n7298_ );
xor  ( new_n7303_, new_n6877_, new_n6873_ );
xnor ( new_n7304_, new_n7303_, new_n6883_ );
nor  ( new_n7305_, new_n7304_, new_n7302_ );
nor  ( new_n7306_, new_n7305_, new_n7301_ );
or   ( new_n7307_, new_n7306_, new_n7296_ );
and  ( new_n7308_, new_n7307_, new_n7295_ );
or   ( new_n7309_, new_n7308_, new_n7279_ );
and  ( new_n7310_, new_n7309_, new_n7278_ );
nor  ( new_n7311_, new_n7310_, new_n7104_ );
and  ( new_n7312_, new_n7310_, new_n7104_ );
xnor ( new_n7313_, new_n6968_, new_n6952_ );
xor  ( new_n7314_, new_n7313_, new_n6938_ );
xnor ( new_n7315_, new_n6901_, new_n6885_ );
xor  ( new_n7316_, new_n7315_, new_n6920_ );
nor  ( new_n7317_, new_n7316_, new_n7314_ );
nand ( new_n7318_, new_n7316_, new_n7314_ );
xor  ( new_n7319_, new_n7005_, new_n6989_ );
xor  ( new_n7320_, new_n7319_, new_n7023_ );
and  ( new_n7321_, new_n7320_, new_n7318_ );
or   ( new_n7322_, new_n7321_, new_n7317_ );
xor  ( new_n7323_, new_n7049_, new_n7047_ );
xor  ( new_n7324_, new_n7323_, new_n7053_ );
and  ( new_n7325_, new_n7324_, new_n7322_ );
nor  ( new_n7326_, new_n7324_, new_n7322_ );
xor  ( new_n7327_, new_n7034_, new_n7032_ );
xor  ( new_n7328_, new_n7327_, new_n7039_ );
not  ( new_n7329_, new_n7328_ );
nor  ( new_n7330_, new_n7329_, new_n7326_ );
nor  ( new_n7331_, new_n7330_, new_n7325_ );
nor  ( new_n7332_, new_n7331_, new_n7312_ );
nor  ( new_n7333_, new_n7332_, new_n7311_ );
nor  ( new_n7334_, new_n7333_, new_n7099_ );
nor  ( new_n7335_, new_n7334_, new_n7098_ );
or   ( new_n7336_, new_n7335_, new_n7086_ );
and  ( new_n7337_, new_n7336_, new_n7085_ );
xor  ( new_n7338_, new_n7069_, new_n7067_ );
xor  ( new_n7339_, new_n7338_, new_n7073_ );
nor  ( new_n7340_, new_n7339_, new_n7337_ );
xor  ( new_n7341_, new_n7077_, new_n7075_ );
and  ( new_n7342_, new_n7341_, new_n7340_ );
xor  ( new_n7343_, new_n7092_, new_n7090_ );
xor  ( new_n7344_, new_n7343_, new_n7095_ );
xor  ( new_n7345_, new_n7277_, new_n7267_ );
xor  ( new_n7346_, new_n7345_, new_n7308_ );
xor  ( new_n7347_, new_n7324_, new_n7322_ );
xor  ( new_n7348_, new_n7347_, new_n7329_ );
or   ( new_n7349_, new_n7348_, new_n7346_ );
and  ( new_n7350_, new_n7348_, new_n7346_ );
xnor ( new_n7351_, new_n7103_, new_n7101_ );
or   ( new_n7352_, new_n7351_, new_n7350_ );
and  ( new_n7353_, new_n7352_, new_n7349_ );
nor  ( new_n7354_, new_n7353_, new_n7344_ );
and  ( new_n7355_, new_n7353_, new_n7344_ );
xor  ( new_n7356_, new_n7294_, new_n7284_ );
xnor ( new_n7357_, new_n7356_, new_n7306_ );
not  ( new_n7358_, new_n7357_ );
xor  ( new_n7359_, new_n7211_, new_n7157_ );
xor  ( new_n7360_, new_n7359_, new_n7265_ );
nor  ( new_n7361_, new_n7360_, new_n7358_ );
xor  ( new_n7362_, new_n7165_, new_n7161_ );
xor  ( new_n7363_, new_n7362_, new_n7171_ );
xnor ( new_n7364_, new_n7221_, new_n7217_ );
xor  ( new_n7365_, new_n7364_, new_n7227_ );
nor  ( new_n7366_, new_n7365_, new_n7363_ );
nand ( new_n7367_, new_n7365_, new_n7363_ );
xor  ( new_n7368_, new_n7201_, new_n7197_ );
xnor ( new_n7369_, new_n7368_, new_n7207_ );
not  ( new_n7370_, new_n7369_ );
and  ( new_n7371_, new_n7370_, new_n7367_ );
or   ( new_n7372_, new_n7371_, new_n7366_ );
not  ( new_n7373_, RIbb2bfb0_117 );
or   ( new_n7374_, new_n7373_, new_n260_ );
xnor ( new_n7375_, new_n7112_, new_n7108_ );
xor  ( new_n7376_, new_n7375_, new_n7118_ );
nand ( new_n7377_, new_n7376_, new_n7374_ );
or   ( new_n7378_, new_n7376_, new_n7374_ );
xor  ( new_n7379_, new_n7146_, new_n7142_ );
xnor ( new_n7380_, new_n7379_, new_n7153_ );
nand ( new_n7381_, new_n7380_, new_n7378_ );
and  ( new_n7382_, new_n7381_, new_n7377_ );
and  ( new_n7383_, new_n7382_, new_n7372_ );
or   ( new_n7384_, new_n7382_, new_n7372_ );
xnor ( new_n7385_, new_n7128_, new_n7124_ );
xor  ( new_n7386_, new_n7385_, new_n7134_ );
xnor ( new_n7387_, new_n7237_, new_n7233_ );
xor  ( new_n7388_, new_n7387_, new_n7243_ );
nor  ( new_n7389_, new_n7388_, new_n7386_ );
nand ( new_n7390_, new_n7388_, new_n7386_ );
xor  ( new_n7391_, new_n7255_, new_n7251_ );
xor  ( new_n7392_, new_n7391_, new_n7261_ );
and  ( new_n7393_, new_n7392_, new_n7390_ );
or   ( new_n7394_, new_n7393_, new_n7389_ );
and  ( new_n7395_, new_n7394_, new_n7384_ );
or   ( new_n7396_, new_n7395_, new_n7383_ );
or   ( new_n7397_, new_n283_, new_n6425_ );
or   ( new_n7398_, new_n286_, new_n6219_ );
and  ( new_n7399_, new_n7398_, new_n7397_ );
xor  ( new_n7400_, new_n7399_, new_n278_ );
or   ( new_n7401_, new_n299_, new_n6943_ );
or   ( new_n7402_, new_n302_, new_n6589_ );
and  ( new_n7403_, new_n7402_, new_n7401_ );
xor  ( new_n7404_, new_n7403_, new_n293_ );
or   ( new_n7405_, new_n7404_, new_n7400_ );
and  ( new_n7406_, new_n7404_, new_n7400_ );
or   ( new_n7407_, new_n268_, new_n7373_ );
or   ( new_n7408_, new_n271_, new_n7149_ );
and  ( new_n7409_, new_n7408_, new_n7407_ );
xor  ( new_n7410_, new_n7409_, new_n263_ );
or   ( new_n7411_, new_n7410_, new_n7406_ );
and  ( new_n7412_, new_n7411_, new_n7405_ );
or   ( new_n7413_, new_n897_, new_n3694_ );
or   ( new_n7414_, new_n899_, new_n3696_ );
and  ( new_n7415_, new_n7414_, new_n7413_ );
xor  ( new_n7416_, new_n7415_, new_n748_ );
or   ( new_n7417_, new_n755_, new_n4069_ );
or   ( new_n7418_, new_n757_, new_n3820_ );
and  ( new_n7419_, new_n7418_, new_n7417_ );
xor  ( new_n7420_, new_n7419_, new_n523_ );
or   ( new_n7421_, new_n7420_, new_n7416_ );
and  ( new_n7422_, new_n7420_, new_n7416_ );
or   ( new_n7423_, new_n524_, new_n4603_ );
or   ( new_n7424_, new_n526_, new_n4267_ );
and  ( new_n7425_, new_n7424_, new_n7423_ );
xor  ( new_n7426_, new_n7425_, new_n403_ );
or   ( new_n7427_, new_n7426_, new_n7422_ );
and  ( new_n7428_, new_n7427_, new_n7421_ );
or   ( new_n7429_, new_n7428_, new_n7412_ );
and  ( new_n7430_, new_n7428_, new_n7412_ );
or   ( new_n7431_, new_n409_, new_n4859_ );
or   ( new_n7432_, new_n411_, new_n4995_ );
and  ( new_n7433_, new_n7432_, new_n7431_ );
xor  ( new_n7434_, new_n7433_, new_n328_ );
or   ( new_n7435_, new_n337_, new_n5428_ );
or   ( new_n7436_, new_n340_, new_n5171_ );
and  ( new_n7437_, new_n7436_, new_n7435_ );
xor  ( new_n7438_, new_n7437_, new_n332_ );
nor  ( new_n7439_, new_n7438_, new_n7434_ );
and  ( new_n7440_, new_n7438_, new_n7434_ );
or   ( new_n7441_, new_n317_, new_n5899_ );
or   ( new_n7442_, new_n320_, new_n5570_ );
and  ( new_n7443_, new_n7442_, new_n7441_ );
xor  ( new_n7444_, new_n7443_, new_n312_ );
nor  ( new_n7445_, new_n7444_, new_n7440_ );
nor  ( new_n7446_, new_n7445_, new_n7439_ );
or   ( new_n7447_, new_n7446_, new_n7430_ );
and  ( new_n7448_, new_n7447_, new_n7429_ );
or   ( new_n7449_, new_n4709_, new_n443_ );
or   ( new_n7450_, new_n4711_, new_n419_ );
and  ( new_n7451_, new_n7450_, new_n7449_ );
xor  ( new_n7452_, new_n7451_, new_n4295_ );
or   ( new_n7453_, new_n4302_, new_n515_ );
or   ( new_n7454_, new_n4304_, new_n509_ );
and  ( new_n7455_, new_n7454_, new_n7453_ );
xor  ( new_n7456_, new_n7455_, new_n3895_ );
or   ( new_n7457_, new_n7456_, new_n7452_ );
and  ( new_n7458_, new_n7456_, new_n7452_ );
or   ( new_n7459_, new_n3896_, new_n805_ );
or   ( new_n7460_, new_n3898_, new_n775_ );
and  ( new_n7461_, new_n7460_, new_n7459_ );
xor  ( new_n7462_, new_n7461_, new_n3460_ );
or   ( new_n7463_, new_n7462_, new_n7458_ );
and  ( new_n7464_, new_n7463_, new_n7457_ );
or   ( new_n7465_, new_n6173_, new_n301_ );
or   ( new_n7466_, new_n6175_, new_n279_ );
and  ( new_n7467_, new_n7466_, new_n7465_ );
xor  ( new_n7468_, new_n7467_, new_n5597_ );
or   ( new_n7469_, new_n5604_, new_n270_ );
or   ( new_n7470_, new_n5606_, new_n294_ );
and  ( new_n7471_, new_n7470_, new_n7469_ );
xor  ( new_n7472_, new_n7471_, new_n5206_ );
or   ( new_n7473_, new_n7472_, new_n7468_ );
and  ( new_n7474_, new_n7472_, new_n7468_ );
or   ( new_n7475_, new_n5207_, new_n348_ );
or   ( new_n7476_, new_n5209_, new_n264_ );
and  ( new_n7477_, new_n7476_, new_n7475_ );
xor  ( new_n7478_, new_n7477_, new_n4708_ );
or   ( new_n7479_, new_n7478_, new_n7474_ );
and  ( new_n7480_, new_n7479_, new_n7473_ );
or   ( new_n7481_, new_n7480_, new_n7464_ );
and  ( new_n7482_, new_n7480_, new_n7464_ );
or   ( new_n7483_, new_n7184_, new_n319_ );
or   ( new_n7484_, new_n7186_, new_n333_ );
and  ( new_n7485_, new_n7484_, new_n7483_ );
xor  ( new_n7486_, new_n7485_, new_n6637_ );
xor  ( new_n7487_, RIbb2dcc0_55, RIbb2dd38_54 );
xor  ( new_n7488_, RIbb2dd38_54, new_n7174_ );
nor  ( new_n7489_, new_n7488_, new_n7487_ );
and  ( new_n7490_, new_n7489_, RIbb2d810_65 );
xor  ( new_n7491_, new_n7490_, new_n7177_ );
and  ( new_n7492_, new_n7491_, new_n7486_ );
nor  ( new_n7493_, new_n7491_, new_n7486_ );
or   ( new_n7494_, new_n6645_, new_n285_ );
or   ( new_n7495_, new_n6647_, new_n313_ );
and  ( new_n7496_, new_n7495_, new_n7494_ );
xor  ( new_n7497_, new_n7496_, new_n6166_ );
nor  ( new_n7498_, new_n7497_, new_n7493_ );
nor  ( new_n7499_, new_n7498_, new_n7492_ );
or   ( new_n7500_, new_n7499_, new_n7482_ );
and  ( new_n7501_, new_n7500_, new_n7481_ );
or   ( new_n7502_, new_n7501_, new_n7448_ );
or   ( new_n7503_, new_n3461_, new_n986_ );
or   ( new_n7504_, new_n3463_, new_n886_ );
and  ( new_n7505_, new_n7504_, new_n7503_ );
xor  ( new_n7506_, new_n7505_, new_n3116_ );
or   ( new_n7507_, new_n3117_, new_n1213_ );
or   ( new_n7508_, new_n3119_, new_n1168_ );
and  ( new_n7509_, new_n7508_, new_n7507_ );
xor  ( new_n7510_, new_n7509_, new_n2800_ );
or   ( new_n7511_, new_n7510_, new_n7506_ );
and  ( new_n7512_, new_n7510_, new_n7506_ );
or   ( new_n7513_, new_n2807_, new_n1525_ );
or   ( new_n7514_, new_n2809_, new_n1318_ );
and  ( new_n7515_, new_n7514_, new_n7513_ );
xor  ( new_n7516_, new_n7515_, new_n2424_ );
or   ( new_n7517_, new_n7516_, new_n7512_ );
and  ( new_n7518_, new_n7517_, new_n7511_ );
or   ( new_n7519_, new_n1593_, new_n2646_ );
or   ( new_n7520_, new_n1595_, new_n2475_ );
and  ( new_n7521_, new_n7520_, new_n7519_ );
xor  ( new_n7522_, new_n7521_, new_n1358_ );
or   ( new_n7523_, new_n1364_, new_n2981_ );
or   ( new_n7524_, new_n1366_, new_n2751_ );
and  ( new_n7525_, new_n7524_, new_n7523_ );
xor  ( new_n7526_, new_n7525_, new_n1129_ );
or   ( new_n7527_, new_n7526_, new_n7522_ );
and  ( new_n7528_, new_n7526_, new_n7522_ );
or   ( new_n7529_, new_n1135_, new_n3306_ );
or   ( new_n7530_, new_n1137_, new_n3178_ );
and  ( new_n7531_, new_n7530_, new_n7529_ );
xor  ( new_n7532_, new_n7531_, new_n896_ );
or   ( new_n7533_, new_n7532_, new_n7528_ );
and  ( new_n7534_, new_n7533_, new_n7527_ );
or   ( new_n7535_, new_n7534_, new_n7518_ );
and  ( new_n7536_, new_n7534_, new_n7518_ );
or   ( new_n7537_, new_n2425_, new_n1754_ );
or   ( new_n7538_, new_n2427_, new_n1523_ );
and  ( new_n7539_, new_n7538_, new_n7537_ );
xor  ( new_n7540_, new_n7539_, new_n2121_ );
or   ( new_n7541_, new_n2122_, new_n2057_ );
or   ( new_n7542_, new_n2124_, new_n1899_ );
and  ( new_n7543_, new_n7542_, new_n7541_ );
xor  ( new_n7544_, new_n7543_, new_n1843_ );
nor  ( new_n7545_, new_n7544_, new_n7540_ );
and  ( new_n7546_, new_n7544_, new_n7540_ );
or   ( new_n7547_, new_n1844_, new_n2291_ );
or   ( new_n7548_, new_n1846_, new_n2178_ );
and  ( new_n7549_, new_n7548_, new_n7547_ );
xor  ( new_n7550_, new_n7549_, new_n1586_ );
nor  ( new_n7551_, new_n7550_, new_n7546_ );
nor  ( new_n7552_, new_n7551_, new_n7545_ );
or   ( new_n7553_, new_n7552_, new_n7536_ );
and  ( new_n7554_, new_n7553_, new_n7535_ );
and  ( new_n7555_, new_n7501_, new_n7448_ );
or   ( new_n7556_, new_n7555_, new_n7554_ );
and  ( new_n7557_, new_n7556_, new_n7502_ );
or   ( new_n7558_, new_n7557_, new_n7396_ );
and  ( new_n7559_, new_n7557_, new_n7396_ );
xor  ( new_n7560_, new_n6912_, new_n6907_ );
xor  ( new_n7561_, new_n7560_, new_n6918_ );
xnor ( new_n7562_, new_n7300_, new_n7298_ );
xor  ( new_n7563_, new_n7562_, new_n7304_ );
and  ( new_n7564_, new_n7563_, new_n7561_ );
or   ( new_n7565_, new_n7563_, new_n7561_ );
xor  ( new_n7566_, new_n7288_, new_n7286_ );
xnor ( new_n7567_, new_n7566_, new_n7292_ );
and  ( new_n7568_, new_n7567_, new_n7565_ );
or   ( new_n7569_, new_n7568_, new_n7564_ );
or   ( new_n7570_, new_n7569_, new_n7559_ );
and  ( new_n7571_, new_n7570_, new_n7558_ );
and  ( new_n7572_, new_n7571_, new_n7361_ );
nor  ( new_n7573_, new_n7571_, new_n7361_ );
xnor ( new_n7574_, new_n7271_, new_n7269_ );
xor  ( new_n7575_, new_n7574_, new_n7275_ );
xor  ( new_n7576_, new_n7316_, new_n7314_ );
xor  ( new_n7577_, new_n7576_, new_n7320_ );
and  ( new_n7578_, new_n7577_, new_n7575_ );
nor  ( new_n7579_, new_n7577_, new_n7575_ );
xor  ( new_n7580_, new_n7245_, new_n7229_ );
xor  ( new_n7581_, new_n7580_, new_n7263_ );
xnor ( new_n7582_, new_n7136_, new_n7120_ );
xor  ( new_n7583_, new_n7582_, new_n7155_ );
nor  ( new_n7584_, new_n7583_, new_n7581_ );
and  ( new_n7585_, new_n7583_, new_n7581_ );
xor  ( new_n7586_, new_n7283_, new_n7281_ );
nor  ( new_n7587_, new_n7586_, new_n7585_ );
nor  ( new_n7588_, new_n7587_, new_n7584_ );
nor  ( new_n7589_, new_n7588_, new_n7579_ );
nor  ( new_n7590_, new_n7589_, new_n7578_ );
nor  ( new_n7591_, new_n7590_, new_n7573_ );
nor  ( new_n7592_, new_n7591_, new_n7572_ );
nor  ( new_n7593_, new_n7592_, new_n7355_ );
or   ( new_n7594_, new_n7593_, new_n7354_ );
xnor ( new_n7595_, new_n7043_, new_n6834_ );
xor  ( new_n7596_, new_n7595_, new_n7063_ );
or   ( new_n7597_, new_n7596_, new_n7594_ );
and  ( new_n7598_, new_n7596_, new_n7594_ );
xor  ( new_n7599_, new_n7097_, new_n7088_ );
xnor ( new_n7600_, new_n7599_, new_n7333_ );
or   ( new_n7601_, new_n7600_, new_n7598_ );
and  ( new_n7602_, new_n7601_, new_n7597_ );
xnor ( new_n7603_, new_n7084_, new_n7082_ );
xor  ( new_n7604_, new_n7603_, new_n7335_ );
and  ( new_n7605_, new_n7604_, new_n7602_ );
xor  ( new_n7606_, new_n7339_, new_n7337_ );
and  ( new_n7607_, new_n7606_, new_n7605_ );
xnor ( new_n7608_, new_n7310_, new_n7104_ );
xor  ( new_n7609_, new_n7608_, new_n7331_ );
xor  ( new_n7610_, new_n7348_, new_n7346_ );
xor  ( new_n7611_, new_n7610_, new_n7351_ );
xor  ( new_n7612_, new_n7557_, new_n7396_ );
xor  ( new_n7613_, new_n7612_, new_n7569_ );
xnor ( new_n7614_, new_n7577_, new_n7575_ );
xor  ( new_n7615_, new_n7614_, new_n7588_ );
nand ( new_n7616_, new_n7615_, new_n7613_ );
or   ( new_n7617_, new_n7615_, new_n7613_ );
xor  ( new_n7618_, new_n7360_, new_n7358_ );
nand ( new_n7619_, new_n7618_, new_n7617_ );
and  ( new_n7620_, new_n7619_, new_n7616_ );
nand ( new_n7621_, new_n7620_, new_n7611_ );
or   ( new_n7622_, new_n7620_, new_n7611_ );
xor  ( new_n7623_, new_n7501_, new_n7448_ );
xor  ( new_n7624_, new_n7623_, new_n7554_ );
xor  ( new_n7625_, new_n7382_, new_n7372_ );
xor  ( new_n7626_, new_n7625_, new_n7394_ );
nand ( new_n7627_, new_n7626_, new_n7624_ );
nor  ( new_n7628_, new_n7626_, new_n7624_ );
xor  ( new_n7629_, new_n7563_, new_n7561_ );
xnor ( new_n7630_, new_n7629_, new_n7567_ );
or   ( new_n7631_, new_n7630_, new_n7628_ );
and  ( new_n7632_, new_n7631_, new_n7627_ );
xnor ( new_n7633_, new_n7191_, new_n7173_ );
xor  ( new_n7634_, new_n7633_, new_n7209_ );
xnor ( new_n7635_, new_n7428_, new_n7412_ );
xor  ( new_n7636_, new_n7635_, new_n7446_ );
xnor ( new_n7637_, new_n7534_, new_n7518_ );
xor  ( new_n7638_, new_n7637_, new_n7552_ );
or   ( new_n7639_, new_n7638_, new_n7636_ );
and  ( new_n7640_, new_n7638_, new_n7636_ );
xor  ( new_n7641_, new_n7376_, new_n7374_ );
xor  ( new_n7642_, new_n7641_, new_n7380_ );
or   ( new_n7643_, new_n7642_, new_n7640_ );
and  ( new_n7644_, new_n7643_, new_n7639_ );
or   ( new_n7645_, new_n7644_, new_n7634_ );
and  ( new_n7646_, new_n7644_, new_n7634_ );
xor  ( new_n7647_, new_n7583_, new_n7581_ );
xor  ( new_n7648_, new_n7647_, new_n7586_ );
or   ( new_n7649_, new_n7648_, new_n7646_ );
and  ( new_n7650_, new_n7649_, new_n7645_ );
nor  ( new_n7651_, new_n7650_, new_n7632_ );
and  ( new_n7652_, new_n7650_, new_n7632_ );
or   ( new_n7653_, new_n317_, new_n6219_ );
or   ( new_n7654_, new_n320_, new_n5899_ );
and  ( new_n7655_, new_n7654_, new_n7653_ );
xor  ( new_n7656_, new_n7655_, new_n312_ );
or   ( new_n7657_, new_n283_, new_n6589_ );
or   ( new_n7658_, new_n286_, new_n6425_ );
and  ( new_n7659_, new_n7658_, new_n7657_ );
xor  ( new_n7660_, new_n7659_, new_n278_ );
or   ( new_n7661_, new_n7660_, new_n7656_ );
and  ( new_n7662_, new_n7660_, new_n7656_ );
or   ( new_n7663_, new_n299_, new_n7149_ );
or   ( new_n7664_, new_n302_, new_n6943_ );
and  ( new_n7665_, new_n7664_, new_n7663_ );
xor  ( new_n7666_, new_n7665_, new_n293_ );
or   ( new_n7667_, new_n7666_, new_n7662_ );
and  ( new_n7668_, new_n7667_, new_n7661_ );
or   ( new_n7669_, new_n524_, new_n4995_ );
or   ( new_n7670_, new_n526_, new_n4603_ );
and  ( new_n7671_, new_n7670_, new_n7669_ );
xor  ( new_n7672_, new_n7671_, new_n403_ );
or   ( new_n7673_, new_n409_, new_n5171_ );
or   ( new_n7674_, new_n411_, new_n4859_ );
and  ( new_n7675_, new_n7674_, new_n7673_ );
xor  ( new_n7676_, new_n7675_, new_n328_ );
or   ( new_n7677_, new_n7676_, new_n7672_ );
and  ( new_n7678_, new_n7676_, new_n7672_ );
or   ( new_n7679_, new_n337_, new_n5570_ );
or   ( new_n7680_, new_n340_, new_n5428_ );
and  ( new_n7681_, new_n7680_, new_n7679_ );
xor  ( new_n7682_, new_n7681_, new_n332_ );
or   ( new_n7683_, new_n7682_, new_n7678_ );
and  ( new_n7684_, new_n7683_, new_n7677_ );
or   ( new_n7685_, new_n7684_, new_n7668_ );
and  ( new_n7686_, new_n7684_, new_n7668_ );
or   ( new_n7687_, new_n1135_, new_n3696_ );
or   ( new_n7688_, new_n1137_, new_n3306_ );
and  ( new_n7689_, new_n7688_, new_n7687_ );
xor  ( new_n7690_, new_n7689_, new_n896_ );
or   ( new_n7691_, new_n897_, new_n3820_ );
or   ( new_n7692_, new_n899_, new_n3694_ );
and  ( new_n7693_, new_n7692_, new_n7691_ );
xor  ( new_n7694_, new_n7693_, new_n748_ );
nor  ( new_n7695_, new_n7694_, new_n7690_ );
and  ( new_n7696_, new_n7694_, new_n7690_ );
or   ( new_n7697_, new_n755_, new_n4267_ );
or   ( new_n7698_, new_n757_, new_n4069_ );
and  ( new_n7699_, new_n7698_, new_n7697_ );
xor  ( new_n7700_, new_n7699_, new_n523_ );
nor  ( new_n7701_, new_n7700_, new_n7696_ );
nor  ( new_n7702_, new_n7701_, new_n7695_ );
or   ( new_n7703_, new_n7702_, new_n7686_ );
and  ( new_n7704_, new_n7703_, new_n7685_ );
or   ( new_n7705_, new_n5207_, new_n419_ );
or   ( new_n7706_, new_n5209_, new_n348_ );
and  ( new_n7707_, new_n7706_, new_n7705_ );
xor  ( new_n7708_, new_n7707_, new_n4708_ );
or   ( new_n7709_, new_n4709_, new_n509_ );
or   ( new_n7710_, new_n4711_, new_n443_ );
and  ( new_n7711_, new_n7710_, new_n7709_ );
xor  ( new_n7712_, new_n7711_, new_n4295_ );
nor  ( new_n7713_, new_n7712_, new_n7708_ );
nand ( new_n7714_, new_n7712_, new_n7708_ );
or   ( new_n7715_, new_n4302_, new_n775_ );
or   ( new_n7716_, new_n4304_, new_n515_ );
and  ( new_n7717_, new_n7716_, new_n7715_ );
xor  ( new_n7718_, new_n7717_, new_n3895_ );
not  ( new_n7719_, new_n7718_ );
and  ( new_n7720_, new_n7719_, new_n7714_ );
or   ( new_n7721_, new_n7720_, new_n7713_ );
not  ( new_n7722_, RIbb2dcc0_55 );
and  ( new_n7723_, RIbb2dbd0_57, RIbb2dc48_56 );
nor  ( new_n7724_, new_n7723_, new_n7722_ );
not  ( new_n7725_, new_n7724_ );
or   ( new_n7726_, new_n7184_, new_n313_ );
or   ( new_n7727_, new_n7186_, new_n319_ );
and  ( new_n7728_, new_n7727_, new_n7726_ );
xor  ( new_n7729_, new_n7728_, new_n6638_ );
nand ( new_n7730_, new_n7729_, new_n7725_ );
or   ( new_n7731_, new_n7729_, new_n7725_ );
not  ( new_n7732_, new_n7489_ );
or   ( new_n7733_, new_n7732_, new_n333_ );
not  ( new_n7734_, new_n7487_ );
or   ( new_n7735_, new_n7734_, new_n339_ );
and  ( new_n7736_, new_n7735_, new_n7733_ );
xor  ( new_n7737_, new_n7736_, new_n7177_ );
nand ( new_n7738_, new_n7737_, new_n7731_ );
and  ( new_n7739_, new_n7738_, new_n7730_ );
nand ( new_n7740_, new_n7739_, new_n7721_ );
nor  ( new_n7741_, new_n7739_, new_n7721_ );
or   ( new_n7742_, new_n6645_, new_n279_ );
or   ( new_n7743_, new_n6647_, new_n285_ );
and  ( new_n7744_, new_n7743_, new_n7742_ );
xor  ( new_n7745_, new_n7744_, new_n6166_ );
or   ( new_n7746_, new_n6173_, new_n294_ );
or   ( new_n7747_, new_n6175_, new_n301_ );
and  ( new_n7748_, new_n7747_, new_n7746_ );
xor  ( new_n7749_, new_n7748_, new_n5597_ );
nor  ( new_n7750_, new_n7749_, new_n7745_ );
and  ( new_n7751_, new_n7749_, new_n7745_ );
or   ( new_n7752_, new_n5604_, new_n264_ );
or   ( new_n7753_, new_n5606_, new_n270_ );
and  ( new_n7754_, new_n7753_, new_n7752_ );
xor  ( new_n7755_, new_n7754_, new_n5206_ );
nor  ( new_n7756_, new_n7755_, new_n7751_ );
nor  ( new_n7757_, new_n7756_, new_n7750_ );
or   ( new_n7758_, new_n7757_, new_n7741_ );
and  ( new_n7759_, new_n7758_, new_n7740_ );
or   ( new_n7760_, new_n7759_, new_n7704_ );
and  ( new_n7761_, new_n7759_, new_n7704_ );
or   ( new_n7762_, new_n3896_, new_n886_ );
or   ( new_n7763_, new_n3898_, new_n805_ );
and  ( new_n7764_, new_n7763_, new_n7762_ );
xor  ( new_n7765_, new_n7764_, new_n3460_ );
or   ( new_n7766_, new_n3461_, new_n1168_ );
or   ( new_n7767_, new_n3463_, new_n986_ );
and  ( new_n7768_, new_n7767_, new_n7766_ );
xor  ( new_n7769_, new_n7768_, new_n3116_ );
or   ( new_n7770_, new_n7769_, new_n7765_ );
and  ( new_n7771_, new_n7769_, new_n7765_ );
or   ( new_n7772_, new_n3117_, new_n1318_ );
or   ( new_n7773_, new_n3119_, new_n1213_ );
and  ( new_n7774_, new_n7773_, new_n7772_ );
xor  ( new_n7775_, new_n7774_, new_n2800_ );
or   ( new_n7776_, new_n7775_, new_n7771_ );
and  ( new_n7777_, new_n7776_, new_n7770_ );
or   ( new_n7778_, new_n1844_, new_n2475_ );
or   ( new_n7779_, new_n1846_, new_n2291_ );
and  ( new_n7780_, new_n7779_, new_n7778_ );
xor  ( new_n7781_, new_n7780_, new_n1586_ );
or   ( new_n7782_, new_n1593_, new_n2751_ );
or   ( new_n7783_, new_n1595_, new_n2646_ );
and  ( new_n7784_, new_n7783_, new_n7782_ );
xor  ( new_n7785_, new_n7784_, new_n1358_ );
or   ( new_n7786_, new_n7785_, new_n7781_ );
and  ( new_n7787_, new_n7785_, new_n7781_ );
or   ( new_n7788_, new_n1364_, new_n3178_ );
or   ( new_n7789_, new_n1366_, new_n2981_ );
and  ( new_n7790_, new_n7789_, new_n7788_ );
xor  ( new_n7791_, new_n7790_, new_n1129_ );
or   ( new_n7792_, new_n7791_, new_n7787_ );
and  ( new_n7793_, new_n7792_, new_n7786_ );
nor  ( new_n7794_, new_n7793_, new_n7777_ );
and  ( new_n7795_, new_n7793_, new_n7777_ );
or   ( new_n7796_, new_n2807_, new_n1523_ );
or   ( new_n7797_, new_n2809_, new_n1525_ );
and  ( new_n7798_, new_n7797_, new_n7796_ );
xor  ( new_n7799_, new_n7798_, new_n2424_ );
or   ( new_n7800_, new_n2425_, new_n1899_ );
or   ( new_n7801_, new_n2427_, new_n1754_ );
and  ( new_n7802_, new_n7801_, new_n7800_ );
xor  ( new_n7803_, new_n7802_, new_n2121_ );
nor  ( new_n7804_, new_n7803_, new_n7799_ );
and  ( new_n7805_, new_n7803_, new_n7799_ );
or   ( new_n7806_, new_n2122_, new_n2178_ );
or   ( new_n7807_, new_n2124_, new_n2057_ );
and  ( new_n7808_, new_n7807_, new_n7806_ );
xor  ( new_n7809_, new_n7808_, new_n1843_ );
nor  ( new_n7810_, new_n7809_, new_n7805_ );
nor  ( new_n7811_, new_n7810_, new_n7804_ );
nor  ( new_n7812_, new_n7811_, new_n7795_ );
nor  ( new_n7813_, new_n7812_, new_n7794_ );
or   ( new_n7814_, new_n7813_, new_n7761_ );
and  ( new_n7815_, new_n7814_, new_n7760_ );
xor  ( new_n7816_, new_n7388_, new_n7386_ );
xor  ( new_n7817_, new_n7816_, new_n7392_ );
xor  ( new_n7818_, new_n7181_, new_n7177_ );
xor  ( new_n7819_, new_n7818_, new_n7189_ );
or   ( new_n7820_, new_n7819_, new_n7817_ );
and  ( new_n7821_, new_n7819_, new_n7817_ );
xor  ( new_n7822_, new_n7365_, new_n7363_ );
xor  ( new_n7823_, new_n7822_, new_n7370_ );
or   ( new_n7824_, new_n7823_, new_n7821_ );
and  ( new_n7825_, new_n7824_, new_n7820_ );
and  ( new_n7826_, new_n7825_, new_n7815_ );
nor  ( new_n7827_, new_n7825_, new_n7815_ );
and  ( new_n7828_, RIbb2bf38_118, RIbb2f610_1 );
not  ( new_n7829_, new_n7828_ );
xnor ( new_n7830_, new_n7404_, new_n7400_ );
xor  ( new_n7831_, new_n7830_, new_n7410_ );
and  ( new_n7832_, new_n7831_, new_n7829_ );
xnor ( new_n7833_, new_n7456_, new_n7452_ );
xor  ( new_n7834_, new_n7833_, new_n7462_ );
xnor ( new_n7835_, new_n7510_, new_n7506_ );
xor  ( new_n7836_, new_n7835_, new_n7516_ );
or   ( new_n7837_, new_n7836_, new_n7834_ );
and  ( new_n7838_, new_n7836_, new_n7834_ );
xor  ( new_n7839_, new_n7544_, new_n7540_ );
xnor ( new_n7840_, new_n7839_, new_n7550_ );
or   ( new_n7841_, new_n7840_, new_n7838_ );
and  ( new_n7842_, new_n7841_, new_n7837_ );
nor  ( new_n7843_, new_n7842_, new_n7832_ );
and  ( new_n7844_, new_n7842_, new_n7832_ );
xnor ( new_n7845_, new_n7420_, new_n7416_ );
xor  ( new_n7846_, new_n7845_, new_n7426_ );
xnor ( new_n7847_, new_n7526_, new_n7522_ );
xor  ( new_n7848_, new_n7847_, new_n7532_ );
nor  ( new_n7849_, new_n7848_, new_n7846_ );
and  ( new_n7850_, new_n7848_, new_n7846_ );
xor  ( new_n7851_, new_n7438_, new_n7434_ );
xnor ( new_n7852_, new_n7851_, new_n7444_ );
nor  ( new_n7853_, new_n7852_, new_n7850_ );
nor  ( new_n7854_, new_n7853_, new_n7849_ );
nor  ( new_n7855_, new_n7854_, new_n7844_ );
nor  ( new_n7856_, new_n7855_, new_n7843_ );
nor  ( new_n7857_, new_n7856_, new_n7827_ );
nor  ( new_n7858_, new_n7857_, new_n7826_ );
nor  ( new_n7859_, new_n7858_, new_n7652_ );
nor  ( new_n7860_, new_n7859_, new_n7651_ );
nand ( new_n7861_, new_n7860_, new_n7622_ );
and  ( new_n7862_, new_n7861_, new_n7621_ );
nor  ( new_n7863_, new_n7862_, new_n7609_ );
nand ( new_n7864_, new_n7862_, new_n7609_ );
xor  ( new_n7865_, new_n7353_, new_n7344_ );
xor  ( new_n7866_, new_n7865_, new_n7592_ );
and  ( new_n7867_, new_n7866_, new_n7864_ );
or   ( new_n7868_, new_n7867_, new_n7863_ );
xnor ( new_n7869_, new_n7596_, new_n7594_ );
xor  ( new_n7870_, new_n7869_, new_n7600_ );
nor  ( new_n7871_, new_n7870_, new_n7868_ );
xor  ( new_n7872_, new_n7604_, new_n7602_ );
and  ( new_n7873_, new_n7872_, new_n7871_ );
xor  ( new_n7874_, new_n7862_, new_n7609_ );
xor  ( new_n7875_, new_n7874_, new_n7866_ );
xor  ( new_n7876_, new_n7571_, new_n7361_ );
xor  ( new_n7877_, new_n7876_, new_n7590_ );
xnor ( new_n7878_, new_n7626_, new_n7624_ );
xor  ( new_n7879_, new_n7878_, new_n7630_ );
xnor ( new_n7880_, new_n7825_, new_n7815_ );
xor  ( new_n7881_, new_n7880_, new_n7856_ );
or   ( new_n7882_, new_n7881_, new_n7879_ );
and  ( new_n7883_, new_n7881_, new_n7879_ );
xor  ( new_n7884_, new_n7644_, new_n7634_ );
xnor ( new_n7885_, new_n7884_, new_n7648_ );
or   ( new_n7886_, new_n7885_, new_n7883_ );
and  ( new_n7887_, new_n7886_, new_n7882_ );
xnor ( new_n7888_, new_n7848_, new_n7846_ );
xor  ( new_n7889_, new_n7888_, new_n7852_ );
xnor ( new_n7890_, new_n7836_, new_n7834_ );
xor  ( new_n7891_, new_n7890_, new_n7840_ );
nor  ( new_n7892_, new_n7891_, new_n7889_ );
nand ( new_n7893_, new_n7891_, new_n7889_ );
xor  ( new_n7894_, new_n7831_, new_n7829_ );
and  ( new_n7895_, new_n7894_, new_n7893_ );
or   ( new_n7896_, new_n7895_, new_n7892_ );
xnor ( new_n7897_, new_n7480_, new_n7464_ );
xor  ( new_n7898_, new_n7897_, new_n7499_ );
nor  ( new_n7899_, new_n7898_, new_n7896_ );
and  ( new_n7900_, new_n7898_, new_n7896_ );
xnor ( new_n7901_, new_n7793_, new_n7777_ );
xor  ( new_n7902_, new_n7901_, new_n7811_ );
xnor ( new_n7903_, new_n7739_, new_n7721_ );
xor  ( new_n7904_, new_n7903_, new_n7757_ );
nor  ( new_n7905_, new_n7904_, new_n7902_ );
and  ( new_n7906_, new_n7904_, new_n7902_ );
xor  ( new_n7907_, new_n7684_, new_n7668_ );
xnor ( new_n7908_, new_n7907_, new_n7702_ );
nor  ( new_n7909_, new_n7908_, new_n7906_ );
nor  ( new_n7910_, new_n7909_, new_n7905_ );
nor  ( new_n7911_, new_n7910_, new_n7900_ );
or   ( new_n7912_, new_n7911_, new_n7899_ );
xor  ( new_n7913_, new_n7749_, new_n7745_ );
xor  ( new_n7914_, new_n7913_, new_n7755_ );
xor  ( new_n7915_, new_n7729_, new_n7725_ );
xor  ( new_n7916_, new_n7915_, new_n7737_ );
nand ( new_n7917_, new_n7916_, new_n7914_ );
nor  ( new_n7918_, new_n7916_, new_n7914_ );
xor  ( new_n7919_, new_n7712_, new_n7708_ );
xor  ( new_n7920_, new_n7919_, new_n7719_ );
or   ( new_n7921_, new_n7920_, new_n7918_ );
and  ( new_n7922_, new_n7921_, new_n7917_ );
xnor ( new_n7923_, new_n7472_, new_n7468_ );
xor  ( new_n7924_, new_n7923_, new_n7478_ );
nor  ( new_n7925_, new_n7924_, new_n7922_ );
and  ( new_n7926_, new_n7924_, new_n7922_ );
xor  ( new_n7927_, new_n7491_, new_n7486_ );
xnor ( new_n7928_, new_n7927_, new_n7497_ );
nor  ( new_n7929_, new_n7928_, new_n7926_ );
or   ( new_n7930_, new_n7929_, new_n7925_ );
or   ( new_n7931_, new_n1844_, new_n2646_ );
or   ( new_n7932_, new_n1846_, new_n2475_ );
and  ( new_n7933_, new_n7932_, new_n7931_ );
xor  ( new_n7934_, new_n7933_, new_n1586_ );
or   ( new_n7935_, new_n1593_, new_n2981_ );
or   ( new_n7936_, new_n1595_, new_n2751_ );
and  ( new_n7937_, new_n7936_, new_n7935_ );
xor  ( new_n7938_, new_n7937_, new_n1358_ );
or   ( new_n7939_, new_n7938_, new_n7934_ );
and  ( new_n7940_, new_n7938_, new_n7934_ );
or   ( new_n7941_, new_n1364_, new_n3306_ );
or   ( new_n7942_, new_n1366_, new_n3178_ );
and  ( new_n7943_, new_n7942_, new_n7941_ );
xor  ( new_n7944_, new_n7943_, new_n1129_ );
or   ( new_n7945_, new_n7944_, new_n7940_ );
and  ( new_n7946_, new_n7945_, new_n7939_ );
or   ( new_n7947_, new_n2807_, new_n1754_ );
or   ( new_n7948_, new_n2809_, new_n1523_ );
and  ( new_n7949_, new_n7948_, new_n7947_ );
xor  ( new_n7950_, new_n7949_, new_n2424_ );
or   ( new_n7951_, new_n2425_, new_n2057_ );
or   ( new_n7952_, new_n2427_, new_n1899_ );
and  ( new_n7953_, new_n7952_, new_n7951_ );
xor  ( new_n7954_, new_n7953_, new_n2121_ );
or   ( new_n7955_, new_n7954_, new_n7950_ );
and  ( new_n7956_, new_n7954_, new_n7950_ );
or   ( new_n7957_, new_n2122_, new_n2291_ );
or   ( new_n7958_, new_n2124_, new_n2178_ );
and  ( new_n7959_, new_n7958_, new_n7957_ );
xor  ( new_n7960_, new_n7959_, new_n1843_ );
or   ( new_n7961_, new_n7960_, new_n7956_ );
and  ( new_n7962_, new_n7961_, new_n7955_ );
or   ( new_n7963_, new_n7962_, new_n7946_ );
and  ( new_n7964_, new_n7962_, new_n7946_ );
or   ( new_n7965_, new_n3896_, new_n986_ );
or   ( new_n7966_, new_n3898_, new_n886_ );
and  ( new_n7967_, new_n7966_, new_n7965_ );
xor  ( new_n7968_, new_n7967_, new_n3460_ );
or   ( new_n7969_, new_n3461_, new_n1213_ );
or   ( new_n7970_, new_n3463_, new_n1168_ );
and  ( new_n7971_, new_n7970_, new_n7969_ );
xor  ( new_n7972_, new_n7971_, new_n3116_ );
nor  ( new_n7973_, new_n7972_, new_n7968_ );
and  ( new_n7974_, new_n7972_, new_n7968_ );
or   ( new_n7975_, new_n3117_, new_n1525_ );
or   ( new_n7976_, new_n3119_, new_n1318_ );
and  ( new_n7977_, new_n7976_, new_n7975_ );
xor  ( new_n7978_, new_n7977_, new_n2800_ );
nor  ( new_n7979_, new_n7978_, new_n7974_ );
nor  ( new_n7980_, new_n7979_, new_n7973_ );
or   ( new_n7981_, new_n7980_, new_n7964_ );
and  ( new_n7982_, new_n7981_, new_n7963_ );
or   ( new_n7983_, new_n1135_, new_n3694_ );
or   ( new_n7984_, new_n1137_, new_n3696_ );
and  ( new_n7985_, new_n7984_, new_n7983_ );
xor  ( new_n7986_, new_n7985_, new_n896_ );
or   ( new_n7987_, new_n897_, new_n4069_ );
or   ( new_n7988_, new_n899_, new_n3820_ );
and  ( new_n7989_, new_n7988_, new_n7987_ );
xor  ( new_n7990_, new_n7989_, new_n748_ );
or   ( new_n7991_, new_n7990_, new_n7986_ );
and  ( new_n7992_, new_n7990_, new_n7986_ );
or   ( new_n7993_, new_n755_, new_n4603_ );
or   ( new_n7994_, new_n757_, new_n4267_ );
and  ( new_n7995_, new_n7994_, new_n7993_ );
xor  ( new_n7996_, new_n7995_, new_n523_ );
or   ( new_n7997_, new_n7996_, new_n7992_ );
and  ( new_n7998_, new_n7997_, new_n7991_ );
or   ( new_n7999_, new_n524_, new_n4859_ );
or   ( new_n8000_, new_n526_, new_n4995_ );
and  ( new_n8001_, new_n8000_, new_n7999_ );
xor  ( new_n8002_, new_n8001_, new_n403_ );
or   ( new_n8003_, new_n409_, new_n5428_ );
or   ( new_n8004_, new_n411_, new_n5171_ );
and  ( new_n8005_, new_n8004_, new_n8003_ );
xor  ( new_n8006_, new_n8005_, new_n328_ );
or   ( new_n8007_, new_n8006_, new_n8002_ );
and  ( new_n8008_, new_n8006_, new_n8002_ );
or   ( new_n8009_, new_n337_, new_n5899_ );
or   ( new_n8010_, new_n340_, new_n5570_ );
and  ( new_n8011_, new_n8010_, new_n8009_ );
xor  ( new_n8012_, new_n8011_, new_n332_ );
or   ( new_n8013_, new_n8012_, new_n8008_ );
and  ( new_n8014_, new_n8013_, new_n8007_ );
or   ( new_n8015_, new_n8014_, new_n7998_ );
and  ( new_n8016_, new_n8014_, new_n7998_ );
or   ( new_n8017_, new_n317_, new_n6425_ );
or   ( new_n8018_, new_n320_, new_n6219_ );
and  ( new_n8019_, new_n8018_, new_n8017_ );
xor  ( new_n8020_, new_n8019_, new_n312_ );
or   ( new_n8021_, new_n283_, new_n6943_ );
or   ( new_n8022_, new_n286_, new_n6589_ );
and  ( new_n8023_, new_n8022_, new_n8021_ );
xor  ( new_n8024_, new_n8023_, new_n278_ );
nor  ( new_n8025_, new_n8024_, new_n8020_ );
and  ( new_n8026_, new_n8024_, new_n8020_ );
or   ( new_n8027_, new_n299_, new_n7373_ );
or   ( new_n8028_, new_n302_, new_n7149_ );
and  ( new_n8029_, new_n8028_, new_n8027_ );
xor  ( new_n8030_, new_n8029_, new_n293_ );
nor  ( new_n8031_, new_n8030_, new_n8026_ );
nor  ( new_n8032_, new_n8031_, new_n8025_ );
or   ( new_n8033_, new_n8032_, new_n8016_ );
and  ( new_n8034_, new_n8033_, new_n8015_ );
or   ( new_n8035_, new_n8034_, new_n7982_ );
or   ( new_n8036_, new_n7732_, new_n319_ );
or   ( new_n8037_, new_n7734_, new_n333_ );
and  ( new_n8038_, new_n8037_, new_n8036_ );
xor  ( new_n8039_, new_n8038_, new_n7176_ );
xor  ( new_n8040_, RIbb2dbd0_57, RIbb2dc48_56 );
xor  ( new_n8041_, RIbb2dc48_56, new_n7722_ );
nor  ( new_n8042_, new_n8041_, new_n8040_ );
and  ( new_n8043_, new_n8042_, RIbb2d810_65 );
xor  ( new_n8044_, new_n8043_, new_n7725_ );
nand ( new_n8045_, new_n8044_, new_n8039_ );
nor  ( new_n8046_, new_n8044_, new_n8039_ );
or   ( new_n8047_, new_n7184_, new_n285_ );
or   ( new_n8048_, new_n7186_, new_n313_ );
and  ( new_n8049_, new_n8048_, new_n8047_ );
xor  ( new_n8050_, new_n8049_, new_n6638_ );
or   ( new_n8051_, new_n8050_, new_n8046_ );
and  ( new_n8052_, new_n8051_, new_n8045_ );
or   ( new_n8053_, new_n5207_, new_n443_ );
or   ( new_n8054_, new_n5209_, new_n419_ );
and  ( new_n8055_, new_n8054_, new_n8053_ );
xor  ( new_n8056_, new_n8055_, new_n4708_ );
or   ( new_n8057_, new_n4709_, new_n515_ );
or   ( new_n8058_, new_n4711_, new_n509_ );
and  ( new_n8059_, new_n8058_, new_n8057_ );
xor  ( new_n8060_, new_n8059_, new_n4295_ );
or   ( new_n8061_, new_n8060_, new_n8056_ );
and  ( new_n8062_, new_n8060_, new_n8056_ );
or   ( new_n8063_, new_n4302_, new_n805_ );
or   ( new_n8064_, new_n4304_, new_n775_ );
and  ( new_n8065_, new_n8064_, new_n8063_ );
xor  ( new_n8066_, new_n8065_, new_n3895_ );
or   ( new_n8067_, new_n8066_, new_n8062_ );
and  ( new_n8068_, new_n8067_, new_n8061_ );
nor  ( new_n8069_, new_n8068_, new_n8052_ );
and  ( new_n8070_, new_n8068_, new_n8052_ );
or   ( new_n8071_, new_n6645_, new_n301_ );
or   ( new_n8072_, new_n6647_, new_n279_ );
and  ( new_n8073_, new_n8072_, new_n8071_ );
xor  ( new_n8074_, new_n8073_, new_n6166_ );
or   ( new_n8075_, new_n6173_, new_n270_ );
or   ( new_n8076_, new_n6175_, new_n294_ );
and  ( new_n8077_, new_n8076_, new_n8075_ );
xor  ( new_n8078_, new_n8077_, new_n5597_ );
nor  ( new_n8079_, new_n8078_, new_n8074_ );
and  ( new_n8080_, new_n8078_, new_n8074_ );
or   ( new_n8081_, new_n5604_, new_n348_ );
or   ( new_n8082_, new_n5606_, new_n264_ );
and  ( new_n8083_, new_n8082_, new_n8081_ );
xor  ( new_n8084_, new_n8083_, new_n5206_ );
nor  ( new_n8085_, new_n8084_, new_n8080_ );
nor  ( new_n8086_, new_n8085_, new_n8079_ );
nor  ( new_n8087_, new_n8086_, new_n8070_ );
nor  ( new_n8088_, new_n8087_, new_n8069_ );
and  ( new_n8089_, new_n8034_, new_n7982_ );
or   ( new_n8090_, new_n8089_, new_n8088_ );
and  ( new_n8091_, new_n8090_, new_n8035_ );
or   ( new_n8092_, new_n8091_, new_n7930_ );
xnor ( new_n8093_, new_n7676_, new_n7672_ );
xor  ( new_n8094_, new_n8093_, new_n7682_ );
xnor ( new_n8095_, new_n7660_, new_n7656_ );
xor  ( new_n8096_, new_n8095_, new_n7666_ );
or   ( new_n8097_, new_n8096_, new_n8094_ );
and  ( new_n8098_, new_n8096_, new_n8094_ );
xor  ( new_n8099_, new_n7694_, new_n7690_ );
xnor ( new_n8100_, new_n8099_, new_n7700_ );
or   ( new_n8101_, new_n8100_, new_n8098_ );
and  ( new_n8102_, new_n8101_, new_n8097_ );
xnor ( new_n8103_, new_n7785_, new_n7781_ );
xor  ( new_n8104_, new_n8103_, new_n7791_ );
xnor ( new_n8105_, new_n7769_, new_n7765_ );
xor  ( new_n8106_, new_n8105_, new_n7775_ );
or   ( new_n8107_, new_n8106_, new_n8104_ );
and  ( new_n8108_, new_n8106_, new_n8104_ );
xor  ( new_n8109_, new_n7803_, new_n7799_ );
xnor ( new_n8110_, new_n8109_, new_n7809_ );
or   ( new_n8111_, new_n8110_, new_n8108_ );
and  ( new_n8112_, new_n8111_, new_n8107_ );
nor  ( new_n8113_, new_n8112_, new_n8102_ );
nand ( new_n8114_, new_n8112_, new_n8102_ );
not  ( new_n8115_, RIbb2bec0_119 );
or   ( new_n8116_, new_n268_, new_n8115_ );
not  ( new_n8117_, RIbb2bf38_118 );
or   ( new_n8118_, new_n271_, new_n8117_ );
and  ( new_n8119_, new_n8118_, new_n8116_ );
xor  ( new_n8120_, new_n8119_, new_n263_ );
and  ( new_n8121_, RIbb2be48_120, RIbb2f610_1 );
or   ( new_n8122_, new_n8121_, new_n8120_ );
or   ( new_n8123_, new_n268_, new_n8117_ );
or   ( new_n8124_, new_n271_, new_n7373_ );
and  ( new_n8125_, new_n8124_, new_n8123_ );
xor  ( new_n8126_, new_n8125_, new_n263_ );
nor  ( new_n8127_, new_n8126_, new_n8122_ );
and  ( new_n8128_, new_n8126_, new_n8122_ );
and  ( new_n8129_, RIbb2bec0_119, RIbb2f610_1 );
nor  ( new_n8130_, new_n8129_, new_n8128_ );
nor  ( new_n8131_, new_n8130_, new_n8127_ );
and  ( new_n8132_, new_n8131_, new_n8114_ );
or   ( new_n8133_, new_n8132_, new_n8113_ );
and  ( new_n8134_, new_n8091_, new_n7930_ );
or   ( new_n8135_, new_n8134_, new_n8133_ );
and  ( new_n8136_, new_n8135_, new_n8092_ );
or   ( new_n8137_, new_n8136_, new_n7912_ );
nand ( new_n8138_, new_n8136_, new_n7912_ );
xnor ( new_n8139_, new_n7842_, new_n7832_ );
xor  ( new_n8140_, new_n8139_, new_n7854_ );
xnor ( new_n8141_, new_n7638_, new_n7636_ );
xor  ( new_n8142_, new_n8141_, new_n7642_ );
and  ( new_n8143_, new_n8142_, new_n8140_ );
nor  ( new_n8144_, new_n8142_, new_n8140_ );
xor  ( new_n8145_, new_n7819_, new_n7817_ );
xnor ( new_n8146_, new_n8145_, new_n7823_ );
nor  ( new_n8147_, new_n8146_, new_n8144_ );
nor  ( new_n8148_, new_n8147_, new_n8143_ );
nand ( new_n8149_, new_n8148_, new_n8138_ );
and  ( new_n8150_, new_n8149_, new_n8137_ );
nand ( new_n8151_, new_n8150_, new_n7887_ );
or   ( new_n8152_, new_n8150_, new_n7887_ );
xor  ( new_n8153_, new_n7615_, new_n7613_ );
xor  ( new_n8154_, new_n8153_, new_n7618_ );
nand ( new_n8155_, new_n8154_, new_n8152_ );
and  ( new_n8156_, new_n8155_, new_n8151_ );
or   ( new_n8157_, new_n8156_, new_n7877_ );
and  ( new_n8158_, new_n8156_, new_n7877_ );
xor  ( new_n8159_, new_n7620_, new_n7611_ );
xor  ( new_n8160_, new_n8159_, new_n7860_ );
or   ( new_n8161_, new_n8160_, new_n8158_ );
and  ( new_n8162_, new_n8161_, new_n8157_ );
nor  ( new_n8163_, new_n8162_, new_n7875_ );
xor  ( new_n8164_, new_n7870_, new_n7868_ );
and  ( new_n8165_, new_n8164_, new_n8163_ );
xor  ( new_n8166_, new_n8150_, new_n7887_ );
xor  ( new_n8167_, new_n8166_, new_n8154_ );
xnor ( new_n8168_, new_n7650_, new_n7632_ );
xor  ( new_n8169_, new_n8168_, new_n7858_ );
and  ( new_n8170_, new_n8169_, new_n8167_ );
or   ( new_n8171_, new_n8169_, new_n8167_ );
xnor ( new_n8172_, new_n7881_, new_n7879_ );
xor  ( new_n8173_, new_n8172_, new_n7885_ );
xor  ( new_n8174_, new_n7898_, new_n7896_ );
xor  ( new_n8175_, new_n8174_, new_n7910_ );
xnor ( new_n8176_, new_n7759_, new_n7704_ );
xor  ( new_n8177_, new_n8176_, new_n7813_ );
or   ( new_n8178_, new_n8177_, new_n8175_ );
and  ( new_n8179_, new_n8177_, new_n8175_ );
xor  ( new_n8180_, new_n8142_, new_n8140_ );
xor  ( new_n8181_, new_n8180_, new_n8146_ );
or   ( new_n8182_, new_n8181_, new_n8179_ );
and  ( new_n8183_, new_n8182_, new_n8178_ );
nor  ( new_n8184_, new_n8183_, new_n8173_ );
nand ( new_n8185_, new_n8183_, new_n8173_ );
or   ( new_n8186_, new_n1364_, new_n3696_ );
or   ( new_n8187_, new_n1366_, new_n3306_ );
and  ( new_n8188_, new_n8187_, new_n8186_ );
xor  ( new_n8189_, new_n8188_, new_n1129_ );
or   ( new_n8190_, new_n1135_, new_n3820_ );
or   ( new_n8191_, new_n1137_, new_n3694_ );
and  ( new_n8192_, new_n8191_, new_n8190_ );
xor  ( new_n8193_, new_n8192_, new_n896_ );
or   ( new_n8194_, new_n8193_, new_n8189_ );
and  ( new_n8195_, new_n8193_, new_n8189_ );
or   ( new_n8196_, new_n897_, new_n4267_ );
or   ( new_n8197_, new_n899_, new_n4069_ );
and  ( new_n8198_, new_n8197_, new_n8196_ );
xor  ( new_n8199_, new_n8198_, new_n748_ );
or   ( new_n8200_, new_n8199_, new_n8195_ );
and  ( new_n8201_, new_n8200_, new_n8194_ );
or   ( new_n8202_, new_n755_, new_n4995_ );
or   ( new_n8203_, new_n757_, new_n4603_ );
and  ( new_n8204_, new_n8203_, new_n8202_ );
xor  ( new_n8205_, new_n8204_, new_n523_ );
or   ( new_n8206_, new_n524_, new_n5171_ );
or   ( new_n8207_, new_n526_, new_n4859_ );
and  ( new_n8208_, new_n8207_, new_n8206_ );
xor  ( new_n8209_, new_n8208_, new_n403_ );
or   ( new_n8210_, new_n8209_, new_n8205_ );
and  ( new_n8211_, new_n8209_, new_n8205_ );
or   ( new_n8212_, new_n409_, new_n5570_ );
or   ( new_n8213_, new_n411_, new_n5428_ );
and  ( new_n8214_, new_n8213_, new_n8212_ );
xor  ( new_n8215_, new_n8214_, new_n328_ );
or   ( new_n8216_, new_n8215_, new_n8211_ );
and  ( new_n8217_, new_n8216_, new_n8210_ );
or   ( new_n8218_, new_n8217_, new_n8201_ );
and  ( new_n8219_, new_n8217_, new_n8201_ );
or   ( new_n8220_, new_n337_, new_n6219_ );
or   ( new_n8221_, new_n340_, new_n5899_ );
and  ( new_n8222_, new_n8221_, new_n8220_ );
xor  ( new_n8223_, new_n8222_, new_n332_ );
or   ( new_n8224_, new_n317_, new_n6589_ );
or   ( new_n8225_, new_n320_, new_n6425_ );
and  ( new_n8226_, new_n8225_, new_n8224_ );
xor  ( new_n8227_, new_n8226_, new_n312_ );
or   ( new_n8228_, new_n8227_, new_n8223_ );
and  ( new_n8229_, new_n8227_, new_n8223_ );
or   ( new_n8230_, new_n283_, new_n7149_ );
or   ( new_n8231_, new_n286_, new_n6943_ );
and  ( new_n8232_, new_n8231_, new_n8230_ );
xor  ( new_n8233_, new_n8232_, new_n278_ );
or   ( new_n8234_, new_n8233_, new_n8229_ );
and  ( new_n8235_, new_n8234_, new_n8228_ );
or   ( new_n8236_, new_n8235_, new_n8219_ );
and  ( new_n8237_, new_n8236_, new_n8218_ );
or   ( new_n8238_, new_n7184_, new_n279_ );
or   ( new_n8239_, new_n7186_, new_n285_ );
and  ( new_n8240_, new_n8239_, new_n8238_ );
xor  ( new_n8241_, new_n8240_, new_n6638_ );
or   ( new_n8242_, new_n6645_, new_n294_ );
or   ( new_n8243_, new_n6647_, new_n301_ );
and  ( new_n8244_, new_n8243_, new_n8242_ );
xor  ( new_n8245_, new_n8244_, new_n6166_ );
nor  ( new_n8246_, new_n8245_, new_n8241_ );
nand ( new_n8247_, new_n8245_, new_n8241_ );
or   ( new_n8248_, new_n6173_, new_n264_ );
or   ( new_n8249_, new_n6175_, new_n270_ );
and  ( new_n8250_, new_n8249_, new_n8248_ );
xor  ( new_n8251_, new_n8250_, new_n5596_ );
and  ( new_n8252_, new_n8251_, new_n8247_ );
or   ( new_n8253_, new_n8252_, new_n8246_ );
not  ( new_n8254_, RIbb2dbd0_57 );
and  ( new_n8255_, RIbb2dae0_59, RIbb2db58_58 );
nor  ( new_n8256_, new_n8255_, new_n8254_ );
not  ( new_n8257_, new_n8256_ );
or   ( new_n8258_, new_n7732_, new_n313_ );
or   ( new_n8259_, new_n7734_, new_n319_ );
and  ( new_n8260_, new_n8259_, new_n8258_ );
xor  ( new_n8261_, new_n8260_, new_n7177_ );
nand ( new_n8262_, new_n8261_, new_n8257_ );
or   ( new_n8263_, new_n8261_, new_n8257_ );
not  ( new_n8264_, new_n8042_ );
or   ( new_n8265_, new_n8264_, new_n333_ );
not  ( new_n8266_, new_n8040_ );
or   ( new_n8267_, new_n8266_, new_n339_ );
and  ( new_n8268_, new_n8267_, new_n8265_ );
xor  ( new_n8269_, new_n8268_, new_n7725_ );
nand ( new_n8270_, new_n8269_, new_n8263_ );
and  ( new_n8271_, new_n8270_, new_n8262_ );
nand ( new_n8272_, new_n8271_, new_n8253_ );
nor  ( new_n8273_, new_n8271_, new_n8253_ );
or   ( new_n8274_, new_n5604_, new_n419_ );
or   ( new_n8275_, new_n5606_, new_n348_ );
and  ( new_n8276_, new_n8275_, new_n8274_ );
xor  ( new_n8277_, new_n8276_, new_n5206_ );
or   ( new_n8278_, new_n5207_, new_n509_ );
or   ( new_n8279_, new_n5209_, new_n443_ );
and  ( new_n8280_, new_n8279_, new_n8278_ );
xor  ( new_n8281_, new_n8280_, new_n4708_ );
nor  ( new_n8282_, new_n8281_, new_n8277_ );
and  ( new_n8283_, new_n8281_, new_n8277_ );
or   ( new_n8284_, new_n4709_, new_n775_ );
or   ( new_n8285_, new_n4711_, new_n515_ );
and  ( new_n8286_, new_n8285_, new_n8284_ );
xor  ( new_n8287_, new_n8286_, new_n4295_ );
nor  ( new_n8288_, new_n8287_, new_n8283_ );
nor  ( new_n8289_, new_n8288_, new_n8282_ );
or   ( new_n8290_, new_n8289_, new_n8273_ );
and  ( new_n8291_, new_n8290_, new_n8272_ );
nor  ( new_n8292_, new_n8291_, new_n8237_ );
and  ( new_n8293_, new_n8291_, new_n8237_ );
or   ( new_n8294_, new_n3117_, new_n1523_ );
or   ( new_n8295_, new_n3119_, new_n1525_ );
and  ( new_n8296_, new_n8295_, new_n8294_ );
xor  ( new_n8297_, new_n8296_, new_n2800_ );
or   ( new_n8298_, new_n2807_, new_n1899_ );
or   ( new_n8299_, new_n2809_, new_n1754_ );
and  ( new_n8300_, new_n8299_, new_n8298_ );
xor  ( new_n8301_, new_n8300_, new_n2424_ );
or   ( new_n8302_, new_n8301_, new_n8297_ );
and  ( new_n8303_, new_n8301_, new_n8297_ );
or   ( new_n8304_, new_n2425_, new_n2178_ );
or   ( new_n8305_, new_n2427_, new_n2057_ );
and  ( new_n8306_, new_n8305_, new_n8304_ );
xor  ( new_n8307_, new_n8306_, new_n2121_ );
or   ( new_n8308_, new_n8307_, new_n8303_ );
and  ( new_n8309_, new_n8308_, new_n8302_ );
or   ( new_n8310_, new_n2122_, new_n2475_ );
or   ( new_n8311_, new_n2124_, new_n2291_ );
and  ( new_n8312_, new_n8311_, new_n8310_ );
xor  ( new_n8313_, new_n8312_, new_n1843_ );
or   ( new_n8314_, new_n1844_, new_n2751_ );
or   ( new_n8315_, new_n1846_, new_n2646_ );
and  ( new_n8316_, new_n8315_, new_n8314_ );
xor  ( new_n8317_, new_n8316_, new_n1586_ );
or   ( new_n8318_, new_n8317_, new_n8313_ );
and  ( new_n8319_, new_n8317_, new_n8313_ );
or   ( new_n8320_, new_n1593_, new_n3178_ );
or   ( new_n8321_, new_n1595_, new_n2981_ );
and  ( new_n8322_, new_n8321_, new_n8320_ );
xor  ( new_n8323_, new_n8322_, new_n1358_ );
or   ( new_n8324_, new_n8323_, new_n8319_ );
and  ( new_n8325_, new_n8324_, new_n8318_ );
nor  ( new_n8326_, new_n8325_, new_n8309_ );
and  ( new_n8327_, new_n8325_, new_n8309_ );
or   ( new_n8328_, new_n4302_, new_n886_ );
or   ( new_n8329_, new_n4304_, new_n805_ );
and  ( new_n8330_, new_n8329_, new_n8328_ );
xor  ( new_n8331_, new_n8330_, new_n3895_ );
or   ( new_n8332_, new_n3896_, new_n1168_ );
or   ( new_n8333_, new_n3898_, new_n986_ );
and  ( new_n8334_, new_n8333_, new_n8332_ );
xor  ( new_n8335_, new_n8334_, new_n3460_ );
nor  ( new_n8336_, new_n8335_, new_n8331_ );
and  ( new_n8337_, new_n8335_, new_n8331_ );
or   ( new_n8338_, new_n3461_, new_n1318_ );
or   ( new_n8339_, new_n3463_, new_n1213_ );
and  ( new_n8340_, new_n8339_, new_n8338_ );
xor  ( new_n8341_, new_n8340_, new_n3116_ );
nor  ( new_n8342_, new_n8341_, new_n8337_ );
nor  ( new_n8343_, new_n8342_, new_n8336_ );
nor  ( new_n8344_, new_n8343_, new_n8327_ );
nor  ( new_n8345_, new_n8344_, new_n8326_ );
nor  ( new_n8346_, new_n8345_, new_n8293_ );
or   ( new_n8347_, new_n8346_, new_n8292_ );
or   ( new_n8348_, new_n299_, new_n8117_ );
or   ( new_n8349_, new_n302_, new_n7373_ );
and  ( new_n8350_, new_n8349_, new_n8348_ );
xor  ( new_n8351_, new_n8350_, new_n293_ );
not  ( new_n8352_, RIbb2be48_120 );
or   ( new_n8353_, new_n268_, new_n8352_ );
or   ( new_n8354_, new_n271_, new_n8115_ );
and  ( new_n8355_, new_n8354_, new_n8353_ );
xor  ( new_n8356_, new_n8355_, new_n263_ );
nor  ( new_n8357_, new_n8356_, new_n8351_ );
and  ( new_n8358_, RIbb2bdd0_121, RIbb2f610_1 );
not  ( new_n8359_, new_n8358_ );
nand ( new_n8360_, new_n8356_, new_n8351_ );
and  ( new_n8361_, new_n8360_, new_n8359_ );
or   ( new_n8362_, new_n8361_, new_n8357_ );
xnor ( new_n8363_, new_n8024_, new_n8020_ );
xor  ( new_n8364_, new_n8363_, new_n8030_ );
or   ( new_n8365_, new_n8364_, new_n8362_ );
and  ( new_n8366_, new_n8364_, new_n8362_ );
xor  ( new_n8367_, new_n8121_, new_n8120_ );
or   ( new_n8368_, new_n8367_, new_n8366_ );
and  ( new_n8369_, new_n8368_, new_n8365_ );
xnor ( new_n8370_, new_n7954_, new_n7950_ );
xor  ( new_n8371_, new_n8370_, new_n7960_ );
xnor ( new_n8372_, new_n8060_, new_n8056_ );
xor  ( new_n8373_, new_n8372_, new_n8066_ );
or   ( new_n8374_, new_n8373_, new_n8371_ );
and  ( new_n8375_, new_n8373_, new_n8371_ );
xor  ( new_n8376_, new_n7972_, new_n7968_ );
xnor ( new_n8377_, new_n8376_, new_n7978_ );
or   ( new_n8378_, new_n8377_, new_n8375_ );
and  ( new_n8379_, new_n8378_, new_n8374_ );
or   ( new_n8380_, new_n8379_, new_n8369_ );
and  ( new_n8381_, new_n8379_, new_n8369_ );
xnor ( new_n8382_, new_n7938_, new_n7934_ );
xor  ( new_n8383_, new_n8382_, new_n7944_ );
xnor ( new_n8384_, new_n8006_, new_n8002_ );
xor  ( new_n8385_, new_n8384_, new_n8012_ );
nor  ( new_n8386_, new_n8385_, new_n8383_ );
and  ( new_n8387_, new_n8385_, new_n8383_ );
xor  ( new_n8388_, new_n7990_, new_n7986_ );
xnor ( new_n8389_, new_n8388_, new_n7996_ );
nor  ( new_n8390_, new_n8389_, new_n8387_ );
nor  ( new_n8391_, new_n8390_, new_n8386_ );
or   ( new_n8392_, new_n8391_, new_n8381_ );
and  ( new_n8393_, new_n8392_, new_n8380_ );
and  ( new_n8394_, new_n8393_, new_n8347_ );
or   ( new_n8395_, new_n8393_, new_n8347_ );
xnor ( new_n8396_, new_n8096_, new_n8094_ );
xor  ( new_n8397_, new_n8396_, new_n8100_ );
xnor ( new_n8398_, new_n8106_, new_n8104_ );
xor  ( new_n8399_, new_n8398_, new_n8110_ );
nor  ( new_n8400_, new_n8399_, new_n8397_ );
nand ( new_n8401_, new_n8399_, new_n8397_ );
xor  ( new_n8402_, new_n7916_, new_n7914_ );
xnor ( new_n8403_, new_n8402_, new_n7920_ );
not  ( new_n8404_, new_n8403_ );
and  ( new_n8405_, new_n8404_, new_n8401_ );
or   ( new_n8406_, new_n8405_, new_n8400_ );
and  ( new_n8407_, new_n8406_, new_n8395_ );
or   ( new_n8408_, new_n8407_, new_n8394_ );
xnor ( new_n8409_, new_n8112_, new_n8102_ );
xor  ( new_n8410_, new_n8409_, new_n8131_ );
xnor ( new_n8411_, new_n8034_, new_n7982_ );
xor  ( new_n8412_, new_n8411_, new_n8088_ );
or   ( new_n8413_, new_n8412_, new_n8410_ );
and  ( new_n8414_, new_n8412_, new_n8410_ );
xor  ( new_n8415_, new_n7924_, new_n7922_ );
xor  ( new_n8416_, new_n8415_, new_n7928_ );
or   ( new_n8417_, new_n8416_, new_n8414_ );
and  ( new_n8418_, new_n8417_, new_n8413_ );
nor  ( new_n8419_, new_n8418_, new_n8408_ );
nand ( new_n8420_, new_n8418_, new_n8408_ );
xnor ( new_n8421_, new_n7891_, new_n7889_ );
xor  ( new_n8422_, new_n8421_, new_n7894_ );
xnor ( new_n8423_, new_n7904_, new_n7902_ );
xor  ( new_n8424_, new_n8423_, new_n7908_ );
and  ( new_n8425_, new_n8424_, new_n8422_ );
nor  ( new_n8426_, new_n8424_, new_n8422_ );
xnor ( new_n8427_, new_n7962_, new_n7946_ );
xor  ( new_n8428_, new_n8427_, new_n7980_ );
xnor ( new_n8429_, new_n8014_, new_n7998_ );
xor  ( new_n8430_, new_n8429_, new_n8032_ );
nor  ( new_n8431_, new_n8430_, new_n8428_ );
and  ( new_n8432_, new_n8430_, new_n8428_ );
xor  ( new_n8433_, new_n8126_, new_n8122_ );
xnor ( new_n8434_, new_n8433_, new_n8129_ );
nor  ( new_n8435_, new_n8434_, new_n8432_ );
nor  ( new_n8436_, new_n8435_, new_n8431_ );
nor  ( new_n8437_, new_n8436_, new_n8426_ );
nor  ( new_n8438_, new_n8437_, new_n8425_ );
not  ( new_n8439_, new_n8438_ );
and  ( new_n8440_, new_n8439_, new_n8420_ );
or   ( new_n8441_, new_n8440_, new_n8419_ );
and  ( new_n8442_, new_n8441_, new_n8185_ );
or   ( new_n8443_, new_n8442_, new_n8184_ );
and  ( new_n8444_, new_n8443_, new_n8171_ );
or   ( new_n8445_, new_n8444_, new_n8170_ );
xnor ( new_n8446_, new_n8156_, new_n7877_ );
xor  ( new_n8447_, new_n8446_, new_n8160_ );
and  ( new_n8448_, new_n8447_, new_n8445_ );
xor  ( new_n8449_, new_n8162_, new_n7875_ );
and  ( new_n8450_, new_n8449_, new_n8448_ );
xor  ( new_n8451_, new_n8418_, new_n8408_ );
xor  ( new_n8452_, new_n8451_, new_n8439_ );
not  ( new_n8453_, new_n8452_ );
xor  ( new_n8454_, new_n8177_, new_n8175_ );
xor  ( new_n8455_, new_n8454_, new_n8181_ );
nor  ( new_n8456_, new_n8455_, new_n8453_ );
xor  ( new_n8457_, new_n8091_, new_n7930_ );
xor  ( new_n8458_, new_n8457_, new_n8133_ );
xnor ( new_n8459_, new_n8068_, new_n8052_ );
xor  ( new_n8460_, new_n8459_, new_n8086_ );
xor  ( new_n8461_, new_n8217_, new_n8201_ );
xor  ( new_n8462_, new_n8461_, new_n8235_ );
xnor ( new_n8463_, new_n8385_, new_n8383_ );
xor  ( new_n8464_, new_n8463_, new_n8389_ );
nand ( new_n8465_, new_n8464_, new_n8462_ );
nor  ( new_n8466_, new_n8464_, new_n8462_ );
xor  ( new_n8467_, new_n8364_, new_n8362_ );
xor  ( new_n8468_, new_n8467_, new_n8367_ );
or   ( new_n8469_, new_n8468_, new_n8466_ );
and  ( new_n8470_, new_n8469_, new_n8465_ );
nor  ( new_n8471_, new_n8470_, new_n8460_ );
nand ( new_n8472_, new_n8470_, new_n8460_ );
xor  ( new_n8473_, new_n8430_, new_n8428_ );
xnor ( new_n8474_, new_n8473_, new_n8434_ );
and  ( new_n8475_, new_n8474_, new_n8472_ );
or   ( new_n8476_, new_n8475_, new_n8471_ );
or   ( new_n8477_, new_n299_, new_n8115_ );
or   ( new_n8478_, new_n302_, new_n8117_ );
and  ( new_n8479_, new_n8478_, new_n8477_ );
xor  ( new_n8480_, new_n8479_, new_n293_ );
not  ( new_n8481_, RIbb2bdd0_121 );
or   ( new_n8482_, new_n268_, new_n8481_ );
or   ( new_n8483_, new_n271_, new_n8352_ );
and  ( new_n8484_, new_n8483_, new_n8482_ );
xor  ( new_n8485_, new_n8484_, new_n263_ );
nor  ( new_n8486_, new_n8485_, new_n8480_ );
and  ( new_n8487_, RIbb2bd58_122, RIbb2f610_1 );
not  ( new_n8488_, new_n8487_ );
nand ( new_n8489_, new_n8485_, new_n8480_ );
and  ( new_n8490_, new_n8489_, new_n8488_ );
or   ( new_n8491_, new_n8490_, new_n8486_ );
xnor ( new_n8492_, new_n8227_, new_n8223_ );
xor  ( new_n8493_, new_n8492_, new_n8233_ );
and  ( new_n8494_, new_n8493_, new_n8491_ );
or   ( new_n8495_, new_n8493_, new_n8491_ );
xor  ( new_n8496_, new_n8356_, new_n8351_ );
xor  ( new_n8497_, new_n8496_, new_n8359_ );
and  ( new_n8498_, new_n8497_, new_n8495_ );
or   ( new_n8499_, new_n8498_, new_n8494_ );
xnor ( new_n8500_, new_n8281_, new_n8277_ );
xor  ( new_n8501_, new_n8500_, new_n8287_ );
xnor ( new_n8502_, new_n8301_, new_n8297_ );
xor  ( new_n8503_, new_n8502_, new_n8307_ );
or   ( new_n8504_, new_n8503_, new_n8501_ );
and  ( new_n8505_, new_n8503_, new_n8501_ );
xor  ( new_n8506_, new_n8335_, new_n8331_ );
xnor ( new_n8507_, new_n8506_, new_n8341_ );
or   ( new_n8508_, new_n8507_, new_n8505_ );
and  ( new_n8509_, new_n8508_, new_n8504_ );
nor  ( new_n8510_, new_n8509_, new_n8499_ );
nand ( new_n8511_, new_n8509_, new_n8499_ );
xnor ( new_n8512_, new_n8317_, new_n8313_ );
xor  ( new_n8513_, new_n8512_, new_n8323_ );
xnor ( new_n8514_, new_n8209_, new_n8205_ );
xor  ( new_n8515_, new_n8514_, new_n8215_ );
nor  ( new_n8516_, new_n8515_, new_n8513_ );
nand ( new_n8517_, new_n8515_, new_n8513_ );
xor  ( new_n8518_, new_n8193_, new_n8189_ );
xor  ( new_n8519_, new_n8518_, new_n8199_ );
and  ( new_n8520_, new_n8519_, new_n8517_ );
or   ( new_n8521_, new_n8520_, new_n8516_ );
and  ( new_n8522_, new_n8521_, new_n8511_ );
or   ( new_n8523_, new_n8522_, new_n8510_ );
or   ( new_n8524_, new_n4302_, new_n986_ );
or   ( new_n8525_, new_n4304_, new_n886_ );
and  ( new_n8526_, new_n8525_, new_n8524_ );
xor  ( new_n8527_, new_n8526_, new_n3895_ );
or   ( new_n8528_, new_n3896_, new_n1213_ );
or   ( new_n8529_, new_n3898_, new_n1168_ );
and  ( new_n8530_, new_n8529_, new_n8528_ );
xor  ( new_n8531_, new_n8530_, new_n3460_ );
or   ( new_n8532_, new_n8531_, new_n8527_ );
and  ( new_n8533_, new_n8531_, new_n8527_ );
or   ( new_n8534_, new_n3461_, new_n1525_ );
or   ( new_n8535_, new_n3463_, new_n1318_ );
and  ( new_n8536_, new_n8535_, new_n8534_ );
xor  ( new_n8537_, new_n8536_, new_n3116_ );
or   ( new_n8538_, new_n8537_, new_n8533_ );
and  ( new_n8539_, new_n8538_, new_n8532_ );
or   ( new_n8540_, new_n2122_, new_n2646_ );
or   ( new_n8541_, new_n2124_, new_n2475_ );
and  ( new_n8542_, new_n8541_, new_n8540_ );
xor  ( new_n8543_, new_n8542_, new_n1843_ );
or   ( new_n8544_, new_n1844_, new_n2981_ );
or   ( new_n8545_, new_n1846_, new_n2751_ );
and  ( new_n8546_, new_n8545_, new_n8544_ );
xor  ( new_n8547_, new_n8546_, new_n1586_ );
or   ( new_n8548_, new_n8547_, new_n8543_ );
and  ( new_n8549_, new_n8547_, new_n8543_ );
or   ( new_n8550_, new_n1593_, new_n3306_ );
or   ( new_n8551_, new_n1595_, new_n3178_ );
and  ( new_n8552_, new_n8551_, new_n8550_ );
xor  ( new_n8553_, new_n8552_, new_n1358_ );
or   ( new_n8554_, new_n8553_, new_n8549_ );
and  ( new_n8555_, new_n8554_, new_n8548_ );
or   ( new_n8556_, new_n8555_, new_n8539_ );
and  ( new_n8557_, new_n8555_, new_n8539_ );
or   ( new_n8558_, new_n3117_, new_n1754_ );
or   ( new_n8559_, new_n3119_, new_n1523_ );
and  ( new_n8560_, new_n8559_, new_n8558_ );
xor  ( new_n8561_, new_n8560_, new_n2800_ );
or   ( new_n8562_, new_n2807_, new_n2057_ );
or   ( new_n8563_, new_n2809_, new_n1899_ );
and  ( new_n8564_, new_n8563_, new_n8562_ );
xor  ( new_n8565_, new_n8564_, new_n2424_ );
nor  ( new_n8566_, new_n8565_, new_n8561_ );
and  ( new_n8567_, new_n8565_, new_n8561_ );
or   ( new_n8568_, new_n2425_, new_n2291_ );
or   ( new_n8569_, new_n2427_, new_n2178_ );
and  ( new_n8570_, new_n8569_, new_n8568_ );
xor  ( new_n8571_, new_n8570_, new_n2121_ );
nor  ( new_n8572_, new_n8571_, new_n8567_ );
nor  ( new_n8573_, new_n8572_, new_n8566_ );
or   ( new_n8574_, new_n8573_, new_n8557_ );
and  ( new_n8575_, new_n8574_, new_n8556_ );
or   ( new_n8576_, new_n755_, new_n4859_ );
or   ( new_n8577_, new_n757_, new_n4995_ );
and  ( new_n8578_, new_n8577_, new_n8576_ );
xor  ( new_n8579_, new_n8578_, new_n523_ );
or   ( new_n8580_, new_n524_, new_n5428_ );
or   ( new_n8581_, new_n526_, new_n5171_ );
and  ( new_n8582_, new_n8581_, new_n8580_ );
xor  ( new_n8583_, new_n8582_, new_n403_ );
or   ( new_n8584_, new_n8583_, new_n8579_ );
and  ( new_n8585_, new_n8583_, new_n8579_ );
or   ( new_n8586_, new_n409_, new_n5899_ );
or   ( new_n8587_, new_n411_, new_n5570_ );
and  ( new_n8588_, new_n8587_, new_n8586_ );
xor  ( new_n8589_, new_n8588_, new_n328_ );
or   ( new_n8590_, new_n8589_, new_n8585_ );
and  ( new_n8591_, new_n8590_, new_n8584_ );
or   ( new_n8592_, new_n337_, new_n6425_ );
or   ( new_n8593_, new_n340_, new_n6219_ );
and  ( new_n8594_, new_n8593_, new_n8592_ );
xor  ( new_n8595_, new_n8594_, new_n332_ );
or   ( new_n8596_, new_n317_, new_n6943_ );
or   ( new_n8597_, new_n320_, new_n6589_ );
and  ( new_n8598_, new_n8597_, new_n8596_ );
xor  ( new_n8599_, new_n8598_, new_n312_ );
or   ( new_n8600_, new_n8599_, new_n8595_ );
and  ( new_n8601_, new_n8599_, new_n8595_ );
or   ( new_n8602_, new_n283_, new_n7373_ );
or   ( new_n8603_, new_n286_, new_n7149_ );
and  ( new_n8604_, new_n8603_, new_n8602_ );
xor  ( new_n8605_, new_n8604_, new_n278_ );
or   ( new_n8606_, new_n8605_, new_n8601_ );
and  ( new_n8607_, new_n8606_, new_n8600_ );
or   ( new_n8608_, new_n8607_, new_n8591_ );
and  ( new_n8609_, new_n8607_, new_n8591_ );
or   ( new_n8610_, new_n1364_, new_n3694_ );
or   ( new_n8611_, new_n1366_, new_n3696_ );
and  ( new_n8612_, new_n8611_, new_n8610_ );
xor  ( new_n8613_, new_n8612_, new_n1129_ );
or   ( new_n8614_, new_n1135_, new_n4069_ );
or   ( new_n8615_, new_n1137_, new_n3820_ );
and  ( new_n8616_, new_n8615_, new_n8614_ );
xor  ( new_n8617_, new_n8616_, new_n896_ );
nor  ( new_n8618_, new_n8617_, new_n8613_ );
and  ( new_n8619_, new_n8617_, new_n8613_ );
or   ( new_n8620_, new_n897_, new_n4603_ );
or   ( new_n8621_, new_n899_, new_n4267_ );
and  ( new_n8622_, new_n8621_, new_n8620_ );
xor  ( new_n8623_, new_n8622_, new_n748_ );
nor  ( new_n8624_, new_n8623_, new_n8619_ );
nor  ( new_n8625_, new_n8624_, new_n8618_ );
or   ( new_n8626_, new_n8625_, new_n8609_ );
and  ( new_n8627_, new_n8626_, new_n8608_ );
or   ( new_n8628_, new_n8627_, new_n8575_ );
or   ( new_n8629_, new_n5604_, new_n443_ );
or   ( new_n8630_, new_n5606_, new_n419_ );
and  ( new_n8631_, new_n8630_, new_n8629_ );
xor  ( new_n8632_, new_n8631_, new_n5206_ );
or   ( new_n8633_, new_n5207_, new_n515_ );
or   ( new_n8634_, new_n5209_, new_n509_ );
and  ( new_n8635_, new_n8634_, new_n8633_ );
xor  ( new_n8636_, new_n8635_, new_n4708_ );
or   ( new_n8637_, new_n8636_, new_n8632_ );
and  ( new_n8638_, new_n8636_, new_n8632_ );
or   ( new_n8639_, new_n4709_, new_n805_ );
or   ( new_n8640_, new_n4711_, new_n775_ );
and  ( new_n8641_, new_n8640_, new_n8639_ );
xor  ( new_n8642_, new_n8641_, new_n4295_ );
or   ( new_n8643_, new_n8642_, new_n8638_ );
and  ( new_n8644_, new_n8643_, new_n8637_ );
or   ( new_n8645_, new_n8264_, new_n319_ );
or   ( new_n8646_, new_n8266_, new_n333_ );
and  ( new_n8647_, new_n8646_, new_n8645_ );
xor  ( new_n8648_, new_n8647_, new_n7724_ );
xor  ( new_n8649_, RIbb2dae0_59, RIbb2db58_58 );
xor  ( new_n8650_, RIbb2db58_58, new_n8254_ );
nor  ( new_n8651_, new_n8650_, new_n8649_ );
and  ( new_n8652_, new_n8651_, RIbb2d810_65 );
xor  ( new_n8653_, new_n8652_, new_n8257_ );
nand ( new_n8654_, new_n8653_, new_n8648_ );
nor  ( new_n8655_, new_n8653_, new_n8648_ );
or   ( new_n8656_, new_n7732_, new_n285_ );
or   ( new_n8657_, new_n7734_, new_n313_ );
and  ( new_n8658_, new_n8657_, new_n8656_ );
xor  ( new_n8659_, new_n8658_, new_n7177_ );
or   ( new_n8660_, new_n8659_, new_n8655_ );
and  ( new_n8661_, new_n8660_, new_n8654_ );
or   ( new_n8662_, new_n8661_, new_n8644_ );
and  ( new_n8663_, new_n8661_, new_n8644_ );
or   ( new_n8664_, new_n7184_, new_n301_ );
or   ( new_n8665_, new_n7186_, new_n279_ );
and  ( new_n8666_, new_n8665_, new_n8664_ );
xor  ( new_n8667_, new_n8666_, new_n6638_ );
or   ( new_n8668_, new_n6645_, new_n270_ );
or   ( new_n8669_, new_n6647_, new_n294_ );
and  ( new_n8670_, new_n8669_, new_n8668_ );
xor  ( new_n8671_, new_n8670_, new_n6166_ );
nor  ( new_n8672_, new_n8671_, new_n8667_ );
and  ( new_n8673_, new_n8671_, new_n8667_ );
or   ( new_n8674_, new_n6173_, new_n348_ );
or   ( new_n8675_, new_n6175_, new_n264_ );
and  ( new_n8676_, new_n8675_, new_n8674_ );
xor  ( new_n8677_, new_n8676_, new_n5597_ );
nor  ( new_n8678_, new_n8677_, new_n8673_ );
nor  ( new_n8679_, new_n8678_, new_n8672_ );
or   ( new_n8680_, new_n8679_, new_n8663_ );
and  ( new_n8681_, new_n8680_, new_n8662_ );
and  ( new_n8682_, new_n8627_, new_n8575_ );
or   ( new_n8683_, new_n8682_, new_n8681_ );
and  ( new_n8684_, new_n8683_, new_n8628_ );
or   ( new_n8685_, new_n8684_, new_n8523_ );
nand ( new_n8686_, new_n8684_, new_n8523_ );
xnor ( new_n8687_, new_n8044_, new_n8039_ );
xor  ( new_n8688_, new_n8687_, new_n8050_ );
xnor ( new_n8689_, new_n8078_, new_n8074_ );
xor  ( new_n8690_, new_n8689_, new_n8084_ );
nor  ( new_n8691_, new_n8690_, new_n8688_ );
and  ( new_n8692_, new_n8690_, new_n8688_ );
xor  ( new_n8693_, new_n8373_, new_n8371_ );
xnor ( new_n8694_, new_n8693_, new_n8377_ );
not  ( new_n8695_, new_n8694_ );
nor  ( new_n8696_, new_n8695_, new_n8692_ );
nor  ( new_n8697_, new_n8696_, new_n8691_ );
nand ( new_n8698_, new_n8697_, new_n8686_ );
and  ( new_n8699_, new_n8698_, new_n8685_ );
or   ( new_n8700_, new_n8699_, new_n8476_ );
nand ( new_n8701_, new_n8699_, new_n8476_ );
xor  ( new_n8702_, new_n8291_, new_n8237_ );
xor  ( new_n8703_, new_n8702_, new_n8345_ );
xnor ( new_n8704_, new_n8379_, new_n8369_ );
xor  ( new_n8705_, new_n8704_, new_n8391_ );
and  ( new_n8706_, new_n8705_, new_n8703_ );
nor  ( new_n8707_, new_n8705_, new_n8703_ );
xor  ( new_n8708_, new_n8399_, new_n8397_ );
xor  ( new_n8709_, new_n8708_, new_n8404_ );
nor  ( new_n8710_, new_n8709_, new_n8707_ );
nor  ( new_n8711_, new_n8710_, new_n8706_ );
nand ( new_n8712_, new_n8711_, new_n8701_ );
and  ( new_n8713_, new_n8712_, new_n8700_ );
or   ( new_n8714_, new_n8713_, new_n8458_ );
nand ( new_n8715_, new_n8713_, new_n8458_ );
xor  ( new_n8716_, new_n8393_, new_n8347_ );
xor  ( new_n8717_, new_n8716_, new_n8406_ );
xor  ( new_n8718_, new_n8412_, new_n8410_ );
xor  ( new_n8719_, new_n8718_, new_n8416_ );
nor  ( new_n8720_, new_n8719_, new_n8717_ );
and  ( new_n8721_, new_n8719_, new_n8717_ );
xor  ( new_n8722_, new_n8424_, new_n8422_ );
xnor ( new_n8723_, new_n8722_, new_n8436_ );
not  ( new_n8724_, new_n8723_ );
nor  ( new_n8725_, new_n8724_, new_n8721_ );
nor  ( new_n8726_, new_n8725_, new_n8720_ );
nand ( new_n8727_, new_n8726_, new_n8715_ );
and  ( new_n8728_, new_n8727_, new_n8714_ );
and  ( new_n8729_, new_n8728_, new_n8456_ );
nor  ( new_n8730_, new_n8728_, new_n8456_ );
xor  ( new_n8731_, new_n8136_, new_n7912_ );
xor  ( new_n8732_, new_n8731_, new_n8148_ );
nor  ( new_n8733_, new_n8732_, new_n8730_ );
nor  ( new_n8734_, new_n8733_, new_n8729_ );
xor  ( new_n8735_, new_n8169_, new_n8167_ );
xnor ( new_n8736_, new_n8735_, new_n8443_ );
nor  ( new_n8737_, new_n8736_, new_n8734_ );
xor  ( new_n8738_, new_n8447_, new_n8445_ );
and  ( new_n8739_, new_n8738_, new_n8737_ );
xnor ( new_n8740_, new_n8736_, new_n8734_ );
xor  ( new_n8741_, new_n8183_, new_n8173_ );
xor  ( new_n8742_, new_n8741_, new_n8441_ );
xnor ( new_n8743_, new_n8728_, new_n8456_ );
xor  ( new_n8744_, new_n8743_, new_n8732_ );
nand ( new_n8745_, new_n8744_, new_n8742_ );
nor  ( new_n8746_, new_n8744_, new_n8742_ );
xor  ( new_n8747_, new_n8719_, new_n8717_ );
xor  ( new_n8748_, new_n8747_, new_n8724_ );
xor  ( new_n8749_, new_n8684_, new_n8523_ );
xor  ( new_n8750_, new_n8749_, new_n8697_ );
xnor ( new_n8751_, new_n8470_, new_n8460_ );
xor  ( new_n8752_, new_n8751_, new_n8474_ );
or   ( new_n8753_, new_n8752_, new_n8750_ );
nand ( new_n8754_, new_n8752_, new_n8750_ );
xor  ( new_n8755_, new_n8705_, new_n8703_ );
xnor ( new_n8756_, new_n8755_, new_n8709_ );
nand ( new_n8757_, new_n8756_, new_n8754_ );
and  ( new_n8758_, new_n8757_, new_n8753_ );
or   ( new_n8759_, new_n8758_, new_n8748_ );
and  ( new_n8760_, new_n8758_, new_n8748_ );
xnor ( new_n8761_, new_n8503_, new_n8501_ );
xor  ( new_n8762_, new_n8761_, new_n8507_ );
xor  ( new_n8763_, new_n8515_, new_n8513_ );
xor  ( new_n8764_, new_n8763_, new_n8519_ );
nor  ( new_n8765_, new_n8764_, new_n8762_ );
and  ( new_n8766_, new_n8764_, new_n8762_ );
xor  ( new_n8767_, new_n8493_, new_n8491_ );
xnor ( new_n8768_, new_n8767_, new_n8497_ );
nor  ( new_n8769_, new_n8768_, new_n8766_ );
or   ( new_n8770_, new_n8769_, new_n8765_ );
xnor ( new_n8771_, new_n8325_, new_n8309_ );
xor  ( new_n8772_, new_n8771_, new_n8343_ );
or   ( new_n8773_, new_n8772_, new_n8770_ );
and  ( new_n8774_, new_n8772_, new_n8770_ );
xnor ( new_n8775_, new_n8555_, new_n8539_ );
xor  ( new_n8776_, new_n8775_, new_n8573_ );
xnor ( new_n8777_, new_n8607_, new_n8591_ );
xor  ( new_n8778_, new_n8777_, new_n8625_ );
nor  ( new_n8779_, new_n8778_, new_n8776_ );
and  ( new_n8780_, new_n8778_, new_n8776_ );
xor  ( new_n8781_, new_n8661_, new_n8644_ );
xnor ( new_n8782_, new_n8781_, new_n8679_ );
nor  ( new_n8783_, new_n8782_, new_n8780_ );
nor  ( new_n8784_, new_n8783_, new_n8779_ );
or   ( new_n8785_, new_n8784_, new_n8774_ );
and  ( new_n8786_, new_n8785_, new_n8773_ );
xnor ( new_n8787_, new_n8271_, new_n8253_ );
xor  ( new_n8788_, new_n8787_, new_n8289_ );
xor  ( new_n8789_, new_n8690_, new_n8688_ );
xor  ( new_n8790_, new_n8789_, new_n8695_ );
or   ( new_n8791_, new_n8790_, new_n8788_ );
and  ( new_n8792_, new_n8790_, new_n8788_ );
xor  ( new_n8793_, new_n8464_, new_n8462_ );
xnor ( new_n8794_, new_n8793_, new_n8468_ );
not  ( new_n8795_, new_n8794_ );
or   ( new_n8796_, new_n8795_, new_n8792_ );
and  ( new_n8797_, new_n8796_, new_n8791_ );
nor  ( new_n8798_, new_n8797_, new_n8786_ );
and  ( new_n8799_, new_n8797_, new_n8786_ );
xor  ( new_n8800_, new_n8245_, new_n8241_ );
xor  ( new_n8801_, new_n8800_, new_n8251_ );
xnor ( new_n8802_, new_n8653_, new_n8648_ );
xor  ( new_n8803_, new_n8802_, new_n8659_ );
xnor ( new_n8804_, new_n8636_, new_n8632_ );
xor  ( new_n8805_, new_n8804_, new_n8642_ );
or   ( new_n8806_, new_n8805_, new_n8803_ );
and  ( new_n8807_, new_n8805_, new_n8803_ );
xnor ( new_n8808_, new_n8671_, new_n8667_ );
xor  ( new_n8809_, new_n8808_, new_n8677_ );
or   ( new_n8810_, new_n8809_, new_n8807_ );
and  ( new_n8811_, new_n8810_, new_n8806_ );
nor  ( new_n8812_, new_n8811_, new_n8801_ );
nand ( new_n8813_, new_n8811_, new_n8801_ );
xor  ( new_n8814_, new_n8261_, new_n8257_ );
xor  ( new_n8815_, new_n8814_, new_n8269_ );
and  ( new_n8816_, new_n8815_, new_n8813_ );
or   ( new_n8817_, new_n8816_, new_n8812_ );
or   ( new_n8818_, new_n2425_, new_n2475_ );
or   ( new_n8819_, new_n2427_, new_n2291_ );
and  ( new_n8820_, new_n8819_, new_n8818_ );
xor  ( new_n8821_, new_n8820_, new_n2121_ );
or   ( new_n8822_, new_n2122_, new_n2751_ );
or   ( new_n8823_, new_n2124_, new_n2646_ );
and  ( new_n8824_, new_n8823_, new_n8822_ );
xor  ( new_n8825_, new_n8824_, new_n1843_ );
or   ( new_n8826_, new_n8825_, new_n8821_ );
and  ( new_n8827_, new_n8825_, new_n8821_ );
or   ( new_n8828_, new_n1844_, new_n3178_ );
or   ( new_n8829_, new_n1846_, new_n2981_ );
and  ( new_n8830_, new_n8829_, new_n8828_ );
xor  ( new_n8831_, new_n8830_, new_n1586_ );
or   ( new_n8832_, new_n8831_, new_n8827_ );
and  ( new_n8833_, new_n8832_, new_n8826_ );
or   ( new_n8834_, new_n3461_, new_n1523_ );
or   ( new_n8835_, new_n3463_, new_n1525_ );
and  ( new_n8836_, new_n8835_, new_n8834_ );
xor  ( new_n8837_, new_n8836_, new_n3116_ );
or   ( new_n8838_, new_n3117_, new_n1899_ );
or   ( new_n8839_, new_n3119_, new_n1754_ );
and  ( new_n8840_, new_n8839_, new_n8838_ );
xor  ( new_n8841_, new_n8840_, new_n2800_ );
or   ( new_n8842_, new_n8841_, new_n8837_ );
and  ( new_n8843_, new_n8841_, new_n8837_ );
or   ( new_n8844_, new_n2807_, new_n2178_ );
or   ( new_n8845_, new_n2809_, new_n2057_ );
and  ( new_n8846_, new_n8845_, new_n8844_ );
xor  ( new_n8847_, new_n8846_, new_n2424_ );
or   ( new_n8848_, new_n8847_, new_n8843_ );
and  ( new_n8849_, new_n8848_, new_n8842_ );
or   ( new_n8850_, new_n8849_, new_n8833_ );
and  ( new_n8851_, new_n8849_, new_n8833_ );
or   ( new_n8852_, new_n4709_, new_n886_ );
or   ( new_n8853_, new_n4711_, new_n805_ );
and  ( new_n8854_, new_n8853_, new_n8852_ );
xor  ( new_n8855_, new_n8854_, new_n4295_ );
or   ( new_n8856_, new_n4302_, new_n1168_ );
or   ( new_n8857_, new_n4304_, new_n986_ );
and  ( new_n8858_, new_n8857_, new_n8856_ );
xor  ( new_n8859_, new_n8858_, new_n3895_ );
nor  ( new_n8860_, new_n8859_, new_n8855_ );
and  ( new_n8861_, new_n8859_, new_n8855_ );
or   ( new_n8862_, new_n3896_, new_n1318_ );
or   ( new_n8863_, new_n3898_, new_n1213_ );
and  ( new_n8864_, new_n8863_, new_n8862_ );
xor  ( new_n8865_, new_n8864_, new_n3460_ );
nor  ( new_n8866_, new_n8865_, new_n8861_ );
nor  ( new_n8867_, new_n8866_, new_n8860_ );
or   ( new_n8868_, new_n8867_, new_n8851_ );
and  ( new_n8869_, new_n8868_, new_n8850_ );
not  ( new_n8870_, RIbb2dae0_59 );
and  ( new_n8871_, RIbb2d9f0_61, RIbb2da68_60 );
nor  ( new_n8872_, new_n8871_, new_n8870_ );
not  ( new_n8873_, new_n8872_ );
not  ( new_n8874_, new_n8651_ );
or   ( new_n8875_, new_n8874_, new_n333_ );
not  ( new_n8876_, new_n8649_ );
or   ( new_n8877_, new_n8876_, new_n339_ );
and  ( new_n8878_, new_n8877_, new_n8875_ );
xor  ( new_n8879_, new_n8878_, new_n8257_ );
and  ( new_n8880_, new_n8879_, new_n8873_ );
or   ( new_n8881_, new_n8879_, new_n8873_ );
or   ( new_n8882_, new_n8264_, new_n313_ );
or   ( new_n8883_, new_n8266_, new_n319_ );
and  ( new_n8884_, new_n8883_, new_n8882_ );
xor  ( new_n8885_, new_n8884_, new_n7725_ );
and  ( new_n8886_, new_n8885_, new_n8881_ );
or   ( new_n8887_, new_n8886_, new_n8880_ );
or   ( new_n8888_, new_n6173_, new_n419_ );
or   ( new_n8889_, new_n6175_, new_n348_ );
and  ( new_n8890_, new_n8889_, new_n8888_ );
xor  ( new_n8891_, new_n8890_, new_n5597_ );
or   ( new_n8892_, new_n5604_, new_n509_ );
or   ( new_n8893_, new_n5606_, new_n443_ );
and  ( new_n8894_, new_n8893_, new_n8892_ );
xor  ( new_n8895_, new_n8894_, new_n5206_ );
or   ( new_n8896_, new_n8895_, new_n8891_ );
and  ( new_n8897_, new_n8895_, new_n8891_ );
or   ( new_n8898_, new_n5207_, new_n775_ );
or   ( new_n8899_, new_n5209_, new_n515_ );
and  ( new_n8900_, new_n8899_, new_n8898_ );
xor  ( new_n8901_, new_n8900_, new_n4708_ );
or   ( new_n8902_, new_n8901_, new_n8897_ );
and  ( new_n8903_, new_n8902_, new_n8896_ );
or   ( new_n8904_, new_n8903_, new_n8887_ );
and  ( new_n8905_, new_n8903_, new_n8887_ );
or   ( new_n8906_, new_n7732_, new_n279_ );
or   ( new_n8907_, new_n7734_, new_n285_ );
and  ( new_n8908_, new_n8907_, new_n8906_ );
xor  ( new_n8909_, new_n8908_, new_n7177_ );
or   ( new_n8910_, new_n7184_, new_n294_ );
or   ( new_n8911_, new_n7186_, new_n301_ );
and  ( new_n8912_, new_n8911_, new_n8910_ );
xor  ( new_n8913_, new_n8912_, new_n6638_ );
nor  ( new_n8914_, new_n8913_, new_n8909_ );
and  ( new_n8915_, new_n8913_, new_n8909_ );
or   ( new_n8916_, new_n6645_, new_n264_ );
or   ( new_n8917_, new_n6647_, new_n270_ );
and  ( new_n8918_, new_n8917_, new_n8916_ );
xor  ( new_n8919_, new_n8918_, new_n6166_ );
nor  ( new_n8920_, new_n8919_, new_n8915_ );
nor  ( new_n8921_, new_n8920_, new_n8914_ );
or   ( new_n8922_, new_n8921_, new_n8905_ );
and  ( new_n8923_, new_n8922_, new_n8904_ );
or   ( new_n8924_, new_n8923_, new_n8869_ );
or   ( new_n8925_, new_n897_, new_n4995_ );
or   ( new_n8926_, new_n899_, new_n4603_ );
and  ( new_n8927_, new_n8926_, new_n8925_ );
xor  ( new_n8928_, new_n8927_, new_n748_ );
or   ( new_n8929_, new_n755_, new_n5171_ );
or   ( new_n8930_, new_n757_, new_n4859_ );
and  ( new_n8931_, new_n8930_, new_n8929_ );
xor  ( new_n8932_, new_n8931_, new_n523_ );
or   ( new_n8933_, new_n8932_, new_n8928_ );
and  ( new_n8934_, new_n8932_, new_n8928_ );
or   ( new_n8935_, new_n524_, new_n5570_ );
or   ( new_n8936_, new_n526_, new_n5428_ );
and  ( new_n8937_, new_n8936_, new_n8935_ );
xor  ( new_n8938_, new_n8937_, new_n403_ );
or   ( new_n8939_, new_n8938_, new_n8934_ );
and  ( new_n8940_, new_n8939_, new_n8933_ );
or   ( new_n8941_, new_n409_, new_n6219_ );
or   ( new_n8942_, new_n411_, new_n5899_ );
and  ( new_n8943_, new_n8942_, new_n8941_ );
xor  ( new_n8944_, new_n8943_, new_n328_ );
or   ( new_n8945_, new_n337_, new_n6589_ );
or   ( new_n8946_, new_n340_, new_n6425_ );
and  ( new_n8947_, new_n8946_, new_n8945_ );
xor  ( new_n8948_, new_n8947_, new_n332_ );
or   ( new_n8949_, new_n8948_, new_n8944_ );
and  ( new_n8950_, new_n8948_, new_n8944_ );
or   ( new_n8951_, new_n317_, new_n7149_ );
or   ( new_n8952_, new_n320_, new_n6943_ );
and  ( new_n8953_, new_n8952_, new_n8951_ );
xor  ( new_n8954_, new_n8953_, new_n312_ );
or   ( new_n8955_, new_n8954_, new_n8950_ );
and  ( new_n8956_, new_n8955_, new_n8949_ );
nor  ( new_n8957_, new_n8956_, new_n8940_ );
and  ( new_n8958_, new_n8956_, new_n8940_ );
or   ( new_n8959_, new_n1593_, new_n3696_ );
or   ( new_n8960_, new_n1595_, new_n3306_ );
and  ( new_n8961_, new_n8960_, new_n8959_ );
xor  ( new_n8962_, new_n8961_, new_n1358_ );
or   ( new_n8963_, new_n1364_, new_n3820_ );
or   ( new_n8964_, new_n1366_, new_n3694_ );
and  ( new_n8965_, new_n8964_, new_n8963_ );
xor  ( new_n8966_, new_n8965_, new_n1129_ );
nor  ( new_n8967_, new_n8966_, new_n8962_ );
and  ( new_n8968_, new_n8966_, new_n8962_ );
or   ( new_n8969_, new_n1135_, new_n4267_ );
or   ( new_n8970_, new_n1137_, new_n4069_ );
and  ( new_n8971_, new_n8970_, new_n8969_ );
xor  ( new_n8972_, new_n8971_, new_n896_ );
nor  ( new_n8973_, new_n8972_, new_n8968_ );
nor  ( new_n8974_, new_n8973_, new_n8967_ );
nor  ( new_n8975_, new_n8974_, new_n8958_ );
nor  ( new_n8976_, new_n8975_, new_n8957_ );
and  ( new_n8977_, new_n8923_, new_n8869_ );
or   ( new_n8978_, new_n8977_, new_n8976_ );
and  ( new_n8979_, new_n8978_, new_n8924_ );
and  ( new_n8980_, new_n8979_, new_n8817_ );
nor  ( new_n8981_, new_n8979_, new_n8817_ );
xor  ( new_n8982_, new_n8485_, new_n8480_ );
xor  ( new_n8983_, new_n8982_, new_n8488_ );
not  ( new_n8984_, new_n8983_ );
or   ( new_n8985_, new_n283_, new_n8117_ );
or   ( new_n8986_, new_n286_, new_n7373_ );
and  ( new_n8987_, new_n8986_, new_n8985_ );
xor  ( new_n8988_, new_n8987_, new_n278_ );
or   ( new_n8989_, new_n299_, new_n8352_ );
or   ( new_n8990_, new_n302_, new_n8115_ );
and  ( new_n8991_, new_n8990_, new_n8989_ );
xor  ( new_n8992_, new_n8991_, new_n293_ );
or   ( new_n8993_, new_n8992_, new_n8988_ );
and  ( new_n8994_, new_n8992_, new_n8988_ );
not  ( new_n8995_, RIbb2bd58_122 );
or   ( new_n8996_, new_n268_, new_n8995_ );
or   ( new_n8997_, new_n271_, new_n8481_ );
and  ( new_n8998_, new_n8997_, new_n8996_ );
xor  ( new_n8999_, new_n8998_, new_n263_ );
or   ( new_n9000_, new_n8999_, new_n8994_ );
and  ( new_n9001_, new_n9000_, new_n8993_ );
nor  ( new_n9002_, new_n9001_, new_n8984_ );
xnor ( new_n9003_, new_n8547_, new_n8543_ );
xor  ( new_n9004_, new_n9003_, new_n8553_ );
xnor ( new_n9005_, new_n8531_, new_n8527_ );
xor  ( new_n9006_, new_n9005_, new_n8537_ );
or   ( new_n9007_, new_n9006_, new_n9004_ );
and  ( new_n9008_, new_n9006_, new_n9004_ );
xor  ( new_n9009_, new_n8565_, new_n8561_ );
xnor ( new_n9010_, new_n9009_, new_n8571_ );
or   ( new_n9011_, new_n9010_, new_n9008_ );
and  ( new_n9012_, new_n9011_, new_n9007_ );
nor  ( new_n9013_, new_n9012_, new_n9002_ );
and  ( new_n9014_, new_n9012_, new_n9002_ );
xnor ( new_n9015_, new_n8599_, new_n8595_ );
xor  ( new_n9016_, new_n9015_, new_n8605_ );
xnor ( new_n9017_, new_n8583_, new_n8579_ );
xor  ( new_n9018_, new_n9017_, new_n8589_ );
nor  ( new_n9019_, new_n9018_, new_n9016_ );
and  ( new_n9020_, new_n9018_, new_n9016_ );
xor  ( new_n9021_, new_n8617_, new_n8613_ );
xnor ( new_n9022_, new_n9021_, new_n8623_ );
nor  ( new_n9023_, new_n9022_, new_n9020_ );
nor  ( new_n9024_, new_n9023_, new_n9019_ );
nor  ( new_n9025_, new_n9024_, new_n9014_ );
nor  ( new_n9026_, new_n9025_, new_n9013_ );
nor  ( new_n9027_, new_n9026_, new_n8981_ );
nor  ( new_n9028_, new_n9027_, new_n8980_ );
nor  ( new_n9029_, new_n9028_, new_n8799_ );
nor  ( new_n9030_, new_n9029_, new_n8798_ );
or   ( new_n9031_, new_n9030_, new_n8760_ );
and  ( new_n9032_, new_n9031_, new_n8759_ );
xor  ( new_n9033_, new_n8713_, new_n8458_ );
xor  ( new_n9034_, new_n9033_, new_n8726_ );
nor  ( new_n9035_, new_n9034_, new_n9032_ );
and  ( new_n9036_, new_n9034_, new_n9032_ );
xor  ( new_n9037_, new_n8455_, new_n8453_ );
not  ( new_n9038_, new_n9037_ );
nor  ( new_n9039_, new_n9038_, new_n9036_ );
nor  ( new_n9040_, new_n9039_, new_n9035_ );
or   ( new_n9041_, new_n9040_, new_n8746_ );
and  ( new_n9042_, new_n9041_, new_n8745_ );
nor  ( new_n9043_, new_n9042_, new_n8740_ );
xor  ( new_n9044_, new_n9034_, new_n9032_ );
xor  ( new_n9045_, new_n9044_, new_n9038_ );
xor  ( new_n9046_, new_n8752_, new_n8750_ );
xor  ( new_n9047_, new_n9046_, new_n8756_ );
xor  ( new_n9048_, new_n8764_, new_n8762_ );
xor  ( new_n9049_, new_n9048_, new_n8768_ );
xnor ( new_n9050_, new_n8778_, new_n8776_ );
xor  ( new_n9051_, new_n9050_, new_n8782_ );
and  ( new_n9052_, new_n9051_, new_n9049_ );
or   ( new_n9053_, new_n9051_, new_n9049_ );
xor  ( new_n9054_, new_n8956_, new_n8940_ );
xor  ( new_n9055_, new_n9054_, new_n8974_ );
xnor ( new_n9056_, new_n9018_, new_n9016_ );
xor  ( new_n9057_, new_n9056_, new_n9022_ );
and  ( new_n9058_, new_n9057_, new_n9055_ );
nor  ( new_n9059_, new_n9057_, new_n9055_ );
xor  ( new_n9060_, new_n9001_, new_n8984_ );
nor  ( new_n9061_, new_n9060_, new_n9059_ );
nor  ( new_n9062_, new_n9061_, new_n9058_ );
not  ( new_n9063_, new_n9062_ );
and  ( new_n9064_, new_n9063_, new_n9053_ );
or   ( new_n9065_, new_n9064_, new_n9052_ );
xnor ( new_n9066_, new_n8992_, new_n8988_ );
xor  ( new_n9067_, new_n9066_, new_n8999_ );
xnor ( new_n9068_, new_n8948_, new_n8944_ );
xor  ( new_n9069_, new_n9068_, new_n8954_ );
or   ( new_n9070_, new_n9069_, new_n9067_ );
and  ( new_n9071_, new_n9069_, new_n9067_ );
xor  ( new_n9072_, new_n8932_, new_n8928_ );
xnor ( new_n9073_, new_n9072_, new_n8938_ );
or   ( new_n9074_, new_n9073_, new_n9071_ );
and  ( new_n9075_, new_n9074_, new_n9070_ );
xnor ( new_n9076_, new_n8966_, new_n8962_ );
xor  ( new_n9077_, new_n9076_, new_n8972_ );
xnor ( new_n9078_, new_n8841_, new_n8837_ );
xor  ( new_n9079_, new_n9078_, new_n8847_ );
or   ( new_n9080_, new_n9079_, new_n9077_ );
and  ( new_n9081_, new_n9079_, new_n9077_ );
xor  ( new_n9082_, new_n8825_, new_n8821_ );
xnor ( new_n9083_, new_n9082_, new_n8831_ );
or   ( new_n9084_, new_n9083_, new_n9081_ );
and  ( new_n9085_, new_n9084_, new_n9080_ );
nor  ( new_n9086_, new_n9085_, new_n9075_ );
nand ( new_n9087_, new_n9085_, new_n9075_ );
and  ( new_n9088_, RIbb2bc68_124, RIbb2f610_1 );
or   ( new_n9089_, new_n283_, new_n8115_ );
or   ( new_n9090_, new_n286_, new_n8117_ );
and  ( new_n9091_, new_n9090_, new_n9089_ );
xor  ( new_n9092_, new_n9091_, new_n278_ );
or   ( new_n9093_, new_n299_, new_n8481_ );
or   ( new_n9094_, new_n302_, new_n8352_ );
and  ( new_n9095_, new_n9094_, new_n9093_ );
xor  ( new_n9096_, new_n9095_, new_n293_ );
or   ( new_n9097_, new_n9096_, new_n9092_ );
and  ( new_n9098_, new_n9096_, new_n9092_ );
not  ( new_n9099_, RIbb2bce0_123 );
or   ( new_n9100_, new_n268_, new_n9099_ );
or   ( new_n9101_, new_n271_, new_n8995_ );
and  ( new_n9102_, new_n9101_, new_n9100_ );
xor  ( new_n9103_, new_n9102_, new_n263_ );
or   ( new_n9104_, new_n9103_, new_n9098_ );
and  ( new_n9105_, new_n9104_, new_n9097_ );
nor  ( new_n9106_, new_n9105_, new_n9088_ );
and  ( new_n9107_, new_n9105_, new_n9088_ );
and  ( new_n9108_, RIbb2bce0_123, RIbb2f610_1 );
nor  ( new_n9109_, new_n9108_, new_n9107_ );
nor  ( new_n9110_, new_n9109_, new_n9106_ );
and  ( new_n9111_, new_n9110_, new_n9087_ );
or   ( new_n9112_, new_n9111_, new_n9086_ );
or   ( new_n9113_, new_n1593_, new_n3694_ );
or   ( new_n9114_, new_n1595_, new_n3696_ );
and  ( new_n9115_, new_n9114_, new_n9113_ );
xor  ( new_n9116_, new_n9115_, new_n1358_ );
or   ( new_n9117_, new_n1364_, new_n4069_ );
or   ( new_n9118_, new_n1366_, new_n3820_ );
and  ( new_n9119_, new_n9118_, new_n9117_ );
xor  ( new_n9120_, new_n9119_, new_n1129_ );
or   ( new_n9121_, new_n9120_, new_n9116_ );
and  ( new_n9122_, new_n9120_, new_n9116_ );
or   ( new_n9123_, new_n1135_, new_n4603_ );
or   ( new_n9124_, new_n1137_, new_n4267_ );
and  ( new_n9125_, new_n9124_, new_n9123_ );
xor  ( new_n9126_, new_n9125_, new_n896_ );
or   ( new_n9127_, new_n9126_, new_n9122_ );
and  ( new_n9128_, new_n9127_, new_n9121_ );
or   ( new_n9129_, new_n897_, new_n4859_ );
or   ( new_n9130_, new_n899_, new_n4995_ );
and  ( new_n9131_, new_n9130_, new_n9129_ );
xor  ( new_n9132_, new_n9131_, new_n748_ );
or   ( new_n9133_, new_n755_, new_n5428_ );
or   ( new_n9134_, new_n757_, new_n5171_ );
and  ( new_n9135_, new_n9134_, new_n9133_ );
xor  ( new_n9136_, new_n9135_, new_n523_ );
or   ( new_n9137_, new_n9136_, new_n9132_ );
and  ( new_n9138_, new_n9136_, new_n9132_ );
or   ( new_n9139_, new_n524_, new_n5899_ );
or   ( new_n9140_, new_n526_, new_n5570_ );
and  ( new_n9141_, new_n9140_, new_n9139_ );
xor  ( new_n9142_, new_n9141_, new_n403_ );
or   ( new_n9143_, new_n9142_, new_n9138_ );
and  ( new_n9144_, new_n9143_, new_n9137_ );
or   ( new_n9145_, new_n9144_, new_n9128_ );
and  ( new_n9146_, new_n9144_, new_n9128_ );
or   ( new_n9147_, new_n409_, new_n6425_ );
or   ( new_n9148_, new_n411_, new_n6219_ );
and  ( new_n9149_, new_n9148_, new_n9147_ );
xor  ( new_n9150_, new_n9149_, new_n328_ );
or   ( new_n9151_, new_n337_, new_n6943_ );
or   ( new_n9152_, new_n340_, new_n6589_ );
and  ( new_n9153_, new_n9152_, new_n9151_ );
xor  ( new_n9154_, new_n9153_, new_n332_ );
nor  ( new_n9155_, new_n9154_, new_n9150_ );
and  ( new_n9156_, new_n9154_, new_n9150_ );
or   ( new_n9157_, new_n317_, new_n7373_ );
or   ( new_n9158_, new_n320_, new_n7149_ );
and  ( new_n9159_, new_n9158_, new_n9157_ );
xor  ( new_n9160_, new_n9159_, new_n312_ );
nor  ( new_n9161_, new_n9160_, new_n9156_ );
nor  ( new_n9162_, new_n9161_, new_n9155_ );
or   ( new_n9163_, new_n9162_, new_n9146_ );
and  ( new_n9164_, new_n9163_, new_n9145_ );
or   ( new_n9165_, new_n6173_, new_n443_ );
or   ( new_n9166_, new_n6175_, new_n419_ );
and  ( new_n9167_, new_n9166_, new_n9165_ );
xor  ( new_n9168_, new_n9167_, new_n5597_ );
or   ( new_n9169_, new_n5604_, new_n515_ );
or   ( new_n9170_, new_n5606_, new_n509_ );
and  ( new_n9171_, new_n9170_, new_n9169_ );
xor  ( new_n9172_, new_n9171_, new_n5206_ );
or   ( new_n9173_, new_n9172_, new_n9168_ );
and  ( new_n9174_, new_n9172_, new_n9168_ );
or   ( new_n9175_, new_n5207_, new_n805_ );
or   ( new_n9176_, new_n5209_, new_n775_ );
and  ( new_n9177_, new_n9176_, new_n9175_ );
xor  ( new_n9178_, new_n9177_, new_n4708_ );
or   ( new_n9179_, new_n9178_, new_n9174_ );
and  ( new_n9180_, new_n9179_, new_n9173_ );
or   ( new_n9181_, new_n8874_, new_n319_ );
or   ( new_n9182_, new_n8876_, new_n333_ );
and  ( new_n9183_, new_n9182_, new_n9181_ );
xor  ( new_n9184_, new_n9183_, new_n8256_ );
xor  ( new_n9185_, RIbb2d9f0_61, RIbb2da68_60 );
xor  ( new_n9186_, RIbb2da68_60, new_n8870_ );
nor  ( new_n9187_, new_n9186_, new_n9185_ );
and  ( new_n9188_, new_n9187_, RIbb2d810_65 );
xor  ( new_n9189_, new_n9188_, new_n8873_ );
nand ( new_n9190_, new_n9189_, new_n9184_ );
nor  ( new_n9191_, new_n9189_, new_n9184_ );
or   ( new_n9192_, new_n8264_, new_n285_ );
or   ( new_n9193_, new_n8266_, new_n313_ );
and  ( new_n9194_, new_n9193_, new_n9192_ );
xor  ( new_n9195_, new_n9194_, new_n7725_ );
or   ( new_n9196_, new_n9195_, new_n9191_ );
and  ( new_n9197_, new_n9196_, new_n9190_ );
or   ( new_n9198_, new_n9197_, new_n9180_ );
and  ( new_n9199_, new_n9197_, new_n9180_ );
or   ( new_n9200_, new_n7732_, new_n301_ );
or   ( new_n9201_, new_n7734_, new_n279_ );
and  ( new_n9202_, new_n9201_, new_n9200_ );
xor  ( new_n9203_, new_n9202_, new_n7177_ );
or   ( new_n9204_, new_n7184_, new_n270_ );
or   ( new_n9205_, new_n7186_, new_n294_ );
and  ( new_n9206_, new_n9205_, new_n9204_ );
xor  ( new_n9207_, new_n9206_, new_n6638_ );
nor  ( new_n9208_, new_n9207_, new_n9203_ );
and  ( new_n9209_, new_n9207_, new_n9203_ );
or   ( new_n9210_, new_n6645_, new_n348_ );
or   ( new_n9211_, new_n6647_, new_n264_ );
and  ( new_n9212_, new_n9211_, new_n9210_ );
xor  ( new_n9213_, new_n9212_, new_n6166_ );
nor  ( new_n9214_, new_n9213_, new_n9209_ );
nor  ( new_n9215_, new_n9214_, new_n9208_ );
or   ( new_n9216_, new_n9215_, new_n9199_ );
and  ( new_n9217_, new_n9216_, new_n9198_ );
or   ( new_n9218_, new_n9217_, new_n9164_ );
or   ( new_n9219_, new_n2425_, new_n2646_ );
or   ( new_n9220_, new_n2427_, new_n2475_ );
and  ( new_n9221_, new_n9220_, new_n9219_ );
xor  ( new_n9222_, new_n9221_, new_n2121_ );
or   ( new_n9223_, new_n2122_, new_n2981_ );
or   ( new_n9224_, new_n2124_, new_n2751_ );
and  ( new_n9225_, new_n9224_, new_n9223_ );
xor  ( new_n9226_, new_n9225_, new_n1843_ );
or   ( new_n9227_, new_n9226_, new_n9222_ );
and  ( new_n9228_, new_n9226_, new_n9222_ );
or   ( new_n9229_, new_n1844_, new_n3306_ );
or   ( new_n9230_, new_n1846_, new_n3178_ );
and  ( new_n9231_, new_n9230_, new_n9229_ );
xor  ( new_n9232_, new_n9231_, new_n1586_ );
or   ( new_n9233_, new_n9232_, new_n9228_ );
and  ( new_n9234_, new_n9233_, new_n9227_ );
or   ( new_n9235_, new_n4709_, new_n986_ );
or   ( new_n9236_, new_n4711_, new_n886_ );
and  ( new_n9237_, new_n9236_, new_n9235_ );
xor  ( new_n9238_, new_n9237_, new_n4295_ );
or   ( new_n9239_, new_n4302_, new_n1213_ );
or   ( new_n9240_, new_n4304_, new_n1168_ );
and  ( new_n9241_, new_n9240_, new_n9239_ );
xor  ( new_n9242_, new_n9241_, new_n3895_ );
or   ( new_n9243_, new_n9242_, new_n9238_ );
and  ( new_n9244_, new_n9242_, new_n9238_ );
or   ( new_n9245_, new_n3896_, new_n1525_ );
or   ( new_n9246_, new_n3898_, new_n1318_ );
and  ( new_n9247_, new_n9246_, new_n9245_ );
xor  ( new_n9248_, new_n9247_, new_n3460_ );
or   ( new_n9249_, new_n9248_, new_n9244_ );
and  ( new_n9250_, new_n9249_, new_n9243_ );
nor  ( new_n9251_, new_n9250_, new_n9234_ );
and  ( new_n9252_, new_n9250_, new_n9234_ );
or   ( new_n9253_, new_n3461_, new_n1754_ );
or   ( new_n9254_, new_n3463_, new_n1523_ );
and  ( new_n9255_, new_n9254_, new_n9253_ );
xor  ( new_n9256_, new_n9255_, new_n3116_ );
or   ( new_n9257_, new_n3117_, new_n2057_ );
or   ( new_n9258_, new_n3119_, new_n1899_ );
and  ( new_n9259_, new_n9258_, new_n9257_ );
xor  ( new_n9260_, new_n9259_, new_n2800_ );
nor  ( new_n9261_, new_n9260_, new_n9256_ );
and  ( new_n9262_, new_n9260_, new_n9256_ );
or   ( new_n9263_, new_n2807_, new_n2291_ );
or   ( new_n9264_, new_n2809_, new_n2178_ );
and  ( new_n9265_, new_n9264_, new_n9263_ );
xor  ( new_n9266_, new_n9265_, new_n2424_ );
nor  ( new_n9267_, new_n9266_, new_n9262_ );
nor  ( new_n9268_, new_n9267_, new_n9261_ );
nor  ( new_n9269_, new_n9268_, new_n9252_ );
nor  ( new_n9270_, new_n9269_, new_n9251_ );
and  ( new_n9271_, new_n9217_, new_n9164_ );
or   ( new_n9272_, new_n9271_, new_n9270_ );
and  ( new_n9273_, new_n9272_, new_n9218_ );
or   ( new_n9274_, new_n9273_, new_n9112_ );
and  ( new_n9275_, new_n9273_, new_n9112_ );
xor  ( new_n9276_, new_n8805_, new_n8803_ );
xor  ( new_n9277_, new_n9276_, new_n8809_ );
xnor ( new_n9278_, new_n8895_, new_n8891_ );
xor  ( new_n9279_, new_n9278_, new_n8901_ );
xnor ( new_n9280_, new_n8913_, new_n8909_ );
xor  ( new_n9281_, new_n9280_, new_n8919_ );
or   ( new_n9282_, new_n9281_, new_n9279_ );
and  ( new_n9283_, new_n9281_, new_n9279_ );
xor  ( new_n9284_, new_n8859_, new_n8855_ );
xnor ( new_n9285_, new_n9284_, new_n8865_ );
or   ( new_n9286_, new_n9285_, new_n9283_ );
and  ( new_n9287_, new_n9286_, new_n9282_ );
nor  ( new_n9288_, new_n9287_, new_n9277_ );
nand ( new_n9289_, new_n9287_, new_n9277_ );
xor  ( new_n9290_, new_n9006_, new_n9004_ );
xnor ( new_n9291_, new_n9290_, new_n9010_ );
and  ( new_n9292_, new_n9291_, new_n9289_ );
or   ( new_n9293_, new_n9292_, new_n9288_ );
or   ( new_n9294_, new_n9293_, new_n9275_ );
and  ( new_n9295_, new_n9294_, new_n9274_ );
or   ( new_n9296_, new_n9295_, new_n9065_ );
nand ( new_n9297_, new_n9295_, new_n9065_ );
xor  ( new_n9298_, new_n9012_, new_n9002_ );
xor  ( new_n9299_, new_n9298_, new_n9024_ );
xnor ( new_n9300_, new_n8923_, new_n8869_ );
xor  ( new_n9301_, new_n9300_, new_n8976_ );
nor  ( new_n9302_, new_n9301_, new_n9299_ );
and  ( new_n9303_, new_n9301_, new_n9299_ );
xor  ( new_n9304_, new_n8811_, new_n8801_ );
xnor ( new_n9305_, new_n9304_, new_n8815_ );
nor  ( new_n9306_, new_n9305_, new_n9303_ );
nor  ( new_n9307_, new_n9306_, new_n9302_ );
nand ( new_n9308_, new_n9307_, new_n9297_ );
and  ( new_n9309_, new_n9308_, new_n9296_ );
nor  ( new_n9310_, new_n9309_, new_n9047_ );
nand ( new_n9311_, new_n9309_, new_n9047_ );
xor  ( new_n9312_, new_n8627_, new_n8575_ );
xor  ( new_n9313_, new_n9312_, new_n8681_ );
xor  ( new_n9314_, new_n8509_, new_n8499_ );
xor  ( new_n9315_, new_n9314_, new_n8521_ );
and  ( new_n9316_, new_n9315_, new_n9313_ );
nor  ( new_n9317_, new_n9315_, new_n9313_ );
xor  ( new_n9318_, new_n8790_, new_n8788_ );
xor  ( new_n9319_, new_n9318_, new_n8795_ );
nor  ( new_n9320_, new_n9319_, new_n9317_ );
nor  ( new_n9321_, new_n9320_, new_n9316_ );
and  ( new_n9322_, new_n9321_, new_n9311_ );
or   ( new_n9323_, new_n9322_, new_n9310_ );
xor  ( new_n9324_, new_n8699_, new_n8476_ );
xor  ( new_n9325_, new_n9324_, new_n8711_ );
or   ( new_n9326_, new_n9325_, new_n9323_ );
and  ( new_n9327_, new_n9325_, new_n9323_ );
xor  ( new_n9328_, new_n8758_, new_n8748_ );
xor  ( new_n9329_, new_n9328_, new_n9030_ );
or   ( new_n9330_, new_n9329_, new_n9327_ );
and  ( new_n9331_, new_n9330_, new_n9326_ );
nor  ( new_n9332_, new_n9331_, new_n9045_ );
xnor ( new_n9333_, new_n8744_, new_n8742_ );
xor  ( new_n9334_, new_n9333_, new_n9040_ );
and  ( new_n9335_, new_n9334_, new_n9332_ );
xor  ( new_n9336_, new_n9325_, new_n9323_ );
xnor ( new_n9337_, new_n9336_, new_n9329_ );
xnor ( new_n9338_, new_n8772_, new_n8770_ );
xor  ( new_n9339_, new_n9338_, new_n8784_ );
xnor ( new_n9340_, new_n8849_, new_n8833_ );
xor  ( new_n9341_, new_n9340_, new_n8867_ );
xor  ( new_n9342_, new_n9105_, new_n9088_ );
xor  ( new_n9343_, new_n9342_, new_n9108_ );
xnor ( new_n9344_, new_n9069_, new_n9067_ );
xor  ( new_n9345_, new_n9344_, new_n9073_ );
nand ( new_n9346_, new_n9345_, new_n9343_ );
or   ( new_n9347_, new_n9345_, new_n9343_ );
xor  ( new_n9348_, new_n9079_, new_n9077_ );
xnor ( new_n9349_, new_n9348_, new_n9083_ );
nand ( new_n9350_, new_n9349_, new_n9347_ );
and  ( new_n9351_, new_n9350_, new_n9346_ );
nor  ( new_n9352_, new_n9351_, new_n9341_ );
and  ( new_n9353_, new_n9351_, new_n9341_ );
xnor ( new_n9354_, new_n9144_, new_n9128_ );
xor  ( new_n9355_, new_n9354_, new_n9162_ );
xnor ( new_n9356_, new_n9197_, new_n9180_ );
xor  ( new_n9357_, new_n9356_, new_n9215_ );
nor  ( new_n9358_, new_n9357_, new_n9355_ );
and  ( new_n9359_, new_n9357_, new_n9355_ );
xor  ( new_n9360_, new_n9250_, new_n9234_ );
xnor ( new_n9361_, new_n9360_, new_n9268_ );
nor  ( new_n9362_, new_n9361_, new_n9359_ );
nor  ( new_n9363_, new_n9362_, new_n9358_ );
nor  ( new_n9364_, new_n9363_, new_n9353_ );
or   ( new_n9365_, new_n9364_, new_n9352_ );
or   ( new_n9366_, new_n1135_, new_n4995_ );
or   ( new_n9367_, new_n1137_, new_n4603_ );
and  ( new_n9368_, new_n9367_, new_n9366_ );
xor  ( new_n9369_, new_n9368_, new_n896_ );
or   ( new_n9370_, new_n897_, new_n5171_ );
or   ( new_n9371_, new_n899_, new_n4859_ );
and  ( new_n9372_, new_n9371_, new_n9370_ );
xor  ( new_n9373_, new_n9372_, new_n748_ );
or   ( new_n9374_, new_n9373_, new_n9369_ );
and  ( new_n9375_, new_n9373_, new_n9369_ );
or   ( new_n9376_, new_n755_, new_n5570_ );
or   ( new_n9377_, new_n757_, new_n5428_ );
and  ( new_n9378_, new_n9377_, new_n9376_ );
xor  ( new_n9379_, new_n9378_, new_n523_ );
or   ( new_n9380_, new_n9379_, new_n9375_ );
and  ( new_n9381_, new_n9380_, new_n9374_ );
or   ( new_n9382_, new_n524_, new_n6219_ );
or   ( new_n9383_, new_n526_, new_n5899_ );
and  ( new_n9384_, new_n9383_, new_n9382_ );
xor  ( new_n9385_, new_n9384_, new_n403_ );
or   ( new_n9386_, new_n409_, new_n6589_ );
or   ( new_n9387_, new_n411_, new_n6425_ );
and  ( new_n9388_, new_n9387_, new_n9386_ );
xor  ( new_n9389_, new_n9388_, new_n328_ );
or   ( new_n9390_, new_n9389_, new_n9385_ );
and  ( new_n9391_, new_n9389_, new_n9385_ );
or   ( new_n9392_, new_n337_, new_n7149_ );
or   ( new_n9393_, new_n340_, new_n6943_ );
and  ( new_n9394_, new_n9393_, new_n9392_ );
xor  ( new_n9395_, new_n9394_, new_n332_ );
or   ( new_n9396_, new_n9395_, new_n9391_ );
and  ( new_n9397_, new_n9396_, new_n9390_ );
or   ( new_n9398_, new_n9397_, new_n9381_ );
and  ( new_n9399_, new_n9397_, new_n9381_ );
or   ( new_n9400_, new_n1844_, new_n3696_ );
or   ( new_n9401_, new_n1846_, new_n3306_ );
and  ( new_n9402_, new_n9401_, new_n9400_ );
xor  ( new_n9403_, new_n9402_, new_n1586_ );
or   ( new_n9404_, new_n1593_, new_n3820_ );
or   ( new_n9405_, new_n1595_, new_n3694_ );
and  ( new_n9406_, new_n9405_, new_n9404_ );
xor  ( new_n9407_, new_n9406_, new_n1358_ );
nor  ( new_n9408_, new_n9407_, new_n9403_ );
and  ( new_n9409_, new_n9407_, new_n9403_ );
or   ( new_n9410_, new_n1364_, new_n4267_ );
or   ( new_n9411_, new_n1366_, new_n4069_ );
and  ( new_n9412_, new_n9411_, new_n9410_ );
xor  ( new_n9413_, new_n9412_, new_n1129_ );
nor  ( new_n9414_, new_n9413_, new_n9409_ );
nor  ( new_n9415_, new_n9414_, new_n9408_ );
or   ( new_n9416_, new_n9415_, new_n9399_ );
and  ( new_n9417_, new_n9416_, new_n9398_ );
not  ( new_n9418_, RIbb2d9f0_61 );
and  ( new_n9419_, RIbb2d900_63, RIbb2d978_62 );
nor  ( new_n9420_, new_n9419_, new_n9418_ );
not  ( new_n9421_, new_n9420_ );
not  ( new_n9422_, new_n9187_ );
or   ( new_n9423_, new_n9422_, new_n333_ );
not  ( new_n9424_, new_n9185_ );
or   ( new_n9425_, new_n9424_, new_n339_ );
and  ( new_n9426_, new_n9425_, new_n9423_ );
xor  ( new_n9427_, new_n9426_, new_n8873_ );
and  ( new_n9428_, new_n9427_, new_n9421_ );
or   ( new_n9429_, new_n9427_, new_n9421_ );
or   ( new_n9430_, new_n8874_, new_n313_ );
or   ( new_n9431_, new_n8876_, new_n319_ );
and  ( new_n9432_, new_n9431_, new_n9430_ );
xor  ( new_n9433_, new_n9432_, new_n8257_ );
and  ( new_n9434_, new_n9433_, new_n9429_ );
or   ( new_n9435_, new_n9434_, new_n9428_ );
or   ( new_n9436_, new_n6645_, new_n419_ );
or   ( new_n9437_, new_n6647_, new_n348_ );
and  ( new_n9438_, new_n9437_, new_n9436_ );
xor  ( new_n9439_, new_n9438_, new_n6166_ );
or   ( new_n9440_, new_n6173_, new_n509_ );
or   ( new_n9441_, new_n6175_, new_n443_ );
and  ( new_n9442_, new_n9441_, new_n9440_ );
xor  ( new_n9443_, new_n9442_, new_n5597_ );
or   ( new_n9444_, new_n9443_, new_n9439_ );
and  ( new_n9445_, new_n9443_, new_n9439_ );
or   ( new_n9446_, new_n5604_, new_n775_ );
or   ( new_n9447_, new_n5606_, new_n515_ );
and  ( new_n9448_, new_n9447_, new_n9446_ );
xor  ( new_n9449_, new_n9448_, new_n5206_ );
or   ( new_n9450_, new_n9449_, new_n9445_ );
and  ( new_n9451_, new_n9450_, new_n9444_ );
or   ( new_n9452_, new_n9451_, new_n9435_ );
and  ( new_n9453_, new_n9451_, new_n9435_ );
or   ( new_n9454_, new_n8264_, new_n279_ );
or   ( new_n9455_, new_n8266_, new_n285_ );
and  ( new_n9456_, new_n9455_, new_n9454_ );
xor  ( new_n9457_, new_n9456_, new_n7725_ );
or   ( new_n9458_, new_n7732_, new_n294_ );
or   ( new_n9459_, new_n7734_, new_n301_ );
and  ( new_n9460_, new_n9459_, new_n9458_ );
xor  ( new_n9461_, new_n9460_, new_n7177_ );
nor  ( new_n9462_, new_n9461_, new_n9457_ );
and  ( new_n9463_, new_n9461_, new_n9457_ );
or   ( new_n9464_, new_n7184_, new_n264_ );
or   ( new_n9465_, new_n7186_, new_n270_ );
and  ( new_n9466_, new_n9465_, new_n9464_ );
xor  ( new_n9467_, new_n9466_, new_n6638_ );
nor  ( new_n9468_, new_n9467_, new_n9463_ );
nor  ( new_n9469_, new_n9468_, new_n9462_ );
or   ( new_n9470_, new_n9469_, new_n9453_ );
and  ( new_n9471_, new_n9470_, new_n9452_ );
nor  ( new_n9472_, new_n9471_, new_n9417_ );
nand ( new_n9473_, new_n9471_, new_n9417_ );
or   ( new_n9474_, new_n3896_, new_n1523_ );
or   ( new_n9475_, new_n3898_, new_n1525_ );
and  ( new_n9476_, new_n9475_, new_n9474_ );
xor  ( new_n9477_, new_n9476_, new_n3460_ );
or   ( new_n9478_, new_n3461_, new_n1899_ );
or   ( new_n9479_, new_n3463_, new_n1754_ );
and  ( new_n9480_, new_n9479_, new_n9478_ );
xor  ( new_n9481_, new_n9480_, new_n3116_ );
or   ( new_n9482_, new_n9481_, new_n9477_ );
and  ( new_n9483_, new_n9481_, new_n9477_ );
or   ( new_n9484_, new_n3117_, new_n2178_ );
or   ( new_n9485_, new_n3119_, new_n2057_ );
and  ( new_n9486_, new_n9485_, new_n9484_ );
xor  ( new_n9487_, new_n9486_, new_n2800_ );
or   ( new_n9488_, new_n9487_, new_n9483_ );
and  ( new_n9489_, new_n9488_, new_n9482_ );
or   ( new_n9490_, new_n2807_, new_n2475_ );
or   ( new_n9491_, new_n2809_, new_n2291_ );
and  ( new_n9492_, new_n9491_, new_n9490_ );
xor  ( new_n9493_, new_n9492_, new_n2424_ );
or   ( new_n9494_, new_n2425_, new_n2751_ );
or   ( new_n9495_, new_n2427_, new_n2646_ );
and  ( new_n9496_, new_n9495_, new_n9494_ );
xor  ( new_n9497_, new_n9496_, new_n2121_ );
or   ( new_n9498_, new_n9497_, new_n9493_ );
and  ( new_n9499_, new_n9497_, new_n9493_ );
or   ( new_n9500_, new_n2122_, new_n3178_ );
or   ( new_n9501_, new_n2124_, new_n2981_ );
and  ( new_n9502_, new_n9501_, new_n9500_ );
xor  ( new_n9503_, new_n9502_, new_n1843_ );
or   ( new_n9504_, new_n9503_, new_n9499_ );
and  ( new_n9505_, new_n9504_, new_n9498_ );
nor  ( new_n9506_, new_n9505_, new_n9489_ );
nand ( new_n9507_, new_n9505_, new_n9489_ );
or   ( new_n9508_, new_n5207_, new_n886_ );
or   ( new_n9509_, new_n5209_, new_n805_ );
and  ( new_n9510_, new_n9509_, new_n9508_ );
xor  ( new_n9511_, new_n9510_, new_n4708_ );
or   ( new_n9512_, new_n4709_, new_n1168_ );
or   ( new_n9513_, new_n4711_, new_n986_ );
and  ( new_n9514_, new_n9513_, new_n9512_ );
xor  ( new_n9515_, new_n9514_, new_n4295_ );
nor  ( new_n9516_, new_n9515_, new_n9511_ );
and  ( new_n9517_, new_n9515_, new_n9511_ );
or   ( new_n9518_, new_n4302_, new_n1318_ );
or   ( new_n9519_, new_n4304_, new_n1213_ );
and  ( new_n9520_, new_n9519_, new_n9518_ );
xor  ( new_n9521_, new_n9520_, new_n3895_ );
nor  ( new_n9522_, new_n9521_, new_n9517_ );
nor  ( new_n9523_, new_n9522_, new_n9516_ );
not  ( new_n9524_, new_n9523_ );
and  ( new_n9525_, new_n9524_, new_n9507_ );
or   ( new_n9526_, new_n9525_, new_n9506_ );
and  ( new_n9527_, new_n9526_, new_n9473_ );
or   ( new_n9528_, new_n9527_, new_n9472_ );
not  ( new_n9529_, new_n9088_ );
or   ( new_n9530_, new_n317_, new_n8117_ );
or   ( new_n9531_, new_n320_, new_n7373_ );
and  ( new_n9532_, new_n9531_, new_n9530_ );
xor  ( new_n9533_, new_n9532_, new_n312_ );
or   ( new_n9534_, new_n283_, new_n8352_ );
or   ( new_n9535_, new_n286_, new_n8115_ );
and  ( new_n9536_, new_n9535_, new_n9534_ );
xor  ( new_n9537_, new_n9536_, new_n278_ );
or   ( new_n9538_, new_n9537_, new_n9533_ );
and  ( new_n9539_, new_n9537_, new_n9533_ );
or   ( new_n9540_, new_n299_, new_n8995_ );
or   ( new_n9541_, new_n302_, new_n8481_ );
and  ( new_n9542_, new_n9541_, new_n9540_ );
xor  ( new_n9543_, new_n9542_, new_n293_ );
or   ( new_n9544_, new_n9543_, new_n9539_ );
and  ( new_n9545_, new_n9544_, new_n9538_ );
nor  ( new_n9546_, new_n9545_, new_n9529_ );
nand ( new_n9547_, new_n9545_, new_n9529_ );
xor  ( new_n9548_, new_n9096_, new_n9092_ );
xnor ( new_n9549_, new_n9548_, new_n9103_ );
and  ( new_n9550_, new_n9549_, new_n9547_ );
or   ( new_n9551_, new_n9550_, new_n9546_ );
xnor ( new_n9552_, new_n9242_, new_n9238_ );
xor  ( new_n9553_, new_n9552_, new_n9248_ );
xnor ( new_n9554_, new_n9226_, new_n9222_ );
xor  ( new_n9555_, new_n9554_, new_n9232_ );
or   ( new_n9556_, new_n9555_, new_n9553_ );
and  ( new_n9557_, new_n9555_, new_n9553_ );
xor  ( new_n9558_, new_n9260_, new_n9256_ );
xnor ( new_n9559_, new_n9558_, new_n9266_ );
or   ( new_n9560_, new_n9559_, new_n9557_ );
and  ( new_n9561_, new_n9560_, new_n9556_ );
or   ( new_n9562_, new_n9561_, new_n9551_ );
and  ( new_n9563_, new_n9561_, new_n9551_ );
xnor ( new_n9564_, new_n9136_, new_n9132_ );
xor  ( new_n9565_, new_n9564_, new_n9142_ );
xnor ( new_n9566_, new_n9120_, new_n9116_ );
xor  ( new_n9567_, new_n9566_, new_n9126_ );
nor  ( new_n9568_, new_n9567_, new_n9565_ );
and  ( new_n9569_, new_n9567_, new_n9565_ );
xor  ( new_n9570_, new_n9154_, new_n9150_ );
xnor ( new_n9571_, new_n9570_, new_n9160_ );
nor  ( new_n9572_, new_n9571_, new_n9569_ );
nor  ( new_n9573_, new_n9572_, new_n9568_ );
or   ( new_n9574_, new_n9573_, new_n9563_ );
and  ( new_n9575_, new_n9574_, new_n9562_ );
nand ( new_n9576_, new_n9575_, new_n9528_ );
or   ( new_n9577_, new_n9575_, new_n9528_ );
xor  ( new_n9578_, new_n8879_, new_n8872_ );
xor  ( new_n9579_, new_n9578_, new_n8885_ );
xnor ( new_n9580_, new_n9189_, new_n9184_ );
xor  ( new_n9581_, new_n9580_, new_n9195_ );
xnor ( new_n9582_, new_n9172_, new_n9168_ );
xor  ( new_n9583_, new_n9582_, new_n9178_ );
or   ( new_n9584_, new_n9583_, new_n9581_ );
and  ( new_n9585_, new_n9583_, new_n9581_ );
xor  ( new_n9586_, new_n9207_, new_n9203_ );
xnor ( new_n9587_, new_n9586_, new_n9213_ );
or   ( new_n9588_, new_n9587_, new_n9585_ );
and  ( new_n9589_, new_n9588_, new_n9584_ );
nor  ( new_n9590_, new_n9589_, new_n9579_ );
and  ( new_n9591_, new_n9589_, new_n9579_ );
xor  ( new_n9592_, new_n9281_, new_n9279_ );
xnor ( new_n9593_, new_n9592_, new_n9285_ );
not  ( new_n9594_, new_n9593_ );
nor  ( new_n9595_, new_n9594_, new_n9591_ );
nor  ( new_n9596_, new_n9595_, new_n9590_ );
nand ( new_n9597_, new_n9596_, new_n9577_ );
and  ( new_n9598_, new_n9597_, new_n9576_ );
or   ( new_n9599_, new_n9598_, new_n9365_ );
nand ( new_n9600_, new_n9598_, new_n9365_ );
xnor ( new_n9601_, new_n8903_, new_n8887_ );
xor  ( new_n9602_, new_n9601_, new_n8921_ );
xnor ( new_n9603_, new_n9287_, new_n9277_ );
xor  ( new_n9604_, new_n9603_, new_n9291_ );
nor  ( new_n9605_, new_n9604_, new_n9602_ );
and  ( new_n9606_, new_n9604_, new_n9602_ );
xor  ( new_n9607_, new_n9057_, new_n9055_ );
xnor ( new_n9608_, new_n9607_, new_n9060_ );
not  ( new_n9609_, new_n9608_ );
nor  ( new_n9610_, new_n9609_, new_n9606_ );
nor  ( new_n9611_, new_n9610_, new_n9605_ );
nand ( new_n9612_, new_n9611_, new_n9600_ );
and  ( new_n9613_, new_n9612_, new_n9599_ );
nor  ( new_n9614_, new_n9613_, new_n9339_ );
nand ( new_n9615_, new_n9613_, new_n9339_ );
xor  ( new_n9616_, new_n9273_, new_n9112_ );
xor  ( new_n9617_, new_n9616_, new_n9293_ );
xnor ( new_n9618_, new_n9301_, new_n9299_ );
xor  ( new_n9619_, new_n9618_, new_n9305_ );
nand ( new_n9620_, new_n9619_, new_n9617_ );
or   ( new_n9621_, new_n9619_, new_n9617_ );
xor  ( new_n9622_, new_n9051_, new_n9049_ );
xor  ( new_n9623_, new_n9622_, new_n9063_ );
nand ( new_n9624_, new_n9623_, new_n9621_ );
and  ( new_n9625_, new_n9624_, new_n9620_ );
and  ( new_n9626_, new_n9625_, new_n9615_ );
or   ( new_n9627_, new_n9626_, new_n9614_ );
xor  ( new_n9628_, new_n8979_, new_n8817_ );
xor  ( new_n9629_, new_n9628_, new_n9026_ );
xor  ( new_n9630_, new_n9295_, new_n9065_ );
xor  ( new_n9631_, new_n9630_, new_n9307_ );
or   ( new_n9632_, new_n9631_, new_n9629_ );
and  ( new_n9633_, new_n9631_, new_n9629_ );
xor  ( new_n9634_, new_n9315_, new_n9313_ );
xnor ( new_n9635_, new_n9634_, new_n9319_ );
not  ( new_n9636_, new_n9635_ );
or   ( new_n9637_, new_n9636_, new_n9633_ );
and  ( new_n9638_, new_n9637_, new_n9632_ );
or   ( new_n9639_, new_n9638_, new_n9627_ );
and  ( new_n9640_, new_n9638_, new_n9627_ );
xor  ( new_n9641_, new_n8797_, new_n8786_ );
xor  ( new_n9642_, new_n9641_, new_n9028_ );
or   ( new_n9643_, new_n9642_, new_n9640_ );
nand ( new_n9644_, new_n9643_, new_n9639_ );
and  ( new_n9645_, new_n9644_, new_n9337_ );
xor  ( new_n9646_, new_n9331_, new_n9045_ );
and  ( new_n9647_, new_n9646_, new_n9645_ );
xnor ( new_n9648_, new_n9644_, new_n9337_ );
xor  ( new_n9649_, new_n9638_, new_n9627_ );
xor  ( new_n9650_, new_n9649_, new_n9642_ );
xor  ( new_n9651_, new_n9619_, new_n9617_ );
xor  ( new_n9652_, new_n9651_, new_n9623_ );
xor  ( new_n9653_, new_n9357_, new_n9355_ );
xor  ( new_n9654_, new_n9653_, new_n9361_ );
xnor ( new_n9655_, new_n9555_, new_n9553_ );
xor  ( new_n9656_, new_n9655_, new_n9559_ );
xnor ( new_n9657_, new_n9567_, new_n9565_ );
xor  ( new_n9658_, new_n9657_, new_n9571_ );
nand ( new_n9659_, new_n9658_, new_n9656_ );
nor  ( new_n9660_, new_n9658_, new_n9656_ );
xor  ( new_n9661_, new_n9545_, new_n9529_ );
xor  ( new_n9662_, new_n9661_, new_n9549_ );
or   ( new_n9663_, new_n9662_, new_n9660_ );
and  ( new_n9664_, new_n9663_, new_n9659_ );
nor  ( new_n9665_, new_n9664_, new_n9654_ );
and  ( new_n9666_, new_n9664_, new_n9654_ );
xnor ( new_n9667_, new_n9397_, new_n9381_ );
xor  ( new_n9668_, new_n9667_, new_n9415_ );
xnor ( new_n9669_, new_n9451_, new_n9435_ );
xor  ( new_n9670_, new_n9669_, new_n9469_ );
nor  ( new_n9671_, new_n9670_, new_n9668_ );
and  ( new_n9672_, new_n9670_, new_n9668_ );
xor  ( new_n9673_, new_n9505_, new_n9489_ );
xor  ( new_n9674_, new_n9673_, new_n9524_ );
nor  ( new_n9675_, new_n9674_, new_n9672_ );
nor  ( new_n9676_, new_n9675_, new_n9671_ );
nor  ( new_n9677_, new_n9676_, new_n9666_ );
or   ( new_n9678_, new_n9677_, new_n9665_ );
not  ( new_n9679_, RIbb2bbf0_125 );
or   ( new_n9680_, new_n268_, new_n9679_ );
not  ( new_n9681_, RIbb2bc68_124 );
or   ( new_n9682_, new_n271_, new_n9681_ );
and  ( new_n9683_, new_n9682_, new_n9680_ );
xor  ( new_n9684_, new_n9683_, new_n263_ );
and  ( new_n9685_, RIbb2bb78_126, RIbb2f610_1 );
or   ( new_n9686_, new_n9685_, new_n9684_ );
or   ( new_n9687_, new_n317_, new_n8115_ );
or   ( new_n9688_, new_n320_, new_n8117_ );
and  ( new_n9689_, new_n9688_, new_n9687_ );
xor  ( new_n9690_, new_n9689_, new_n312_ );
or   ( new_n9691_, new_n283_, new_n8481_ );
or   ( new_n9692_, new_n286_, new_n8352_ );
and  ( new_n9693_, new_n9692_, new_n9691_ );
xor  ( new_n9694_, new_n9693_, new_n278_ );
or   ( new_n9695_, new_n9694_, new_n9690_ );
and  ( new_n9696_, new_n9694_, new_n9690_ );
or   ( new_n9697_, new_n299_, new_n9099_ );
or   ( new_n9698_, new_n302_, new_n8995_ );
and  ( new_n9699_, new_n9698_, new_n9697_ );
xor  ( new_n9700_, new_n9699_, new_n293_ );
or   ( new_n9701_, new_n9700_, new_n9696_ );
and  ( new_n9702_, new_n9701_, new_n9695_ );
and  ( new_n9703_, new_n9702_, new_n9686_ );
or   ( new_n9704_, new_n9702_, new_n9686_ );
or   ( new_n9705_, new_n268_, new_n9681_ );
or   ( new_n9706_, new_n271_, new_n9099_ );
and  ( new_n9707_, new_n9706_, new_n9705_ );
xor  ( new_n9708_, new_n9707_, new_n263_ );
and  ( new_n9709_, new_n9708_, new_n9704_ );
or   ( new_n9710_, new_n9709_, new_n9703_ );
or   ( new_n9711_, new_n9679_, new_n260_ );
xnor ( new_n9712_, new_n9389_, new_n9385_ );
xor  ( new_n9713_, new_n9712_, new_n9395_ );
nand ( new_n9714_, new_n9713_, new_n9711_ );
or   ( new_n9715_, new_n9713_, new_n9711_ );
xor  ( new_n9716_, new_n9537_, new_n9533_ );
xnor ( new_n9717_, new_n9716_, new_n9543_ );
nand ( new_n9718_, new_n9717_, new_n9715_ );
and  ( new_n9719_, new_n9718_, new_n9714_ );
and  ( new_n9720_, new_n9719_, new_n9710_ );
nor  ( new_n9721_, new_n9719_, new_n9710_ );
xnor ( new_n9722_, new_n9497_, new_n9493_ );
xor  ( new_n9723_, new_n9722_, new_n9503_ );
xnor ( new_n9724_, new_n9373_, new_n9369_ );
xor  ( new_n9725_, new_n9724_, new_n9379_ );
nor  ( new_n9726_, new_n9725_, new_n9723_ );
and  ( new_n9727_, new_n9725_, new_n9723_ );
xor  ( new_n9728_, new_n9407_, new_n9403_ );
xnor ( new_n9729_, new_n9728_, new_n9413_ );
nor  ( new_n9730_, new_n9729_, new_n9727_ );
nor  ( new_n9731_, new_n9730_, new_n9726_ );
nor  ( new_n9732_, new_n9731_, new_n9721_ );
or   ( new_n9733_, new_n9732_, new_n9720_ );
or   ( new_n9734_, new_n9422_, new_n319_ );
or   ( new_n9735_, new_n9424_, new_n333_ );
and  ( new_n9736_, new_n9735_, new_n9734_ );
xor  ( new_n9737_, new_n9736_, new_n8872_ );
xor  ( new_n9738_, RIbb2d900_63, RIbb2d978_62 );
xor  ( new_n9739_, RIbb2d978_62, new_n9418_ );
nor  ( new_n9740_, new_n9739_, new_n9738_ );
and  ( new_n9741_, new_n9740_, RIbb2d810_65 );
xor  ( new_n9742_, new_n9741_, new_n9421_ );
nand ( new_n9743_, new_n9742_, new_n9737_ );
nor  ( new_n9744_, new_n9742_, new_n9737_ );
or   ( new_n9745_, new_n8874_, new_n285_ );
or   ( new_n9746_, new_n8876_, new_n313_ );
and  ( new_n9747_, new_n9746_, new_n9745_ );
xor  ( new_n9748_, new_n9747_, new_n8257_ );
or   ( new_n9749_, new_n9748_, new_n9744_ );
and  ( new_n9750_, new_n9749_, new_n9743_ );
or   ( new_n9751_, new_n6645_, new_n443_ );
or   ( new_n9752_, new_n6647_, new_n419_ );
and  ( new_n9753_, new_n9752_, new_n9751_ );
xor  ( new_n9754_, new_n9753_, new_n6166_ );
or   ( new_n9755_, new_n6173_, new_n515_ );
or   ( new_n9756_, new_n6175_, new_n509_ );
and  ( new_n9757_, new_n9756_, new_n9755_ );
xor  ( new_n9758_, new_n9757_, new_n5597_ );
or   ( new_n9759_, new_n9758_, new_n9754_ );
and  ( new_n9760_, new_n9758_, new_n9754_ );
or   ( new_n9761_, new_n5604_, new_n805_ );
or   ( new_n9762_, new_n5606_, new_n775_ );
and  ( new_n9763_, new_n9762_, new_n9761_ );
xor  ( new_n9764_, new_n9763_, new_n5206_ );
or   ( new_n9765_, new_n9764_, new_n9760_ );
and  ( new_n9766_, new_n9765_, new_n9759_ );
or   ( new_n9767_, new_n9766_, new_n9750_ );
and  ( new_n9768_, new_n9766_, new_n9750_ );
or   ( new_n9769_, new_n8264_, new_n301_ );
or   ( new_n9770_, new_n8266_, new_n279_ );
and  ( new_n9771_, new_n9770_, new_n9769_ );
xor  ( new_n9772_, new_n9771_, new_n7725_ );
or   ( new_n9773_, new_n7732_, new_n270_ );
or   ( new_n9774_, new_n7734_, new_n294_ );
and  ( new_n9775_, new_n9774_, new_n9773_ );
xor  ( new_n9776_, new_n9775_, new_n7177_ );
nor  ( new_n9777_, new_n9776_, new_n9772_ );
and  ( new_n9778_, new_n9776_, new_n9772_ );
or   ( new_n9779_, new_n7184_, new_n348_ );
or   ( new_n9780_, new_n7186_, new_n264_ );
and  ( new_n9781_, new_n9780_, new_n9779_ );
xor  ( new_n9782_, new_n9781_, new_n6638_ );
nor  ( new_n9783_, new_n9782_, new_n9778_ );
nor  ( new_n9784_, new_n9783_, new_n9777_ );
or   ( new_n9785_, new_n9784_, new_n9768_ );
and  ( new_n9786_, new_n9785_, new_n9767_ );
or   ( new_n9787_, new_n1844_, new_n3694_ );
or   ( new_n9788_, new_n1846_, new_n3696_ );
and  ( new_n9789_, new_n9788_, new_n9787_ );
xor  ( new_n9790_, new_n9789_, new_n1586_ );
or   ( new_n9791_, new_n1593_, new_n4069_ );
or   ( new_n9792_, new_n1595_, new_n3820_ );
and  ( new_n9793_, new_n9792_, new_n9791_ );
xor  ( new_n9794_, new_n9793_, new_n1358_ );
or   ( new_n9795_, new_n9794_, new_n9790_ );
and  ( new_n9796_, new_n9794_, new_n9790_ );
or   ( new_n9797_, new_n1364_, new_n4603_ );
or   ( new_n9798_, new_n1366_, new_n4267_ );
and  ( new_n9799_, new_n9798_, new_n9797_ );
xor  ( new_n9800_, new_n9799_, new_n1129_ );
or   ( new_n9801_, new_n9800_, new_n9796_ );
and  ( new_n9802_, new_n9801_, new_n9795_ );
or   ( new_n9803_, new_n524_, new_n6425_ );
or   ( new_n9804_, new_n526_, new_n6219_ );
and  ( new_n9805_, new_n9804_, new_n9803_ );
xor  ( new_n9806_, new_n9805_, new_n403_ );
or   ( new_n9807_, new_n409_, new_n6943_ );
or   ( new_n9808_, new_n411_, new_n6589_ );
and  ( new_n9809_, new_n9808_, new_n9807_ );
xor  ( new_n9810_, new_n9809_, new_n328_ );
or   ( new_n9811_, new_n9810_, new_n9806_ );
and  ( new_n9812_, new_n9810_, new_n9806_ );
or   ( new_n9813_, new_n337_, new_n7373_ );
or   ( new_n9814_, new_n340_, new_n7149_ );
and  ( new_n9815_, new_n9814_, new_n9813_ );
xor  ( new_n9816_, new_n9815_, new_n332_ );
or   ( new_n9817_, new_n9816_, new_n9812_ );
and  ( new_n9818_, new_n9817_, new_n9811_ );
or   ( new_n9819_, new_n9818_, new_n9802_ );
and  ( new_n9820_, new_n9818_, new_n9802_ );
or   ( new_n9821_, new_n1135_, new_n4859_ );
or   ( new_n9822_, new_n1137_, new_n4995_ );
and  ( new_n9823_, new_n9822_, new_n9821_ );
xor  ( new_n9824_, new_n9823_, new_n896_ );
or   ( new_n9825_, new_n897_, new_n5428_ );
or   ( new_n9826_, new_n899_, new_n5171_ );
and  ( new_n9827_, new_n9826_, new_n9825_ );
xor  ( new_n9828_, new_n9827_, new_n748_ );
nor  ( new_n9829_, new_n9828_, new_n9824_ );
and  ( new_n9830_, new_n9828_, new_n9824_ );
or   ( new_n9831_, new_n755_, new_n5899_ );
or   ( new_n9832_, new_n757_, new_n5570_ );
and  ( new_n9833_, new_n9832_, new_n9831_ );
xor  ( new_n9834_, new_n9833_, new_n523_ );
nor  ( new_n9835_, new_n9834_, new_n9830_ );
nor  ( new_n9836_, new_n9835_, new_n9829_ );
or   ( new_n9837_, new_n9836_, new_n9820_ );
and  ( new_n9838_, new_n9837_, new_n9819_ );
or   ( new_n9839_, new_n9838_, new_n9786_ );
or   ( new_n9840_, new_n2807_, new_n2646_ );
or   ( new_n9841_, new_n2809_, new_n2475_ );
and  ( new_n9842_, new_n9841_, new_n9840_ );
xor  ( new_n9843_, new_n9842_, new_n2424_ );
or   ( new_n9844_, new_n2425_, new_n2981_ );
or   ( new_n9845_, new_n2427_, new_n2751_ );
and  ( new_n9846_, new_n9845_, new_n9844_ );
xor  ( new_n9847_, new_n9846_, new_n2121_ );
or   ( new_n9848_, new_n9847_, new_n9843_ );
and  ( new_n9849_, new_n9847_, new_n9843_ );
or   ( new_n9850_, new_n2122_, new_n3306_ );
or   ( new_n9851_, new_n2124_, new_n3178_ );
and  ( new_n9852_, new_n9851_, new_n9850_ );
xor  ( new_n9853_, new_n9852_, new_n1843_ );
or   ( new_n9854_, new_n9853_, new_n9849_ );
and  ( new_n9855_, new_n9854_, new_n9848_ );
or   ( new_n9856_, new_n5207_, new_n986_ );
or   ( new_n9857_, new_n5209_, new_n886_ );
and  ( new_n9858_, new_n9857_, new_n9856_ );
xor  ( new_n9859_, new_n9858_, new_n4708_ );
or   ( new_n9860_, new_n4709_, new_n1213_ );
or   ( new_n9861_, new_n4711_, new_n1168_ );
and  ( new_n9862_, new_n9861_, new_n9860_ );
xor  ( new_n9863_, new_n9862_, new_n4295_ );
or   ( new_n9864_, new_n9863_, new_n9859_ );
and  ( new_n9865_, new_n9863_, new_n9859_ );
or   ( new_n9866_, new_n4302_, new_n1525_ );
or   ( new_n9867_, new_n4304_, new_n1318_ );
and  ( new_n9868_, new_n9867_, new_n9866_ );
xor  ( new_n9869_, new_n9868_, new_n3895_ );
or   ( new_n9870_, new_n9869_, new_n9865_ );
and  ( new_n9871_, new_n9870_, new_n9864_ );
or   ( new_n9872_, new_n9871_, new_n9855_ );
and  ( new_n9873_, new_n9871_, new_n9855_ );
or   ( new_n9874_, new_n3896_, new_n1754_ );
or   ( new_n9875_, new_n3898_, new_n1523_ );
and  ( new_n9876_, new_n9875_, new_n9874_ );
xor  ( new_n9877_, new_n9876_, new_n3460_ );
or   ( new_n9878_, new_n3461_, new_n2057_ );
or   ( new_n9879_, new_n3463_, new_n1899_ );
and  ( new_n9880_, new_n9879_, new_n9878_ );
xor  ( new_n9881_, new_n9880_, new_n3116_ );
nor  ( new_n9882_, new_n9881_, new_n9877_ );
and  ( new_n9883_, new_n9881_, new_n9877_ );
or   ( new_n9884_, new_n3117_, new_n2291_ );
or   ( new_n9885_, new_n3119_, new_n2178_ );
and  ( new_n9886_, new_n9885_, new_n9884_ );
xor  ( new_n9887_, new_n9886_, new_n2800_ );
nor  ( new_n9888_, new_n9887_, new_n9883_ );
nor  ( new_n9889_, new_n9888_, new_n9882_ );
or   ( new_n9890_, new_n9889_, new_n9873_ );
and  ( new_n9891_, new_n9890_, new_n9872_ );
and  ( new_n9892_, new_n9838_, new_n9786_ );
or   ( new_n9893_, new_n9892_, new_n9891_ );
and  ( new_n9894_, new_n9893_, new_n9839_ );
or   ( new_n9895_, new_n9894_, new_n9733_ );
nand ( new_n9896_, new_n9894_, new_n9733_ );
xor  ( new_n9897_, new_n9461_, new_n9457_ );
xnor ( new_n9898_, new_n9897_, new_n9467_ );
not  ( new_n9899_, new_n9898_ );
xor  ( new_n9900_, new_n9427_, new_n9421_ );
xor  ( new_n9901_, new_n9900_, new_n9433_ );
nand ( new_n9902_, new_n9901_, new_n9899_ );
xnor ( new_n9903_, new_n9443_, new_n9439_ );
xor  ( new_n9904_, new_n9903_, new_n9449_ );
xnor ( new_n9905_, new_n9481_, new_n9477_ );
xor  ( new_n9906_, new_n9905_, new_n9487_ );
or   ( new_n9907_, new_n9906_, new_n9904_ );
and  ( new_n9908_, new_n9906_, new_n9904_ );
xnor ( new_n9909_, new_n9515_, new_n9511_ );
xor  ( new_n9910_, new_n9909_, new_n9521_ );
or   ( new_n9911_, new_n9910_, new_n9908_ );
and  ( new_n9912_, new_n9911_, new_n9907_ );
nor  ( new_n9913_, new_n9912_, new_n9902_ );
and  ( new_n9914_, new_n9912_, new_n9902_ );
xor  ( new_n9915_, new_n9583_, new_n9581_ );
xnor ( new_n9916_, new_n9915_, new_n9587_ );
not  ( new_n9917_, new_n9916_ );
nor  ( new_n9918_, new_n9917_, new_n9914_ );
nor  ( new_n9919_, new_n9918_, new_n9913_ );
nand ( new_n9920_, new_n9919_, new_n9896_ );
and  ( new_n9921_, new_n9920_, new_n9895_ );
or   ( new_n9922_, new_n9921_, new_n9678_ );
nand ( new_n9923_, new_n9921_, new_n9678_ );
xor  ( new_n9924_, new_n9345_, new_n9343_ );
xor  ( new_n9925_, new_n9924_, new_n9349_ );
xnor ( new_n9926_, new_n9561_, new_n9551_ );
xor  ( new_n9927_, new_n9926_, new_n9573_ );
and  ( new_n9928_, new_n9927_, new_n9925_ );
nor  ( new_n9929_, new_n9927_, new_n9925_ );
xor  ( new_n9930_, new_n9589_, new_n9579_ );
xor  ( new_n9931_, new_n9930_, new_n9594_ );
nor  ( new_n9932_, new_n9931_, new_n9929_ );
nor  ( new_n9933_, new_n9932_, new_n9928_ );
nand ( new_n9934_, new_n9933_, new_n9923_ );
and  ( new_n9935_, new_n9934_, new_n9922_ );
nor  ( new_n9936_, new_n9935_, new_n9652_ );
nand ( new_n9937_, new_n9935_, new_n9652_ );
xnor ( new_n9938_, new_n9085_, new_n9075_ );
xor  ( new_n9939_, new_n9938_, new_n9110_ );
xnor ( new_n9940_, new_n9217_, new_n9164_ );
xor  ( new_n9941_, new_n9940_, new_n9270_ );
or   ( new_n9942_, new_n9941_, new_n9939_ );
and  ( new_n9943_, new_n9941_, new_n9939_ );
xor  ( new_n9944_, new_n9604_, new_n9602_ );
xor  ( new_n9945_, new_n9944_, new_n9609_ );
or   ( new_n9946_, new_n9945_, new_n9943_ );
and  ( new_n9947_, new_n9946_, new_n9942_ );
and  ( new_n9948_, new_n9947_, new_n9937_ );
or   ( new_n9949_, new_n9948_, new_n9936_ );
xor  ( new_n9950_, new_n9613_, new_n9339_ );
xor  ( new_n9951_, new_n9950_, new_n9625_ );
or   ( new_n9952_, new_n9951_, new_n9949_ );
and  ( new_n9953_, new_n9951_, new_n9949_ );
xor  ( new_n9954_, new_n9631_, new_n9629_ );
xor  ( new_n9955_, new_n9954_, new_n9636_ );
or   ( new_n9956_, new_n9955_, new_n9953_ );
and  ( new_n9957_, new_n9956_, new_n9952_ );
or   ( new_n9958_, new_n9957_, new_n9650_ );
and  ( new_n9959_, new_n9957_, new_n9650_ );
xor  ( new_n9960_, new_n9309_, new_n9047_ );
xor  ( new_n9961_, new_n9960_, new_n9321_ );
or   ( new_n9962_, new_n9961_, new_n9959_ );
and  ( new_n9963_, new_n9962_, new_n9958_ );
nor  ( new_n9964_, new_n9963_, new_n9648_ );
xor  ( new_n9965_, new_n9351_, new_n9341_ );
xor  ( new_n9966_, new_n9965_, new_n9363_ );
xor  ( new_n9967_, new_n9664_, new_n9654_ );
xor  ( new_n9968_, new_n9967_, new_n9676_ );
xor  ( new_n9969_, new_n9471_, new_n9417_ );
xor  ( new_n9970_, new_n9969_, new_n9526_ );
or   ( new_n9971_, new_n9970_, new_n9968_ );
and  ( new_n9972_, new_n9970_, new_n9968_ );
xor  ( new_n9973_, new_n9927_, new_n9925_ );
xnor ( new_n9974_, new_n9973_, new_n9931_ );
not  ( new_n9975_, new_n9974_ );
or   ( new_n9976_, new_n9975_, new_n9972_ );
and  ( new_n9977_, new_n9976_, new_n9971_ );
or   ( new_n9978_, new_n9977_, new_n9966_ );
and  ( new_n9979_, new_n9977_, new_n9966_ );
xnor ( new_n9980_, new_n9702_, new_n9686_ );
xor  ( new_n9981_, new_n9980_, new_n9708_ );
xor  ( new_n9982_, new_n9713_, new_n9711_ );
xor  ( new_n9983_, new_n9982_, new_n9717_ );
nor  ( new_n9984_, new_n9983_, new_n9981_ );
nand ( new_n9985_, new_n9983_, new_n9981_ );
xnor ( new_n9986_, new_n9725_, new_n9723_ );
xor  ( new_n9987_, new_n9986_, new_n9729_ );
and  ( new_n9988_, new_n9987_, new_n9985_ );
or   ( new_n9989_, new_n9988_, new_n9984_ );
xnor ( new_n9990_, new_n9670_, new_n9668_ );
xor  ( new_n9991_, new_n9990_, new_n9674_ );
nand ( new_n9992_, new_n9991_, new_n9989_ );
nor  ( new_n9993_, new_n9991_, new_n9989_ );
xnor ( new_n9994_, new_n9766_, new_n9750_ );
xor  ( new_n9995_, new_n9994_, new_n9784_ );
xnor ( new_n9996_, new_n9818_, new_n9802_ );
xor  ( new_n9997_, new_n9996_, new_n9836_ );
nor  ( new_n9998_, new_n9997_, new_n9995_ );
and  ( new_n9999_, new_n9997_, new_n9995_ );
xor  ( new_n10000_, new_n9871_, new_n9855_ );
xnor ( new_n10001_, new_n10000_, new_n9889_ );
nor  ( new_n10002_, new_n10001_, new_n9999_ );
nor  ( new_n10003_, new_n10002_, new_n9998_ );
or   ( new_n10004_, new_n10003_, new_n9993_ );
and  ( new_n10005_, new_n10004_, new_n9992_ );
xor  ( new_n10006_, new_n9719_, new_n9710_ );
xor  ( new_n10007_, new_n10006_, new_n9731_ );
xor  ( new_n10008_, new_n9912_, new_n9902_ );
xor  ( new_n10009_, new_n10008_, new_n9917_ );
or   ( new_n10010_, new_n10009_, new_n10007_ );
and  ( new_n10011_, new_n10009_, new_n10007_ );
xor  ( new_n10012_, new_n9658_, new_n9656_ );
xnor ( new_n10013_, new_n10012_, new_n9662_ );
not  ( new_n10014_, new_n10013_ );
or   ( new_n10015_, new_n10014_, new_n10011_ );
and  ( new_n10016_, new_n10015_, new_n10010_ );
or   ( new_n10017_, new_n10016_, new_n10005_ );
and  ( new_n10018_, new_n10016_, new_n10005_ );
xor  ( new_n10019_, new_n9906_, new_n9904_ );
xor  ( new_n10020_, new_n10019_, new_n9910_ );
xnor ( new_n10021_, new_n9863_, new_n9859_ );
xor  ( new_n10022_, new_n10021_, new_n9869_ );
xnor ( new_n10023_, new_n9758_, new_n9754_ );
xor  ( new_n10024_, new_n10023_, new_n9764_ );
or   ( new_n10025_, new_n10024_, new_n10022_ );
and  ( new_n10026_, new_n10024_, new_n10022_ );
xor  ( new_n10027_, new_n9776_, new_n9772_ );
xnor ( new_n10028_, new_n10027_, new_n9782_ );
or   ( new_n10029_, new_n10028_, new_n10026_ );
and  ( new_n10030_, new_n10029_, new_n10025_ );
nor  ( new_n10031_, new_n10030_, new_n10020_ );
nand ( new_n10032_, new_n10030_, new_n10020_ );
xor  ( new_n10033_, new_n9901_, new_n9899_ );
and  ( new_n10034_, new_n10033_, new_n10032_ );
or   ( new_n10035_, new_n10034_, new_n10031_ );
or   ( new_n10036_, new_n8874_, new_n279_ );
or   ( new_n10037_, new_n8876_, new_n285_ );
and  ( new_n10038_, new_n10037_, new_n10036_ );
xor  ( new_n10039_, new_n10038_, new_n8257_ );
or   ( new_n10040_, new_n8264_, new_n294_ );
or   ( new_n10041_, new_n8266_, new_n301_ );
and  ( new_n10042_, new_n10041_, new_n10040_ );
xor  ( new_n10043_, new_n10042_, new_n7725_ );
or   ( new_n10044_, new_n10043_, new_n10039_ );
and  ( new_n10045_, new_n10043_, new_n10039_ );
or   ( new_n10046_, new_n7732_, new_n264_ );
or   ( new_n10047_, new_n7734_, new_n270_ );
and  ( new_n10048_, new_n10047_, new_n10046_ );
xor  ( new_n10049_, new_n10048_, new_n7177_ );
or   ( new_n10050_, new_n10049_, new_n10045_ );
and  ( new_n10051_, new_n10050_, new_n10044_ );
not  ( new_n10052_, RIbb2d900_63 );
or   ( new_n10053_, new_n9422_, new_n313_ );
or   ( new_n10054_, new_n9424_, new_n319_ );
and  ( new_n10055_, new_n10054_, new_n10053_ );
xor  ( new_n10056_, new_n10055_, new_n8873_ );
or   ( new_n10057_, new_n10056_, new_n10052_ );
and  ( new_n10058_, new_n10056_, new_n10052_ );
not  ( new_n10059_, new_n9740_ );
or   ( new_n10060_, new_n10059_, new_n333_ );
not  ( new_n10061_, new_n9738_ );
or   ( new_n10062_, new_n10061_, new_n339_ );
and  ( new_n10063_, new_n10062_, new_n10060_ );
xor  ( new_n10064_, new_n10063_, new_n9421_ );
or   ( new_n10065_, new_n10064_, new_n10058_ );
and  ( new_n10066_, new_n10065_, new_n10057_ );
or   ( new_n10067_, new_n10066_, new_n10051_ );
and  ( new_n10068_, new_n10066_, new_n10051_ );
or   ( new_n10069_, new_n7184_, new_n419_ );
or   ( new_n10070_, new_n7186_, new_n348_ );
and  ( new_n10071_, new_n10070_, new_n10069_ );
xor  ( new_n10072_, new_n10071_, new_n6638_ );
or   ( new_n10073_, new_n6645_, new_n509_ );
or   ( new_n10074_, new_n6647_, new_n443_ );
and  ( new_n10075_, new_n10074_, new_n10073_ );
xor  ( new_n10076_, new_n10075_, new_n6166_ );
nor  ( new_n10077_, new_n10076_, new_n10072_ );
and  ( new_n10078_, new_n10076_, new_n10072_ );
or   ( new_n10079_, new_n6173_, new_n775_ );
or   ( new_n10080_, new_n6175_, new_n515_ );
and  ( new_n10081_, new_n10080_, new_n10079_ );
xor  ( new_n10082_, new_n10081_, new_n5597_ );
nor  ( new_n10083_, new_n10082_, new_n10078_ );
nor  ( new_n10084_, new_n10083_, new_n10077_ );
or   ( new_n10085_, new_n10084_, new_n10068_ );
and  ( new_n10086_, new_n10085_, new_n10067_ );
or   ( new_n10087_, new_n2122_, new_n3696_ );
or   ( new_n10088_, new_n2124_, new_n3306_ );
and  ( new_n10089_, new_n10088_, new_n10087_ );
xor  ( new_n10090_, new_n10089_, new_n1843_ );
or   ( new_n10091_, new_n1844_, new_n3820_ );
or   ( new_n10092_, new_n1846_, new_n3694_ );
and  ( new_n10093_, new_n10092_, new_n10091_ );
xor  ( new_n10094_, new_n10093_, new_n1586_ );
or   ( new_n10095_, new_n10094_, new_n10090_ );
and  ( new_n10096_, new_n10094_, new_n10090_ );
or   ( new_n10097_, new_n1593_, new_n4267_ );
or   ( new_n10098_, new_n1595_, new_n4069_ );
and  ( new_n10099_, new_n10098_, new_n10097_ );
xor  ( new_n10100_, new_n10099_, new_n1358_ );
or   ( new_n10101_, new_n10100_, new_n10096_ );
and  ( new_n10102_, new_n10101_, new_n10095_ );
or   ( new_n10103_, new_n1364_, new_n4995_ );
or   ( new_n10104_, new_n1366_, new_n4603_ );
and  ( new_n10105_, new_n10104_, new_n10103_ );
xor  ( new_n10106_, new_n10105_, new_n1129_ );
or   ( new_n10107_, new_n1135_, new_n5171_ );
or   ( new_n10108_, new_n1137_, new_n4859_ );
and  ( new_n10109_, new_n10108_, new_n10107_ );
xor  ( new_n10110_, new_n10109_, new_n896_ );
or   ( new_n10111_, new_n10110_, new_n10106_ );
and  ( new_n10112_, new_n10110_, new_n10106_ );
or   ( new_n10113_, new_n897_, new_n5570_ );
or   ( new_n10114_, new_n899_, new_n5428_ );
and  ( new_n10115_, new_n10114_, new_n10113_ );
xor  ( new_n10116_, new_n10115_, new_n748_ );
or   ( new_n10117_, new_n10116_, new_n10112_ );
and  ( new_n10118_, new_n10117_, new_n10111_ );
or   ( new_n10119_, new_n10118_, new_n10102_ );
and  ( new_n10120_, new_n10118_, new_n10102_ );
or   ( new_n10121_, new_n755_, new_n6219_ );
or   ( new_n10122_, new_n757_, new_n5899_ );
and  ( new_n10123_, new_n10122_, new_n10121_ );
xor  ( new_n10124_, new_n10123_, new_n523_ );
or   ( new_n10125_, new_n524_, new_n6589_ );
or   ( new_n10126_, new_n526_, new_n6425_ );
and  ( new_n10127_, new_n10126_, new_n10125_ );
xor  ( new_n10128_, new_n10127_, new_n403_ );
nor  ( new_n10129_, new_n10128_, new_n10124_ );
and  ( new_n10130_, new_n10128_, new_n10124_ );
or   ( new_n10131_, new_n409_, new_n7149_ );
or   ( new_n10132_, new_n411_, new_n6943_ );
and  ( new_n10133_, new_n10132_, new_n10131_ );
xor  ( new_n10134_, new_n10133_, new_n328_ );
nor  ( new_n10135_, new_n10134_, new_n10130_ );
nor  ( new_n10136_, new_n10135_, new_n10129_ );
or   ( new_n10137_, new_n10136_, new_n10120_ );
and  ( new_n10138_, new_n10137_, new_n10119_ );
or   ( new_n10139_, new_n10138_, new_n10086_ );
or   ( new_n10140_, new_n3117_, new_n2475_ );
or   ( new_n10141_, new_n3119_, new_n2291_ );
and  ( new_n10142_, new_n10141_, new_n10140_ );
xor  ( new_n10143_, new_n10142_, new_n2800_ );
or   ( new_n10144_, new_n2807_, new_n2751_ );
or   ( new_n10145_, new_n2809_, new_n2646_ );
and  ( new_n10146_, new_n10145_, new_n10144_ );
xor  ( new_n10147_, new_n10146_, new_n2424_ );
or   ( new_n10148_, new_n10147_, new_n10143_ );
and  ( new_n10149_, new_n10147_, new_n10143_ );
or   ( new_n10150_, new_n2425_, new_n3178_ );
or   ( new_n10151_, new_n2427_, new_n2981_ );
and  ( new_n10152_, new_n10151_, new_n10150_ );
xor  ( new_n10153_, new_n10152_, new_n2121_ );
or   ( new_n10154_, new_n10153_, new_n10149_ );
and  ( new_n10155_, new_n10154_, new_n10148_ );
or   ( new_n10156_, new_n4302_, new_n1523_ );
or   ( new_n10157_, new_n4304_, new_n1525_ );
and  ( new_n10158_, new_n10157_, new_n10156_ );
xor  ( new_n10159_, new_n10158_, new_n3895_ );
or   ( new_n10160_, new_n3896_, new_n1899_ );
or   ( new_n10161_, new_n3898_, new_n1754_ );
and  ( new_n10162_, new_n10161_, new_n10160_ );
xor  ( new_n10163_, new_n10162_, new_n3460_ );
or   ( new_n10164_, new_n10163_, new_n10159_ );
and  ( new_n10165_, new_n10163_, new_n10159_ );
or   ( new_n10166_, new_n3461_, new_n2178_ );
or   ( new_n10167_, new_n3463_, new_n2057_ );
and  ( new_n10168_, new_n10167_, new_n10166_ );
xor  ( new_n10169_, new_n10168_, new_n3116_ );
or   ( new_n10170_, new_n10169_, new_n10165_ );
and  ( new_n10171_, new_n10170_, new_n10164_ );
nor  ( new_n10172_, new_n10171_, new_n10155_ );
and  ( new_n10173_, new_n10171_, new_n10155_ );
or   ( new_n10174_, new_n5604_, new_n886_ );
or   ( new_n10175_, new_n5606_, new_n805_ );
and  ( new_n10176_, new_n10175_, new_n10174_ );
xor  ( new_n10177_, new_n10176_, new_n5206_ );
or   ( new_n10178_, new_n5207_, new_n1168_ );
or   ( new_n10179_, new_n5209_, new_n986_ );
and  ( new_n10180_, new_n10179_, new_n10178_ );
xor  ( new_n10181_, new_n10180_, new_n4708_ );
nor  ( new_n10182_, new_n10181_, new_n10177_ );
and  ( new_n10183_, new_n10181_, new_n10177_ );
or   ( new_n10184_, new_n4709_, new_n1318_ );
or   ( new_n10185_, new_n4711_, new_n1213_ );
and  ( new_n10186_, new_n10185_, new_n10184_ );
xor  ( new_n10187_, new_n10186_, new_n4295_ );
nor  ( new_n10188_, new_n10187_, new_n10183_ );
nor  ( new_n10189_, new_n10188_, new_n10182_ );
nor  ( new_n10190_, new_n10189_, new_n10173_ );
nor  ( new_n10191_, new_n10190_, new_n10172_ );
and  ( new_n10192_, new_n10138_, new_n10086_ );
or   ( new_n10193_, new_n10192_, new_n10191_ );
and  ( new_n10194_, new_n10193_, new_n10139_ );
and  ( new_n10195_, new_n10194_, new_n10035_ );
nor  ( new_n10196_, new_n10194_, new_n10035_ );
xnor ( new_n10197_, new_n9685_, new_n9684_ );
or   ( new_n10198_, new_n337_, new_n8117_ );
or   ( new_n10199_, new_n340_, new_n7373_ );
and  ( new_n10200_, new_n10199_, new_n10198_ );
xor  ( new_n10201_, new_n10200_, new_n332_ );
or   ( new_n10202_, new_n317_, new_n8352_ );
or   ( new_n10203_, new_n320_, new_n8115_ );
and  ( new_n10204_, new_n10203_, new_n10202_ );
xor  ( new_n10205_, new_n10204_, new_n312_ );
or   ( new_n10206_, new_n10205_, new_n10201_ );
and  ( new_n10207_, new_n10205_, new_n10201_ );
or   ( new_n10208_, new_n283_, new_n8995_ );
or   ( new_n10209_, new_n286_, new_n8481_ );
and  ( new_n10210_, new_n10209_, new_n10208_ );
xor  ( new_n10211_, new_n10210_, new_n278_ );
or   ( new_n10212_, new_n10211_, new_n10207_ );
and  ( new_n10213_, new_n10212_, new_n10206_ );
nor  ( new_n10214_, new_n10213_, new_n10197_ );
and  ( new_n10215_, new_n10213_, new_n10197_ );
or   ( new_n10216_, new_n299_, new_n9681_ );
or   ( new_n10217_, new_n302_, new_n9099_ );
and  ( new_n10218_, new_n10217_, new_n10216_ );
xor  ( new_n10219_, new_n10218_, new_n293_ );
not  ( new_n10220_, RIbb2bb78_126 );
or   ( new_n10221_, new_n268_, new_n10220_ );
or   ( new_n10222_, new_n271_, new_n9679_ );
and  ( new_n10223_, new_n10222_, new_n10221_ );
xor  ( new_n10224_, new_n10223_, new_n263_ );
nor  ( new_n10225_, new_n10224_, new_n10219_ );
and  ( new_n10226_, RIbb31500_127, RIbb2f610_1 );
and  ( new_n10227_, new_n10224_, new_n10219_ );
nor  ( new_n10228_, new_n10227_, new_n10226_ );
nor  ( new_n10229_, new_n10228_, new_n10225_ );
nor  ( new_n10230_, new_n10229_, new_n10215_ );
or   ( new_n10231_, new_n10230_, new_n10214_ );
xnor ( new_n10232_, new_n9847_, new_n9843_ );
xor  ( new_n10233_, new_n10232_, new_n9853_ );
xnor ( new_n10234_, new_n9881_, new_n9877_ );
xor  ( new_n10235_, new_n10234_, new_n9887_ );
or   ( new_n10236_, new_n10235_, new_n10233_ );
and  ( new_n10237_, new_n10235_, new_n10233_ );
xor  ( new_n10238_, new_n9794_, new_n9790_ );
xnor ( new_n10239_, new_n10238_, new_n9800_ );
or   ( new_n10240_, new_n10239_, new_n10237_ );
and  ( new_n10241_, new_n10240_, new_n10236_ );
nor  ( new_n10242_, new_n10241_, new_n10231_ );
and  ( new_n10243_, new_n10241_, new_n10231_ );
xnor ( new_n10244_, new_n9810_, new_n9806_ );
xor  ( new_n10245_, new_n10244_, new_n9816_ );
xnor ( new_n10246_, new_n9694_, new_n9690_ );
xor  ( new_n10247_, new_n10246_, new_n9700_ );
nor  ( new_n10248_, new_n10247_, new_n10245_ );
and  ( new_n10249_, new_n10247_, new_n10245_ );
xor  ( new_n10250_, new_n9828_, new_n9824_ );
xnor ( new_n10251_, new_n10250_, new_n9834_ );
nor  ( new_n10252_, new_n10251_, new_n10249_ );
nor  ( new_n10253_, new_n10252_, new_n10248_ );
nor  ( new_n10254_, new_n10253_, new_n10243_ );
nor  ( new_n10255_, new_n10254_, new_n10242_ );
nor  ( new_n10256_, new_n10255_, new_n10196_ );
nor  ( new_n10257_, new_n10256_, new_n10195_ );
or   ( new_n10258_, new_n10257_, new_n10018_ );
and  ( new_n10259_, new_n10258_, new_n10017_ );
or   ( new_n10260_, new_n10259_, new_n9979_ );
and  ( new_n10261_, new_n10260_, new_n9978_ );
xor  ( new_n10262_, new_n9575_, new_n9528_ );
xor  ( new_n10263_, new_n10262_, new_n9596_ );
xor  ( new_n10264_, new_n9921_, new_n9678_ );
xor  ( new_n10265_, new_n10264_, new_n9933_ );
or   ( new_n10266_, new_n10265_, new_n10263_ );
and  ( new_n10267_, new_n10265_, new_n10263_ );
xor  ( new_n10268_, new_n9941_, new_n9939_ );
xnor ( new_n10269_, new_n10268_, new_n9945_ );
not  ( new_n10270_, new_n10269_ );
or   ( new_n10271_, new_n10270_, new_n10267_ );
and  ( new_n10272_, new_n10271_, new_n10266_ );
nor  ( new_n10273_, new_n10272_, new_n10261_ );
and  ( new_n10274_, new_n10272_, new_n10261_ );
xor  ( new_n10275_, new_n9598_, new_n9365_ );
xor  ( new_n10276_, new_n10275_, new_n9611_ );
nor  ( new_n10277_, new_n10276_, new_n10274_ );
nor  ( new_n10278_, new_n10277_, new_n10273_ );
xnor ( new_n10279_, new_n9951_, new_n9949_ );
xnor ( new_n10280_, new_n10279_, new_n9955_ );
nor  ( new_n10281_, new_n10280_, new_n10278_ );
xnor ( new_n10282_, new_n9957_, new_n9650_ );
xor  ( new_n10283_, new_n10282_, new_n9961_ );
and  ( new_n10284_, new_n10283_, new_n10281_ );
xnor ( new_n10285_, new_n10280_, new_n10278_ );
xor  ( new_n10286_, new_n10272_, new_n10261_ );
xor  ( new_n10287_, new_n10286_, new_n10276_ );
xor  ( new_n10288_, new_n9894_, new_n9733_ );
xor  ( new_n10289_, new_n10288_, new_n9919_ );
xor  ( new_n10290_, new_n9838_, new_n9786_ );
xor  ( new_n10291_, new_n10290_, new_n9891_ );
xnor ( new_n10292_, new_n9991_, new_n9989_ );
xor  ( new_n10293_, new_n10292_, new_n10003_ );
nand ( new_n10294_, new_n10293_, new_n10291_ );
nor  ( new_n10295_, new_n10293_, new_n10291_ );
xor  ( new_n10296_, new_n10009_, new_n10007_ );
xor  ( new_n10297_, new_n10296_, new_n10014_ );
or   ( new_n10298_, new_n10297_, new_n10295_ );
and  ( new_n10299_, new_n10298_, new_n10294_ );
or   ( new_n10300_, new_n10299_, new_n10289_ );
and  ( new_n10301_, new_n10299_, new_n10289_ );
xor  ( new_n10302_, new_n9983_, new_n9981_ );
xor  ( new_n10303_, new_n10302_, new_n9987_ );
xnor ( new_n10304_, new_n10241_, new_n10231_ );
xor  ( new_n10305_, new_n10304_, new_n10253_ );
or   ( new_n10306_, new_n10305_, new_n10303_ );
and  ( new_n10307_, new_n10305_, new_n10303_ );
xor  ( new_n10308_, new_n10030_, new_n10020_ );
xor  ( new_n10309_, new_n10308_, new_n10033_ );
or   ( new_n10310_, new_n10309_, new_n10307_ );
and  ( new_n10311_, new_n10310_, new_n10306_ );
xnor ( new_n10312_, new_n10024_, new_n10022_ );
xor  ( new_n10313_, new_n10312_, new_n10028_ );
xnor ( new_n10314_, new_n10235_, new_n10233_ );
xor  ( new_n10315_, new_n10314_, new_n10239_ );
or   ( new_n10316_, new_n10315_, new_n10313_ );
and  ( new_n10317_, new_n10315_, new_n10313_ );
xor  ( new_n10318_, new_n10247_, new_n10245_ );
xnor ( new_n10319_, new_n10318_, new_n10251_ );
or   ( new_n10320_, new_n10319_, new_n10317_ );
and  ( new_n10321_, new_n10320_, new_n10316_ );
xnor ( new_n10322_, new_n9997_, new_n9995_ );
xor  ( new_n10323_, new_n10322_, new_n10001_ );
or   ( new_n10324_, new_n10323_, new_n10321_ );
nand ( new_n10325_, new_n10323_, new_n10321_ );
xnor ( new_n10326_, new_n10118_, new_n10102_ );
xor  ( new_n10327_, new_n10326_, new_n10136_ );
xnor ( new_n10328_, new_n10171_, new_n10155_ );
xor  ( new_n10329_, new_n10328_, new_n10189_ );
nor  ( new_n10330_, new_n10329_, new_n10327_ );
and  ( new_n10331_, new_n10329_, new_n10327_ );
xor  ( new_n10332_, new_n10213_, new_n10197_ );
xor  ( new_n10333_, new_n10332_, new_n10229_ );
not  ( new_n10334_, new_n10333_ );
nor  ( new_n10335_, new_n10334_, new_n10331_ );
nor  ( new_n10336_, new_n10335_, new_n10330_ );
nand ( new_n10337_, new_n10336_, new_n10325_ );
and  ( new_n10338_, new_n10337_, new_n10324_ );
and  ( new_n10339_, new_n10338_, new_n10311_ );
nor  ( new_n10340_, new_n10338_, new_n10311_ );
xor  ( new_n10341_, new_n10043_, new_n10039_ );
xnor ( new_n10342_, new_n10341_, new_n10049_ );
xor  ( new_n10343_, new_n10056_, RIbb2d900_63 );
xor  ( new_n10344_, new_n10343_, new_n10064_ );
or   ( new_n10345_, new_n10344_, new_n10342_ );
xnor ( new_n10346_, new_n10163_, new_n10159_ );
xor  ( new_n10347_, new_n10346_, new_n10169_ );
xnor ( new_n10348_, new_n10076_, new_n10072_ );
xor  ( new_n10349_, new_n10348_, new_n10082_ );
or   ( new_n10350_, new_n10349_, new_n10347_ );
and  ( new_n10351_, new_n10349_, new_n10347_ );
xnor ( new_n10352_, new_n10181_, new_n10177_ );
xor  ( new_n10353_, new_n10352_, new_n10187_ );
or   ( new_n10354_, new_n10353_, new_n10351_ );
and  ( new_n10355_, new_n10354_, new_n10350_ );
nor  ( new_n10356_, new_n10355_, new_n10345_ );
and  ( new_n10357_, new_n10355_, new_n10345_ );
xor  ( new_n10358_, new_n9742_, new_n9737_ );
xnor ( new_n10359_, new_n10358_, new_n9748_ );
nor  ( new_n10360_, new_n10359_, new_n10357_ );
or   ( new_n10361_, new_n10360_, new_n10356_ );
or   ( new_n10362_, new_n897_, new_n5899_ );
or   ( new_n10363_, new_n899_, new_n5570_ );
and  ( new_n10364_, new_n10363_, new_n10362_ );
xor  ( new_n10365_, new_n10364_, new_n748_ );
or   ( new_n10366_, new_n755_, new_n6425_ );
or   ( new_n10367_, new_n757_, new_n6219_ );
and  ( new_n10368_, new_n10367_, new_n10366_ );
xor  ( new_n10369_, new_n10368_, new_n523_ );
or   ( new_n10370_, new_n10369_, new_n10365_ );
and  ( new_n10371_, new_n10369_, new_n10365_ );
or   ( new_n10372_, new_n524_, new_n6943_ );
or   ( new_n10373_, new_n526_, new_n6589_ );
and  ( new_n10374_, new_n10373_, new_n10372_ );
xor  ( new_n10375_, new_n10374_, new_n403_ );
or   ( new_n10376_, new_n10375_, new_n10371_ );
and  ( new_n10377_, new_n10376_, new_n10370_ );
or   ( new_n10378_, new_n1593_, new_n4603_ );
or   ( new_n10379_, new_n1595_, new_n4267_ );
and  ( new_n10380_, new_n10379_, new_n10378_ );
xor  ( new_n10381_, new_n10380_, new_n1358_ );
or   ( new_n10382_, new_n1364_, new_n4859_ );
or   ( new_n10383_, new_n1366_, new_n4995_ );
and  ( new_n10384_, new_n10383_, new_n10382_ );
xor  ( new_n10385_, new_n10384_, new_n1129_ );
or   ( new_n10386_, new_n10385_, new_n10381_ );
and  ( new_n10387_, new_n10385_, new_n10381_ );
or   ( new_n10388_, new_n1135_, new_n5428_ );
or   ( new_n10389_, new_n1137_, new_n5171_ );
and  ( new_n10390_, new_n10389_, new_n10388_ );
xor  ( new_n10391_, new_n10390_, new_n896_ );
or   ( new_n10392_, new_n10391_, new_n10387_ );
and  ( new_n10393_, new_n10392_, new_n10386_ );
or   ( new_n10394_, new_n10393_, new_n10377_ );
and  ( new_n10395_, new_n10393_, new_n10377_ );
or   ( new_n10396_, new_n2425_, new_n3306_ );
or   ( new_n10397_, new_n2427_, new_n3178_ );
and  ( new_n10398_, new_n10397_, new_n10396_ );
xor  ( new_n10399_, new_n10398_, new_n2121_ );
or   ( new_n10400_, new_n2122_, new_n3694_ );
or   ( new_n10401_, new_n2124_, new_n3696_ );
and  ( new_n10402_, new_n10401_, new_n10400_ );
xor  ( new_n10403_, new_n10402_, new_n1843_ );
nor  ( new_n10404_, new_n10403_, new_n10399_ );
and  ( new_n10405_, new_n10403_, new_n10399_ );
or   ( new_n10406_, new_n1844_, new_n4069_ );
or   ( new_n10407_, new_n1846_, new_n3820_ );
and  ( new_n10408_, new_n10407_, new_n10406_ );
xor  ( new_n10409_, new_n10408_, new_n1586_ );
nor  ( new_n10410_, new_n10409_, new_n10405_ );
nor  ( new_n10411_, new_n10410_, new_n10404_ );
or   ( new_n10412_, new_n10411_, new_n10395_ );
and  ( new_n10413_, new_n10412_, new_n10394_ );
or   ( new_n10414_, new_n3461_, new_n2291_ );
or   ( new_n10415_, new_n3463_, new_n2178_ );
and  ( new_n10416_, new_n10415_, new_n10414_ );
xor  ( new_n10417_, new_n10416_, new_n3116_ );
or   ( new_n10418_, new_n3117_, new_n2646_ );
or   ( new_n10419_, new_n3119_, new_n2475_ );
and  ( new_n10420_, new_n10419_, new_n10418_ );
xor  ( new_n10421_, new_n10420_, new_n2800_ );
or   ( new_n10422_, new_n10421_, new_n10417_ );
and  ( new_n10423_, new_n10421_, new_n10417_ );
or   ( new_n10424_, new_n2807_, new_n2981_ );
or   ( new_n10425_, new_n2809_, new_n2751_ );
and  ( new_n10426_, new_n10425_, new_n10424_ );
xor  ( new_n10427_, new_n10426_, new_n2424_ );
or   ( new_n10428_, new_n10427_, new_n10423_ );
and  ( new_n10429_, new_n10428_, new_n10422_ );
or   ( new_n10430_, new_n4709_, new_n1525_ );
or   ( new_n10431_, new_n4711_, new_n1318_ );
and  ( new_n10432_, new_n10431_, new_n10430_ );
xor  ( new_n10433_, new_n10432_, new_n4295_ );
or   ( new_n10434_, new_n4302_, new_n1754_ );
or   ( new_n10435_, new_n4304_, new_n1523_ );
and  ( new_n10436_, new_n10435_, new_n10434_ );
xor  ( new_n10437_, new_n10436_, new_n3895_ );
or   ( new_n10438_, new_n10437_, new_n10433_ );
and  ( new_n10439_, new_n10437_, new_n10433_ );
or   ( new_n10440_, new_n3896_, new_n2057_ );
or   ( new_n10441_, new_n3898_, new_n1899_ );
and  ( new_n10442_, new_n10441_, new_n10440_ );
xor  ( new_n10443_, new_n10442_, new_n3460_ );
or   ( new_n10444_, new_n10443_, new_n10439_ );
and  ( new_n10445_, new_n10444_, new_n10438_ );
or   ( new_n10446_, new_n10445_, new_n10429_ );
and  ( new_n10447_, new_n10445_, new_n10429_ );
or   ( new_n10448_, new_n6173_, new_n805_ );
or   ( new_n10449_, new_n6175_, new_n775_ );
and  ( new_n10450_, new_n10449_, new_n10448_ );
xor  ( new_n10451_, new_n10450_, new_n5597_ );
or   ( new_n10452_, new_n5604_, new_n986_ );
or   ( new_n10453_, new_n5606_, new_n886_ );
and  ( new_n10454_, new_n10453_, new_n10452_ );
xor  ( new_n10455_, new_n10454_, new_n5206_ );
nor  ( new_n10456_, new_n10455_, new_n10451_ );
and  ( new_n10457_, new_n10455_, new_n10451_ );
or   ( new_n10458_, new_n5207_, new_n1213_ );
or   ( new_n10459_, new_n5209_, new_n1168_ );
and  ( new_n10460_, new_n10459_, new_n10458_ );
xor  ( new_n10461_, new_n10460_, new_n4708_ );
nor  ( new_n10462_, new_n10461_, new_n10457_ );
nor  ( new_n10463_, new_n10462_, new_n10456_ );
or   ( new_n10464_, new_n10463_, new_n10447_ );
and  ( new_n10465_, new_n10464_, new_n10446_ );
or   ( new_n10466_, new_n10465_, new_n10413_ );
and  ( new_n10467_, new_n10465_, new_n10413_ );
or   ( new_n10468_, new_n9422_, new_n285_ );
or   ( new_n10469_, new_n9424_, new_n313_ );
and  ( new_n10470_, new_n10469_, new_n10468_ );
xor  ( new_n10471_, new_n10470_, new_n8873_ );
or   ( new_n10472_, new_n8874_, new_n301_ );
or   ( new_n10473_, new_n8876_, new_n279_ );
and  ( new_n10474_, new_n10473_, new_n10472_ );
xor  ( new_n10475_, new_n10474_, new_n8257_ );
nor  ( new_n10476_, new_n10475_, new_n10471_ );
and  ( new_n10477_, new_n10475_, new_n10471_ );
or   ( new_n10478_, new_n8264_, new_n270_ );
or   ( new_n10479_, new_n8266_, new_n294_ );
and  ( new_n10480_, new_n10479_, new_n10478_ );
xor  ( new_n10481_, new_n10480_, new_n7725_ );
nor  ( new_n10482_, new_n10481_, new_n10477_ );
nor  ( new_n10483_, new_n10482_, new_n10476_ );
or   ( new_n10484_, new_n10059_, new_n319_ );
or   ( new_n10485_, new_n10061_, new_n333_ );
and  ( new_n10486_, new_n10485_, new_n10484_ );
xor  ( new_n10487_, new_n10486_, new_n9421_ );
or   ( new_n10488_, RIbb2d888_64, new_n339_ );
and  ( new_n10489_, new_n10488_, RIbb2d900_63 );
and  ( new_n10490_, new_n10489_, new_n10487_ );
or   ( new_n10491_, new_n7732_, new_n348_ );
or   ( new_n10492_, new_n7734_, new_n264_ );
and  ( new_n10493_, new_n10492_, new_n10491_ );
xor  ( new_n10494_, new_n10493_, new_n7177_ );
or   ( new_n10495_, new_n7184_, new_n443_ );
or   ( new_n10496_, new_n7186_, new_n419_ );
and  ( new_n10497_, new_n10496_, new_n10495_ );
xor  ( new_n10498_, new_n10497_, new_n6638_ );
nor  ( new_n10499_, new_n10498_, new_n10494_ );
and  ( new_n10500_, new_n10498_, new_n10494_ );
or   ( new_n10501_, new_n6645_, new_n515_ );
or   ( new_n10502_, new_n6647_, new_n509_ );
and  ( new_n10503_, new_n10502_, new_n10501_ );
xor  ( new_n10504_, new_n10503_, new_n6166_ );
nor  ( new_n10505_, new_n10504_, new_n10500_ );
nor  ( new_n10506_, new_n10505_, new_n10499_ );
and  ( new_n10507_, new_n10506_, new_n10490_ );
nor  ( new_n10508_, new_n10507_, new_n10483_ );
nor  ( new_n10509_, new_n10506_, new_n10490_ );
nor  ( new_n10510_, new_n10509_, new_n10508_ );
or   ( new_n10511_, new_n10510_, new_n10467_ );
and  ( new_n10512_, new_n10511_, new_n10466_ );
and  ( new_n10513_, new_n10512_, new_n10361_ );
nor  ( new_n10514_, new_n10512_, new_n10361_ );
or   ( new_n10515_, new_n409_, new_n7373_ );
or   ( new_n10516_, new_n411_, new_n7149_ );
and  ( new_n10517_, new_n10516_, new_n10515_ );
xor  ( new_n10518_, new_n10517_, new_n328_ );
or   ( new_n10519_, new_n337_, new_n8115_ );
or   ( new_n10520_, new_n340_, new_n8117_ );
and  ( new_n10521_, new_n10520_, new_n10519_ );
xor  ( new_n10522_, new_n10521_, new_n332_ );
or   ( new_n10523_, new_n10522_, new_n10518_ );
and  ( new_n10524_, new_n10522_, new_n10518_ );
or   ( new_n10525_, new_n317_, new_n8481_ );
or   ( new_n10526_, new_n320_, new_n8352_ );
and  ( new_n10527_, new_n10526_, new_n10525_ );
xor  ( new_n10528_, new_n10527_, new_n312_ );
or   ( new_n10529_, new_n10528_, new_n10524_ );
and  ( new_n10530_, new_n10529_, new_n10523_ );
or   ( new_n10531_, new_n283_, new_n9099_ );
or   ( new_n10532_, new_n286_, new_n8995_ );
and  ( new_n10533_, new_n10532_, new_n10531_ );
xor  ( new_n10534_, new_n10533_, new_n278_ );
or   ( new_n10535_, new_n299_, new_n9679_ );
or   ( new_n10536_, new_n302_, new_n9681_ );
and  ( new_n10537_, new_n10536_, new_n10535_ );
xor  ( new_n10538_, new_n10537_, new_n293_ );
or   ( new_n10539_, new_n10538_, new_n10534_ );
and  ( new_n10540_, new_n10538_, new_n10534_ );
not  ( new_n10541_, RIbb31500_127 );
or   ( new_n10542_, new_n268_, new_n10541_ );
or   ( new_n10543_, new_n271_, new_n10220_ );
and  ( new_n10544_, new_n10543_, new_n10542_ );
xor  ( new_n10545_, new_n10544_, new_n263_ );
or   ( new_n10546_, new_n10545_, new_n10540_ );
and  ( new_n10547_, new_n10546_, new_n10539_ );
nor  ( new_n10548_, new_n10547_, new_n10530_ );
xnor ( new_n10549_, new_n10205_, new_n10201_ );
xor  ( new_n10550_, new_n10549_, new_n10211_ );
xnor ( new_n10551_, new_n10224_, new_n10219_ );
xor  ( new_n10552_, new_n10551_, new_n10226_ );
or   ( new_n10553_, new_n10552_, new_n10550_ );
and  ( new_n10554_, new_n10552_, new_n10550_ );
xor  ( new_n10555_, new_n10128_, new_n10124_ );
xnor ( new_n10556_, new_n10555_, new_n10134_ );
or   ( new_n10557_, new_n10556_, new_n10554_ );
and  ( new_n10558_, new_n10557_, new_n10553_ );
nor  ( new_n10559_, new_n10558_, new_n10548_ );
and  ( new_n10560_, new_n10558_, new_n10548_ );
xnor ( new_n10561_, new_n10110_, new_n10106_ );
xor  ( new_n10562_, new_n10561_, new_n10116_ );
xnor ( new_n10563_, new_n10094_, new_n10090_ );
xor  ( new_n10564_, new_n10563_, new_n10100_ );
nor  ( new_n10565_, new_n10564_, new_n10562_ );
and  ( new_n10566_, new_n10564_, new_n10562_ );
xor  ( new_n10567_, new_n10147_, new_n10143_ );
xnor ( new_n10568_, new_n10567_, new_n10153_ );
nor  ( new_n10569_, new_n10568_, new_n10566_ );
nor  ( new_n10570_, new_n10569_, new_n10565_ );
nor  ( new_n10571_, new_n10570_, new_n10560_ );
nor  ( new_n10572_, new_n10571_, new_n10559_ );
nor  ( new_n10573_, new_n10572_, new_n10514_ );
nor  ( new_n10574_, new_n10573_, new_n10513_ );
nor  ( new_n10575_, new_n10574_, new_n10340_ );
nor  ( new_n10576_, new_n10575_, new_n10339_ );
or   ( new_n10577_, new_n10576_, new_n10301_ );
and  ( new_n10578_, new_n10577_, new_n10300_ );
xor  ( new_n10579_, new_n9977_, new_n9966_ );
xor  ( new_n10580_, new_n10579_, new_n10259_ );
or   ( new_n10581_, new_n10580_, new_n10578_ );
and  ( new_n10582_, new_n10580_, new_n10578_ );
xor  ( new_n10583_, new_n10265_, new_n10263_ );
xor  ( new_n10584_, new_n10583_, new_n10270_ );
or   ( new_n10585_, new_n10584_, new_n10582_ );
and  ( new_n10586_, new_n10585_, new_n10581_ );
or   ( new_n10587_, new_n10586_, new_n10287_ );
and  ( new_n10588_, new_n10586_, new_n10287_ );
xor  ( new_n10589_, new_n9935_, new_n9652_ );
xor  ( new_n10590_, new_n10589_, new_n9947_ );
or   ( new_n10591_, new_n10590_, new_n10588_ );
and  ( new_n10592_, new_n10591_, new_n10587_ );
nor  ( new_n10593_, new_n10592_, new_n10285_ );
xor  ( new_n10594_, new_n10586_, new_n10287_ );
xor  ( new_n10595_, new_n10594_, new_n10590_ );
xor  ( new_n10596_, new_n10016_, new_n10005_ );
xnor ( new_n10597_, new_n10596_, new_n10257_ );
xnor ( new_n10598_, new_n10299_, new_n10289_ );
xor  ( new_n10599_, new_n10598_, new_n10576_ );
nand ( new_n10600_, new_n10599_, new_n10597_ );
xor  ( new_n10601_, new_n10338_, new_n10311_ );
xnor ( new_n10602_, new_n10601_, new_n10574_ );
xnor ( new_n10603_, new_n10293_, new_n10291_ );
xor  ( new_n10604_, new_n10603_, new_n10297_ );
and  ( new_n10605_, new_n10604_, new_n10602_ );
xor  ( new_n10606_, new_n10194_, new_n10035_ );
xor  ( new_n10607_, new_n10606_, new_n10255_ );
xnor ( new_n10608_, new_n10138_, new_n10086_ );
xor  ( new_n10609_, new_n10608_, new_n10191_ );
xor  ( new_n10610_, new_n10323_, new_n10321_ );
xor  ( new_n10611_, new_n10610_, new_n10336_ );
or   ( new_n10612_, new_n10611_, new_n10609_ );
and  ( new_n10613_, new_n10611_, new_n10609_ );
xnor ( new_n10614_, new_n10305_, new_n10303_ );
xor  ( new_n10615_, new_n10614_, new_n10309_ );
or   ( new_n10616_, new_n10615_, new_n10613_ );
and  ( new_n10617_, new_n10616_, new_n10612_ );
nand ( new_n10618_, new_n10617_, new_n10607_ );
or   ( new_n10619_, new_n10617_, new_n10607_ );
xnor ( new_n10620_, new_n10564_, new_n10562_ );
xor  ( new_n10621_, new_n10620_, new_n10568_ );
xnor ( new_n10622_, new_n10552_, new_n10550_ );
xor  ( new_n10623_, new_n10622_, new_n10556_ );
nor  ( new_n10624_, new_n10623_, new_n10621_ );
nand ( new_n10625_, new_n10623_, new_n10621_ );
xor  ( new_n10626_, new_n10547_, new_n10530_ );
and  ( new_n10627_, new_n10626_, new_n10625_ );
or   ( new_n10628_, new_n10627_, new_n10624_ );
xnor ( new_n10629_, new_n10066_, new_n10051_ );
xor  ( new_n10630_, new_n10629_, new_n10084_ );
or   ( new_n10631_, new_n10630_, new_n10628_ );
and  ( new_n10632_, new_n10630_, new_n10628_ );
xnor ( new_n10633_, new_n10393_, new_n10377_ );
xor  ( new_n10634_, new_n10633_, new_n10411_ );
xnor ( new_n10635_, new_n10445_, new_n10429_ );
xor  ( new_n10636_, new_n10635_, new_n10463_ );
nor  ( new_n10637_, new_n10636_, new_n10634_ );
and  ( new_n10638_, new_n10636_, new_n10634_ );
xnor ( new_n10639_, new_n10506_, new_n10490_ );
xnor ( new_n10640_, new_n10639_, new_n10483_ );
not  ( new_n10641_, new_n10640_ );
nor  ( new_n10642_, new_n10641_, new_n10638_ );
nor  ( new_n10643_, new_n10642_, new_n10637_ );
or   ( new_n10644_, new_n10643_, new_n10632_ );
and  ( new_n10645_, new_n10644_, new_n10631_ );
xor  ( new_n10646_, new_n10355_, new_n10345_ );
xor  ( new_n10647_, new_n10646_, new_n10359_ );
xnor ( new_n10648_, new_n10315_, new_n10313_ );
xor  ( new_n10649_, new_n10648_, new_n10319_ );
or   ( new_n10650_, new_n10649_, new_n10647_ );
and  ( new_n10651_, new_n10649_, new_n10647_ );
xor  ( new_n10652_, new_n10329_, new_n10327_ );
xor  ( new_n10653_, new_n10652_, new_n10334_ );
or   ( new_n10654_, new_n10653_, new_n10651_ );
and  ( new_n10655_, new_n10654_, new_n10650_ );
nor  ( new_n10656_, new_n10655_, new_n10645_ );
and  ( new_n10657_, new_n10655_, new_n10645_ );
xor  ( new_n10658_, new_n10349_, new_n10347_ );
xor  ( new_n10659_, new_n10658_, new_n10353_ );
xnor ( new_n10660_, new_n10475_, new_n10471_ );
xor  ( new_n10661_, new_n10660_, new_n10481_ );
xnor ( new_n10662_, new_n10498_, new_n10494_ );
xor  ( new_n10663_, new_n10662_, new_n10504_ );
or   ( new_n10664_, new_n10663_, new_n10661_ );
and  ( new_n10665_, new_n10663_, new_n10661_ );
xor  ( new_n10666_, new_n10455_, new_n10451_ );
xnor ( new_n10667_, new_n10666_, new_n10461_ );
or   ( new_n10668_, new_n10667_, new_n10665_ );
and  ( new_n10669_, new_n10668_, new_n10664_ );
nor  ( new_n10670_, new_n10669_, new_n10659_ );
nand ( new_n10671_, new_n10669_, new_n10659_ );
xor  ( new_n10672_, new_n10344_, new_n10342_ );
and  ( new_n10673_, new_n10672_, new_n10671_ );
or   ( new_n10674_, new_n10673_, new_n10670_ );
or   ( new_n10675_, new_n5604_, new_n1168_ );
or   ( new_n10676_, new_n5606_, new_n986_ );
and  ( new_n10677_, new_n10676_, new_n10675_ );
xor  ( new_n10678_, new_n10677_, new_n5206_ );
or   ( new_n10679_, new_n5207_, new_n1318_ );
or   ( new_n10680_, new_n5209_, new_n1213_ );
and  ( new_n10681_, new_n10680_, new_n10679_ );
xor  ( new_n10682_, new_n10681_, new_n4708_ );
or   ( new_n10683_, new_n10682_, new_n10678_ );
and  ( new_n10684_, new_n10682_, new_n10678_ );
or   ( new_n10685_, new_n4709_, new_n1523_ );
or   ( new_n10686_, new_n4711_, new_n1525_ );
and  ( new_n10687_, new_n10686_, new_n10685_ );
xor  ( new_n10688_, new_n10687_, new_n4295_ );
or   ( new_n10689_, new_n10688_, new_n10684_ );
and  ( new_n10690_, new_n10689_, new_n10683_ );
or   ( new_n10691_, new_n4302_, new_n1899_ );
or   ( new_n10692_, new_n4304_, new_n1754_ );
and  ( new_n10693_, new_n10692_, new_n10691_ );
xor  ( new_n10694_, new_n10693_, new_n3895_ );
or   ( new_n10695_, new_n3896_, new_n2178_ );
or   ( new_n10696_, new_n3898_, new_n2057_ );
and  ( new_n10697_, new_n10696_, new_n10695_ );
xor  ( new_n10698_, new_n10697_, new_n3460_ );
or   ( new_n10699_, new_n10698_, new_n10694_ );
and  ( new_n10700_, new_n10698_, new_n10694_ );
or   ( new_n10701_, new_n3461_, new_n2475_ );
or   ( new_n10702_, new_n3463_, new_n2291_ );
and  ( new_n10703_, new_n10702_, new_n10701_ );
xor  ( new_n10704_, new_n10703_, new_n3116_ );
or   ( new_n10705_, new_n10704_, new_n10700_ );
and  ( new_n10706_, new_n10705_, new_n10699_ );
or   ( new_n10707_, new_n10706_, new_n10690_ );
and  ( new_n10708_, new_n10706_, new_n10690_ );
or   ( new_n10709_, new_n3117_, new_n2751_ );
or   ( new_n10710_, new_n3119_, new_n2646_ );
and  ( new_n10711_, new_n10710_, new_n10709_ );
xor  ( new_n10712_, new_n10711_, new_n2800_ );
or   ( new_n10713_, new_n2807_, new_n3178_ );
or   ( new_n10714_, new_n2809_, new_n2981_ );
and  ( new_n10715_, new_n10714_, new_n10713_ );
xor  ( new_n10716_, new_n10715_, new_n2424_ );
nor  ( new_n10717_, new_n10716_, new_n10712_ );
and  ( new_n10718_, new_n10716_, new_n10712_ );
or   ( new_n10719_, new_n2425_, new_n3696_ );
or   ( new_n10720_, new_n2427_, new_n3306_ );
and  ( new_n10721_, new_n10720_, new_n10719_ );
xor  ( new_n10722_, new_n10721_, new_n2121_ );
nor  ( new_n10723_, new_n10722_, new_n10718_ );
nor  ( new_n10724_, new_n10723_, new_n10717_ );
or   ( new_n10725_, new_n10724_, new_n10708_ );
and  ( new_n10726_, new_n10725_, new_n10707_ );
or   ( new_n10727_, new_n8874_, new_n294_ );
or   ( new_n10728_, new_n8876_, new_n301_ );
and  ( new_n10729_, new_n10728_, new_n10727_ );
xor  ( new_n10730_, new_n10729_, new_n8257_ );
or   ( new_n10731_, new_n8264_, new_n264_ );
or   ( new_n10732_, new_n8266_, new_n270_ );
and  ( new_n10733_, new_n10732_, new_n10731_ );
xor  ( new_n10734_, new_n10733_, new_n7725_ );
or   ( new_n10735_, new_n10734_, new_n10730_ );
and  ( new_n10736_, new_n10734_, new_n10730_ );
or   ( new_n10737_, new_n7732_, new_n419_ );
or   ( new_n10738_, new_n7734_, new_n348_ );
and  ( new_n10739_, new_n10738_, new_n10737_ );
xor  ( new_n10740_, new_n10739_, new_n7177_ );
or   ( new_n10741_, new_n10740_, new_n10736_ );
and  ( new_n10742_, new_n10741_, new_n10735_ );
or   ( new_n10743_, new_n7184_, new_n509_ );
or   ( new_n10744_, new_n7186_, new_n443_ );
and  ( new_n10745_, new_n10744_, new_n10743_ );
xor  ( new_n10746_, new_n10745_, new_n6638_ );
or   ( new_n10747_, new_n6645_, new_n775_ );
or   ( new_n10748_, new_n6647_, new_n515_ );
and  ( new_n10749_, new_n10748_, new_n10747_ );
xor  ( new_n10750_, new_n10749_, new_n6166_ );
or   ( new_n10751_, new_n10750_, new_n10746_ );
and  ( new_n10752_, new_n10750_, new_n10746_ );
or   ( new_n10753_, new_n6173_, new_n886_ );
or   ( new_n10754_, new_n6175_, new_n805_ );
and  ( new_n10755_, new_n10754_, new_n10753_ );
xor  ( new_n10756_, new_n10755_, new_n5597_ );
or   ( new_n10757_, new_n10756_, new_n10752_ );
and  ( new_n10758_, new_n10757_, new_n10751_ );
or   ( new_n10759_, new_n10758_, new_n10742_ );
and  ( new_n10760_, new_n10758_, new_n10742_ );
or   ( new_n10761_, new_n10059_, new_n313_ );
or   ( new_n10762_, new_n10061_, new_n319_ );
and  ( new_n10763_, new_n10762_, new_n10761_ );
xor  ( new_n10764_, new_n10763_, new_n9421_ );
and  ( new_n10765_, RIbb2d888_64, RIbb2d810_65 );
or   ( new_n10766_, RIbb2d888_64, new_n333_ );
and  ( new_n10767_, new_n10766_, RIbb2d900_63 );
or   ( new_n10768_, new_n10767_, new_n10765_ );
and  ( new_n10769_, RIbb2d888_64, RIbb2d900_63 );
not  ( new_n10770_, new_n10769_ );
or   ( new_n10771_, new_n10770_, new_n339_ );
and  ( new_n10772_, new_n10771_, new_n10768_ );
nor  ( new_n10773_, new_n10772_, new_n10764_ );
and  ( new_n10774_, new_n10772_, new_n10764_ );
or   ( new_n10775_, new_n9422_, new_n279_ );
or   ( new_n10776_, new_n9424_, new_n285_ );
and  ( new_n10777_, new_n10776_, new_n10775_ );
xor  ( new_n10778_, new_n10777_, new_n8873_ );
nor  ( new_n10779_, new_n10778_, new_n10774_ );
nor  ( new_n10780_, new_n10779_, new_n10773_ );
or   ( new_n10781_, new_n10780_, new_n10760_ );
and  ( new_n10782_, new_n10781_, new_n10759_ );
or   ( new_n10783_, new_n10782_, new_n10726_ );
or   ( new_n10784_, new_n2122_, new_n3820_ );
or   ( new_n10785_, new_n2124_, new_n3694_ );
and  ( new_n10786_, new_n10785_, new_n10784_ );
xor  ( new_n10787_, new_n10786_, new_n1843_ );
or   ( new_n10788_, new_n1844_, new_n4267_ );
or   ( new_n10789_, new_n1846_, new_n4069_ );
and  ( new_n10790_, new_n10789_, new_n10788_ );
xor  ( new_n10791_, new_n10790_, new_n1586_ );
or   ( new_n10792_, new_n10791_, new_n10787_ );
and  ( new_n10793_, new_n10791_, new_n10787_ );
or   ( new_n10794_, new_n1593_, new_n4995_ );
or   ( new_n10795_, new_n1595_, new_n4603_ );
and  ( new_n10796_, new_n10795_, new_n10794_ );
xor  ( new_n10797_, new_n10796_, new_n1358_ );
or   ( new_n10798_, new_n10797_, new_n10793_ );
and  ( new_n10799_, new_n10798_, new_n10792_ );
or   ( new_n10800_, new_n1364_, new_n5171_ );
or   ( new_n10801_, new_n1366_, new_n4859_ );
and  ( new_n10802_, new_n10801_, new_n10800_ );
xor  ( new_n10803_, new_n10802_, new_n1129_ );
or   ( new_n10804_, new_n1135_, new_n5570_ );
or   ( new_n10805_, new_n1137_, new_n5428_ );
and  ( new_n10806_, new_n10805_, new_n10804_ );
xor  ( new_n10807_, new_n10806_, new_n896_ );
or   ( new_n10808_, new_n10807_, new_n10803_ );
and  ( new_n10809_, new_n10807_, new_n10803_ );
or   ( new_n10810_, new_n897_, new_n6219_ );
or   ( new_n10811_, new_n899_, new_n5899_ );
and  ( new_n10812_, new_n10811_, new_n10810_ );
xor  ( new_n10813_, new_n10812_, new_n748_ );
or   ( new_n10814_, new_n10813_, new_n10809_ );
and  ( new_n10815_, new_n10814_, new_n10808_ );
or   ( new_n10816_, new_n10815_, new_n10799_ );
and  ( new_n10817_, new_n10815_, new_n10799_ );
or   ( new_n10818_, new_n755_, new_n6589_ );
or   ( new_n10819_, new_n757_, new_n6425_ );
and  ( new_n10820_, new_n10819_, new_n10818_ );
xor  ( new_n10821_, new_n10820_, new_n523_ );
or   ( new_n10822_, new_n524_, new_n7149_ );
or   ( new_n10823_, new_n526_, new_n6943_ );
and  ( new_n10824_, new_n10823_, new_n10822_ );
xor  ( new_n10825_, new_n10824_, new_n403_ );
nor  ( new_n10826_, new_n10825_, new_n10821_ );
and  ( new_n10827_, new_n10825_, new_n10821_ );
or   ( new_n10828_, new_n409_, new_n8117_ );
or   ( new_n10829_, new_n411_, new_n7373_ );
and  ( new_n10830_, new_n10829_, new_n10828_ );
xor  ( new_n10831_, new_n10830_, new_n328_ );
nor  ( new_n10832_, new_n10831_, new_n10827_ );
nor  ( new_n10833_, new_n10832_, new_n10826_ );
or   ( new_n10834_, new_n10833_, new_n10817_ );
and  ( new_n10835_, new_n10834_, new_n10816_ );
and  ( new_n10836_, new_n10782_, new_n10726_ );
or   ( new_n10837_, new_n10836_, new_n10835_ );
and  ( new_n10838_, new_n10837_, new_n10783_ );
and  ( new_n10839_, new_n10838_, new_n10674_ );
nor  ( new_n10840_, new_n10838_, new_n10674_ );
not  ( new_n10841_, RIbb31578_128 );
or   ( new_n10842_, new_n10841_, new_n260_ );
xnor ( new_n10843_, new_n10538_, new_n10534_ );
xor  ( new_n10844_, new_n10843_, new_n10545_ );
or   ( new_n10845_, new_n10844_, new_n10842_ );
and  ( new_n10846_, new_n10844_, new_n10842_ );
or   ( new_n10847_, new_n337_, new_n8352_ );
or   ( new_n10848_, new_n340_, new_n8115_ );
and  ( new_n10849_, new_n10848_, new_n10847_ );
xor  ( new_n10850_, new_n10849_, new_n332_ );
or   ( new_n10851_, new_n317_, new_n8995_ );
or   ( new_n10852_, new_n320_, new_n8481_ );
and  ( new_n10853_, new_n10852_, new_n10851_ );
xor  ( new_n10854_, new_n10853_, new_n312_ );
nor  ( new_n10855_, new_n10854_, new_n10850_ );
and  ( new_n10856_, new_n10854_, new_n10850_ );
or   ( new_n10857_, new_n283_, new_n9681_ );
or   ( new_n10858_, new_n286_, new_n9099_ );
and  ( new_n10859_, new_n10858_, new_n10857_ );
xor  ( new_n10860_, new_n10859_, new_n278_ );
nor  ( new_n10861_, new_n10860_, new_n10856_ );
nor  ( new_n10862_, new_n10861_, new_n10855_ );
not  ( new_n10863_, new_n10862_ );
or   ( new_n10864_, new_n10863_, new_n10846_ );
and  ( new_n10865_, new_n10864_, new_n10845_ );
xnor ( new_n10866_, new_n10437_, new_n10433_ );
xor  ( new_n10867_, new_n10866_, new_n10443_ );
xnor ( new_n10868_, new_n10421_, new_n10417_ );
xor  ( new_n10869_, new_n10868_, new_n10427_ );
or   ( new_n10870_, new_n10869_, new_n10867_ );
and  ( new_n10871_, new_n10869_, new_n10867_ );
xnor ( new_n10872_, new_n10403_, new_n10399_ );
xor  ( new_n10873_, new_n10872_, new_n10409_ );
or   ( new_n10874_, new_n10873_, new_n10871_ );
and  ( new_n10875_, new_n10874_, new_n10870_ );
nor  ( new_n10876_, new_n10875_, new_n10865_ );
and  ( new_n10877_, new_n10875_, new_n10865_ );
xnor ( new_n10878_, new_n10385_, new_n10381_ );
xor  ( new_n10879_, new_n10878_, new_n10391_ );
xnor ( new_n10880_, new_n10522_, new_n10518_ );
xor  ( new_n10881_, new_n10880_, new_n10528_ );
nor  ( new_n10882_, new_n10881_, new_n10879_ );
and  ( new_n10883_, new_n10881_, new_n10879_ );
xor  ( new_n10884_, new_n10369_, new_n10365_ );
xnor ( new_n10885_, new_n10884_, new_n10375_ );
nor  ( new_n10886_, new_n10885_, new_n10883_ );
nor  ( new_n10887_, new_n10886_, new_n10882_ );
nor  ( new_n10888_, new_n10887_, new_n10877_ );
nor  ( new_n10889_, new_n10888_, new_n10876_ );
nor  ( new_n10890_, new_n10889_, new_n10840_ );
nor  ( new_n10891_, new_n10890_, new_n10839_ );
nor  ( new_n10892_, new_n10891_, new_n10657_ );
nor  ( new_n10893_, new_n10892_, new_n10656_ );
nand ( new_n10894_, new_n10893_, new_n10619_ );
and  ( new_n10895_, new_n10894_, new_n10618_ );
nand ( new_n10896_, new_n10895_, new_n10605_ );
nor  ( new_n10897_, new_n10895_, new_n10605_ );
xor  ( new_n10898_, new_n9970_, new_n9968_ );
xor  ( new_n10899_, new_n10898_, new_n9975_ );
or   ( new_n10900_, new_n10899_, new_n10897_ );
and  ( new_n10901_, new_n10900_, new_n10896_ );
or   ( new_n10902_, new_n10901_, new_n10600_ );
nand ( new_n10903_, new_n10901_, new_n10600_ );
xor  ( new_n10904_, new_n10580_, new_n10578_ );
xnor ( new_n10905_, new_n10904_, new_n10584_ );
nand ( new_n10906_, new_n10905_, new_n10903_ );
and  ( new_n10907_, new_n10906_, new_n10902_ );
nor  ( new_n10908_, new_n10907_, new_n10595_ );
xor  ( new_n10909_, new_n10901_, new_n10600_ );
xor  ( new_n10910_, new_n10909_, new_n10905_ );
xnor ( new_n10911_, new_n10663_, new_n10661_ );
xor  ( new_n10912_, new_n10911_, new_n10667_ );
xnor ( new_n10913_, new_n10881_, new_n10879_ );
xor  ( new_n10914_, new_n10913_, new_n10885_ );
nor  ( new_n10915_, new_n10914_, new_n10912_ );
nand ( new_n10916_, new_n10914_, new_n10912_ );
xor  ( new_n10917_, new_n10869_, new_n10867_ );
xor  ( new_n10918_, new_n10917_, new_n10873_ );
and  ( new_n10919_, new_n10918_, new_n10916_ );
or   ( new_n10920_, new_n10919_, new_n10915_ );
xor  ( new_n10921_, new_n10636_, new_n10634_ );
xor  ( new_n10922_, new_n10921_, new_n10641_ );
nor  ( new_n10923_, new_n10922_, new_n10920_ );
nand ( new_n10924_, new_n10922_, new_n10920_ );
xnor ( new_n10925_, new_n10706_, new_n10690_ );
xor  ( new_n10926_, new_n10925_, new_n10724_ );
xnor ( new_n10927_, new_n10815_, new_n10799_ );
xor  ( new_n10928_, new_n10927_, new_n10833_ );
nor  ( new_n10929_, new_n10928_, new_n10926_ );
and  ( new_n10930_, new_n10928_, new_n10926_ );
xor  ( new_n10931_, new_n10844_, new_n10842_ );
xor  ( new_n10932_, new_n10931_, new_n10863_ );
nor  ( new_n10933_, new_n10932_, new_n10930_ );
or   ( new_n10934_, new_n10933_, new_n10929_ );
and  ( new_n10935_, new_n10934_, new_n10924_ );
or   ( new_n10936_, new_n10935_, new_n10923_ );
xor  ( new_n10937_, new_n10734_, new_n10730_ );
xnor ( new_n10938_, new_n10937_, new_n10740_ );
xnor ( new_n10939_, new_n10772_, new_n10764_ );
xor  ( new_n10940_, new_n10939_, new_n10778_ );
or   ( new_n10941_, new_n10940_, new_n10938_ );
xnor ( new_n10942_, new_n10698_, new_n10694_ );
xor  ( new_n10943_, new_n10942_, new_n10704_ );
xnor ( new_n10944_, new_n10682_, new_n10678_ );
xor  ( new_n10945_, new_n10944_, new_n10688_ );
or   ( new_n10946_, new_n10945_, new_n10943_ );
and  ( new_n10947_, new_n10945_, new_n10943_ );
xnor ( new_n10948_, new_n10750_, new_n10746_ );
xor  ( new_n10949_, new_n10948_, new_n10756_ );
or   ( new_n10950_, new_n10949_, new_n10947_ );
and  ( new_n10951_, new_n10950_, new_n10946_ );
nor  ( new_n10952_, new_n10951_, new_n10941_ );
nand ( new_n10953_, new_n10951_, new_n10941_ );
xor  ( new_n10954_, new_n10489_, new_n10487_ );
and  ( new_n10955_, new_n10954_, new_n10953_ );
or   ( new_n10956_, new_n10955_, new_n10952_ );
xnor ( new_n10957_, new_n10807_, new_n10803_ );
xor  ( new_n10958_, new_n10957_, new_n10813_ );
xnor ( new_n10959_, new_n10791_, new_n10787_ );
xor  ( new_n10960_, new_n10959_, new_n10797_ );
nor  ( new_n10961_, new_n10960_, new_n10958_ );
and  ( new_n10962_, new_n10960_, new_n10958_ );
xor  ( new_n10963_, new_n10716_, new_n10712_ );
xnor ( new_n10964_, new_n10963_, new_n10722_ );
nor  ( new_n10965_, new_n10964_, new_n10962_ );
or   ( new_n10966_, new_n10965_, new_n10961_ );
or   ( new_n10967_, new_n299_, new_n10220_ );
or   ( new_n10968_, new_n302_, new_n9679_ );
and  ( new_n10969_, new_n10968_, new_n10967_ );
xor  ( new_n10970_, new_n10969_, new_n293_ );
or   ( new_n10971_, new_n283_, new_n9679_ );
or   ( new_n10972_, new_n286_, new_n9681_ );
and  ( new_n10973_, new_n10972_, new_n10971_ );
xor  ( new_n10974_, new_n10973_, new_n278_ );
or   ( new_n10975_, new_n299_, new_n10541_ );
or   ( new_n10976_, new_n302_, new_n10220_ );
and  ( new_n10977_, new_n10976_, new_n10975_ );
xor  ( new_n10978_, new_n10977_, new_n293_ );
or   ( new_n10979_, new_n10978_, new_n10974_ );
and  ( new_n10980_, new_n10978_, new_n10974_ );
and  ( new_n10981_, new_n265_, RIbb31578_128 );
nor  ( new_n10982_, new_n10981_, new_n262_ );
and  ( new_n10983_, new_n10981_, RIbb2f610_1 );
nor  ( new_n10984_, new_n10983_, new_n10982_ );
or   ( new_n10985_, new_n10984_, new_n10980_ );
and  ( new_n10986_, new_n10985_, new_n10979_ );
or   ( new_n10987_, new_n10986_, new_n10970_ );
and  ( new_n10988_, new_n10986_, new_n10970_ );
or   ( new_n10989_, new_n409_, new_n8115_ );
or   ( new_n10990_, new_n411_, new_n8117_ );
and  ( new_n10991_, new_n10990_, new_n10989_ );
xor  ( new_n10992_, new_n10991_, new_n328_ );
or   ( new_n10993_, new_n337_, new_n8481_ );
or   ( new_n10994_, new_n340_, new_n8352_ );
and  ( new_n10995_, new_n10994_, new_n10993_ );
xor  ( new_n10996_, new_n10995_, new_n332_ );
nor  ( new_n10997_, new_n10996_, new_n10992_ );
and  ( new_n10998_, new_n10996_, new_n10992_ );
or   ( new_n10999_, new_n317_, new_n9099_ );
or   ( new_n11000_, new_n320_, new_n8995_ );
and  ( new_n11001_, new_n11000_, new_n10999_ );
xor  ( new_n11002_, new_n11001_, new_n312_ );
nor  ( new_n11003_, new_n11002_, new_n10998_ );
nor  ( new_n11004_, new_n11003_, new_n10997_ );
or   ( new_n11005_, new_n11004_, new_n10988_ );
and  ( new_n11006_, new_n11005_, new_n10987_ );
or   ( new_n11007_, new_n11006_, new_n10966_ );
and  ( new_n11008_, new_n11006_, new_n10966_ );
or   ( new_n11009_, new_n268_, new_n10841_ );
or   ( new_n11010_, new_n271_, new_n10541_ );
and  ( new_n11011_, new_n11010_, new_n11009_ );
xor  ( new_n11012_, new_n11011_, new_n262_ );
xnor ( new_n11013_, new_n10825_, new_n10821_ );
xor  ( new_n11014_, new_n11013_, new_n10831_ );
and  ( new_n11015_, new_n11014_, new_n11012_ );
nor  ( new_n11016_, new_n11014_, new_n11012_ );
xor  ( new_n11017_, new_n10854_, new_n10850_ );
xnor ( new_n11018_, new_n11017_, new_n10860_ );
not  ( new_n11019_, new_n11018_ );
nor  ( new_n11020_, new_n11019_, new_n11016_ );
nor  ( new_n11021_, new_n11020_, new_n11015_ );
or   ( new_n11022_, new_n11021_, new_n11008_ );
and  ( new_n11023_, new_n11022_, new_n11007_ );
or   ( new_n11024_, new_n11023_, new_n10956_ );
and  ( new_n11025_, new_n11023_, new_n10956_ );
or   ( new_n11026_, new_n2425_, new_n3694_ );
or   ( new_n11027_, new_n2427_, new_n3696_ );
and  ( new_n11028_, new_n11027_, new_n11026_ );
xor  ( new_n11029_, new_n11028_, new_n2121_ );
or   ( new_n11030_, new_n2122_, new_n4069_ );
or   ( new_n11031_, new_n2124_, new_n3820_ );
and  ( new_n11032_, new_n11031_, new_n11030_ );
xor  ( new_n11033_, new_n11032_, new_n1843_ );
or   ( new_n11034_, new_n11033_, new_n11029_ );
and  ( new_n11035_, new_n11033_, new_n11029_ );
or   ( new_n11036_, new_n1844_, new_n4603_ );
or   ( new_n11037_, new_n1846_, new_n4267_ );
and  ( new_n11038_, new_n11037_, new_n11036_ );
xor  ( new_n11039_, new_n11038_, new_n1586_ );
or   ( new_n11040_, new_n11039_, new_n11035_ );
and  ( new_n11041_, new_n11040_, new_n11034_ );
or   ( new_n11042_, new_n1593_, new_n4859_ );
or   ( new_n11043_, new_n1595_, new_n4995_ );
and  ( new_n11044_, new_n11043_, new_n11042_ );
xor  ( new_n11045_, new_n11044_, new_n1358_ );
or   ( new_n11046_, new_n1364_, new_n5428_ );
or   ( new_n11047_, new_n1366_, new_n5171_ );
and  ( new_n11048_, new_n11047_, new_n11046_ );
xor  ( new_n11049_, new_n11048_, new_n1129_ );
or   ( new_n11050_, new_n11049_, new_n11045_ );
and  ( new_n11051_, new_n11049_, new_n11045_ );
or   ( new_n11052_, new_n1135_, new_n5899_ );
or   ( new_n11053_, new_n1137_, new_n5570_ );
and  ( new_n11054_, new_n11053_, new_n11052_ );
xor  ( new_n11055_, new_n11054_, new_n896_ );
or   ( new_n11056_, new_n11055_, new_n11051_ );
and  ( new_n11057_, new_n11056_, new_n11050_ );
or   ( new_n11058_, new_n11057_, new_n11041_ );
and  ( new_n11059_, new_n11057_, new_n11041_ );
or   ( new_n11060_, new_n897_, new_n6425_ );
or   ( new_n11061_, new_n899_, new_n6219_ );
and  ( new_n11062_, new_n11061_, new_n11060_ );
xor  ( new_n11063_, new_n11062_, new_n748_ );
or   ( new_n11064_, new_n755_, new_n6943_ );
or   ( new_n11065_, new_n757_, new_n6589_ );
and  ( new_n11066_, new_n11065_, new_n11064_ );
xor  ( new_n11067_, new_n11066_, new_n523_ );
or   ( new_n11068_, new_n11067_, new_n11063_ );
and  ( new_n11069_, new_n11067_, new_n11063_ );
or   ( new_n11070_, new_n524_, new_n7373_ );
or   ( new_n11071_, new_n526_, new_n7149_ );
and  ( new_n11072_, new_n11071_, new_n11070_ );
xor  ( new_n11073_, new_n11072_, new_n403_ );
or   ( new_n11074_, new_n11073_, new_n11069_ );
and  ( new_n11075_, new_n11074_, new_n11068_ );
or   ( new_n11076_, new_n11075_, new_n11059_ );
and  ( new_n11077_, new_n11076_, new_n11058_ );
or   ( new_n11078_, new_n7732_, new_n443_ );
or   ( new_n11079_, new_n7734_, new_n419_ );
and  ( new_n11080_, new_n11079_, new_n11078_ );
xor  ( new_n11081_, new_n11080_, new_n7177_ );
or   ( new_n11082_, new_n7184_, new_n515_ );
or   ( new_n11083_, new_n7186_, new_n509_ );
and  ( new_n11084_, new_n11083_, new_n11082_ );
xor  ( new_n11085_, new_n11084_, new_n6638_ );
nor  ( new_n11086_, new_n11085_, new_n11081_ );
and  ( new_n11087_, new_n11085_, new_n11081_ );
or   ( new_n11088_, new_n6645_, new_n805_ );
or   ( new_n11089_, new_n6647_, new_n775_ );
and  ( new_n11090_, new_n11089_, new_n11088_ );
xor  ( new_n11091_, new_n11090_, new_n6166_ );
nor  ( new_n11092_, new_n11091_, new_n11087_ );
nor  ( new_n11093_, new_n11092_, new_n11086_ );
or   ( new_n11094_, new_n10059_, new_n285_ );
or   ( new_n11095_, new_n10061_, new_n313_ );
and  ( new_n11096_, new_n11095_, new_n11094_ );
xor  ( new_n11097_, new_n11096_, new_n9421_ );
and  ( new_n11098_, RIbb2d888_64, RIbb2d798_66 );
or   ( new_n11099_, RIbb2d888_64, new_n319_ );
and  ( new_n11100_, new_n11099_, RIbb2d900_63 );
or   ( new_n11101_, new_n11100_, new_n11098_ );
or   ( new_n11102_, new_n10770_, new_n333_ );
and  ( new_n11103_, new_n11102_, new_n11101_ );
nor  ( new_n11104_, new_n11103_, new_n11097_ );
and  ( new_n11105_, new_n11103_, new_n11097_ );
nor  ( new_n11106_, new_n11105_, new_n262_ );
nor  ( new_n11107_, new_n11106_, new_n11104_ );
or   ( new_n11108_, new_n9422_, new_n301_ );
or   ( new_n11109_, new_n9424_, new_n279_ );
and  ( new_n11110_, new_n11109_, new_n11108_ );
xor  ( new_n11111_, new_n11110_, new_n8873_ );
or   ( new_n11112_, new_n8874_, new_n270_ );
or   ( new_n11113_, new_n8876_, new_n294_ );
and  ( new_n11114_, new_n11113_, new_n11112_ );
xor  ( new_n11115_, new_n11114_, new_n8257_ );
or   ( new_n11116_, new_n11115_, new_n11111_ );
and  ( new_n11117_, new_n11115_, new_n11111_ );
or   ( new_n11118_, new_n8264_, new_n348_ );
or   ( new_n11119_, new_n8266_, new_n264_ );
and  ( new_n11120_, new_n11119_, new_n11118_ );
xor  ( new_n11121_, new_n11120_, new_n7725_ );
or   ( new_n11122_, new_n11121_, new_n11117_ );
and  ( new_n11123_, new_n11122_, new_n11116_ );
and  ( new_n11124_, new_n11123_, new_n11107_ );
or   ( new_n11125_, new_n11124_, new_n11093_ );
or   ( new_n11126_, new_n11123_, new_n11107_ );
and  ( new_n11127_, new_n11126_, new_n11125_ );
nor  ( new_n11128_, new_n11127_, new_n11077_ );
or   ( new_n11129_, new_n6173_, new_n986_ );
or   ( new_n11130_, new_n6175_, new_n886_ );
and  ( new_n11131_, new_n11130_, new_n11129_ );
xor  ( new_n11132_, new_n11131_, new_n5597_ );
or   ( new_n11133_, new_n5604_, new_n1213_ );
or   ( new_n11134_, new_n5606_, new_n1168_ );
and  ( new_n11135_, new_n11134_, new_n11133_ );
xor  ( new_n11136_, new_n11135_, new_n5206_ );
or   ( new_n11137_, new_n11136_, new_n11132_ );
and  ( new_n11138_, new_n11136_, new_n11132_ );
or   ( new_n11139_, new_n5207_, new_n1525_ );
or   ( new_n11140_, new_n5209_, new_n1318_ );
and  ( new_n11141_, new_n11140_, new_n11139_ );
xor  ( new_n11142_, new_n11141_, new_n4708_ );
or   ( new_n11143_, new_n11142_, new_n11138_ );
and  ( new_n11144_, new_n11143_, new_n11137_ );
or   ( new_n11145_, new_n4709_, new_n1754_ );
or   ( new_n11146_, new_n4711_, new_n1523_ );
and  ( new_n11147_, new_n11146_, new_n11145_ );
xor  ( new_n11148_, new_n11147_, new_n4295_ );
or   ( new_n11149_, new_n4302_, new_n2057_ );
or   ( new_n11150_, new_n4304_, new_n1899_ );
and  ( new_n11151_, new_n11150_, new_n11149_ );
xor  ( new_n11152_, new_n11151_, new_n3895_ );
or   ( new_n11153_, new_n11152_, new_n11148_ );
and  ( new_n11154_, new_n11152_, new_n11148_ );
or   ( new_n11155_, new_n3896_, new_n2291_ );
or   ( new_n11156_, new_n3898_, new_n2178_ );
and  ( new_n11157_, new_n11156_, new_n11155_ );
xor  ( new_n11158_, new_n11157_, new_n3460_ );
or   ( new_n11159_, new_n11158_, new_n11154_ );
and  ( new_n11160_, new_n11159_, new_n11153_ );
nor  ( new_n11161_, new_n11160_, new_n11144_ );
and  ( new_n11162_, new_n11160_, new_n11144_ );
or   ( new_n11163_, new_n3461_, new_n2646_ );
or   ( new_n11164_, new_n3463_, new_n2475_ );
and  ( new_n11165_, new_n11164_, new_n11163_ );
xor  ( new_n11166_, new_n11165_, new_n3116_ );
or   ( new_n11167_, new_n3117_, new_n2981_ );
or   ( new_n11168_, new_n3119_, new_n2751_ );
and  ( new_n11169_, new_n11168_, new_n11167_ );
xor  ( new_n11170_, new_n11169_, new_n2800_ );
nor  ( new_n11171_, new_n11170_, new_n11166_ );
and  ( new_n11172_, new_n11170_, new_n11166_ );
or   ( new_n11173_, new_n2807_, new_n3306_ );
or   ( new_n11174_, new_n2809_, new_n3178_ );
and  ( new_n11175_, new_n11174_, new_n11173_ );
xor  ( new_n11176_, new_n11175_, new_n2424_ );
nor  ( new_n11177_, new_n11176_, new_n11172_ );
nor  ( new_n11178_, new_n11177_, new_n11171_ );
nor  ( new_n11179_, new_n11178_, new_n11162_ );
nor  ( new_n11180_, new_n11179_, new_n11161_ );
and  ( new_n11181_, new_n11127_, new_n11077_ );
nor  ( new_n11182_, new_n11181_, new_n11180_ );
nor  ( new_n11183_, new_n11182_, new_n11128_ );
or   ( new_n11184_, new_n11183_, new_n11025_ );
and  ( new_n11185_, new_n11184_, new_n11024_ );
nor  ( new_n11186_, new_n11185_, new_n10936_ );
nand ( new_n11187_, new_n11185_, new_n10936_ );
xor  ( new_n11188_, new_n10875_, new_n10865_ );
xor  ( new_n11189_, new_n11188_, new_n10887_ );
xor  ( new_n11190_, new_n10623_, new_n10621_ );
xor  ( new_n11191_, new_n11190_, new_n10626_ );
or   ( new_n11192_, new_n11191_, new_n11189_ );
nand ( new_n11193_, new_n11191_, new_n11189_ );
xor  ( new_n11194_, new_n10669_, new_n10659_ );
xor  ( new_n11195_, new_n11194_, new_n10672_ );
nand ( new_n11196_, new_n11195_, new_n11193_ );
and  ( new_n11197_, new_n11196_, new_n11192_ );
and  ( new_n11198_, new_n11197_, new_n11187_ );
or   ( new_n11199_, new_n11198_, new_n11186_ );
xor  ( new_n11200_, new_n10558_, new_n10548_ );
xor  ( new_n11201_, new_n11200_, new_n10570_ );
xnor ( new_n11202_, new_n10465_, new_n10413_ );
xor  ( new_n11203_, new_n11202_, new_n10510_ );
or   ( new_n11204_, new_n11203_, new_n11201_ );
and  ( new_n11205_, new_n11203_, new_n11201_ );
xor  ( new_n11206_, new_n10649_, new_n10647_ );
xnor ( new_n11207_, new_n11206_, new_n10653_ );
not  ( new_n11208_, new_n11207_ );
or   ( new_n11209_, new_n11208_, new_n11205_ );
and  ( new_n11210_, new_n11209_, new_n11204_ );
or   ( new_n11211_, new_n11210_, new_n11199_ );
nand ( new_n11212_, new_n11210_, new_n11199_ );
xor  ( new_n11213_, new_n10512_, new_n10361_ );
xnor ( new_n11214_, new_n11213_, new_n10572_ );
nand ( new_n11215_, new_n11214_, new_n11212_ );
and  ( new_n11216_, new_n11215_, new_n11211_ );
xor  ( new_n11217_, new_n10617_, new_n10607_ );
xor  ( new_n11218_, new_n11217_, new_n10893_ );
nor  ( new_n11219_, new_n11218_, new_n11216_ );
nand ( new_n11220_, new_n11218_, new_n11216_ );
xor  ( new_n11221_, new_n10604_, new_n10602_ );
and  ( new_n11222_, new_n11221_, new_n11220_ );
or   ( new_n11223_, new_n11222_, new_n11219_ );
xnor ( new_n11224_, new_n10895_, new_n10605_ );
xor  ( new_n11225_, new_n11224_, new_n10899_ );
or   ( new_n11226_, new_n11225_, new_n11223_ );
and  ( new_n11227_, new_n11225_, new_n11223_ );
xor  ( new_n11228_, new_n10599_, new_n10597_ );
or   ( new_n11229_, new_n11228_, new_n11227_ );
and  ( new_n11230_, new_n11229_, new_n11226_ );
and  ( new_n11231_, new_n11230_, new_n10910_ );
xnor ( new_n11232_, new_n11225_, new_n11223_ );
xor  ( new_n11233_, new_n11232_, new_n11228_ );
xor  ( new_n11234_, new_n10655_, new_n10645_ );
xnor ( new_n11235_, new_n11234_, new_n10891_ );
xor  ( new_n11236_, new_n11210_, new_n11199_ );
xor  ( new_n11237_, new_n11236_, new_n11214_ );
nand ( new_n11238_, new_n11237_, new_n11235_ );
xor  ( new_n11239_, new_n10838_, new_n10674_ );
xor  ( new_n11240_, new_n11239_, new_n10889_ );
xor  ( new_n11241_, new_n11185_, new_n10936_ );
xor  ( new_n11242_, new_n11241_, new_n11197_ );
nor  ( new_n11243_, new_n11242_, new_n11240_ );
and  ( new_n11244_, new_n11242_, new_n11240_ );
xor  ( new_n11245_, new_n11203_, new_n11201_ );
xor  ( new_n11246_, new_n11245_, new_n11208_ );
nor  ( new_n11247_, new_n11246_, new_n11244_ );
or   ( new_n11248_, new_n11247_, new_n11243_ );
xor  ( new_n11249_, new_n10782_, new_n10726_ );
xor  ( new_n11250_, new_n11249_, new_n10835_ );
xor  ( new_n11251_, new_n10922_, new_n10920_ );
xor  ( new_n11252_, new_n11251_, new_n10934_ );
or   ( new_n11253_, new_n11252_, new_n11250_ );
and  ( new_n11254_, new_n11252_, new_n11250_ );
xor  ( new_n11255_, new_n11191_, new_n11189_ );
xor  ( new_n11256_, new_n11255_, new_n11195_ );
or   ( new_n11257_, new_n11256_, new_n11254_ );
and  ( new_n11258_, new_n11257_, new_n11253_ );
xor  ( new_n11259_, new_n10960_, new_n10958_ );
xor  ( new_n11260_, new_n11259_, new_n10964_ );
xnor ( new_n11261_, new_n10986_, new_n10970_ );
xor  ( new_n11262_, new_n11261_, new_n11004_ );
or   ( new_n11263_, new_n11262_, new_n11260_ );
and  ( new_n11264_, new_n11262_, new_n11260_ );
xor  ( new_n11265_, new_n11014_, new_n11012_ );
xor  ( new_n11266_, new_n11265_, new_n11018_ );
or   ( new_n11267_, new_n11266_, new_n11264_ );
and  ( new_n11268_, new_n11267_, new_n11263_ );
xor  ( new_n11269_, new_n11057_, new_n11041_ );
xor  ( new_n11270_, new_n11269_, new_n11075_ );
xor  ( new_n11271_, new_n11123_, new_n11107_ );
xor  ( new_n11272_, new_n11271_, new_n11093_ );
nand ( new_n11273_, new_n11272_, new_n11270_ );
nor  ( new_n11274_, new_n11272_, new_n11270_ );
xor  ( new_n11275_, new_n11160_, new_n11144_ );
xnor ( new_n11276_, new_n11275_, new_n11178_ );
or   ( new_n11277_, new_n11276_, new_n11274_ );
and  ( new_n11278_, new_n11277_, new_n11273_ );
nor  ( new_n11279_, new_n11278_, new_n11268_ );
and  ( new_n11280_, new_n11278_, new_n11268_ );
xor  ( new_n11281_, new_n10758_, new_n10742_ );
xnor ( new_n11282_, new_n11281_, new_n10780_ );
nor  ( new_n11283_, new_n11282_, new_n11280_ );
or   ( new_n11284_, new_n11283_, new_n11279_ );
xnor ( new_n11285_, new_n11152_, new_n11148_ );
xor  ( new_n11286_, new_n11285_, new_n11158_ );
xnor ( new_n11287_, new_n11136_, new_n11132_ );
xor  ( new_n11288_, new_n11287_, new_n11142_ );
nor  ( new_n11289_, new_n11288_, new_n11286_ );
nand ( new_n11290_, new_n11288_, new_n11286_ );
xor  ( new_n11291_, new_n11170_, new_n11166_ );
xnor ( new_n11292_, new_n11291_, new_n11176_ );
not  ( new_n11293_, new_n11292_ );
and  ( new_n11294_, new_n11293_, new_n11290_ );
or   ( new_n11295_, new_n11294_, new_n11289_ );
xor  ( new_n11296_, new_n10996_, new_n10992_ );
xor  ( new_n11297_, new_n11296_, new_n11002_ );
or   ( new_n11298_, new_n337_, new_n8995_ );
or   ( new_n11299_, new_n340_, new_n8481_ );
and  ( new_n11300_, new_n11299_, new_n11298_ );
xor  ( new_n11301_, new_n11300_, new_n332_ );
or   ( new_n11302_, new_n317_, new_n9681_ );
or   ( new_n11303_, new_n320_, new_n9099_ );
and  ( new_n11304_, new_n11303_, new_n11302_ );
xor  ( new_n11305_, new_n11304_, new_n312_ );
or   ( new_n11306_, new_n11305_, new_n11301_ );
and  ( new_n11307_, new_n11305_, new_n11301_ );
or   ( new_n11308_, new_n283_, new_n10220_ );
or   ( new_n11309_, new_n286_, new_n9679_ );
and  ( new_n11310_, new_n11309_, new_n11308_ );
xor  ( new_n11311_, new_n11310_, new_n278_ );
or   ( new_n11312_, new_n11311_, new_n11307_ );
and  ( new_n11313_, new_n11312_, new_n11306_ );
or   ( new_n11314_, new_n11313_, new_n11297_ );
nand ( new_n11315_, new_n11313_, new_n11297_ );
xor  ( new_n11316_, new_n10978_, new_n10974_ );
xnor ( new_n11317_, new_n11316_, new_n10984_ );
nand ( new_n11318_, new_n11317_, new_n11315_ );
and  ( new_n11319_, new_n11318_, new_n11314_ );
and  ( new_n11320_, new_n11319_, new_n11295_ );
or   ( new_n11321_, new_n11319_, new_n11295_ );
xnor ( new_n11322_, new_n11049_, new_n11045_ );
xor  ( new_n11323_, new_n11322_, new_n11055_ );
xnor ( new_n11324_, new_n11033_, new_n11029_ );
xor  ( new_n11325_, new_n11324_, new_n11039_ );
nor  ( new_n11326_, new_n11325_, new_n11323_ );
nand ( new_n11327_, new_n11325_, new_n11323_ );
xor  ( new_n11328_, new_n11067_, new_n11063_ );
xnor ( new_n11329_, new_n11328_, new_n11073_ );
not  ( new_n11330_, new_n11329_ );
and  ( new_n11331_, new_n11330_, new_n11327_ );
or   ( new_n11332_, new_n11331_, new_n11326_ );
and  ( new_n11333_, new_n11332_, new_n11321_ );
or   ( new_n11334_, new_n11333_, new_n11320_ );
or   ( new_n11335_, new_n10059_, new_n279_ );
or   ( new_n11336_, new_n10061_, new_n285_ );
and  ( new_n11337_, new_n11336_, new_n11335_ );
xor  ( new_n11338_, new_n11337_, new_n9421_ );
and  ( new_n11339_, RIbb2d888_64, RIbb2d720_67 );
or   ( new_n11340_, RIbb2d888_64, new_n313_ );
and  ( new_n11341_, new_n11340_, RIbb2d900_63 );
or   ( new_n11342_, new_n11341_, new_n11339_ );
or   ( new_n11343_, new_n10770_, new_n319_ );
and  ( new_n11344_, new_n11343_, new_n11342_ );
or   ( new_n11345_, new_n11344_, new_n11338_ );
and  ( new_n11346_, new_n11344_, new_n11338_ );
or   ( new_n11347_, new_n9422_, new_n294_ );
or   ( new_n11348_, new_n9424_, new_n301_ );
and  ( new_n11349_, new_n11348_, new_n11347_ );
xor  ( new_n11350_, new_n11349_, new_n8873_ );
or   ( new_n11351_, new_n11350_, new_n11346_ );
and  ( new_n11352_, new_n11351_, new_n11345_ );
or   ( new_n11353_, new_n8874_, new_n264_ );
or   ( new_n11354_, new_n8876_, new_n270_ );
and  ( new_n11355_, new_n11354_, new_n11353_ );
xor  ( new_n11356_, new_n11355_, new_n8257_ );
or   ( new_n11357_, new_n8264_, new_n419_ );
or   ( new_n11358_, new_n8266_, new_n348_ );
and  ( new_n11359_, new_n11358_, new_n11357_ );
xor  ( new_n11360_, new_n11359_, new_n7725_ );
or   ( new_n11361_, new_n11360_, new_n11356_ );
and  ( new_n11362_, new_n11360_, new_n11356_ );
or   ( new_n11363_, new_n7732_, new_n509_ );
or   ( new_n11364_, new_n7734_, new_n443_ );
and  ( new_n11365_, new_n11364_, new_n11363_ );
xor  ( new_n11366_, new_n11365_, new_n7177_ );
or   ( new_n11367_, new_n11366_, new_n11362_ );
and  ( new_n11368_, new_n11367_, new_n11361_ );
or   ( new_n11369_, new_n11368_, new_n11352_ );
and  ( new_n11370_, new_n11368_, new_n11352_ );
or   ( new_n11371_, new_n7184_, new_n775_ );
or   ( new_n11372_, new_n7186_, new_n515_ );
and  ( new_n11373_, new_n11372_, new_n11371_ );
xor  ( new_n11374_, new_n11373_, new_n6638_ );
or   ( new_n11375_, new_n6645_, new_n886_ );
or   ( new_n11376_, new_n6647_, new_n805_ );
and  ( new_n11377_, new_n11376_, new_n11375_ );
xor  ( new_n11378_, new_n11377_, new_n6166_ );
nor  ( new_n11379_, new_n11378_, new_n11374_ );
and  ( new_n11380_, new_n11378_, new_n11374_ );
or   ( new_n11381_, new_n6173_, new_n1168_ );
or   ( new_n11382_, new_n6175_, new_n986_ );
and  ( new_n11383_, new_n11382_, new_n11381_ );
xor  ( new_n11384_, new_n11383_, new_n5597_ );
nor  ( new_n11385_, new_n11384_, new_n11380_ );
nor  ( new_n11386_, new_n11385_, new_n11379_ );
or   ( new_n11387_, new_n11386_, new_n11370_ );
and  ( new_n11388_, new_n11387_, new_n11369_ );
or   ( new_n11389_, new_n755_, new_n7149_ );
or   ( new_n11390_, new_n757_, new_n6943_ );
and  ( new_n11391_, new_n11390_, new_n11389_ );
xor  ( new_n11392_, new_n11391_, new_n523_ );
or   ( new_n11393_, new_n524_, new_n8117_ );
or   ( new_n11394_, new_n526_, new_n7373_ );
and  ( new_n11395_, new_n11394_, new_n11393_ );
xor  ( new_n11396_, new_n11395_, new_n403_ );
or   ( new_n11397_, new_n11396_, new_n11392_ );
and  ( new_n11398_, new_n11396_, new_n11392_ );
or   ( new_n11399_, new_n409_, new_n8352_ );
or   ( new_n11400_, new_n411_, new_n8115_ );
and  ( new_n11401_, new_n11400_, new_n11399_ );
xor  ( new_n11402_, new_n11401_, new_n328_ );
or   ( new_n11403_, new_n11402_, new_n11398_ );
and  ( new_n11404_, new_n11403_, new_n11397_ );
or   ( new_n11405_, new_n1364_, new_n5570_ );
or   ( new_n11406_, new_n1366_, new_n5428_ );
and  ( new_n11407_, new_n11406_, new_n11405_ );
xor  ( new_n11408_, new_n11407_, new_n1129_ );
or   ( new_n11409_, new_n1135_, new_n6219_ );
or   ( new_n11410_, new_n1137_, new_n5899_ );
and  ( new_n11411_, new_n11410_, new_n11409_ );
xor  ( new_n11412_, new_n11411_, new_n896_ );
or   ( new_n11413_, new_n11412_, new_n11408_ );
and  ( new_n11414_, new_n11412_, new_n11408_ );
or   ( new_n11415_, new_n897_, new_n6589_ );
or   ( new_n11416_, new_n899_, new_n6425_ );
and  ( new_n11417_, new_n11416_, new_n11415_ );
xor  ( new_n11418_, new_n11417_, new_n748_ );
or   ( new_n11419_, new_n11418_, new_n11414_ );
and  ( new_n11420_, new_n11419_, new_n11413_ );
or   ( new_n11421_, new_n11420_, new_n11404_ );
and  ( new_n11422_, new_n11420_, new_n11404_ );
or   ( new_n11423_, new_n2122_, new_n4267_ );
or   ( new_n11424_, new_n2124_, new_n4069_ );
and  ( new_n11425_, new_n11424_, new_n11423_ );
xor  ( new_n11426_, new_n11425_, new_n1843_ );
or   ( new_n11427_, new_n1844_, new_n4995_ );
or   ( new_n11428_, new_n1846_, new_n4603_ );
and  ( new_n11429_, new_n11428_, new_n11427_ );
xor  ( new_n11430_, new_n11429_, new_n1586_ );
nor  ( new_n11431_, new_n11430_, new_n11426_ );
and  ( new_n11432_, new_n11430_, new_n11426_ );
or   ( new_n11433_, new_n1593_, new_n5171_ );
or   ( new_n11434_, new_n1595_, new_n4859_ );
and  ( new_n11435_, new_n11434_, new_n11433_ );
xor  ( new_n11436_, new_n11435_, new_n1358_ );
nor  ( new_n11437_, new_n11436_, new_n11432_ );
nor  ( new_n11438_, new_n11437_, new_n11431_ );
or   ( new_n11439_, new_n11438_, new_n11422_ );
and  ( new_n11440_, new_n11439_, new_n11421_ );
or   ( new_n11441_, new_n11440_, new_n11388_ );
or   ( new_n11442_, new_n3117_, new_n3178_ );
or   ( new_n11443_, new_n3119_, new_n2981_ );
and  ( new_n11444_, new_n11443_, new_n11442_ );
xor  ( new_n11445_, new_n11444_, new_n2800_ );
or   ( new_n11446_, new_n2807_, new_n3696_ );
or   ( new_n11447_, new_n2809_, new_n3306_ );
and  ( new_n11448_, new_n11447_, new_n11446_ );
xor  ( new_n11449_, new_n11448_, new_n2424_ );
or   ( new_n11450_, new_n11449_, new_n11445_ );
and  ( new_n11451_, new_n11449_, new_n11445_ );
or   ( new_n11452_, new_n2425_, new_n3820_ );
or   ( new_n11453_, new_n2427_, new_n3694_ );
and  ( new_n11454_, new_n11453_, new_n11452_ );
xor  ( new_n11455_, new_n11454_, new_n2121_ );
or   ( new_n11456_, new_n11455_, new_n11451_ );
and  ( new_n11457_, new_n11456_, new_n11450_ );
or   ( new_n11458_, new_n5604_, new_n1318_ );
or   ( new_n11459_, new_n5606_, new_n1213_ );
and  ( new_n11460_, new_n11459_, new_n11458_ );
xor  ( new_n11461_, new_n11460_, new_n5206_ );
or   ( new_n11462_, new_n5207_, new_n1523_ );
or   ( new_n11463_, new_n5209_, new_n1525_ );
and  ( new_n11464_, new_n11463_, new_n11462_ );
xor  ( new_n11465_, new_n11464_, new_n4708_ );
or   ( new_n11466_, new_n11465_, new_n11461_ );
and  ( new_n11467_, new_n11465_, new_n11461_ );
or   ( new_n11468_, new_n4709_, new_n1899_ );
or   ( new_n11469_, new_n4711_, new_n1754_ );
and  ( new_n11470_, new_n11469_, new_n11468_ );
xor  ( new_n11471_, new_n11470_, new_n4295_ );
or   ( new_n11472_, new_n11471_, new_n11467_ );
and  ( new_n11473_, new_n11472_, new_n11466_ );
or   ( new_n11474_, new_n11473_, new_n11457_ );
and  ( new_n11475_, new_n11473_, new_n11457_ );
or   ( new_n11476_, new_n4302_, new_n2178_ );
or   ( new_n11477_, new_n4304_, new_n2057_ );
and  ( new_n11478_, new_n11477_, new_n11476_ );
xor  ( new_n11479_, new_n11478_, new_n3895_ );
or   ( new_n11480_, new_n3896_, new_n2475_ );
or   ( new_n11481_, new_n3898_, new_n2291_ );
and  ( new_n11482_, new_n11481_, new_n11480_ );
xor  ( new_n11483_, new_n11482_, new_n3460_ );
nor  ( new_n11484_, new_n11483_, new_n11479_ );
and  ( new_n11485_, new_n11483_, new_n11479_ );
or   ( new_n11486_, new_n3461_, new_n2751_ );
or   ( new_n11487_, new_n3463_, new_n2646_ );
and  ( new_n11488_, new_n11487_, new_n11486_ );
xor  ( new_n11489_, new_n11488_, new_n3116_ );
nor  ( new_n11490_, new_n11489_, new_n11485_ );
nor  ( new_n11491_, new_n11490_, new_n11484_ );
or   ( new_n11492_, new_n11491_, new_n11475_ );
and  ( new_n11493_, new_n11492_, new_n11474_ );
and  ( new_n11494_, new_n11440_, new_n11388_ );
or   ( new_n11495_, new_n11494_, new_n11493_ );
and  ( new_n11496_, new_n11495_, new_n11441_ );
or   ( new_n11497_, new_n11496_, new_n11334_ );
and  ( new_n11498_, new_n11496_, new_n11334_ );
xor  ( new_n11499_, new_n10945_, new_n10943_ );
xor  ( new_n11500_, new_n11499_, new_n10949_ );
xnor ( new_n11501_, new_n11085_, new_n11081_ );
xor  ( new_n11502_, new_n11501_, new_n11091_ );
xor  ( new_n11503_, new_n11103_, new_n11097_ );
xor  ( new_n11504_, new_n11503_, new_n263_ );
or   ( new_n11505_, new_n11504_, new_n11502_ );
and  ( new_n11506_, new_n11504_, new_n11502_ );
xnor ( new_n11507_, new_n11115_, new_n11111_ );
xor  ( new_n11508_, new_n11507_, new_n11121_ );
or   ( new_n11509_, new_n11508_, new_n11506_ );
and  ( new_n11510_, new_n11509_, new_n11505_ );
nor  ( new_n11511_, new_n11510_, new_n11500_ );
nand ( new_n11512_, new_n11510_, new_n11500_ );
xor  ( new_n11513_, new_n10940_, new_n10938_ );
and  ( new_n11514_, new_n11513_, new_n11512_ );
or   ( new_n11515_, new_n11514_, new_n11511_ );
or   ( new_n11516_, new_n11515_, new_n11498_ );
and  ( new_n11517_, new_n11516_, new_n11497_ );
or   ( new_n11518_, new_n11517_, new_n11284_ );
nand ( new_n11519_, new_n11517_, new_n11284_ );
xor  ( new_n11520_, new_n10928_, new_n10926_ );
xor  ( new_n11521_, new_n11520_, new_n10932_ );
xor  ( new_n11522_, new_n10914_, new_n10912_ );
xor  ( new_n11523_, new_n11522_, new_n10918_ );
nor  ( new_n11524_, new_n11523_, new_n11521_ );
and  ( new_n11525_, new_n11523_, new_n11521_ );
xor  ( new_n11526_, new_n10951_, new_n10941_ );
xor  ( new_n11527_, new_n11526_, new_n10954_ );
not  ( new_n11528_, new_n11527_ );
nor  ( new_n11529_, new_n11528_, new_n11525_ );
nor  ( new_n11530_, new_n11529_, new_n11524_ );
nand ( new_n11531_, new_n11530_, new_n11519_ );
and  ( new_n11532_, new_n11531_, new_n11518_ );
or   ( new_n11533_, new_n11532_, new_n11258_ );
and  ( new_n11534_, new_n11532_, new_n11258_ );
xor  ( new_n11535_, new_n10630_, new_n10628_ );
xnor ( new_n11536_, new_n11535_, new_n10643_ );
or   ( new_n11537_, new_n11536_, new_n11534_ );
and  ( new_n11538_, new_n11537_, new_n11533_ );
nand ( new_n11539_, new_n11538_, new_n11248_ );
nor  ( new_n11540_, new_n11538_, new_n11248_ );
xor  ( new_n11541_, new_n10611_, new_n10609_ );
xor  ( new_n11542_, new_n11541_, new_n10615_ );
or   ( new_n11543_, new_n11542_, new_n11540_ );
and  ( new_n11544_, new_n11543_, new_n11539_ );
or   ( new_n11545_, new_n11544_, new_n11238_ );
and  ( new_n11546_, new_n11544_, new_n11238_ );
xnor ( new_n11547_, new_n11218_, new_n11216_ );
xor  ( new_n11548_, new_n11547_, new_n11221_ );
or   ( new_n11549_, new_n11548_, new_n11546_ );
and  ( new_n11550_, new_n11549_, new_n11545_ );
nor  ( new_n11551_, new_n11550_, new_n11233_ );
xor  ( new_n11552_, new_n11544_, new_n11238_ );
xor  ( new_n11553_, new_n11552_, new_n11548_ );
xor  ( new_n11554_, new_n11538_, new_n11248_ );
xor  ( new_n11555_, new_n11554_, new_n11542_ );
xnor ( new_n11556_, new_n11532_, new_n11258_ );
xor  ( new_n11557_, new_n11556_, new_n11536_ );
xor  ( new_n11558_, new_n11523_, new_n11521_ );
xor  ( new_n11559_, new_n11558_, new_n11528_ );
xnor ( new_n11560_, new_n11006_, new_n10966_ );
xor  ( new_n11561_, new_n11560_, new_n11021_ );
or   ( new_n11562_, new_n11561_, new_n11559_ );
and  ( new_n11563_, new_n11561_, new_n11559_ );
xor  ( new_n11564_, new_n11127_, new_n11077_ );
xnor ( new_n11565_, new_n11564_, new_n11180_ );
or   ( new_n11566_, new_n11565_, new_n11563_ );
and  ( new_n11567_, new_n11566_, new_n11562_ );
xor  ( new_n11568_, new_n11440_, new_n11388_ );
xor  ( new_n11569_, new_n11568_, new_n11493_ );
xor  ( new_n11570_, new_n11319_, new_n11295_ );
xor  ( new_n11571_, new_n11570_, new_n11332_ );
nor  ( new_n11572_, new_n11571_, new_n11569_ );
nand ( new_n11573_, new_n11571_, new_n11569_ );
xnor ( new_n11574_, new_n11510_, new_n11500_ );
xor  ( new_n11575_, new_n11574_, new_n11513_ );
and  ( new_n11576_, new_n11575_, new_n11573_ );
or   ( new_n11577_, new_n11576_, new_n11572_ );
xnor ( new_n11578_, new_n11272_, new_n11270_ );
xor  ( new_n11579_, new_n11578_, new_n11276_ );
xnor ( new_n11580_, new_n11262_, new_n11260_ );
xor  ( new_n11581_, new_n11580_, new_n11266_ );
nand ( new_n11582_, new_n11581_, new_n11579_ );
nor  ( new_n11583_, new_n11581_, new_n11579_ );
xnor ( new_n11584_, new_n11420_, new_n11404_ );
xor  ( new_n11585_, new_n11584_, new_n11438_ );
xor  ( new_n11586_, new_n11313_, new_n11297_ );
xor  ( new_n11587_, new_n11586_, new_n11317_ );
nor  ( new_n11588_, new_n11587_, new_n11585_ );
and  ( new_n11589_, new_n11587_, new_n11585_ );
xor  ( new_n11590_, new_n11325_, new_n11323_ );
xor  ( new_n11591_, new_n11590_, new_n11330_ );
not  ( new_n11592_, new_n11591_ );
nor  ( new_n11593_, new_n11592_, new_n11589_ );
nor  ( new_n11594_, new_n11593_, new_n11588_ );
or   ( new_n11595_, new_n11594_, new_n11583_ );
and  ( new_n11596_, new_n11595_, new_n11582_ );
or   ( new_n11597_, new_n11596_, new_n11577_ );
and  ( new_n11598_, new_n11596_, new_n11577_ );
or   ( new_n11599_, new_n283_, new_n10541_ );
or   ( new_n11600_, new_n286_, new_n10220_ );
and  ( new_n11601_, new_n11600_, new_n11599_ );
xor  ( new_n11602_, new_n11601_, new_n278_ );
and  ( new_n11603_, new_n295_, RIbb31578_128 );
or   ( new_n11604_, new_n11603_, new_n292_ );
nand ( new_n11605_, new_n11603_, RIbb2f520_3 );
and  ( new_n11606_, new_n11605_, new_n11604_ );
and  ( new_n11607_, new_n11606_, new_n11602_ );
or   ( new_n11608_, new_n299_, new_n10841_ );
or   ( new_n11609_, new_n302_, new_n10541_ );
and  ( new_n11610_, new_n11609_, new_n11608_ );
xor  ( new_n11611_, new_n11610_, new_n293_ );
nor  ( new_n11612_, new_n11611_, new_n11607_ );
nand ( new_n11613_, new_n11611_, new_n11607_ );
or   ( new_n11614_, new_n409_, new_n8481_ );
or   ( new_n11615_, new_n411_, new_n8352_ );
and  ( new_n11616_, new_n11615_, new_n11614_ );
xor  ( new_n11617_, new_n11616_, new_n328_ );
or   ( new_n11618_, new_n337_, new_n9099_ );
or   ( new_n11619_, new_n340_, new_n8995_ );
and  ( new_n11620_, new_n11619_, new_n11618_ );
xor  ( new_n11621_, new_n11620_, new_n332_ );
nor  ( new_n11622_, new_n11621_, new_n11617_ );
and  ( new_n11623_, new_n11621_, new_n11617_ );
or   ( new_n11624_, new_n317_, new_n9679_ );
or   ( new_n11625_, new_n320_, new_n9681_ );
and  ( new_n11626_, new_n11625_, new_n11624_ );
xor  ( new_n11627_, new_n11626_, new_n312_ );
nor  ( new_n11628_, new_n11627_, new_n11623_ );
or   ( new_n11629_, new_n11628_, new_n11622_ );
and  ( new_n11630_, new_n11629_, new_n11613_ );
or   ( new_n11631_, new_n11630_, new_n11612_ );
xnor ( new_n11632_, new_n11430_, new_n11426_ );
xor  ( new_n11633_, new_n11632_, new_n11436_ );
xnor ( new_n11634_, new_n11449_, new_n11445_ );
xor  ( new_n11635_, new_n11634_, new_n11455_ );
or   ( new_n11636_, new_n11635_, new_n11633_ );
and  ( new_n11637_, new_n11635_, new_n11633_ );
xor  ( new_n11638_, new_n11483_, new_n11479_ );
xnor ( new_n11639_, new_n11638_, new_n11489_ );
or   ( new_n11640_, new_n11639_, new_n11637_ );
and  ( new_n11641_, new_n11640_, new_n11636_ );
nor  ( new_n11642_, new_n11641_, new_n11631_ );
nand ( new_n11643_, new_n11641_, new_n11631_ );
xnor ( new_n11644_, new_n11412_, new_n11408_ );
xor  ( new_n11645_, new_n11644_, new_n11418_ );
xnor ( new_n11646_, new_n11396_, new_n11392_ );
xor  ( new_n11647_, new_n11646_, new_n11402_ );
nor  ( new_n11648_, new_n11647_, new_n11645_ );
and  ( new_n11649_, new_n11647_, new_n11645_ );
xor  ( new_n11650_, new_n11305_, new_n11301_ );
xnor ( new_n11651_, new_n11650_, new_n11311_ );
nor  ( new_n11652_, new_n11651_, new_n11649_ );
or   ( new_n11653_, new_n11652_, new_n11648_ );
and  ( new_n11654_, new_n11653_, new_n11643_ );
or   ( new_n11655_, new_n11654_, new_n11642_ );
or   ( new_n11656_, new_n2425_, new_n4069_ );
or   ( new_n11657_, new_n2427_, new_n3820_ );
and  ( new_n11658_, new_n11657_, new_n11656_ );
xor  ( new_n11659_, new_n11658_, new_n2121_ );
or   ( new_n11660_, new_n2122_, new_n4603_ );
or   ( new_n11661_, new_n2124_, new_n4267_ );
and  ( new_n11662_, new_n11661_, new_n11660_ );
xor  ( new_n11663_, new_n11662_, new_n1843_ );
or   ( new_n11664_, new_n11663_, new_n11659_ );
and  ( new_n11665_, new_n11663_, new_n11659_ );
or   ( new_n11666_, new_n1844_, new_n4859_ );
or   ( new_n11667_, new_n1846_, new_n4995_ );
and  ( new_n11668_, new_n11667_, new_n11666_ );
xor  ( new_n11669_, new_n11668_, new_n1586_ );
or   ( new_n11670_, new_n11669_, new_n11665_ );
and  ( new_n11671_, new_n11670_, new_n11664_ );
or   ( new_n11672_, new_n897_, new_n6943_ );
or   ( new_n11673_, new_n899_, new_n6589_ );
and  ( new_n11674_, new_n11673_, new_n11672_ );
xor  ( new_n11675_, new_n11674_, new_n748_ );
or   ( new_n11676_, new_n755_, new_n7373_ );
or   ( new_n11677_, new_n757_, new_n7149_ );
and  ( new_n11678_, new_n11677_, new_n11676_ );
xor  ( new_n11679_, new_n11678_, new_n523_ );
or   ( new_n11680_, new_n11679_, new_n11675_ );
and  ( new_n11681_, new_n11679_, new_n11675_ );
or   ( new_n11682_, new_n524_, new_n8115_ );
or   ( new_n11683_, new_n526_, new_n8117_ );
and  ( new_n11684_, new_n11683_, new_n11682_ );
xor  ( new_n11685_, new_n11684_, new_n403_ );
or   ( new_n11686_, new_n11685_, new_n11681_ );
and  ( new_n11687_, new_n11686_, new_n11680_ );
or   ( new_n11688_, new_n11687_, new_n11671_ );
and  ( new_n11689_, new_n11687_, new_n11671_ );
or   ( new_n11690_, new_n1593_, new_n5428_ );
or   ( new_n11691_, new_n1595_, new_n5171_ );
and  ( new_n11692_, new_n11691_, new_n11690_ );
xor  ( new_n11693_, new_n11692_, new_n1358_ );
or   ( new_n11694_, new_n1364_, new_n5899_ );
or   ( new_n11695_, new_n1366_, new_n5570_ );
and  ( new_n11696_, new_n11695_, new_n11694_ );
xor  ( new_n11697_, new_n11696_, new_n1129_ );
or   ( new_n11698_, new_n11697_, new_n11693_ );
and  ( new_n11699_, new_n11697_, new_n11693_ );
or   ( new_n11700_, new_n1135_, new_n6425_ );
or   ( new_n11701_, new_n1137_, new_n6219_ );
and  ( new_n11702_, new_n11701_, new_n11700_ );
xor  ( new_n11703_, new_n11702_, new_n896_ );
or   ( new_n11704_, new_n11703_, new_n11699_ );
and  ( new_n11705_, new_n11704_, new_n11698_ );
or   ( new_n11706_, new_n11705_, new_n11689_ );
and  ( new_n11707_, new_n11706_, new_n11688_ );
or   ( new_n11708_, new_n7732_, new_n515_ );
or   ( new_n11709_, new_n7734_, new_n509_ );
and  ( new_n11710_, new_n11709_, new_n11708_ );
xor  ( new_n11711_, new_n11710_, new_n7177_ );
or   ( new_n11712_, new_n7184_, new_n805_ );
or   ( new_n11713_, new_n7186_, new_n775_ );
and  ( new_n11714_, new_n11713_, new_n11712_ );
xor  ( new_n11715_, new_n11714_, new_n6638_ );
nor  ( new_n11716_, new_n11715_, new_n11711_ );
and  ( new_n11717_, new_n11715_, new_n11711_ );
or   ( new_n11718_, new_n6645_, new_n986_ );
or   ( new_n11719_, new_n6647_, new_n886_ );
and  ( new_n11720_, new_n11719_, new_n11718_ );
xor  ( new_n11721_, new_n11720_, new_n6166_ );
nor  ( new_n11722_, new_n11721_, new_n11717_ );
nor  ( new_n11723_, new_n11722_, new_n11716_ );
or   ( new_n11724_, new_n10059_, new_n301_ );
or   ( new_n11725_, new_n10061_, new_n279_ );
and  ( new_n11726_, new_n11725_, new_n11724_ );
xor  ( new_n11727_, new_n11726_, new_n9421_ );
and  ( new_n11728_, RIbb2d888_64, RIbb2d6a8_68 );
or   ( new_n11729_, RIbb2d888_64, new_n285_ );
and  ( new_n11730_, new_n11729_, RIbb2d900_63 );
or   ( new_n11731_, new_n11730_, new_n11728_ );
or   ( new_n11732_, new_n10770_, new_n313_ );
and  ( new_n11733_, new_n11732_, new_n11731_ );
nor  ( new_n11734_, new_n11733_, new_n11727_ );
and  ( new_n11735_, new_n11733_, new_n11727_ );
nor  ( new_n11736_, new_n11735_, new_n292_ );
nor  ( new_n11737_, new_n11736_, new_n11734_ );
or   ( new_n11738_, new_n9422_, new_n270_ );
or   ( new_n11739_, new_n9424_, new_n294_ );
and  ( new_n11740_, new_n11739_, new_n11738_ );
xor  ( new_n11741_, new_n11740_, new_n8873_ );
or   ( new_n11742_, new_n8874_, new_n348_ );
or   ( new_n11743_, new_n8876_, new_n264_ );
and  ( new_n11744_, new_n11743_, new_n11742_ );
xor  ( new_n11745_, new_n11744_, new_n8257_ );
or   ( new_n11746_, new_n11745_, new_n11741_ );
and  ( new_n11747_, new_n11745_, new_n11741_ );
or   ( new_n11748_, new_n8264_, new_n443_ );
or   ( new_n11749_, new_n8266_, new_n419_ );
and  ( new_n11750_, new_n11749_, new_n11748_ );
xor  ( new_n11751_, new_n11750_, new_n7725_ );
or   ( new_n11752_, new_n11751_, new_n11747_ );
and  ( new_n11753_, new_n11752_, new_n11746_ );
and  ( new_n11754_, new_n11753_, new_n11737_ );
or   ( new_n11755_, new_n11754_, new_n11723_ );
or   ( new_n11756_, new_n11753_, new_n11737_ );
and  ( new_n11757_, new_n11756_, new_n11755_ );
or   ( new_n11758_, new_n11757_, new_n11707_ );
or   ( new_n11759_, new_n4709_, new_n2057_ );
or   ( new_n11760_, new_n4711_, new_n1899_ );
and  ( new_n11761_, new_n11760_, new_n11759_ );
xor  ( new_n11762_, new_n11761_, new_n4295_ );
or   ( new_n11763_, new_n4302_, new_n2291_ );
or   ( new_n11764_, new_n4304_, new_n2178_ );
and  ( new_n11765_, new_n11764_, new_n11763_ );
xor  ( new_n11766_, new_n11765_, new_n3895_ );
or   ( new_n11767_, new_n11766_, new_n11762_ );
and  ( new_n11768_, new_n11766_, new_n11762_ );
or   ( new_n11769_, new_n3896_, new_n2646_ );
or   ( new_n11770_, new_n3898_, new_n2475_ );
and  ( new_n11771_, new_n11770_, new_n11769_ );
xor  ( new_n11772_, new_n11771_, new_n3460_ );
or   ( new_n11773_, new_n11772_, new_n11768_ );
and  ( new_n11774_, new_n11773_, new_n11767_ );
or   ( new_n11775_, new_n6173_, new_n1213_ );
or   ( new_n11776_, new_n6175_, new_n1168_ );
and  ( new_n11777_, new_n11776_, new_n11775_ );
xor  ( new_n11778_, new_n11777_, new_n5597_ );
or   ( new_n11779_, new_n5604_, new_n1525_ );
or   ( new_n11780_, new_n5606_, new_n1318_ );
and  ( new_n11781_, new_n11780_, new_n11779_ );
xor  ( new_n11782_, new_n11781_, new_n5206_ );
or   ( new_n11783_, new_n11782_, new_n11778_ );
and  ( new_n11784_, new_n11782_, new_n11778_ );
or   ( new_n11785_, new_n5207_, new_n1754_ );
or   ( new_n11786_, new_n5209_, new_n1523_ );
and  ( new_n11787_, new_n11786_, new_n11785_ );
xor  ( new_n11788_, new_n11787_, new_n4708_ );
or   ( new_n11789_, new_n11788_, new_n11784_ );
and  ( new_n11790_, new_n11789_, new_n11783_ );
or   ( new_n11791_, new_n11790_, new_n11774_ );
and  ( new_n11792_, new_n11790_, new_n11774_ );
or   ( new_n11793_, new_n3461_, new_n2981_ );
or   ( new_n11794_, new_n3463_, new_n2751_ );
and  ( new_n11795_, new_n11794_, new_n11793_ );
xor  ( new_n11796_, new_n11795_, new_n3116_ );
or   ( new_n11797_, new_n3117_, new_n3306_ );
or   ( new_n11798_, new_n3119_, new_n3178_ );
and  ( new_n11799_, new_n11798_, new_n11797_ );
xor  ( new_n11800_, new_n11799_, new_n2800_ );
nor  ( new_n11801_, new_n11800_, new_n11796_ );
and  ( new_n11802_, new_n11800_, new_n11796_ );
or   ( new_n11803_, new_n2807_, new_n3694_ );
or   ( new_n11804_, new_n2809_, new_n3696_ );
and  ( new_n11805_, new_n11804_, new_n11803_ );
xor  ( new_n11806_, new_n11805_, new_n2424_ );
nor  ( new_n11807_, new_n11806_, new_n11802_ );
nor  ( new_n11808_, new_n11807_, new_n11801_ );
or   ( new_n11809_, new_n11808_, new_n11792_ );
and  ( new_n11810_, new_n11809_, new_n11791_ );
and  ( new_n11811_, new_n11757_, new_n11707_ );
or   ( new_n11812_, new_n11811_, new_n11810_ );
and  ( new_n11813_, new_n11812_, new_n11758_ );
and  ( new_n11814_, new_n11813_, new_n11655_ );
nor  ( new_n11815_, new_n11813_, new_n11655_ );
xor  ( new_n11816_, new_n11504_, new_n11502_ );
xor  ( new_n11817_, new_n11816_, new_n11508_ );
xnor ( new_n11818_, new_n11360_, new_n11356_ );
xor  ( new_n11819_, new_n11818_, new_n11366_ );
xnor ( new_n11820_, new_n11465_, new_n11461_ );
xor  ( new_n11821_, new_n11820_, new_n11471_ );
or   ( new_n11822_, new_n11821_, new_n11819_ );
and  ( new_n11823_, new_n11821_, new_n11819_ );
xor  ( new_n11824_, new_n11378_, new_n11374_ );
xnor ( new_n11825_, new_n11824_, new_n11384_ );
or   ( new_n11826_, new_n11825_, new_n11823_ );
and  ( new_n11827_, new_n11826_, new_n11822_ );
nor  ( new_n11828_, new_n11827_, new_n11817_ );
and  ( new_n11829_, new_n11827_, new_n11817_ );
xor  ( new_n11830_, new_n11288_, new_n11286_ );
xor  ( new_n11831_, new_n11830_, new_n11293_ );
not  ( new_n11832_, new_n11831_ );
nor  ( new_n11833_, new_n11832_, new_n11829_ );
nor  ( new_n11834_, new_n11833_, new_n11828_ );
nor  ( new_n11835_, new_n11834_, new_n11815_ );
nor  ( new_n11836_, new_n11835_, new_n11814_ );
or   ( new_n11837_, new_n11836_, new_n11598_ );
and  ( new_n11838_, new_n11837_, new_n11597_ );
or   ( new_n11839_, new_n11838_, new_n11567_ );
and  ( new_n11840_, new_n11838_, new_n11567_ );
xor  ( new_n11841_, new_n11023_, new_n10956_ );
xnor ( new_n11842_, new_n11841_, new_n11183_ );
or   ( new_n11843_, new_n11842_, new_n11840_ );
and  ( new_n11844_, new_n11843_, new_n11839_ );
or   ( new_n11845_, new_n11844_, new_n11557_ );
and  ( new_n11846_, new_n11844_, new_n11557_ );
xor  ( new_n11847_, new_n11242_, new_n11240_ );
xor  ( new_n11848_, new_n11847_, new_n11246_ );
or   ( new_n11849_, new_n11848_, new_n11846_ );
and  ( new_n11850_, new_n11849_, new_n11845_ );
or   ( new_n11851_, new_n11850_, new_n11555_ );
and  ( new_n11852_, new_n11850_, new_n11555_ );
xnor ( new_n11853_, new_n11237_, new_n11235_ );
or   ( new_n11854_, new_n11853_, new_n11852_ );
and  ( new_n11855_, new_n11854_, new_n11851_ );
nor  ( new_n11856_, new_n11855_, new_n11553_ );
xor  ( new_n11857_, new_n11850_, new_n11555_ );
xor  ( new_n11858_, new_n11857_, new_n11853_ );
xor  ( new_n11859_, new_n11517_, new_n11284_ );
xor  ( new_n11860_, new_n11859_, new_n11530_ );
not  ( new_n11861_, new_n11860_ );
xnor ( new_n11862_, new_n11838_, new_n11567_ );
xor  ( new_n11863_, new_n11862_, new_n11842_ );
nand ( new_n11864_, new_n11863_, new_n11861_ );
xnor ( new_n11865_, new_n11252_, new_n11250_ );
xor  ( new_n11866_, new_n11865_, new_n11256_ );
xor  ( new_n11867_, new_n11496_, new_n11334_ );
xor  ( new_n11868_, new_n11867_, new_n11515_ );
xnor ( new_n11869_, new_n11596_, new_n11577_ );
xor  ( new_n11870_, new_n11869_, new_n11836_ );
nand ( new_n11871_, new_n11870_, new_n11868_ );
or   ( new_n11872_, new_n11870_, new_n11868_ );
xor  ( new_n11873_, new_n11561_, new_n11559_ );
xnor ( new_n11874_, new_n11873_, new_n11565_ );
nand ( new_n11875_, new_n11874_, new_n11872_ );
and  ( new_n11876_, new_n11875_, new_n11871_ );
or   ( new_n11877_, new_n11876_, new_n11866_ );
and  ( new_n11878_, new_n11876_, new_n11866_ );
xor  ( new_n11879_, new_n11278_, new_n11268_ );
xor  ( new_n11880_, new_n11879_, new_n11282_ );
xnor ( new_n11881_, new_n11581_, new_n11579_ );
xor  ( new_n11882_, new_n11881_, new_n11594_ );
xnor ( new_n11883_, new_n11813_, new_n11655_ );
xor  ( new_n11884_, new_n11883_, new_n11834_ );
nand ( new_n11885_, new_n11884_, new_n11882_ );
nor  ( new_n11886_, new_n11884_, new_n11882_ );
xor  ( new_n11887_, new_n11571_, new_n11569_ );
xor  ( new_n11888_, new_n11887_, new_n11575_ );
or   ( new_n11889_, new_n11888_, new_n11886_ );
and  ( new_n11890_, new_n11889_, new_n11885_ );
or   ( new_n11891_, new_n11890_, new_n11880_ );
and  ( new_n11892_, new_n11890_, new_n11880_ );
xor  ( new_n11893_, new_n11687_, new_n11671_ );
xor  ( new_n11894_, new_n11893_, new_n11705_ );
xor  ( new_n11895_, new_n11753_, new_n11737_ );
xor  ( new_n11896_, new_n11895_, new_n11723_ );
and  ( new_n11897_, new_n11896_, new_n11894_ );
nor  ( new_n11898_, new_n11896_, new_n11894_ );
xor  ( new_n11899_, new_n11790_, new_n11774_ );
xnor ( new_n11900_, new_n11899_, new_n11808_ );
nor  ( new_n11901_, new_n11900_, new_n11898_ );
or   ( new_n11902_, new_n11901_, new_n11897_ );
xor  ( new_n11903_, new_n11647_, new_n11645_ );
xor  ( new_n11904_, new_n11903_, new_n11651_ );
xor  ( new_n11905_, new_n11611_, new_n11607_ );
xor  ( new_n11906_, new_n11905_, new_n11629_ );
nand ( new_n11907_, new_n11906_, new_n11904_ );
nor  ( new_n11908_, new_n11906_, new_n11904_ );
xor  ( new_n11909_, new_n11635_, new_n11633_ );
xnor ( new_n11910_, new_n11909_, new_n11639_ );
or   ( new_n11911_, new_n11910_, new_n11908_ );
and  ( new_n11912_, new_n11911_, new_n11907_ );
nand ( new_n11913_, new_n11912_, new_n11902_ );
nor  ( new_n11914_, new_n11912_, new_n11902_ );
xor  ( new_n11915_, new_n11473_, new_n11457_ );
xnor ( new_n11916_, new_n11915_, new_n11491_ );
or   ( new_n11917_, new_n11916_, new_n11914_ );
and  ( new_n11918_, new_n11917_, new_n11913_ );
xnor ( new_n11919_, new_n11368_, new_n11352_ );
xor  ( new_n11920_, new_n11919_, new_n11386_ );
xor  ( new_n11921_, new_n11587_, new_n11585_ );
xor  ( new_n11922_, new_n11921_, new_n11592_ );
or   ( new_n11923_, new_n11922_, new_n11920_ );
and  ( new_n11924_, new_n11922_, new_n11920_ );
xor  ( new_n11925_, new_n11827_, new_n11817_ );
xor  ( new_n11926_, new_n11925_, new_n11832_ );
or   ( new_n11927_, new_n11926_, new_n11924_ );
and  ( new_n11928_, new_n11927_, new_n11923_ );
or   ( new_n11929_, new_n11928_, new_n11918_ );
and  ( new_n11930_, new_n11928_, new_n11918_ );
xnor ( new_n11931_, new_n11344_, new_n11338_ );
xor  ( new_n11932_, new_n11931_, new_n11350_ );
xnor ( new_n11933_, new_n11715_, new_n11711_ );
xor  ( new_n11934_, new_n11933_, new_n11721_ );
xnor ( new_n11935_, new_n11745_, new_n11741_ );
xor  ( new_n11936_, new_n11935_, new_n11751_ );
or   ( new_n11937_, new_n11936_, new_n11934_ );
and  ( new_n11938_, new_n11936_, new_n11934_ );
xor  ( new_n11939_, new_n11733_, new_n11727_ );
xor  ( new_n11940_, new_n11939_, new_n293_ );
or   ( new_n11941_, new_n11940_, new_n11938_ );
and  ( new_n11942_, new_n11941_, new_n11937_ );
nor  ( new_n11943_, new_n11942_, new_n11932_ );
nand ( new_n11944_, new_n11942_, new_n11932_ );
xor  ( new_n11945_, new_n11821_, new_n11819_ );
xnor ( new_n11946_, new_n11945_, new_n11825_ );
and  ( new_n11947_, new_n11946_, new_n11944_ );
or   ( new_n11948_, new_n11947_, new_n11943_ );
or   ( new_n11949_, new_n5604_, new_n1523_ );
or   ( new_n11950_, new_n5606_, new_n1525_ );
and  ( new_n11951_, new_n11950_, new_n11949_ );
xor  ( new_n11952_, new_n11951_, new_n5206_ );
or   ( new_n11953_, new_n5207_, new_n1899_ );
or   ( new_n11954_, new_n5209_, new_n1754_ );
and  ( new_n11955_, new_n11954_, new_n11953_ );
xor  ( new_n11956_, new_n11955_, new_n4708_ );
or   ( new_n11957_, new_n11956_, new_n11952_ );
and  ( new_n11958_, new_n11956_, new_n11952_ );
or   ( new_n11959_, new_n4709_, new_n2178_ );
or   ( new_n11960_, new_n4711_, new_n2057_ );
and  ( new_n11961_, new_n11960_, new_n11959_ );
xor  ( new_n11962_, new_n11961_, new_n4295_ );
or   ( new_n11963_, new_n11962_, new_n11958_ );
and  ( new_n11964_, new_n11963_, new_n11957_ );
or   ( new_n11965_, new_n3117_, new_n3696_ );
or   ( new_n11966_, new_n3119_, new_n3306_ );
and  ( new_n11967_, new_n11966_, new_n11965_ );
xor  ( new_n11968_, new_n11967_, new_n2800_ );
or   ( new_n11969_, new_n2807_, new_n3820_ );
or   ( new_n11970_, new_n2809_, new_n3694_ );
and  ( new_n11971_, new_n11970_, new_n11969_ );
xor  ( new_n11972_, new_n11971_, new_n2424_ );
or   ( new_n11973_, new_n11972_, new_n11968_ );
and  ( new_n11974_, new_n11972_, new_n11968_ );
or   ( new_n11975_, new_n2425_, new_n4267_ );
or   ( new_n11976_, new_n2427_, new_n4069_ );
and  ( new_n11977_, new_n11976_, new_n11975_ );
xor  ( new_n11978_, new_n11977_, new_n2121_ );
or   ( new_n11979_, new_n11978_, new_n11974_ );
and  ( new_n11980_, new_n11979_, new_n11973_ );
or   ( new_n11981_, new_n11980_, new_n11964_ );
and  ( new_n11982_, new_n11980_, new_n11964_ );
or   ( new_n11983_, new_n4302_, new_n2475_ );
or   ( new_n11984_, new_n4304_, new_n2291_ );
and  ( new_n11985_, new_n11984_, new_n11983_ );
xor  ( new_n11986_, new_n11985_, new_n3895_ );
or   ( new_n11987_, new_n3896_, new_n2751_ );
or   ( new_n11988_, new_n3898_, new_n2646_ );
and  ( new_n11989_, new_n11988_, new_n11987_ );
xor  ( new_n11990_, new_n11989_, new_n3460_ );
nor  ( new_n11991_, new_n11990_, new_n11986_ );
and  ( new_n11992_, new_n11990_, new_n11986_ );
or   ( new_n11993_, new_n3461_, new_n3178_ );
or   ( new_n11994_, new_n3463_, new_n2981_ );
and  ( new_n11995_, new_n11994_, new_n11993_ );
xor  ( new_n11996_, new_n11995_, new_n3116_ );
nor  ( new_n11997_, new_n11996_, new_n11992_ );
nor  ( new_n11998_, new_n11997_, new_n11991_ );
or   ( new_n11999_, new_n11998_, new_n11982_ );
and  ( new_n12000_, new_n11999_, new_n11981_ );
or   ( new_n12001_, new_n10059_, new_n294_ );
or   ( new_n12002_, new_n10061_, new_n301_ );
and  ( new_n12003_, new_n12002_, new_n12001_ );
xor  ( new_n12004_, new_n12003_, new_n9421_ );
and  ( new_n12005_, RIbb2d888_64, RIbb2d630_69 );
or   ( new_n12006_, RIbb2d888_64, new_n279_ );
and  ( new_n12007_, new_n12006_, RIbb2d900_63 );
or   ( new_n12008_, new_n12007_, new_n12005_ );
or   ( new_n12009_, new_n10770_, new_n285_ );
and  ( new_n12010_, new_n12009_, new_n12008_ );
or   ( new_n12011_, new_n12010_, new_n12004_ );
and  ( new_n12012_, new_n12010_, new_n12004_ );
or   ( new_n12013_, new_n9422_, new_n264_ );
or   ( new_n12014_, new_n9424_, new_n270_ );
and  ( new_n12015_, new_n12014_, new_n12013_ );
xor  ( new_n12016_, new_n12015_, new_n8873_ );
or   ( new_n12017_, new_n12016_, new_n12012_ );
and  ( new_n12018_, new_n12017_, new_n12011_ );
or   ( new_n12019_, new_n7184_, new_n886_ );
or   ( new_n12020_, new_n7186_, new_n805_ );
and  ( new_n12021_, new_n12020_, new_n12019_ );
xor  ( new_n12022_, new_n12021_, new_n6638_ );
or   ( new_n12023_, new_n6645_, new_n1168_ );
or   ( new_n12024_, new_n6647_, new_n986_ );
and  ( new_n12025_, new_n12024_, new_n12023_ );
xor  ( new_n12026_, new_n12025_, new_n6166_ );
or   ( new_n12027_, new_n12026_, new_n12022_ );
and  ( new_n12028_, new_n12026_, new_n12022_ );
or   ( new_n12029_, new_n6173_, new_n1318_ );
or   ( new_n12030_, new_n6175_, new_n1213_ );
and  ( new_n12031_, new_n12030_, new_n12029_ );
xor  ( new_n12032_, new_n12031_, new_n5597_ );
or   ( new_n12033_, new_n12032_, new_n12028_ );
and  ( new_n12034_, new_n12033_, new_n12027_ );
or   ( new_n12035_, new_n12034_, new_n12018_ );
and  ( new_n12036_, new_n12034_, new_n12018_ );
or   ( new_n12037_, new_n8874_, new_n419_ );
or   ( new_n12038_, new_n8876_, new_n348_ );
and  ( new_n12039_, new_n12038_, new_n12037_ );
xor  ( new_n12040_, new_n12039_, new_n8257_ );
or   ( new_n12041_, new_n8264_, new_n509_ );
or   ( new_n12042_, new_n8266_, new_n443_ );
and  ( new_n12043_, new_n12042_, new_n12041_ );
xor  ( new_n12044_, new_n12043_, new_n7725_ );
nor  ( new_n12045_, new_n12044_, new_n12040_ );
and  ( new_n12046_, new_n12044_, new_n12040_ );
or   ( new_n12047_, new_n7732_, new_n775_ );
or   ( new_n12048_, new_n7734_, new_n515_ );
and  ( new_n12049_, new_n12048_, new_n12047_ );
xor  ( new_n12050_, new_n12049_, new_n7177_ );
nor  ( new_n12051_, new_n12050_, new_n12046_ );
nor  ( new_n12052_, new_n12051_, new_n12045_ );
or   ( new_n12053_, new_n12052_, new_n12036_ );
and  ( new_n12054_, new_n12053_, new_n12035_ );
or   ( new_n12055_, new_n12054_, new_n12000_ );
or   ( new_n12056_, new_n755_, new_n8117_ );
or   ( new_n12057_, new_n757_, new_n7373_ );
and  ( new_n12058_, new_n12057_, new_n12056_ );
xor  ( new_n12059_, new_n12058_, new_n523_ );
or   ( new_n12060_, new_n524_, new_n8352_ );
or   ( new_n12061_, new_n526_, new_n8115_ );
and  ( new_n12062_, new_n12061_, new_n12060_ );
xor  ( new_n12063_, new_n12062_, new_n403_ );
or   ( new_n12064_, new_n12063_, new_n12059_ );
and  ( new_n12065_, new_n12063_, new_n12059_ );
or   ( new_n12066_, new_n409_, new_n8995_ );
or   ( new_n12067_, new_n411_, new_n8481_ );
and  ( new_n12068_, new_n12067_, new_n12066_ );
xor  ( new_n12069_, new_n12068_, new_n328_ );
or   ( new_n12070_, new_n12069_, new_n12065_ );
and  ( new_n12071_, new_n12070_, new_n12064_ );
or   ( new_n12072_, new_n2122_, new_n4995_ );
or   ( new_n12073_, new_n2124_, new_n4603_ );
and  ( new_n12074_, new_n12073_, new_n12072_ );
xor  ( new_n12075_, new_n12074_, new_n1843_ );
or   ( new_n12076_, new_n1844_, new_n5171_ );
or   ( new_n12077_, new_n1846_, new_n4859_ );
and  ( new_n12078_, new_n12077_, new_n12076_ );
xor  ( new_n12079_, new_n12078_, new_n1586_ );
or   ( new_n12080_, new_n12079_, new_n12075_ );
and  ( new_n12081_, new_n12079_, new_n12075_ );
or   ( new_n12082_, new_n1593_, new_n5570_ );
or   ( new_n12083_, new_n1595_, new_n5428_ );
and  ( new_n12084_, new_n12083_, new_n12082_ );
xor  ( new_n12085_, new_n12084_, new_n1358_ );
or   ( new_n12086_, new_n12085_, new_n12081_ );
and  ( new_n12087_, new_n12086_, new_n12080_ );
or   ( new_n12088_, new_n12087_, new_n12071_ );
and  ( new_n12089_, new_n12087_, new_n12071_ );
or   ( new_n12090_, new_n1364_, new_n6219_ );
or   ( new_n12091_, new_n1366_, new_n5899_ );
and  ( new_n12092_, new_n12091_, new_n12090_ );
xor  ( new_n12093_, new_n12092_, new_n1129_ );
or   ( new_n12094_, new_n1135_, new_n6589_ );
or   ( new_n12095_, new_n1137_, new_n6425_ );
and  ( new_n12096_, new_n12095_, new_n12094_ );
xor  ( new_n12097_, new_n12096_, new_n896_ );
nor  ( new_n12098_, new_n12097_, new_n12093_ );
and  ( new_n12099_, new_n12097_, new_n12093_ );
or   ( new_n12100_, new_n897_, new_n7149_ );
or   ( new_n12101_, new_n899_, new_n6943_ );
and  ( new_n12102_, new_n12101_, new_n12100_ );
xor  ( new_n12103_, new_n12102_, new_n748_ );
nor  ( new_n12104_, new_n12103_, new_n12099_ );
nor  ( new_n12105_, new_n12104_, new_n12098_ );
or   ( new_n12106_, new_n12105_, new_n12089_ );
and  ( new_n12107_, new_n12106_, new_n12088_ );
and  ( new_n12108_, new_n12054_, new_n12000_ );
or   ( new_n12109_, new_n12108_, new_n12107_ );
and  ( new_n12110_, new_n12109_, new_n12055_ );
nand ( new_n12111_, new_n12110_, new_n11948_ );
nor  ( new_n12112_, new_n12110_, new_n11948_ );
xor  ( new_n12113_, new_n11621_, new_n11617_ );
xor  ( new_n12114_, new_n12113_, new_n11627_ );
or   ( new_n12115_, new_n337_, new_n9681_ );
or   ( new_n12116_, new_n340_, new_n9099_ );
and  ( new_n12117_, new_n12116_, new_n12115_ );
xor  ( new_n12118_, new_n12117_, new_n332_ );
or   ( new_n12119_, new_n317_, new_n10220_ );
or   ( new_n12120_, new_n320_, new_n9679_ );
and  ( new_n12121_, new_n12120_, new_n12119_ );
xor  ( new_n12122_, new_n12121_, new_n312_ );
or   ( new_n12123_, new_n12122_, new_n12118_ );
and  ( new_n12124_, new_n12122_, new_n12118_ );
or   ( new_n12125_, new_n283_, new_n10841_ );
or   ( new_n12126_, new_n286_, new_n10541_ );
and  ( new_n12127_, new_n12126_, new_n12125_ );
xor  ( new_n12128_, new_n12127_, new_n278_ );
or   ( new_n12129_, new_n12128_, new_n12124_ );
and  ( new_n12130_, new_n12129_, new_n12123_ );
nor  ( new_n12131_, new_n12130_, new_n12114_ );
nand ( new_n12132_, new_n12130_, new_n12114_ );
xor  ( new_n12133_, new_n11606_, new_n11602_ );
not  ( new_n12134_, new_n12133_ );
and  ( new_n12135_, new_n12134_, new_n12132_ );
or   ( new_n12136_, new_n12135_, new_n12131_ );
xnor ( new_n12137_, new_n11679_, new_n11675_ );
xor  ( new_n12138_, new_n12137_, new_n11685_ );
xnor ( new_n12139_, new_n11663_, new_n11659_ );
xor  ( new_n12140_, new_n12139_, new_n11669_ );
or   ( new_n12141_, new_n12140_, new_n12138_ );
and  ( new_n12142_, new_n12140_, new_n12138_ );
xor  ( new_n12143_, new_n11697_, new_n11693_ );
xnor ( new_n12144_, new_n12143_, new_n11703_ );
or   ( new_n12145_, new_n12144_, new_n12142_ );
and  ( new_n12146_, new_n12145_, new_n12141_ );
or   ( new_n12147_, new_n12146_, new_n12136_ );
and  ( new_n12148_, new_n12146_, new_n12136_ );
xnor ( new_n12149_, new_n11782_, new_n11778_ );
xor  ( new_n12150_, new_n12149_, new_n11788_ );
xnor ( new_n12151_, new_n11766_, new_n11762_ );
xor  ( new_n12152_, new_n12151_, new_n11772_ );
nor  ( new_n12153_, new_n12152_, new_n12150_ );
and  ( new_n12154_, new_n12152_, new_n12150_ );
xor  ( new_n12155_, new_n11800_, new_n11796_ );
xnor ( new_n12156_, new_n12155_, new_n11806_ );
nor  ( new_n12157_, new_n12156_, new_n12154_ );
nor  ( new_n12158_, new_n12157_, new_n12153_ );
or   ( new_n12159_, new_n12158_, new_n12148_ );
and  ( new_n12160_, new_n12159_, new_n12147_ );
or   ( new_n12161_, new_n12160_, new_n12112_ );
and  ( new_n12162_, new_n12161_, new_n12111_ );
or   ( new_n12163_, new_n12162_, new_n11930_ );
and  ( new_n12164_, new_n12163_, new_n11929_ );
or   ( new_n12165_, new_n12164_, new_n11892_ );
and  ( new_n12166_, new_n12165_, new_n11891_ );
or   ( new_n12167_, new_n12166_, new_n11878_ );
and  ( new_n12168_, new_n12167_, new_n11877_ );
or   ( new_n12169_, new_n12168_, new_n11864_ );
and  ( new_n12170_, new_n12168_, new_n11864_ );
xor  ( new_n12171_, new_n11844_, new_n11557_ );
xor  ( new_n12172_, new_n12171_, new_n11848_ );
or   ( new_n12173_, new_n12172_, new_n12170_ );
and  ( new_n12174_, new_n12173_, new_n12169_ );
nor  ( new_n12175_, new_n12174_, new_n11858_ );
xor  ( new_n12176_, new_n12168_, new_n11864_ );
xor  ( new_n12177_, new_n12176_, new_n12172_ );
xor  ( new_n12178_, new_n11876_, new_n11866_ );
xor  ( new_n12179_, new_n12178_, new_n12166_ );
xor  ( new_n12180_, new_n11884_, new_n11882_ );
xor  ( new_n12181_, new_n12180_, new_n11888_ );
xor  ( new_n12182_, new_n11757_, new_n11707_ );
xor  ( new_n12183_, new_n12182_, new_n11810_ );
xor  ( new_n12184_, new_n11641_, new_n11631_ );
xor  ( new_n12185_, new_n12184_, new_n11653_ );
nand ( new_n12186_, new_n12185_, new_n12183_ );
nor  ( new_n12187_, new_n12185_, new_n12183_ );
xor  ( new_n12188_, new_n11922_, new_n11920_ );
xor  ( new_n12189_, new_n12188_, new_n11926_ );
or   ( new_n12190_, new_n12189_, new_n12187_ );
and  ( new_n12191_, new_n12190_, new_n12186_ );
or   ( new_n12192_, new_n12191_, new_n12181_ );
and  ( new_n12193_, new_n12191_, new_n12181_ );
xor  ( new_n12194_, new_n11896_, new_n11894_ );
xor  ( new_n12195_, new_n12194_, new_n11900_ );
xnor ( new_n12196_, new_n11906_, new_n11904_ );
xor  ( new_n12197_, new_n12196_, new_n11910_ );
or   ( new_n12198_, new_n12197_, new_n12195_ );
and  ( new_n12199_, new_n12197_, new_n12195_ );
xnor ( new_n12200_, new_n11980_, new_n11964_ );
xor  ( new_n12201_, new_n12200_, new_n11998_ );
xnor ( new_n12202_, new_n12087_, new_n12071_ );
xor  ( new_n12203_, new_n12202_, new_n12105_ );
nor  ( new_n12204_, new_n12203_, new_n12201_ );
and  ( new_n12205_, new_n12203_, new_n12201_ );
xor  ( new_n12206_, new_n12130_, new_n12114_ );
xor  ( new_n12207_, new_n12206_, new_n12134_ );
nor  ( new_n12208_, new_n12207_, new_n12205_ );
nor  ( new_n12209_, new_n12208_, new_n12204_ );
or   ( new_n12210_, new_n12209_, new_n12199_ );
and  ( new_n12211_, new_n12210_, new_n12198_ );
xor  ( new_n12212_, new_n12054_, new_n12000_ );
xor  ( new_n12213_, new_n12212_, new_n12107_ );
xnor ( new_n12214_, new_n12146_, new_n12136_ );
xor  ( new_n12215_, new_n12214_, new_n12158_ );
nand ( new_n12216_, new_n12215_, new_n12213_ );
nor  ( new_n12217_, new_n12215_, new_n12213_ );
xnor ( new_n12218_, new_n11942_, new_n11932_ );
xor  ( new_n12219_, new_n12218_, new_n11946_ );
or   ( new_n12220_, new_n12219_, new_n12217_ );
and  ( new_n12221_, new_n12220_, new_n12216_ );
and  ( new_n12222_, new_n12221_, new_n12211_ );
nor  ( new_n12223_, new_n12221_, new_n12211_ );
xnor ( new_n12224_, new_n11936_, new_n11934_ );
xor  ( new_n12225_, new_n12224_, new_n11940_ );
xnor ( new_n12226_, new_n12140_, new_n12138_ );
xor  ( new_n12227_, new_n12226_, new_n12144_ );
or   ( new_n12228_, new_n12227_, new_n12225_ );
and  ( new_n12229_, new_n12227_, new_n12225_ );
xnor ( new_n12230_, new_n12152_, new_n12150_ );
xor  ( new_n12231_, new_n12230_, new_n12156_ );
or   ( new_n12232_, new_n12231_, new_n12229_ );
and  ( new_n12233_, new_n12232_, new_n12228_ );
or   ( new_n12234_, new_n4709_, new_n2291_ );
or   ( new_n12235_, new_n4711_, new_n2178_ );
and  ( new_n12236_, new_n12235_, new_n12234_ );
xor  ( new_n12237_, new_n12236_, new_n4295_ );
or   ( new_n12238_, new_n4302_, new_n2646_ );
or   ( new_n12239_, new_n4304_, new_n2475_ );
and  ( new_n12240_, new_n12239_, new_n12238_ );
xor  ( new_n12241_, new_n12240_, new_n3895_ );
or   ( new_n12242_, new_n12241_, new_n12237_ );
and  ( new_n12243_, new_n12241_, new_n12237_ );
or   ( new_n12244_, new_n3896_, new_n2981_ );
or   ( new_n12245_, new_n3898_, new_n2751_ );
and  ( new_n12246_, new_n12245_, new_n12244_ );
xor  ( new_n12247_, new_n12246_, new_n3460_ );
or   ( new_n12248_, new_n12247_, new_n12243_ );
and  ( new_n12249_, new_n12248_, new_n12242_ );
or   ( new_n12250_, new_n3461_, new_n3306_ );
or   ( new_n12251_, new_n3463_, new_n3178_ );
and  ( new_n12252_, new_n12251_, new_n12250_ );
xor  ( new_n12253_, new_n12252_, new_n3116_ );
or   ( new_n12254_, new_n3117_, new_n3694_ );
or   ( new_n12255_, new_n3119_, new_n3696_ );
and  ( new_n12256_, new_n12255_, new_n12254_ );
xor  ( new_n12257_, new_n12256_, new_n2800_ );
or   ( new_n12258_, new_n12257_, new_n12253_ );
and  ( new_n12259_, new_n12257_, new_n12253_ );
or   ( new_n12260_, new_n2807_, new_n4069_ );
or   ( new_n12261_, new_n2809_, new_n3820_ );
and  ( new_n12262_, new_n12261_, new_n12260_ );
xor  ( new_n12263_, new_n12262_, new_n2424_ );
or   ( new_n12264_, new_n12263_, new_n12259_ );
and  ( new_n12265_, new_n12264_, new_n12258_ );
or   ( new_n12266_, new_n12265_, new_n12249_ );
and  ( new_n12267_, new_n12265_, new_n12249_ );
or   ( new_n12268_, new_n6173_, new_n1525_ );
or   ( new_n12269_, new_n6175_, new_n1318_ );
and  ( new_n12270_, new_n12269_, new_n12268_ );
xor  ( new_n12271_, new_n12270_, new_n5597_ );
or   ( new_n12272_, new_n5604_, new_n1754_ );
or   ( new_n12273_, new_n5606_, new_n1523_ );
and  ( new_n12274_, new_n12273_, new_n12272_ );
xor  ( new_n12275_, new_n12274_, new_n5206_ );
nor  ( new_n12276_, new_n12275_, new_n12271_ );
and  ( new_n12277_, new_n12275_, new_n12271_ );
or   ( new_n12278_, new_n5207_, new_n2057_ );
or   ( new_n12279_, new_n5209_, new_n1899_ );
and  ( new_n12280_, new_n12279_, new_n12278_ );
xor  ( new_n12281_, new_n12280_, new_n4708_ );
nor  ( new_n12282_, new_n12281_, new_n12277_ );
nor  ( new_n12283_, new_n12282_, new_n12276_ );
or   ( new_n12284_, new_n12283_, new_n12267_ );
and  ( new_n12285_, new_n12284_, new_n12266_ );
or   ( new_n12286_, new_n7732_, new_n805_ );
or   ( new_n12287_, new_n7734_, new_n775_ );
and  ( new_n12288_, new_n12287_, new_n12286_ );
xor  ( new_n12289_, new_n12288_, new_n7177_ );
or   ( new_n12290_, new_n7184_, new_n986_ );
or   ( new_n12291_, new_n7186_, new_n886_ );
and  ( new_n12292_, new_n12291_, new_n12290_ );
xor  ( new_n12293_, new_n12292_, new_n6638_ );
or   ( new_n12294_, new_n12293_, new_n12289_ );
and  ( new_n12295_, new_n12293_, new_n12289_ );
or   ( new_n12296_, new_n6645_, new_n1213_ );
or   ( new_n12297_, new_n6647_, new_n1168_ );
and  ( new_n12298_, new_n12297_, new_n12296_ );
xor  ( new_n12299_, new_n12298_, new_n6166_ );
or   ( new_n12300_, new_n12299_, new_n12295_ );
and  ( new_n12301_, new_n12300_, new_n12294_ );
or   ( new_n12302_, new_n10059_, new_n270_ );
or   ( new_n12303_, new_n10061_, new_n294_ );
and  ( new_n12304_, new_n12303_, new_n12302_ );
xor  ( new_n12305_, new_n12304_, new_n9421_ );
and  ( new_n12306_, RIbb2d888_64, RIbb2d5b8_70 );
or   ( new_n12307_, RIbb2d888_64, new_n301_ );
and  ( new_n12308_, new_n12307_, RIbb2d900_63 );
or   ( new_n12309_, new_n12308_, new_n12306_ );
or   ( new_n12310_, new_n10770_, new_n279_ );
and  ( new_n12311_, new_n12310_, new_n12309_ );
nor  ( new_n12312_, new_n12311_, new_n12305_ );
and  ( new_n12313_, new_n12311_, new_n12305_ );
nor  ( new_n12314_, new_n12313_, new_n277_ );
nor  ( new_n12315_, new_n12314_, new_n12312_ );
or   ( new_n12316_, new_n9422_, new_n348_ );
or   ( new_n12317_, new_n9424_, new_n264_ );
and  ( new_n12318_, new_n12317_, new_n12316_ );
xor  ( new_n12319_, new_n12318_, new_n8873_ );
or   ( new_n12320_, new_n8874_, new_n443_ );
or   ( new_n12321_, new_n8876_, new_n419_ );
and  ( new_n12322_, new_n12321_, new_n12320_ );
xor  ( new_n12323_, new_n12322_, new_n8257_ );
or   ( new_n12324_, new_n12323_, new_n12319_ );
and  ( new_n12325_, new_n12323_, new_n12319_ );
or   ( new_n12326_, new_n8264_, new_n515_ );
or   ( new_n12327_, new_n8266_, new_n509_ );
and  ( new_n12328_, new_n12327_, new_n12326_ );
xor  ( new_n12329_, new_n12328_, new_n7725_ );
or   ( new_n12330_, new_n12329_, new_n12325_ );
and  ( new_n12331_, new_n12330_, new_n12324_ );
and  ( new_n12332_, new_n12331_, new_n12315_ );
or   ( new_n12333_, new_n12332_, new_n12301_ );
or   ( new_n12334_, new_n12331_, new_n12315_ );
and  ( new_n12335_, new_n12334_, new_n12333_ );
or   ( new_n12336_, new_n12335_, new_n12285_ );
or   ( new_n12337_, new_n1593_, new_n5899_ );
or   ( new_n12338_, new_n1595_, new_n5570_ );
and  ( new_n12339_, new_n12338_, new_n12337_ );
xor  ( new_n12340_, new_n12339_, new_n1358_ );
or   ( new_n12341_, new_n1364_, new_n6425_ );
or   ( new_n12342_, new_n1366_, new_n6219_ );
and  ( new_n12343_, new_n12342_, new_n12341_ );
xor  ( new_n12344_, new_n12343_, new_n1129_ );
or   ( new_n12345_, new_n12344_, new_n12340_ );
and  ( new_n12346_, new_n12344_, new_n12340_ );
or   ( new_n12347_, new_n1135_, new_n6943_ );
or   ( new_n12348_, new_n1137_, new_n6589_ );
and  ( new_n12349_, new_n12348_, new_n12347_ );
xor  ( new_n12350_, new_n12349_, new_n896_ );
or   ( new_n12351_, new_n12350_, new_n12346_ );
and  ( new_n12352_, new_n12351_, new_n12345_ );
or   ( new_n12353_, new_n2425_, new_n4603_ );
or   ( new_n12354_, new_n2427_, new_n4267_ );
and  ( new_n12355_, new_n12354_, new_n12353_ );
xor  ( new_n12356_, new_n12355_, new_n2121_ );
or   ( new_n12357_, new_n2122_, new_n4859_ );
or   ( new_n12358_, new_n2124_, new_n4995_ );
and  ( new_n12359_, new_n12358_, new_n12357_ );
xor  ( new_n12360_, new_n12359_, new_n1843_ );
or   ( new_n12361_, new_n12360_, new_n12356_ );
and  ( new_n12362_, new_n12360_, new_n12356_ );
or   ( new_n12363_, new_n1844_, new_n5428_ );
or   ( new_n12364_, new_n1846_, new_n5171_ );
and  ( new_n12365_, new_n12364_, new_n12363_ );
xor  ( new_n12366_, new_n12365_, new_n1586_ );
or   ( new_n12367_, new_n12366_, new_n12362_ );
and  ( new_n12368_, new_n12367_, new_n12361_ );
nor  ( new_n12369_, new_n12368_, new_n12352_ );
and  ( new_n12370_, new_n12368_, new_n12352_ );
or   ( new_n12371_, new_n897_, new_n7373_ );
or   ( new_n12372_, new_n899_, new_n7149_ );
and  ( new_n12373_, new_n12372_, new_n12371_ );
xor  ( new_n12374_, new_n12373_, new_n748_ );
or   ( new_n12375_, new_n755_, new_n8115_ );
or   ( new_n12376_, new_n757_, new_n8117_ );
and  ( new_n12377_, new_n12376_, new_n12375_ );
xor  ( new_n12378_, new_n12377_, new_n523_ );
nor  ( new_n12379_, new_n12378_, new_n12374_ );
and  ( new_n12380_, new_n12378_, new_n12374_ );
or   ( new_n12381_, new_n524_, new_n8481_ );
or   ( new_n12382_, new_n526_, new_n8352_ );
and  ( new_n12383_, new_n12382_, new_n12381_ );
xor  ( new_n12384_, new_n12383_, new_n403_ );
nor  ( new_n12385_, new_n12384_, new_n12380_ );
nor  ( new_n12386_, new_n12385_, new_n12379_ );
nor  ( new_n12387_, new_n12386_, new_n12370_ );
nor  ( new_n12388_, new_n12387_, new_n12369_ );
and  ( new_n12389_, new_n12335_, new_n12285_ );
or   ( new_n12390_, new_n12389_, new_n12388_ );
and  ( new_n12391_, new_n12390_, new_n12336_ );
nor  ( new_n12392_, new_n12391_, new_n12233_ );
and  ( new_n12393_, new_n12391_, new_n12233_ );
xnor ( new_n12394_, new_n11972_, new_n11968_ );
xor  ( new_n12395_, new_n12394_, new_n11978_ );
xnor ( new_n12396_, new_n12079_, new_n12075_ );
xor  ( new_n12397_, new_n12396_, new_n12085_ );
nor  ( new_n12398_, new_n12397_, new_n12395_ );
nand ( new_n12399_, new_n12397_, new_n12395_ );
xor  ( new_n12400_, new_n12097_, new_n12093_ );
xor  ( new_n12401_, new_n12400_, new_n12103_ );
and  ( new_n12402_, new_n12401_, new_n12399_ );
or   ( new_n12403_, new_n12402_, new_n12398_ );
xor  ( new_n12404_, new_n12122_, new_n12118_ );
xor  ( new_n12405_, new_n12404_, new_n12128_ );
or   ( new_n12406_, new_n409_, new_n9099_ );
or   ( new_n12407_, new_n411_, new_n8995_ );
and  ( new_n12408_, new_n12407_, new_n12406_ );
xor  ( new_n12409_, new_n12408_, new_n328_ );
or   ( new_n12410_, new_n337_, new_n9679_ );
or   ( new_n12411_, new_n340_, new_n9681_ );
and  ( new_n12412_, new_n12411_, new_n12410_ );
xor  ( new_n12413_, new_n12412_, new_n332_ );
or   ( new_n12414_, new_n12413_, new_n12409_ );
and  ( new_n12415_, new_n12413_, new_n12409_ );
or   ( new_n12416_, new_n317_, new_n10541_ );
or   ( new_n12417_, new_n320_, new_n10220_ );
and  ( new_n12418_, new_n12417_, new_n12416_ );
xor  ( new_n12419_, new_n12418_, new_n312_ );
or   ( new_n12420_, new_n12419_, new_n12415_ );
and  ( new_n12421_, new_n12420_, new_n12414_ );
or   ( new_n12422_, new_n12421_, new_n12405_ );
nand ( new_n12423_, new_n12421_, new_n12405_ );
xor  ( new_n12424_, new_n12063_, new_n12059_ );
xnor ( new_n12425_, new_n12424_, new_n12069_ );
nand ( new_n12426_, new_n12425_, new_n12423_ );
and  ( new_n12427_, new_n12426_, new_n12422_ );
and  ( new_n12428_, new_n12427_, new_n12403_ );
nor  ( new_n12429_, new_n12427_, new_n12403_ );
xnor ( new_n12430_, new_n12026_, new_n12022_ );
xor  ( new_n12431_, new_n12430_, new_n12032_ );
xnor ( new_n12432_, new_n11956_, new_n11952_ );
xor  ( new_n12433_, new_n12432_, new_n11962_ );
nor  ( new_n12434_, new_n12433_, new_n12431_ );
and  ( new_n12435_, new_n12433_, new_n12431_ );
xor  ( new_n12436_, new_n11990_, new_n11986_ );
xnor ( new_n12437_, new_n12436_, new_n11996_ );
nor  ( new_n12438_, new_n12437_, new_n12435_ );
nor  ( new_n12439_, new_n12438_, new_n12434_ );
nor  ( new_n12440_, new_n12439_, new_n12429_ );
nor  ( new_n12441_, new_n12440_, new_n12428_ );
not  ( new_n12442_, new_n12441_ );
nor  ( new_n12443_, new_n12442_, new_n12393_ );
nor  ( new_n12444_, new_n12443_, new_n12392_ );
nor  ( new_n12445_, new_n12444_, new_n12223_ );
nor  ( new_n12446_, new_n12445_, new_n12222_ );
not  ( new_n12447_, new_n12446_ );
or   ( new_n12448_, new_n12447_, new_n12193_ );
and  ( new_n12449_, new_n12448_, new_n12192_ );
xor  ( new_n12450_, new_n11890_, new_n11880_ );
xor  ( new_n12451_, new_n12450_, new_n12164_ );
or   ( new_n12452_, new_n12451_, new_n12449_ );
and  ( new_n12453_, new_n12451_, new_n12449_ );
xor  ( new_n12454_, new_n11870_, new_n11868_ );
xor  ( new_n12455_, new_n12454_, new_n11874_ );
not  ( new_n12456_, new_n12455_ );
or   ( new_n12457_, new_n12456_, new_n12453_ );
and  ( new_n12458_, new_n12457_, new_n12452_ );
or   ( new_n12459_, new_n12458_, new_n12179_ );
nand ( new_n12460_, new_n12458_, new_n12179_ );
xor  ( new_n12461_, new_n11863_, new_n11861_ );
nand ( new_n12462_, new_n12461_, new_n12460_ );
and  ( new_n12463_, new_n12462_, new_n12459_ );
nor  ( new_n12464_, new_n12463_, new_n12177_ );
xor  ( new_n12465_, new_n12451_, new_n12449_ );
xor  ( new_n12466_, new_n12465_, new_n12456_ );
xor  ( new_n12467_, new_n11928_, new_n11918_ );
xor  ( new_n12468_, new_n12467_, new_n12162_ );
xnor ( new_n12469_, new_n11912_, new_n11902_ );
xor  ( new_n12470_, new_n12469_, new_n11916_ );
xor  ( new_n12471_, new_n12427_, new_n12403_ );
xor  ( new_n12472_, new_n12471_, new_n12439_ );
xnor ( new_n12473_, new_n12335_, new_n12285_ );
xor  ( new_n12474_, new_n12473_, new_n12388_ );
nor  ( new_n12475_, new_n12474_, new_n12472_ );
nand ( new_n12476_, new_n12474_, new_n12472_ );
xor  ( new_n12477_, new_n12227_, new_n12225_ );
xor  ( new_n12478_, new_n12477_, new_n12231_ );
and  ( new_n12479_, new_n12478_, new_n12476_ );
or   ( new_n12480_, new_n12479_, new_n12475_ );
xor  ( new_n12481_, new_n12413_, new_n12409_ );
xor  ( new_n12482_, new_n12481_, new_n12419_ );
and  ( new_n12483_, new_n280_, RIbb31578_128 );
or   ( new_n12484_, new_n12483_, new_n277_ );
nand ( new_n12485_, new_n12483_, RIbb2f430_5 );
and  ( new_n12486_, new_n12485_, new_n12484_ );
nor  ( new_n12487_, new_n12486_, new_n12482_ );
nand ( new_n12488_, new_n12486_, new_n12482_ );
xor  ( new_n12489_, new_n12378_, new_n12374_ );
xnor ( new_n12490_, new_n12489_, new_n12384_ );
and  ( new_n12491_, new_n12490_, new_n12488_ );
or   ( new_n12492_, new_n12491_, new_n12487_ );
xnor ( new_n12493_, new_n12293_, new_n12289_ );
xor  ( new_n12494_, new_n12493_, new_n12299_ );
xnor ( new_n12495_, new_n12241_, new_n12237_ );
xor  ( new_n12496_, new_n12495_, new_n12247_ );
or   ( new_n12497_, new_n12496_, new_n12494_ );
and  ( new_n12498_, new_n12496_, new_n12494_ );
xor  ( new_n12499_, new_n12275_, new_n12271_ );
xnor ( new_n12500_, new_n12499_, new_n12281_ );
or   ( new_n12501_, new_n12500_, new_n12498_ );
and  ( new_n12502_, new_n12501_, new_n12497_ );
nor  ( new_n12503_, new_n12502_, new_n12492_ );
nand ( new_n12504_, new_n12502_, new_n12492_ );
xnor ( new_n12505_, new_n12257_, new_n12253_ );
xor  ( new_n12506_, new_n12505_, new_n12263_ );
xnor ( new_n12507_, new_n12360_, new_n12356_ );
xor  ( new_n12508_, new_n12507_, new_n12366_ );
nor  ( new_n12509_, new_n12508_, new_n12506_ );
nand ( new_n12510_, new_n12508_, new_n12506_ );
xor  ( new_n12511_, new_n12344_, new_n12340_ );
xor  ( new_n12512_, new_n12511_, new_n12350_ );
and  ( new_n12513_, new_n12512_, new_n12510_ );
or   ( new_n12514_, new_n12513_, new_n12509_ );
and  ( new_n12515_, new_n12514_, new_n12504_ );
or   ( new_n12516_, new_n12515_, new_n12503_ );
or   ( new_n12517_, new_n3117_, new_n3820_ );
or   ( new_n12518_, new_n3119_, new_n3694_ );
and  ( new_n12519_, new_n12518_, new_n12517_ );
xor  ( new_n12520_, new_n12519_, new_n2800_ );
or   ( new_n12521_, new_n2807_, new_n4267_ );
or   ( new_n12522_, new_n2809_, new_n4069_ );
and  ( new_n12523_, new_n12522_, new_n12521_ );
xor  ( new_n12524_, new_n12523_, new_n2424_ );
or   ( new_n12525_, new_n12524_, new_n12520_ );
and  ( new_n12526_, new_n12524_, new_n12520_ );
or   ( new_n12527_, new_n2425_, new_n4995_ );
or   ( new_n12528_, new_n2427_, new_n4603_ );
and  ( new_n12529_, new_n12528_, new_n12527_ );
xor  ( new_n12530_, new_n12529_, new_n2121_ );
or   ( new_n12531_, new_n12530_, new_n12526_ );
and  ( new_n12532_, new_n12531_, new_n12525_ );
or   ( new_n12533_, new_n4302_, new_n2751_ );
or   ( new_n12534_, new_n4304_, new_n2646_ );
and  ( new_n12535_, new_n12534_, new_n12533_ );
xor  ( new_n12536_, new_n12535_, new_n3895_ );
or   ( new_n12537_, new_n3896_, new_n3178_ );
or   ( new_n12538_, new_n3898_, new_n2981_ );
and  ( new_n12539_, new_n12538_, new_n12537_ );
xor  ( new_n12540_, new_n12539_, new_n3460_ );
or   ( new_n12541_, new_n12540_, new_n12536_ );
and  ( new_n12542_, new_n12540_, new_n12536_ );
or   ( new_n12543_, new_n3461_, new_n3696_ );
or   ( new_n12544_, new_n3463_, new_n3306_ );
and  ( new_n12545_, new_n12544_, new_n12543_ );
xor  ( new_n12546_, new_n12545_, new_n3116_ );
or   ( new_n12547_, new_n12546_, new_n12542_ );
and  ( new_n12548_, new_n12547_, new_n12541_ );
or   ( new_n12549_, new_n12548_, new_n12532_ );
and  ( new_n12550_, new_n12548_, new_n12532_ );
or   ( new_n12551_, new_n5604_, new_n1899_ );
or   ( new_n12552_, new_n5606_, new_n1754_ );
and  ( new_n12553_, new_n12552_, new_n12551_ );
xor  ( new_n12554_, new_n12553_, new_n5206_ );
or   ( new_n12555_, new_n5207_, new_n2178_ );
or   ( new_n12556_, new_n5209_, new_n2057_ );
and  ( new_n12557_, new_n12556_, new_n12555_ );
xor  ( new_n12558_, new_n12557_, new_n4708_ );
nor  ( new_n12559_, new_n12558_, new_n12554_ );
and  ( new_n12560_, new_n12558_, new_n12554_ );
or   ( new_n12561_, new_n4709_, new_n2475_ );
or   ( new_n12562_, new_n4711_, new_n2291_ );
and  ( new_n12563_, new_n12562_, new_n12561_ );
xor  ( new_n12564_, new_n12563_, new_n4295_ );
nor  ( new_n12565_, new_n12564_, new_n12560_ );
nor  ( new_n12566_, new_n12565_, new_n12559_ );
or   ( new_n12567_, new_n12566_, new_n12550_ );
and  ( new_n12568_, new_n12567_, new_n12549_ );
or   ( new_n12569_, new_n755_, new_n8352_ );
or   ( new_n12570_, new_n757_, new_n8115_ );
and  ( new_n12571_, new_n12570_, new_n12569_ );
xor  ( new_n12572_, new_n12571_, new_n523_ );
or   ( new_n12573_, new_n524_, new_n8995_ );
or   ( new_n12574_, new_n526_, new_n8481_ );
and  ( new_n12575_, new_n12574_, new_n12573_ );
xor  ( new_n12576_, new_n12575_, new_n403_ );
or   ( new_n12577_, new_n12576_, new_n12572_ );
and  ( new_n12578_, new_n12576_, new_n12572_ );
or   ( new_n12579_, new_n409_, new_n9681_ );
or   ( new_n12580_, new_n411_, new_n9099_ );
and  ( new_n12581_, new_n12580_, new_n12579_ );
xor  ( new_n12582_, new_n12581_, new_n328_ );
or   ( new_n12583_, new_n12582_, new_n12578_ );
and  ( new_n12584_, new_n12583_, new_n12577_ );
or   ( new_n12585_, new_n1364_, new_n6589_ );
or   ( new_n12586_, new_n1366_, new_n6425_ );
and  ( new_n12587_, new_n12586_, new_n12585_ );
xor  ( new_n12588_, new_n12587_, new_n1129_ );
or   ( new_n12589_, new_n1135_, new_n7149_ );
or   ( new_n12590_, new_n1137_, new_n6943_ );
and  ( new_n12591_, new_n12590_, new_n12589_ );
xor  ( new_n12592_, new_n12591_, new_n896_ );
or   ( new_n12593_, new_n12592_, new_n12588_ );
and  ( new_n12594_, new_n12592_, new_n12588_ );
or   ( new_n12595_, new_n897_, new_n8117_ );
or   ( new_n12596_, new_n899_, new_n7373_ );
and  ( new_n12597_, new_n12596_, new_n12595_ );
xor  ( new_n12598_, new_n12597_, new_n748_ );
or   ( new_n12599_, new_n12598_, new_n12594_ );
and  ( new_n12600_, new_n12599_, new_n12593_ );
or   ( new_n12601_, new_n12600_, new_n12584_ );
and  ( new_n12602_, new_n12600_, new_n12584_ );
or   ( new_n12603_, new_n2122_, new_n5171_ );
or   ( new_n12604_, new_n2124_, new_n4859_ );
and  ( new_n12605_, new_n12604_, new_n12603_ );
xor  ( new_n12606_, new_n12605_, new_n1843_ );
or   ( new_n12607_, new_n1844_, new_n5570_ );
or   ( new_n12608_, new_n1846_, new_n5428_ );
and  ( new_n12609_, new_n12608_, new_n12607_ );
xor  ( new_n12610_, new_n12609_, new_n1586_ );
nor  ( new_n12611_, new_n12610_, new_n12606_ );
and  ( new_n12612_, new_n12610_, new_n12606_ );
or   ( new_n12613_, new_n1593_, new_n6219_ );
or   ( new_n12614_, new_n1595_, new_n5899_ );
and  ( new_n12615_, new_n12614_, new_n12613_ );
xor  ( new_n12616_, new_n12615_, new_n1358_ );
nor  ( new_n12617_, new_n12616_, new_n12612_ );
nor  ( new_n12618_, new_n12617_, new_n12611_ );
or   ( new_n12619_, new_n12618_, new_n12602_ );
and  ( new_n12620_, new_n12619_, new_n12601_ );
or   ( new_n12621_, new_n12620_, new_n12568_ );
or   ( new_n12622_, new_n8874_, new_n509_ );
or   ( new_n12623_, new_n8876_, new_n443_ );
and  ( new_n12624_, new_n12623_, new_n12622_ );
xor  ( new_n12625_, new_n12624_, new_n8257_ );
or   ( new_n12626_, new_n8264_, new_n775_ );
or   ( new_n12627_, new_n8266_, new_n515_ );
and  ( new_n12628_, new_n12627_, new_n12626_ );
xor  ( new_n12629_, new_n12628_, new_n7725_ );
or   ( new_n12630_, new_n12629_, new_n12625_ );
and  ( new_n12631_, new_n12629_, new_n12625_ );
or   ( new_n12632_, new_n7732_, new_n886_ );
or   ( new_n12633_, new_n7734_, new_n805_ );
and  ( new_n12634_, new_n12633_, new_n12632_ );
xor  ( new_n12635_, new_n12634_, new_n7177_ );
or   ( new_n12636_, new_n12635_, new_n12631_ );
and  ( new_n12637_, new_n12636_, new_n12630_ );
or   ( new_n12638_, new_n10059_, new_n264_ );
or   ( new_n12639_, new_n10061_, new_n270_ );
and  ( new_n12640_, new_n12639_, new_n12638_ );
xor  ( new_n12641_, new_n12640_, new_n9421_ );
and  ( new_n12642_, RIbb2d888_64, RIbb2d540_71 );
or   ( new_n12643_, RIbb2d888_64, new_n294_ );
and  ( new_n12644_, new_n12643_, RIbb2d900_63 );
or   ( new_n12645_, new_n12644_, new_n12642_ );
or   ( new_n12646_, new_n10770_, new_n301_ );
and  ( new_n12647_, new_n12646_, new_n12645_ );
or   ( new_n12648_, new_n12647_, new_n12641_ );
and  ( new_n12649_, new_n12647_, new_n12641_ );
or   ( new_n12650_, new_n9422_, new_n419_ );
or   ( new_n12651_, new_n9424_, new_n348_ );
and  ( new_n12652_, new_n12651_, new_n12650_ );
xor  ( new_n12653_, new_n12652_, new_n8873_ );
or   ( new_n12654_, new_n12653_, new_n12649_ );
and  ( new_n12655_, new_n12654_, new_n12648_ );
or   ( new_n12656_, new_n12655_, new_n12637_ );
and  ( new_n12657_, new_n12655_, new_n12637_ );
or   ( new_n12658_, new_n7184_, new_n1168_ );
or   ( new_n12659_, new_n7186_, new_n986_ );
and  ( new_n12660_, new_n12659_, new_n12658_ );
xor  ( new_n12661_, new_n12660_, new_n6638_ );
or   ( new_n12662_, new_n6645_, new_n1318_ );
or   ( new_n12663_, new_n6647_, new_n1213_ );
and  ( new_n12664_, new_n12663_, new_n12662_ );
xor  ( new_n12665_, new_n12664_, new_n6166_ );
nor  ( new_n12666_, new_n12665_, new_n12661_ );
and  ( new_n12667_, new_n12665_, new_n12661_ );
or   ( new_n12668_, new_n6173_, new_n1523_ );
or   ( new_n12669_, new_n6175_, new_n1525_ );
and  ( new_n12670_, new_n12669_, new_n12668_ );
xor  ( new_n12671_, new_n12670_, new_n5597_ );
nor  ( new_n12672_, new_n12671_, new_n12667_ );
nor  ( new_n12673_, new_n12672_, new_n12666_ );
or   ( new_n12674_, new_n12673_, new_n12657_ );
and  ( new_n12675_, new_n12674_, new_n12656_ );
and  ( new_n12676_, new_n12620_, new_n12568_ );
or   ( new_n12677_, new_n12676_, new_n12675_ );
and  ( new_n12678_, new_n12677_, new_n12621_ );
or   ( new_n12679_, new_n12678_, new_n12516_ );
and  ( new_n12680_, new_n12678_, new_n12516_ );
xnor ( new_n12681_, new_n12010_, new_n12004_ );
xor  ( new_n12682_, new_n12681_, new_n12016_ );
xnor ( new_n12683_, new_n12044_, new_n12040_ );
xor  ( new_n12684_, new_n12683_, new_n12050_ );
nor  ( new_n12685_, new_n12684_, new_n12682_ );
nand ( new_n12686_, new_n12684_, new_n12682_ );
xor  ( new_n12687_, new_n12433_, new_n12431_ );
xnor ( new_n12688_, new_n12687_, new_n12437_ );
and  ( new_n12689_, new_n12688_, new_n12686_ );
or   ( new_n12690_, new_n12689_, new_n12685_ );
or   ( new_n12691_, new_n12690_, new_n12680_ );
and  ( new_n12692_, new_n12691_, new_n12679_ );
or   ( new_n12693_, new_n12692_, new_n12480_ );
nand ( new_n12694_, new_n12692_, new_n12480_ );
xnor ( new_n12695_, new_n12034_, new_n12018_ );
xor  ( new_n12696_, new_n12695_, new_n12052_ );
xor  ( new_n12697_, new_n12368_, new_n12352_ );
xor  ( new_n12698_, new_n12697_, new_n12386_ );
xor  ( new_n12699_, new_n12397_, new_n12395_ );
xor  ( new_n12700_, new_n12699_, new_n12401_ );
nand ( new_n12701_, new_n12700_, new_n12698_ );
nor  ( new_n12702_, new_n12700_, new_n12698_ );
xor  ( new_n12703_, new_n12421_, new_n12405_ );
xor  ( new_n12704_, new_n12703_, new_n12425_ );
or   ( new_n12705_, new_n12704_, new_n12702_ );
and  ( new_n12706_, new_n12705_, new_n12701_ );
nor  ( new_n12707_, new_n12706_, new_n12696_ );
and  ( new_n12708_, new_n12706_, new_n12696_ );
xor  ( new_n12709_, new_n12203_, new_n12201_ );
xnor ( new_n12710_, new_n12709_, new_n12207_ );
not  ( new_n12711_, new_n12710_ );
nor  ( new_n12712_, new_n12711_, new_n12708_ );
nor  ( new_n12713_, new_n12712_, new_n12707_ );
nand ( new_n12714_, new_n12713_, new_n12694_ );
and  ( new_n12715_, new_n12714_, new_n12693_ );
nor  ( new_n12716_, new_n12715_, new_n12470_ );
xor  ( new_n12717_, new_n12391_, new_n12233_ );
xor  ( new_n12718_, new_n12717_, new_n12442_ );
xnor ( new_n12719_, new_n12197_, new_n12195_ );
xor  ( new_n12720_, new_n12719_, new_n12209_ );
nor  ( new_n12721_, new_n12720_, new_n12718_ );
nand ( new_n12722_, new_n12720_, new_n12718_ );
xor  ( new_n12723_, new_n12215_, new_n12213_ );
xor  ( new_n12724_, new_n12723_, new_n12219_ );
and  ( new_n12725_, new_n12724_, new_n12722_ );
or   ( new_n12726_, new_n12725_, new_n12721_ );
nand ( new_n12727_, new_n12715_, new_n12470_ );
and  ( new_n12728_, new_n12727_, new_n12726_ );
or   ( new_n12729_, new_n12728_, new_n12716_ );
or   ( new_n12730_, new_n12729_, new_n12468_ );
and  ( new_n12731_, new_n12729_, new_n12468_ );
xor  ( new_n12732_, new_n12110_, new_n11948_ );
xor  ( new_n12733_, new_n12732_, new_n12160_ );
xnor ( new_n12734_, new_n12221_, new_n12211_ );
xor  ( new_n12735_, new_n12734_, new_n12444_ );
or   ( new_n12736_, new_n12735_, new_n12733_ );
and  ( new_n12737_, new_n12735_, new_n12733_ );
xor  ( new_n12738_, new_n12185_, new_n12183_ );
xor  ( new_n12739_, new_n12738_, new_n12189_ );
or   ( new_n12740_, new_n12739_, new_n12737_ );
and  ( new_n12741_, new_n12740_, new_n12736_ );
or   ( new_n12742_, new_n12741_, new_n12731_ );
and  ( new_n12743_, new_n12742_, new_n12730_ );
nor  ( new_n12744_, new_n12743_, new_n12466_ );
xor  ( new_n12745_, new_n12458_, new_n12179_ );
xor  ( new_n12746_, new_n12745_, new_n12461_ );
and  ( new_n12747_, new_n12746_, new_n12744_ );
xnor ( new_n12748_, new_n12743_, new_n12466_ );
xor  ( new_n12749_, new_n12741_, new_n12468_ );
xor  ( new_n12750_, new_n12749_, new_n12729_ );
xor  ( new_n12751_, new_n12720_, new_n12718_ );
xor  ( new_n12752_, new_n12751_, new_n12724_ );
xor  ( new_n12753_, new_n12678_, new_n12516_ );
xor  ( new_n12754_, new_n12753_, new_n12690_ );
xor  ( new_n12755_, new_n12474_, new_n12472_ );
xor  ( new_n12756_, new_n12755_, new_n12478_ );
nand ( new_n12757_, new_n12756_, new_n12754_ );
nor  ( new_n12758_, new_n12756_, new_n12754_ );
xor  ( new_n12759_, new_n12706_, new_n12696_ );
xor  ( new_n12760_, new_n12759_, new_n12711_ );
or   ( new_n12761_, new_n12760_, new_n12758_ );
and  ( new_n12762_, new_n12761_, new_n12757_ );
or   ( new_n12763_, new_n12762_, new_n12752_ );
and  ( new_n12764_, new_n12762_, new_n12752_ );
xnor ( new_n12765_, new_n12265_, new_n12249_ );
xor  ( new_n12766_, new_n12765_, new_n12283_ );
xnor ( new_n12767_, new_n12496_, new_n12494_ );
xor  ( new_n12768_, new_n12767_, new_n12500_ );
xor  ( new_n12769_, new_n12508_, new_n12506_ );
xor  ( new_n12770_, new_n12769_, new_n12512_ );
nand ( new_n12771_, new_n12770_, new_n12768_ );
nor  ( new_n12772_, new_n12770_, new_n12768_ );
xor  ( new_n12773_, new_n12486_, new_n12482_ );
xor  ( new_n12774_, new_n12773_, new_n12490_ );
or   ( new_n12775_, new_n12774_, new_n12772_ );
and  ( new_n12776_, new_n12775_, new_n12771_ );
or   ( new_n12777_, new_n12776_, new_n12766_ );
and  ( new_n12778_, new_n12776_, new_n12766_ );
xnor ( new_n12779_, new_n12548_, new_n12532_ );
xor  ( new_n12780_, new_n12779_, new_n12566_ );
xnor ( new_n12781_, new_n12600_, new_n12584_ );
xor  ( new_n12782_, new_n12781_, new_n12618_ );
or   ( new_n12783_, new_n12782_, new_n12780_ );
and  ( new_n12784_, new_n12782_, new_n12780_ );
xor  ( new_n12785_, new_n12655_, new_n12637_ );
xnor ( new_n12786_, new_n12785_, new_n12673_ );
or   ( new_n12787_, new_n12786_, new_n12784_ );
and  ( new_n12788_, new_n12787_, new_n12783_ );
or   ( new_n12789_, new_n12788_, new_n12778_ );
and  ( new_n12790_, new_n12789_, new_n12777_ );
xnor ( new_n12791_, new_n12331_, new_n12315_ );
xor  ( new_n12792_, new_n12791_, new_n12301_ );
xnor ( new_n12793_, new_n12684_, new_n12682_ );
xor  ( new_n12794_, new_n12793_, new_n12688_ );
or   ( new_n12795_, new_n12794_, new_n12792_ );
and  ( new_n12796_, new_n12794_, new_n12792_ );
xor  ( new_n12797_, new_n12700_, new_n12698_ );
xor  ( new_n12798_, new_n12797_, new_n12704_ );
or   ( new_n12799_, new_n12798_, new_n12796_ );
and  ( new_n12800_, new_n12799_, new_n12795_ );
nor  ( new_n12801_, new_n12800_, new_n12790_ );
and  ( new_n12802_, new_n12800_, new_n12790_ );
xor  ( new_n12803_, new_n12311_, new_n12305_ );
xor  ( new_n12804_, new_n12803_, new_n278_ );
xnor ( new_n12805_, new_n12647_, new_n12641_ );
xor  ( new_n12806_, new_n12805_, new_n12653_ );
xnor ( new_n12807_, new_n12629_, new_n12625_ );
xor  ( new_n12808_, new_n12807_, new_n12635_ );
or   ( new_n12809_, new_n12808_, new_n12806_ );
and  ( new_n12810_, new_n12808_, new_n12806_ );
xor  ( new_n12811_, new_n12665_, new_n12661_ );
xnor ( new_n12812_, new_n12811_, new_n12671_ );
or   ( new_n12813_, new_n12812_, new_n12810_ );
and  ( new_n12814_, new_n12813_, new_n12809_ );
nor  ( new_n12815_, new_n12814_, new_n12804_ );
and  ( new_n12816_, new_n12814_, new_n12804_ );
xor  ( new_n12817_, new_n12323_, new_n12319_ );
xnor ( new_n12818_, new_n12817_, new_n12329_ );
nor  ( new_n12819_, new_n12818_, new_n12816_ );
or   ( new_n12820_, new_n12819_, new_n12815_ );
or   ( new_n12821_, new_n6173_, new_n1754_ );
or   ( new_n12822_, new_n6175_, new_n1523_ );
and  ( new_n12823_, new_n12822_, new_n12821_ );
xor  ( new_n12824_, new_n12823_, new_n5597_ );
or   ( new_n12825_, new_n5604_, new_n2057_ );
or   ( new_n12826_, new_n5606_, new_n1899_ );
and  ( new_n12827_, new_n12826_, new_n12825_ );
xor  ( new_n12828_, new_n12827_, new_n5206_ );
or   ( new_n12829_, new_n12828_, new_n12824_ );
and  ( new_n12830_, new_n12828_, new_n12824_ );
or   ( new_n12831_, new_n5207_, new_n2291_ );
or   ( new_n12832_, new_n5209_, new_n2178_ );
and  ( new_n12833_, new_n12832_, new_n12831_ );
xor  ( new_n12834_, new_n12833_, new_n4708_ );
or   ( new_n12835_, new_n12834_, new_n12830_ );
and  ( new_n12836_, new_n12835_, new_n12829_ );
or   ( new_n12837_, new_n3461_, new_n3694_ );
or   ( new_n12838_, new_n3463_, new_n3696_ );
and  ( new_n12839_, new_n12838_, new_n12837_ );
xor  ( new_n12840_, new_n12839_, new_n3116_ );
or   ( new_n12841_, new_n3117_, new_n4069_ );
or   ( new_n12842_, new_n3119_, new_n3820_ );
and  ( new_n12843_, new_n12842_, new_n12841_ );
xor  ( new_n12844_, new_n12843_, new_n2800_ );
or   ( new_n12845_, new_n12844_, new_n12840_ );
and  ( new_n12846_, new_n12844_, new_n12840_ );
or   ( new_n12847_, new_n2807_, new_n4603_ );
or   ( new_n12848_, new_n2809_, new_n4267_ );
and  ( new_n12849_, new_n12848_, new_n12847_ );
xor  ( new_n12850_, new_n12849_, new_n2424_ );
or   ( new_n12851_, new_n12850_, new_n12846_ );
and  ( new_n12852_, new_n12851_, new_n12845_ );
or   ( new_n12853_, new_n12852_, new_n12836_ );
and  ( new_n12854_, new_n12852_, new_n12836_ );
or   ( new_n12855_, new_n4709_, new_n2646_ );
or   ( new_n12856_, new_n4711_, new_n2475_ );
and  ( new_n12857_, new_n12856_, new_n12855_ );
xor  ( new_n12858_, new_n12857_, new_n4295_ );
or   ( new_n12859_, new_n4302_, new_n2981_ );
or   ( new_n12860_, new_n4304_, new_n2751_ );
and  ( new_n12861_, new_n12860_, new_n12859_ );
xor  ( new_n12862_, new_n12861_, new_n3895_ );
nor  ( new_n12863_, new_n12862_, new_n12858_ );
and  ( new_n12864_, new_n12862_, new_n12858_ );
or   ( new_n12865_, new_n3896_, new_n3306_ );
or   ( new_n12866_, new_n3898_, new_n3178_ );
and  ( new_n12867_, new_n12866_, new_n12865_ );
xor  ( new_n12868_, new_n12867_, new_n3460_ );
nor  ( new_n12869_, new_n12868_, new_n12864_ );
nor  ( new_n12870_, new_n12869_, new_n12863_ );
or   ( new_n12871_, new_n12870_, new_n12854_ );
and  ( new_n12872_, new_n12871_, new_n12853_ );
or   ( new_n12873_, new_n9422_, new_n443_ );
or   ( new_n12874_, new_n9424_, new_n419_ );
and  ( new_n12875_, new_n12874_, new_n12873_ );
xor  ( new_n12876_, new_n12875_, new_n8873_ );
or   ( new_n12877_, new_n8874_, new_n515_ );
or   ( new_n12878_, new_n8876_, new_n509_ );
and  ( new_n12879_, new_n12878_, new_n12877_ );
xor  ( new_n12880_, new_n12879_, new_n8257_ );
or   ( new_n12881_, new_n12880_, new_n12876_ );
and  ( new_n12882_, new_n12880_, new_n12876_ );
or   ( new_n12883_, new_n8264_, new_n805_ );
or   ( new_n12884_, new_n8266_, new_n775_ );
and  ( new_n12885_, new_n12884_, new_n12883_ );
xor  ( new_n12886_, new_n12885_, new_n7725_ );
or   ( new_n12887_, new_n12886_, new_n12882_ );
and  ( new_n12888_, new_n12887_, new_n12881_ );
or   ( new_n12889_, new_n10059_, new_n348_ );
or   ( new_n12890_, new_n10061_, new_n264_ );
and  ( new_n12891_, new_n12890_, new_n12889_ );
xor  ( new_n12892_, new_n12891_, new_n9421_ );
and  ( new_n12893_, RIbb2d888_64, RIbb2d4c8_72 );
or   ( new_n12894_, RIbb2d888_64, new_n270_ );
and  ( new_n12895_, new_n12894_, RIbb2d900_63 );
or   ( new_n12896_, new_n12895_, new_n12893_ );
or   ( new_n12897_, new_n10770_, new_n294_ );
and  ( new_n12898_, new_n12897_, new_n12896_ );
nor  ( new_n12899_, new_n12898_, new_n12892_ );
and  ( new_n12900_, new_n12898_, new_n12892_ );
nor  ( new_n12901_, new_n12900_, new_n311_ );
nor  ( new_n12902_, new_n12901_, new_n12899_ );
or   ( new_n12903_, new_n7732_, new_n986_ );
or   ( new_n12904_, new_n7734_, new_n886_ );
and  ( new_n12905_, new_n12904_, new_n12903_ );
xor  ( new_n12906_, new_n12905_, new_n7177_ );
or   ( new_n12907_, new_n7184_, new_n1213_ );
or   ( new_n12908_, new_n7186_, new_n1168_ );
and  ( new_n12909_, new_n12908_, new_n12907_ );
xor  ( new_n12910_, new_n12909_, new_n6638_ );
or   ( new_n12911_, new_n12910_, new_n12906_ );
and  ( new_n12912_, new_n12910_, new_n12906_ );
or   ( new_n12913_, new_n6645_, new_n1525_ );
or   ( new_n12914_, new_n6647_, new_n1318_ );
and  ( new_n12915_, new_n12914_, new_n12913_ );
xor  ( new_n12916_, new_n12915_, new_n6166_ );
or   ( new_n12917_, new_n12916_, new_n12912_ );
and  ( new_n12918_, new_n12917_, new_n12911_ );
and  ( new_n12919_, new_n12918_, new_n12902_ );
or   ( new_n12920_, new_n12919_, new_n12888_ );
or   ( new_n12921_, new_n12918_, new_n12902_ );
and  ( new_n12922_, new_n12921_, new_n12920_ );
or   ( new_n12923_, new_n12922_, new_n12872_ );
or   ( new_n12924_, new_n897_, new_n8115_ );
or   ( new_n12925_, new_n899_, new_n8117_ );
and  ( new_n12926_, new_n12925_, new_n12924_ );
xor  ( new_n12927_, new_n12926_, new_n748_ );
or   ( new_n12928_, new_n755_, new_n8481_ );
or   ( new_n12929_, new_n757_, new_n8352_ );
and  ( new_n12930_, new_n12929_, new_n12928_ );
xor  ( new_n12931_, new_n12930_, new_n523_ );
or   ( new_n12932_, new_n12931_, new_n12927_ );
and  ( new_n12933_, new_n12931_, new_n12927_ );
or   ( new_n12934_, new_n524_, new_n9099_ );
or   ( new_n12935_, new_n526_, new_n8995_ );
and  ( new_n12936_, new_n12935_, new_n12934_ );
xor  ( new_n12937_, new_n12936_, new_n403_ );
or   ( new_n12938_, new_n12937_, new_n12933_ );
and  ( new_n12939_, new_n12938_, new_n12932_ );
or   ( new_n12940_, new_n1593_, new_n6425_ );
or   ( new_n12941_, new_n1595_, new_n6219_ );
and  ( new_n12942_, new_n12941_, new_n12940_ );
xor  ( new_n12943_, new_n12942_, new_n1358_ );
or   ( new_n12944_, new_n1364_, new_n6943_ );
or   ( new_n12945_, new_n1366_, new_n6589_ );
and  ( new_n12946_, new_n12945_, new_n12944_ );
xor  ( new_n12947_, new_n12946_, new_n1129_ );
or   ( new_n12948_, new_n12947_, new_n12943_ );
and  ( new_n12949_, new_n12947_, new_n12943_ );
or   ( new_n12950_, new_n1135_, new_n7373_ );
or   ( new_n12951_, new_n1137_, new_n7149_ );
and  ( new_n12952_, new_n12951_, new_n12950_ );
xor  ( new_n12953_, new_n12952_, new_n896_ );
or   ( new_n12954_, new_n12953_, new_n12949_ );
and  ( new_n12955_, new_n12954_, new_n12948_ );
nor  ( new_n12956_, new_n12955_, new_n12939_ );
and  ( new_n12957_, new_n12955_, new_n12939_ );
or   ( new_n12958_, new_n2425_, new_n4859_ );
or   ( new_n12959_, new_n2427_, new_n4995_ );
and  ( new_n12960_, new_n12959_, new_n12958_ );
xor  ( new_n12961_, new_n12960_, new_n2121_ );
or   ( new_n12962_, new_n2122_, new_n5428_ );
or   ( new_n12963_, new_n2124_, new_n5171_ );
and  ( new_n12964_, new_n12963_, new_n12962_ );
xor  ( new_n12965_, new_n12964_, new_n1843_ );
nor  ( new_n12966_, new_n12965_, new_n12961_ );
and  ( new_n12967_, new_n12965_, new_n12961_ );
or   ( new_n12968_, new_n1844_, new_n5899_ );
or   ( new_n12969_, new_n1846_, new_n5570_ );
and  ( new_n12970_, new_n12969_, new_n12968_ );
xor  ( new_n12971_, new_n12970_, new_n1586_ );
nor  ( new_n12972_, new_n12971_, new_n12967_ );
nor  ( new_n12973_, new_n12972_, new_n12966_ );
nor  ( new_n12974_, new_n12973_, new_n12957_ );
nor  ( new_n12975_, new_n12974_, new_n12956_ );
and  ( new_n12976_, new_n12922_, new_n12872_ );
or   ( new_n12977_, new_n12976_, new_n12975_ );
and  ( new_n12978_, new_n12977_, new_n12923_ );
and  ( new_n12979_, new_n12978_, new_n12820_ );
nor  ( new_n12980_, new_n12978_, new_n12820_ );
xnor ( new_n12981_, new_n12592_, new_n12588_ );
xor  ( new_n12982_, new_n12981_, new_n12598_ );
xnor ( new_n12983_, new_n12576_, new_n12572_ );
xor  ( new_n12984_, new_n12983_, new_n12582_ );
or   ( new_n12985_, new_n12984_, new_n12982_ );
and  ( new_n12986_, new_n12984_, new_n12982_ );
xor  ( new_n12987_, new_n12610_, new_n12606_ );
xnor ( new_n12988_, new_n12987_, new_n12616_ );
or   ( new_n12989_, new_n12988_, new_n12986_ );
and  ( new_n12990_, new_n12989_, new_n12985_ );
xnor ( new_n12991_, new_n12540_, new_n12536_ );
xor  ( new_n12992_, new_n12991_, new_n12546_ );
xnor ( new_n12993_, new_n12524_, new_n12520_ );
xor  ( new_n12994_, new_n12993_, new_n12530_ );
or   ( new_n12995_, new_n12994_, new_n12992_ );
and  ( new_n12996_, new_n12994_, new_n12992_ );
xor  ( new_n12997_, new_n12558_, new_n12554_ );
xnor ( new_n12998_, new_n12997_, new_n12564_ );
or   ( new_n12999_, new_n12998_, new_n12996_ );
and  ( new_n13000_, new_n12999_, new_n12995_ );
nor  ( new_n13001_, new_n13000_, new_n12990_ );
and  ( new_n13002_, new_n13000_, new_n12990_ );
or   ( new_n13003_, new_n337_, new_n10220_ );
or   ( new_n13004_, new_n340_, new_n9679_ );
and  ( new_n13005_, new_n13004_, new_n13003_ );
xor  ( new_n13006_, new_n13005_, new_n332_ );
or   ( new_n13007_, new_n409_, new_n9679_ );
or   ( new_n13008_, new_n411_, new_n9681_ );
and  ( new_n13009_, new_n13008_, new_n13007_ );
xor  ( new_n13010_, new_n13009_, new_n328_ );
or   ( new_n13011_, new_n337_, new_n10541_ );
or   ( new_n13012_, new_n340_, new_n10220_ );
and  ( new_n13013_, new_n13012_, new_n13011_ );
xor  ( new_n13014_, new_n13013_, new_n332_ );
or   ( new_n13015_, new_n13014_, new_n13010_ );
and  ( new_n13016_, new_n13014_, new_n13010_ );
and  ( new_n13017_, new_n314_, RIbb31578_128 );
nor  ( new_n13018_, new_n13017_, new_n311_ );
and  ( new_n13019_, new_n13017_, RIbb2f340_7 );
nor  ( new_n13020_, new_n13019_, new_n13018_ );
or   ( new_n13021_, new_n13020_, new_n13016_ );
and  ( new_n13022_, new_n13021_, new_n13015_ );
and  ( new_n13023_, new_n13022_, new_n13006_ );
nor  ( new_n13024_, new_n13022_, new_n13006_ );
or   ( new_n13025_, new_n317_, new_n10841_ );
or   ( new_n13026_, new_n320_, new_n10541_ );
and  ( new_n13027_, new_n13026_, new_n13025_ );
xor  ( new_n13028_, new_n13027_, new_n312_ );
not  ( new_n13029_, new_n13028_ );
nor  ( new_n13030_, new_n13029_, new_n13024_ );
nor  ( new_n13031_, new_n13030_, new_n13023_ );
nor  ( new_n13032_, new_n13031_, new_n13002_ );
nor  ( new_n13033_, new_n13032_, new_n13001_ );
nor  ( new_n13034_, new_n13033_, new_n12980_ );
nor  ( new_n13035_, new_n13034_, new_n12979_ );
nor  ( new_n13036_, new_n13035_, new_n12802_ );
nor  ( new_n13037_, new_n13036_, new_n12801_ );
or   ( new_n13038_, new_n13037_, new_n12764_ );
and  ( new_n13039_, new_n13038_, new_n12763_ );
xor  ( new_n13040_, new_n12715_, new_n12470_ );
xor  ( new_n13041_, new_n13040_, new_n12726_ );
or   ( new_n13042_, new_n13041_, new_n13039_ );
and  ( new_n13043_, new_n13041_, new_n13039_ );
xor  ( new_n13044_, new_n12735_, new_n12733_ );
xor  ( new_n13045_, new_n13044_, new_n12739_ );
or   ( new_n13046_, new_n13045_, new_n13043_ );
and  ( new_n13047_, new_n13046_, new_n13042_ );
or   ( new_n13048_, new_n13047_, new_n12750_ );
and  ( new_n13049_, new_n13047_, new_n12750_ );
xor  ( new_n13050_, new_n12191_, new_n12181_ );
xor  ( new_n13051_, new_n13050_, new_n12447_ );
or   ( new_n13052_, new_n13051_, new_n13049_ );
and  ( new_n13053_, new_n13052_, new_n13048_ );
nor  ( new_n13054_, new_n13053_, new_n12748_ );
xor  ( new_n13055_, new_n13041_, new_n13039_ );
xor  ( new_n13056_, new_n13055_, new_n13045_ );
xor  ( new_n13057_, new_n12756_, new_n12754_ );
xor  ( new_n13058_, new_n13057_, new_n12760_ );
xor  ( new_n13059_, new_n12620_, new_n12568_ );
xor  ( new_n13060_, new_n13059_, new_n12675_ );
xor  ( new_n13061_, new_n12502_, new_n12492_ );
xor  ( new_n13062_, new_n13061_, new_n12514_ );
nand ( new_n13063_, new_n13062_, new_n13060_ );
nor  ( new_n13064_, new_n13062_, new_n13060_ );
xor  ( new_n13065_, new_n12794_, new_n12792_ );
xor  ( new_n13066_, new_n13065_, new_n12798_ );
or   ( new_n13067_, new_n13066_, new_n13064_ );
and  ( new_n13068_, new_n13067_, new_n13063_ );
or   ( new_n13069_, new_n13068_, new_n13058_ );
and  ( new_n13070_, new_n13068_, new_n13058_ );
xnor ( new_n13071_, new_n12770_, new_n12768_ );
xor  ( new_n13072_, new_n13071_, new_n12774_ );
xnor ( new_n13073_, new_n12782_, new_n12780_ );
xor  ( new_n13074_, new_n13073_, new_n12786_ );
nand ( new_n13075_, new_n13074_, new_n13072_ );
nor  ( new_n13076_, new_n13074_, new_n13072_ );
xor  ( new_n13077_, new_n13022_, new_n13006_ );
xor  ( new_n13078_, new_n13077_, new_n13029_ );
xnor ( new_n13079_, new_n12852_, new_n12836_ );
xor  ( new_n13080_, new_n13079_, new_n12870_ );
or   ( new_n13081_, new_n13080_, new_n13078_ );
and  ( new_n13082_, new_n13080_, new_n13078_ );
xnor ( new_n13083_, new_n12955_, new_n12939_ );
xor  ( new_n13084_, new_n13083_, new_n12973_ );
or   ( new_n13085_, new_n13084_, new_n13082_ );
and  ( new_n13086_, new_n13085_, new_n13081_ );
or   ( new_n13087_, new_n13086_, new_n13076_ );
and  ( new_n13088_, new_n13087_, new_n13075_ );
xor  ( new_n13089_, new_n13000_, new_n12990_ );
xor  ( new_n13090_, new_n13089_, new_n13031_ );
xnor ( new_n13091_, new_n12922_, new_n12872_ );
xor  ( new_n13092_, new_n13091_, new_n12975_ );
or   ( new_n13093_, new_n13092_, new_n13090_ );
and  ( new_n13094_, new_n13092_, new_n13090_ );
xor  ( new_n13095_, new_n12814_, new_n12804_ );
xor  ( new_n13096_, new_n13095_, new_n12818_ );
or   ( new_n13097_, new_n13096_, new_n13094_ );
and  ( new_n13098_, new_n13097_, new_n13093_ );
and  ( new_n13099_, new_n13098_, new_n13088_ );
nor  ( new_n13100_, new_n13098_, new_n13088_ );
xnor ( new_n13101_, new_n12984_, new_n12982_ );
xor  ( new_n13102_, new_n13101_, new_n12988_ );
xnor ( new_n13103_, new_n12808_, new_n12806_ );
xor  ( new_n13104_, new_n13103_, new_n12812_ );
or   ( new_n13105_, new_n13104_, new_n13102_ );
and  ( new_n13106_, new_n13104_, new_n13102_ );
xor  ( new_n13107_, new_n12994_, new_n12992_ );
xnor ( new_n13108_, new_n13107_, new_n12998_ );
or   ( new_n13109_, new_n13108_, new_n13106_ );
and  ( new_n13110_, new_n13109_, new_n13105_ );
or   ( new_n13111_, new_n3117_, new_n4267_ );
or   ( new_n13112_, new_n3119_, new_n4069_ );
and  ( new_n13113_, new_n13112_, new_n13111_ );
xor  ( new_n13114_, new_n13113_, new_n2800_ );
or   ( new_n13115_, new_n2807_, new_n4995_ );
or   ( new_n13116_, new_n2809_, new_n4603_ );
and  ( new_n13117_, new_n13116_, new_n13115_ );
xor  ( new_n13118_, new_n13117_, new_n2424_ );
or   ( new_n13119_, new_n13118_, new_n13114_ );
and  ( new_n13120_, new_n13118_, new_n13114_ );
or   ( new_n13121_, new_n2425_, new_n5171_ );
or   ( new_n13122_, new_n2427_, new_n4859_ );
and  ( new_n13123_, new_n13122_, new_n13121_ );
xor  ( new_n13124_, new_n13123_, new_n2121_ );
or   ( new_n13125_, new_n13124_, new_n13120_ );
and  ( new_n13126_, new_n13125_, new_n13119_ );
or   ( new_n13127_, new_n5604_, new_n2178_ );
or   ( new_n13128_, new_n5606_, new_n2057_ );
and  ( new_n13129_, new_n13128_, new_n13127_ );
xor  ( new_n13130_, new_n13129_, new_n5206_ );
or   ( new_n13131_, new_n5207_, new_n2475_ );
or   ( new_n13132_, new_n5209_, new_n2291_ );
and  ( new_n13133_, new_n13132_, new_n13131_ );
xor  ( new_n13134_, new_n13133_, new_n4708_ );
or   ( new_n13135_, new_n13134_, new_n13130_ );
and  ( new_n13136_, new_n13134_, new_n13130_ );
or   ( new_n13137_, new_n4709_, new_n2751_ );
or   ( new_n13138_, new_n4711_, new_n2646_ );
and  ( new_n13139_, new_n13138_, new_n13137_ );
xor  ( new_n13140_, new_n13139_, new_n4295_ );
or   ( new_n13141_, new_n13140_, new_n13136_ );
and  ( new_n13142_, new_n13141_, new_n13135_ );
or   ( new_n13143_, new_n13142_, new_n13126_ );
and  ( new_n13144_, new_n13142_, new_n13126_ );
or   ( new_n13145_, new_n4302_, new_n3178_ );
or   ( new_n13146_, new_n4304_, new_n2981_ );
and  ( new_n13147_, new_n13146_, new_n13145_ );
xor  ( new_n13148_, new_n13147_, new_n3895_ );
or   ( new_n13149_, new_n3896_, new_n3696_ );
or   ( new_n13150_, new_n3898_, new_n3306_ );
and  ( new_n13151_, new_n13150_, new_n13149_ );
xor  ( new_n13152_, new_n13151_, new_n3460_ );
nor  ( new_n13153_, new_n13152_, new_n13148_ );
and  ( new_n13154_, new_n13152_, new_n13148_ );
or   ( new_n13155_, new_n3461_, new_n3820_ );
or   ( new_n13156_, new_n3463_, new_n3694_ );
and  ( new_n13157_, new_n13156_, new_n13155_ );
xor  ( new_n13158_, new_n13157_, new_n3116_ );
nor  ( new_n13159_, new_n13158_, new_n13154_ );
nor  ( new_n13160_, new_n13159_, new_n13153_ );
or   ( new_n13161_, new_n13160_, new_n13144_ );
and  ( new_n13162_, new_n13161_, new_n13143_ );
or   ( new_n13163_, new_n1364_, new_n7149_ );
or   ( new_n13164_, new_n1366_, new_n6943_ );
and  ( new_n13165_, new_n13164_, new_n13163_ );
xor  ( new_n13166_, new_n13165_, new_n1129_ );
or   ( new_n13167_, new_n1135_, new_n8117_ );
or   ( new_n13168_, new_n1137_, new_n7373_ );
and  ( new_n13169_, new_n13168_, new_n13167_ );
xor  ( new_n13170_, new_n13169_, new_n896_ );
or   ( new_n13171_, new_n13170_, new_n13166_ );
and  ( new_n13172_, new_n13170_, new_n13166_ );
or   ( new_n13173_, new_n897_, new_n8352_ );
or   ( new_n13174_, new_n899_, new_n8115_ );
and  ( new_n13175_, new_n13174_, new_n13173_ );
xor  ( new_n13176_, new_n13175_, new_n748_ );
or   ( new_n13177_, new_n13176_, new_n13172_ );
and  ( new_n13178_, new_n13177_, new_n13171_ );
or   ( new_n13179_, new_n755_, new_n8995_ );
or   ( new_n13180_, new_n757_, new_n8481_ );
and  ( new_n13181_, new_n13180_, new_n13179_ );
xor  ( new_n13182_, new_n13181_, new_n523_ );
or   ( new_n13183_, new_n524_, new_n9681_ );
or   ( new_n13184_, new_n526_, new_n9099_ );
and  ( new_n13185_, new_n13184_, new_n13183_ );
xor  ( new_n13186_, new_n13185_, new_n403_ );
or   ( new_n13187_, new_n13186_, new_n13182_ );
and  ( new_n13188_, new_n13186_, new_n13182_ );
or   ( new_n13189_, new_n409_, new_n10220_ );
or   ( new_n13190_, new_n411_, new_n9679_ );
and  ( new_n13191_, new_n13190_, new_n13189_ );
xor  ( new_n13192_, new_n13191_, new_n328_ );
or   ( new_n13193_, new_n13192_, new_n13188_ );
and  ( new_n13194_, new_n13193_, new_n13187_ );
or   ( new_n13195_, new_n13194_, new_n13178_ );
and  ( new_n13196_, new_n13194_, new_n13178_ );
or   ( new_n13197_, new_n2122_, new_n5570_ );
or   ( new_n13198_, new_n2124_, new_n5428_ );
and  ( new_n13199_, new_n13198_, new_n13197_ );
xor  ( new_n13200_, new_n13199_, new_n1843_ );
or   ( new_n13201_, new_n1844_, new_n6219_ );
or   ( new_n13202_, new_n1846_, new_n5899_ );
and  ( new_n13203_, new_n13202_, new_n13201_ );
xor  ( new_n13204_, new_n13203_, new_n1586_ );
nor  ( new_n13205_, new_n13204_, new_n13200_ );
and  ( new_n13206_, new_n13204_, new_n13200_ );
or   ( new_n13207_, new_n1593_, new_n6589_ );
or   ( new_n13208_, new_n1595_, new_n6425_ );
and  ( new_n13209_, new_n13208_, new_n13207_ );
xor  ( new_n13210_, new_n13209_, new_n1358_ );
nor  ( new_n13211_, new_n13210_, new_n13206_ );
nor  ( new_n13212_, new_n13211_, new_n13205_ );
or   ( new_n13213_, new_n13212_, new_n13196_ );
and  ( new_n13214_, new_n13213_, new_n13195_ );
or   ( new_n13215_, new_n13214_, new_n13162_ );
or   ( new_n13216_, new_n10059_, new_n419_ );
or   ( new_n13217_, new_n10061_, new_n348_ );
and  ( new_n13218_, new_n13217_, new_n13216_ );
xor  ( new_n13219_, new_n13218_, new_n9421_ );
and  ( new_n13220_, RIbb2d888_64, RIbb2d450_73 );
or   ( new_n13221_, RIbb2d888_64, new_n264_ );
and  ( new_n13222_, new_n13221_, RIbb2d900_63 );
or   ( new_n13223_, new_n13222_, new_n13220_ );
or   ( new_n13224_, new_n10770_, new_n270_ );
and  ( new_n13225_, new_n13224_, new_n13223_ );
or   ( new_n13226_, new_n13225_, new_n13219_ );
and  ( new_n13227_, new_n13225_, new_n13219_ );
or   ( new_n13228_, new_n9422_, new_n509_ );
or   ( new_n13229_, new_n9424_, new_n443_ );
and  ( new_n13230_, new_n13229_, new_n13228_ );
xor  ( new_n13231_, new_n13230_, new_n8873_ );
or   ( new_n13232_, new_n13231_, new_n13227_ );
and  ( new_n13233_, new_n13232_, new_n13226_ );
or   ( new_n13234_, new_n7184_, new_n1318_ );
or   ( new_n13235_, new_n7186_, new_n1213_ );
and  ( new_n13236_, new_n13235_, new_n13234_ );
xor  ( new_n13237_, new_n13236_, new_n6638_ );
or   ( new_n13238_, new_n6645_, new_n1523_ );
or   ( new_n13239_, new_n6647_, new_n1525_ );
and  ( new_n13240_, new_n13239_, new_n13238_ );
xor  ( new_n13241_, new_n13240_, new_n6166_ );
or   ( new_n13242_, new_n13241_, new_n13237_ );
and  ( new_n13243_, new_n13241_, new_n13237_ );
or   ( new_n13244_, new_n6173_, new_n1899_ );
or   ( new_n13245_, new_n6175_, new_n1754_ );
and  ( new_n13246_, new_n13245_, new_n13244_ );
xor  ( new_n13247_, new_n13246_, new_n5597_ );
or   ( new_n13248_, new_n13247_, new_n13243_ );
and  ( new_n13249_, new_n13248_, new_n13242_ );
nor  ( new_n13250_, new_n13249_, new_n13233_ );
and  ( new_n13251_, new_n13249_, new_n13233_ );
or   ( new_n13252_, new_n8874_, new_n775_ );
or   ( new_n13253_, new_n8876_, new_n515_ );
and  ( new_n13254_, new_n13253_, new_n13252_ );
xor  ( new_n13255_, new_n13254_, new_n8257_ );
or   ( new_n13256_, new_n8264_, new_n886_ );
or   ( new_n13257_, new_n8266_, new_n805_ );
and  ( new_n13258_, new_n13257_, new_n13256_ );
xor  ( new_n13259_, new_n13258_, new_n7725_ );
nor  ( new_n13260_, new_n13259_, new_n13255_ );
and  ( new_n13261_, new_n13259_, new_n13255_ );
or   ( new_n13262_, new_n7732_, new_n1168_ );
or   ( new_n13263_, new_n7734_, new_n986_ );
and  ( new_n13264_, new_n13263_, new_n13262_ );
xor  ( new_n13265_, new_n13264_, new_n7177_ );
nor  ( new_n13266_, new_n13265_, new_n13261_ );
nor  ( new_n13267_, new_n13266_, new_n13260_ );
nor  ( new_n13268_, new_n13267_, new_n13251_ );
nor  ( new_n13269_, new_n13268_, new_n13250_ );
and  ( new_n13270_, new_n13214_, new_n13162_ );
or   ( new_n13271_, new_n13270_, new_n13269_ );
and  ( new_n13272_, new_n13271_, new_n13215_ );
nor  ( new_n13273_, new_n13272_, new_n13110_ );
and  ( new_n13274_, new_n13272_, new_n13110_ );
not  ( new_n13275_, new_n13274_ );
xnor ( new_n13276_, new_n12844_, new_n12840_ );
xor  ( new_n13277_, new_n13276_, new_n12850_ );
xnor ( new_n13278_, new_n12862_, new_n12858_ );
xor  ( new_n13279_, new_n13278_, new_n12868_ );
or   ( new_n13280_, new_n13279_, new_n13277_ );
and  ( new_n13281_, new_n13279_, new_n13277_ );
xor  ( new_n13282_, new_n12965_, new_n12961_ );
xnor ( new_n13283_, new_n13282_, new_n12971_ );
or   ( new_n13284_, new_n13283_, new_n13281_ );
and  ( new_n13285_, new_n13284_, new_n13280_ );
xnor ( new_n13286_, new_n12947_, new_n12943_ );
xor  ( new_n13287_, new_n13286_, new_n12953_ );
xnor ( new_n13288_, new_n13014_, new_n13010_ );
xor  ( new_n13289_, new_n13288_, new_n13020_ );
or   ( new_n13290_, new_n13289_, new_n13287_ );
and  ( new_n13291_, new_n13289_, new_n13287_ );
xor  ( new_n13292_, new_n12931_, new_n12927_ );
xnor ( new_n13293_, new_n13292_, new_n12937_ );
or   ( new_n13294_, new_n13293_, new_n13291_ );
and  ( new_n13295_, new_n13294_, new_n13290_ );
nor  ( new_n13296_, new_n13295_, new_n13285_ );
and  ( new_n13297_, new_n13295_, new_n13285_ );
xnor ( new_n13298_, new_n12880_, new_n12876_ );
xor  ( new_n13299_, new_n13298_, new_n12886_ );
xnor ( new_n13300_, new_n12910_, new_n12906_ );
xor  ( new_n13301_, new_n13300_, new_n12916_ );
nor  ( new_n13302_, new_n13301_, new_n13299_ );
and  ( new_n13303_, new_n13301_, new_n13299_ );
xor  ( new_n13304_, new_n12828_, new_n12824_ );
xnor ( new_n13305_, new_n13304_, new_n12834_ );
nor  ( new_n13306_, new_n13305_, new_n13303_ );
nor  ( new_n13307_, new_n13306_, new_n13302_ );
nor  ( new_n13308_, new_n13307_, new_n13297_ );
nor  ( new_n13309_, new_n13308_, new_n13296_ );
and  ( new_n13310_, new_n13309_, new_n13275_ );
nor  ( new_n13311_, new_n13310_, new_n13273_ );
nor  ( new_n13312_, new_n13311_, new_n13100_ );
nor  ( new_n13313_, new_n13312_, new_n13099_ );
not  ( new_n13314_, new_n13313_ );
or   ( new_n13315_, new_n13314_, new_n13070_ );
and  ( new_n13316_, new_n13315_, new_n13069_ );
xor  ( new_n13317_, new_n12692_, new_n12480_ );
xor  ( new_n13318_, new_n13317_, new_n12713_ );
or   ( new_n13319_, new_n13318_, new_n13316_ );
and  ( new_n13320_, new_n13318_, new_n13316_ );
xor  ( new_n13321_, new_n12762_, new_n12752_ );
xor  ( new_n13322_, new_n13321_, new_n13037_ );
or   ( new_n13323_, new_n13322_, new_n13320_ );
and  ( new_n13324_, new_n13323_, new_n13319_ );
nor  ( new_n13325_, new_n13324_, new_n13056_ );
xnor ( new_n13326_, new_n13047_, new_n12750_ );
xor  ( new_n13327_, new_n13326_, new_n13051_ );
and  ( new_n13328_, new_n13327_, new_n13325_ );
xor  ( new_n13329_, new_n12800_, new_n12790_ );
xor  ( new_n13330_, new_n13329_, new_n13035_ );
xor  ( new_n13331_, new_n12978_, new_n12820_ );
xor  ( new_n13332_, new_n13331_, new_n13033_ );
xnor ( new_n13333_, new_n13098_, new_n13088_ );
xor  ( new_n13334_, new_n13333_, new_n13311_ );
or   ( new_n13335_, new_n13334_, new_n13332_ );
and  ( new_n13336_, new_n13334_, new_n13332_ );
xor  ( new_n13337_, new_n13062_, new_n13060_ );
xor  ( new_n13338_, new_n13337_, new_n13066_ );
or   ( new_n13339_, new_n13338_, new_n13336_ );
and  ( new_n13340_, new_n13339_, new_n13335_ );
nor  ( new_n13341_, new_n13340_, new_n13330_ );
and  ( new_n13342_, new_n13340_, new_n13330_ );
xor  ( new_n13343_, new_n12776_, new_n12766_ );
xor  ( new_n13344_, new_n13343_, new_n12788_ );
xor  ( new_n13345_, new_n13272_, new_n13110_ );
xor  ( new_n13346_, new_n13345_, new_n13309_ );
xor  ( new_n13347_, new_n13092_, new_n13090_ );
xor  ( new_n13348_, new_n13347_, new_n13096_ );
or   ( new_n13349_, new_n13348_, new_n13346_ );
and  ( new_n13350_, new_n13348_, new_n13346_ );
xor  ( new_n13351_, new_n13074_, new_n13072_ );
xor  ( new_n13352_, new_n13351_, new_n13086_ );
or   ( new_n13353_, new_n13352_, new_n13350_ );
and  ( new_n13354_, new_n13353_, new_n13349_ );
nor  ( new_n13355_, new_n13354_, new_n13344_ );
and  ( new_n13356_, new_n13354_, new_n13344_ );
xnor ( new_n13357_, new_n12918_, new_n12902_ );
xor  ( new_n13358_, new_n13357_, new_n12888_ );
xnor ( new_n13359_, new_n13142_, new_n13126_ );
xor  ( new_n13360_, new_n13359_, new_n13160_ );
xnor ( new_n13361_, new_n13194_, new_n13178_ );
xor  ( new_n13362_, new_n13361_, new_n13212_ );
or   ( new_n13363_, new_n13362_, new_n13360_ );
and  ( new_n13364_, new_n13362_, new_n13360_ );
xor  ( new_n13365_, new_n13289_, new_n13287_ );
xnor ( new_n13366_, new_n13365_, new_n13293_ );
not  ( new_n13367_, new_n13366_ );
or   ( new_n13368_, new_n13367_, new_n13364_ );
and  ( new_n13369_, new_n13368_, new_n13363_ );
or   ( new_n13370_, new_n13369_, new_n13358_ );
and  ( new_n13371_, new_n13369_, new_n13358_ );
xor  ( new_n13372_, new_n13080_, new_n13078_ );
xor  ( new_n13373_, new_n13372_, new_n13084_ );
or   ( new_n13374_, new_n13373_, new_n13371_ );
and  ( new_n13375_, new_n13374_, new_n13370_ );
xor  ( new_n13376_, new_n13295_, new_n13285_ );
xor  ( new_n13377_, new_n13376_, new_n13307_ );
xnor ( new_n13378_, new_n13214_, new_n13162_ );
xor  ( new_n13379_, new_n13378_, new_n13269_ );
or   ( new_n13380_, new_n13379_, new_n13377_ );
and  ( new_n13381_, new_n13379_, new_n13377_ );
xnor ( new_n13382_, new_n13104_, new_n13102_ );
xor  ( new_n13383_, new_n13382_, new_n13108_ );
or   ( new_n13384_, new_n13383_, new_n13381_ );
and  ( new_n13385_, new_n13384_, new_n13380_ );
nor  ( new_n13386_, new_n13385_, new_n13375_ );
and  ( new_n13387_, new_n13385_, new_n13375_ );
xor  ( new_n13388_, new_n12898_, new_n12892_ );
xor  ( new_n13389_, new_n13388_, new_n311_ );
xnor ( new_n13390_, new_n13301_, new_n13299_ );
xor  ( new_n13391_, new_n13390_, new_n13305_ );
and  ( new_n13392_, new_n13391_, new_n13389_ );
or   ( new_n13393_, new_n13391_, new_n13389_ );
xor  ( new_n13394_, new_n13279_, new_n13277_ );
xnor ( new_n13395_, new_n13394_, new_n13283_ );
and  ( new_n13396_, new_n13395_, new_n13393_ );
or   ( new_n13397_, new_n13396_, new_n13392_ );
or   ( new_n13398_, new_n2425_, new_n5428_ );
or   ( new_n13399_, new_n2427_, new_n5171_ );
and  ( new_n13400_, new_n13399_, new_n13398_ );
xor  ( new_n13401_, new_n13400_, new_n2121_ );
or   ( new_n13402_, new_n2122_, new_n5899_ );
or   ( new_n13403_, new_n2124_, new_n5570_ );
and  ( new_n13404_, new_n13403_, new_n13402_ );
xor  ( new_n13405_, new_n13404_, new_n1843_ );
or   ( new_n13406_, new_n13405_, new_n13401_ );
and  ( new_n13407_, new_n13405_, new_n13401_ );
or   ( new_n13408_, new_n1844_, new_n6425_ );
or   ( new_n13409_, new_n1846_, new_n6219_ );
and  ( new_n13410_, new_n13409_, new_n13408_ );
xor  ( new_n13411_, new_n13410_, new_n1586_ );
or   ( new_n13412_, new_n13411_, new_n13407_ );
and  ( new_n13413_, new_n13412_, new_n13406_ );
or   ( new_n13414_, new_n897_, new_n8481_ );
or   ( new_n13415_, new_n899_, new_n8352_ );
and  ( new_n13416_, new_n13415_, new_n13414_ );
xor  ( new_n13417_, new_n13416_, new_n748_ );
or   ( new_n13418_, new_n755_, new_n9099_ );
or   ( new_n13419_, new_n757_, new_n8995_ );
and  ( new_n13420_, new_n13419_, new_n13418_ );
xor  ( new_n13421_, new_n13420_, new_n523_ );
or   ( new_n13422_, new_n13421_, new_n13417_ );
and  ( new_n13423_, new_n13421_, new_n13417_ );
or   ( new_n13424_, new_n524_, new_n9679_ );
or   ( new_n13425_, new_n526_, new_n9681_ );
and  ( new_n13426_, new_n13425_, new_n13424_ );
xor  ( new_n13427_, new_n13426_, new_n403_ );
or   ( new_n13428_, new_n13427_, new_n13423_ );
and  ( new_n13429_, new_n13428_, new_n13422_ );
or   ( new_n13430_, new_n13429_, new_n13413_ );
and  ( new_n13431_, new_n13429_, new_n13413_ );
or   ( new_n13432_, new_n1593_, new_n6943_ );
or   ( new_n13433_, new_n1595_, new_n6589_ );
and  ( new_n13434_, new_n13433_, new_n13432_ );
xor  ( new_n13435_, new_n13434_, new_n1358_ );
or   ( new_n13436_, new_n1364_, new_n7373_ );
or   ( new_n13437_, new_n1366_, new_n7149_ );
and  ( new_n13438_, new_n13437_, new_n13436_ );
xor  ( new_n13439_, new_n13438_, new_n1129_ );
nor  ( new_n13440_, new_n13439_, new_n13435_ );
and  ( new_n13441_, new_n13439_, new_n13435_ );
or   ( new_n13442_, new_n1135_, new_n8115_ );
or   ( new_n13443_, new_n1137_, new_n8117_ );
and  ( new_n13444_, new_n13443_, new_n13442_ );
xor  ( new_n13445_, new_n13444_, new_n896_ );
nor  ( new_n13446_, new_n13445_, new_n13441_ );
nor  ( new_n13447_, new_n13446_, new_n13440_ );
or   ( new_n13448_, new_n13447_, new_n13431_ );
and  ( new_n13449_, new_n13448_, new_n13430_ );
or   ( new_n13450_, new_n7732_, new_n1213_ );
or   ( new_n13451_, new_n7734_, new_n1168_ );
and  ( new_n13452_, new_n13451_, new_n13450_ );
xor  ( new_n13453_, new_n13452_, new_n7177_ );
or   ( new_n13454_, new_n7184_, new_n1525_ );
or   ( new_n13455_, new_n7186_, new_n1318_ );
and  ( new_n13456_, new_n13455_, new_n13454_ );
xor  ( new_n13457_, new_n13456_, new_n6638_ );
or   ( new_n13458_, new_n13457_, new_n13453_ );
and  ( new_n13459_, new_n13457_, new_n13453_ );
or   ( new_n13460_, new_n6645_, new_n1754_ );
or   ( new_n13461_, new_n6647_, new_n1523_ );
and  ( new_n13462_, new_n13461_, new_n13460_ );
xor  ( new_n13463_, new_n13462_, new_n6166_ );
or   ( new_n13464_, new_n13463_, new_n13459_ );
and  ( new_n13465_, new_n13464_, new_n13458_ );
or   ( new_n13466_, new_n10059_, new_n443_ );
or   ( new_n13467_, new_n10061_, new_n419_ );
and  ( new_n13468_, new_n13467_, new_n13466_ );
xor  ( new_n13469_, new_n13468_, new_n9421_ );
and  ( new_n13470_, RIbb2d888_64, RIbb2d3d8_74 );
or   ( new_n13471_, RIbb2d888_64, new_n348_ );
and  ( new_n13472_, new_n13471_, RIbb2d900_63 );
or   ( new_n13473_, new_n13472_, new_n13470_ );
or   ( new_n13474_, new_n10770_, new_n264_ );
and  ( new_n13475_, new_n13474_, new_n13473_ );
nor  ( new_n13476_, new_n13475_, new_n13469_ );
and  ( new_n13477_, new_n13475_, new_n13469_ );
nor  ( new_n13478_, new_n13477_, new_n331_ );
nor  ( new_n13479_, new_n13478_, new_n13476_ );
or   ( new_n13480_, new_n9422_, new_n515_ );
or   ( new_n13481_, new_n9424_, new_n509_ );
and  ( new_n13482_, new_n13481_, new_n13480_ );
xor  ( new_n13483_, new_n13482_, new_n8873_ );
or   ( new_n13484_, new_n8874_, new_n805_ );
or   ( new_n13485_, new_n8876_, new_n775_ );
and  ( new_n13486_, new_n13485_, new_n13484_ );
xor  ( new_n13487_, new_n13486_, new_n8257_ );
or   ( new_n13488_, new_n13487_, new_n13483_ );
and  ( new_n13489_, new_n13487_, new_n13483_ );
or   ( new_n13490_, new_n8264_, new_n986_ );
or   ( new_n13491_, new_n8266_, new_n886_ );
and  ( new_n13492_, new_n13491_, new_n13490_ );
xor  ( new_n13493_, new_n13492_, new_n7725_ );
or   ( new_n13494_, new_n13493_, new_n13489_ );
and  ( new_n13495_, new_n13494_, new_n13488_ );
and  ( new_n13496_, new_n13495_, new_n13479_ );
or   ( new_n13497_, new_n13496_, new_n13465_ );
or   ( new_n13498_, new_n13495_, new_n13479_ );
and  ( new_n13499_, new_n13498_, new_n13497_ );
or   ( new_n13500_, new_n13499_, new_n13449_ );
or   ( new_n13501_, new_n4709_, new_n2981_ );
or   ( new_n13502_, new_n4711_, new_n2751_ );
and  ( new_n13503_, new_n13502_, new_n13501_ );
xor  ( new_n13504_, new_n13503_, new_n4295_ );
or   ( new_n13505_, new_n4302_, new_n3306_ );
or   ( new_n13506_, new_n4304_, new_n3178_ );
and  ( new_n13507_, new_n13506_, new_n13505_ );
xor  ( new_n13508_, new_n13507_, new_n3895_ );
or   ( new_n13509_, new_n13508_, new_n13504_ );
and  ( new_n13510_, new_n13508_, new_n13504_ );
or   ( new_n13511_, new_n3896_, new_n3694_ );
or   ( new_n13512_, new_n3898_, new_n3696_ );
and  ( new_n13513_, new_n13512_, new_n13511_ );
xor  ( new_n13514_, new_n13513_, new_n3460_ );
or   ( new_n13515_, new_n13514_, new_n13510_ );
and  ( new_n13516_, new_n13515_, new_n13509_ );
or   ( new_n13517_, new_n3461_, new_n4069_ );
or   ( new_n13518_, new_n3463_, new_n3820_ );
and  ( new_n13519_, new_n13518_, new_n13517_ );
xor  ( new_n13520_, new_n13519_, new_n3116_ );
or   ( new_n13521_, new_n3117_, new_n4603_ );
or   ( new_n13522_, new_n3119_, new_n4267_ );
and  ( new_n13523_, new_n13522_, new_n13521_ );
xor  ( new_n13524_, new_n13523_, new_n2800_ );
or   ( new_n13525_, new_n13524_, new_n13520_ );
and  ( new_n13526_, new_n13524_, new_n13520_ );
or   ( new_n13527_, new_n2807_, new_n4859_ );
or   ( new_n13528_, new_n2809_, new_n4995_ );
and  ( new_n13529_, new_n13528_, new_n13527_ );
xor  ( new_n13530_, new_n13529_, new_n2424_ );
or   ( new_n13531_, new_n13530_, new_n13526_ );
and  ( new_n13532_, new_n13531_, new_n13525_ );
or   ( new_n13533_, new_n13532_, new_n13516_ );
and  ( new_n13534_, new_n13532_, new_n13516_ );
or   ( new_n13535_, new_n6173_, new_n2057_ );
or   ( new_n13536_, new_n6175_, new_n1899_ );
and  ( new_n13537_, new_n13536_, new_n13535_ );
xor  ( new_n13538_, new_n13537_, new_n5597_ );
or   ( new_n13539_, new_n5604_, new_n2291_ );
or   ( new_n13540_, new_n5606_, new_n2178_ );
and  ( new_n13541_, new_n13540_, new_n13539_ );
xor  ( new_n13542_, new_n13541_, new_n5206_ );
nor  ( new_n13543_, new_n13542_, new_n13538_ );
and  ( new_n13544_, new_n13542_, new_n13538_ );
or   ( new_n13545_, new_n5207_, new_n2646_ );
or   ( new_n13546_, new_n5209_, new_n2475_ );
and  ( new_n13547_, new_n13546_, new_n13545_ );
xor  ( new_n13548_, new_n13547_, new_n4708_ );
nor  ( new_n13549_, new_n13548_, new_n13544_ );
nor  ( new_n13550_, new_n13549_, new_n13543_ );
or   ( new_n13551_, new_n13550_, new_n13534_ );
and  ( new_n13552_, new_n13551_, new_n13533_ );
and  ( new_n13553_, new_n13499_, new_n13449_ );
or   ( new_n13554_, new_n13553_, new_n13552_ );
and  ( new_n13555_, new_n13554_, new_n13500_ );
and  ( new_n13556_, new_n13555_, new_n13397_ );
nor  ( new_n13557_, new_n13555_, new_n13397_ );
or   ( new_n13558_, new_n337_, new_n10841_ );
or   ( new_n13559_, new_n340_, new_n10541_ );
and  ( new_n13560_, new_n13559_, new_n13558_ );
xor  ( new_n13561_, new_n13560_, new_n331_ );
xnor ( new_n13562_, new_n13186_, new_n13182_ );
xor  ( new_n13563_, new_n13562_, new_n13192_ );
and  ( new_n13564_, new_n13563_, new_n13561_ );
or   ( new_n13565_, new_n13563_, new_n13561_ );
xor  ( new_n13566_, new_n13170_, new_n13166_ );
xnor ( new_n13567_, new_n13566_, new_n13176_ );
and  ( new_n13568_, new_n13567_, new_n13565_ );
or   ( new_n13569_, new_n13568_, new_n13564_ );
xnor ( new_n13570_, new_n13118_, new_n13114_ );
xor  ( new_n13571_, new_n13570_, new_n13124_ );
xnor ( new_n13572_, new_n13152_, new_n13148_ );
xor  ( new_n13573_, new_n13572_, new_n13158_ );
or   ( new_n13574_, new_n13573_, new_n13571_ );
and  ( new_n13575_, new_n13573_, new_n13571_ );
xor  ( new_n13576_, new_n13204_, new_n13200_ );
xnor ( new_n13577_, new_n13576_, new_n13210_ );
or   ( new_n13578_, new_n13577_, new_n13575_ );
and  ( new_n13579_, new_n13578_, new_n13574_ );
nor  ( new_n13580_, new_n13579_, new_n13569_ );
and  ( new_n13581_, new_n13579_, new_n13569_ );
xnor ( new_n13582_, new_n13134_, new_n13130_ );
xor  ( new_n13583_, new_n13582_, new_n13140_ );
xnor ( new_n13584_, new_n13241_, new_n13237_ );
xor  ( new_n13585_, new_n13584_, new_n13247_ );
nor  ( new_n13586_, new_n13585_, new_n13583_ );
and  ( new_n13587_, new_n13585_, new_n13583_ );
xor  ( new_n13588_, new_n13259_, new_n13255_ );
xnor ( new_n13589_, new_n13588_, new_n13265_ );
nor  ( new_n13590_, new_n13589_, new_n13587_ );
nor  ( new_n13591_, new_n13590_, new_n13586_ );
nor  ( new_n13592_, new_n13591_, new_n13581_ );
nor  ( new_n13593_, new_n13592_, new_n13580_ );
nor  ( new_n13594_, new_n13593_, new_n13557_ );
nor  ( new_n13595_, new_n13594_, new_n13556_ );
nor  ( new_n13596_, new_n13595_, new_n13387_ );
nor  ( new_n13597_, new_n13596_, new_n13386_ );
nor  ( new_n13598_, new_n13597_, new_n13356_ );
nor  ( new_n13599_, new_n13598_, new_n13355_ );
nor  ( new_n13600_, new_n13599_, new_n13342_ );
nor  ( new_n13601_, new_n13600_, new_n13341_ );
xnor ( new_n13602_, new_n13318_, new_n13316_ );
xnor ( new_n13603_, new_n13602_, new_n13322_ );
nor  ( new_n13604_, new_n13603_, new_n13601_ );
xor  ( new_n13605_, new_n13324_, new_n13056_ );
and  ( new_n13606_, new_n13605_, new_n13604_ );
xnor ( new_n13607_, new_n13603_, new_n13601_ );
xor  ( new_n13608_, new_n13340_, new_n13330_ );
xor  ( new_n13609_, new_n13608_, new_n13599_ );
xor  ( new_n13610_, new_n13348_, new_n13346_ );
xor  ( new_n13611_, new_n13610_, new_n13352_ );
xor  ( new_n13612_, new_n13555_, new_n13397_ );
xor  ( new_n13613_, new_n13612_, new_n13593_ );
xor  ( new_n13614_, new_n13369_, new_n13358_ );
xor  ( new_n13615_, new_n13614_, new_n13373_ );
or   ( new_n13616_, new_n13615_, new_n13613_ );
and  ( new_n13617_, new_n13615_, new_n13613_ );
xor  ( new_n13618_, new_n13379_, new_n13377_ );
xor  ( new_n13619_, new_n13618_, new_n13383_ );
or   ( new_n13620_, new_n13619_, new_n13617_ );
and  ( new_n13621_, new_n13620_, new_n13616_ );
or   ( new_n13622_, new_n13621_, new_n13611_ );
and  ( new_n13623_, new_n13621_, new_n13611_ );
xnor ( new_n13624_, new_n13249_, new_n13233_ );
xor  ( new_n13625_, new_n13624_, new_n13267_ );
xnor ( new_n13626_, new_n13429_, new_n13413_ );
xor  ( new_n13627_, new_n13626_, new_n13447_ );
xnor ( new_n13628_, new_n13532_, new_n13516_ );
xor  ( new_n13629_, new_n13628_, new_n13550_ );
or   ( new_n13630_, new_n13629_, new_n13627_ );
and  ( new_n13631_, new_n13629_, new_n13627_ );
xor  ( new_n13632_, new_n13563_, new_n13561_ );
xor  ( new_n13633_, new_n13632_, new_n13567_ );
or   ( new_n13634_, new_n13633_, new_n13631_ );
and  ( new_n13635_, new_n13634_, new_n13630_ );
or   ( new_n13636_, new_n13635_, new_n13625_ );
and  ( new_n13637_, new_n13635_, new_n13625_ );
xor  ( new_n13638_, new_n13362_, new_n13360_ );
xor  ( new_n13639_, new_n13638_, new_n13367_ );
or   ( new_n13640_, new_n13639_, new_n13637_ );
and  ( new_n13641_, new_n13640_, new_n13636_ );
xor  ( new_n13642_, new_n13499_, new_n13449_ );
xor  ( new_n13643_, new_n13642_, new_n13552_ );
xnor ( new_n13644_, new_n13579_, new_n13569_ );
xor  ( new_n13645_, new_n13644_, new_n13591_ );
nand ( new_n13646_, new_n13645_, new_n13643_ );
nor  ( new_n13647_, new_n13645_, new_n13643_ );
xnor ( new_n13648_, new_n13391_, new_n13389_ );
xor  ( new_n13649_, new_n13648_, new_n13395_ );
or   ( new_n13650_, new_n13649_, new_n13647_ );
and  ( new_n13651_, new_n13650_, new_n13646_ );
or   ( new_n13652_, new_n13651_, new_n13641_ );
and  ( new_n13653_, new_n13651_, new_n13641_ );
xor  ( new_n13654_, new_n13225_, new_n13219_ );
xor  ( new_n13655_, new_n13654_, new_n13231_ );
xnor ( new_n13656_, new_n13573_, new_n13571_ );
xor  ( new_n13657_, new_n13656_, new_n13577_ );
and  ( new_n13658_, new_n13657_, new_n13655_ );
or   ( new_n13659_, new_n13657_, new_n13655_ );
xor  ( new_n13660_, new_n13585_, new_n13583_ );
xnor ( new_n13661_, new_n13660_, new_n13589_ );
and  ( new_n13662_, new_n13661_, new_n13659_ );
or   ( new_n13663_, new_n13662_, new_n13658_ );
or   ( new_n13664_, new_n2122_, new_n6219_ );
or   ( new_n13665_, new_n2124_, new_n5899_ );
and  ( new_n13666_, new_n13665_, new_n13664_ );
xor  ( new_n13667_, new_n13666_, new_n1843_ );
or   ( new_n13668_, new_n1844_, new_n6589_ );
or   ( new_n13669_, new_n1846_, new_n6425_ );
and  ( new_n13670_, new_n13669_, new_n13668_ );
xor  ( new_n13671_, new_n13670_, new_n1586_ );
or   ( new_n13672_, new_n13671_, new_n13667_ );
and  ( new_n13673_, new_n13671_, new_n13667_ );
or   ( new_n13674_, new_n1593_, new_n7149_ );
or   ( new_n13675_, new_n1595_, new_n6943_ );
and  ( new_n13676_, new_n13675_, new_n13674_ );
xor  ( new_n13677_, new_n13676_, new_n1358_ );
or   ( new_n13678_, new_n13677_, new_n13673_ );
and  ( new_n13679_, new_n13678_, new_n13672_ );
or   ( new_n13680_, new_n755_, new_n9681_ );
or   ( new_n13681_, new_n757_, new_n9099_ );
and  ( new_n13682_, new_n13681_, new_n13680_ );
xor  ( new_n13683_, new_n13682_, new_n523_ );
or   ( new_n13684_, new_n524_, new_n10220_ );
or   ( new_n13685_, new_n526_, new_n9679_ );
and  ( new_n13686_, new_n13685_, new_n13684_ );
xor  ( new_n13687_, new_n13686_, new_n403_ );
or   ( new_n13688_, new_n13687_, new_n13683_ );
and  ( new_n13689_, new_n13687_, new_n13683_ );
or   ( new_n13690_, new_n409_, new_n10841_ );
or   ( new_n13691_, new_n411_, new_n10541_ );
and  ( new_n13692_, new_n13691_, new_n13690_ );
xor  ( new_n13693_, new_n13692_, new_n328_ );
or   ( new_n13694_, new_n13693_, new_n13689_ );
and  ( new_n13695_, new_n13694_, new_n13688_ );
or   ( new_n13696_, new_n13695_, new_n13679_ );
and  ( new_n13697_, new_n13695_, new_n13679_ );
or   ( new_n13698_, new_n1364_, new_n8117_ );
or   ( new_n13699_, new_n1366_, new_n7373_ );
and  ( new_n13700_, new_n13699_, new_n13698_ );
xor  ( new_n13701_, new_n13700_, new_n1129_ );
or   ( new_n13702_, new_n1135_, new_n8352_ );
or   ( new_n13703_, new_n1137_, new_n8115_ );
and  ( new_n13704_, new_n13703_, new_n13702_ );
xor  ( new_n13705_, new_n13704_, new_n896_ );
or   ( new_n13706_, new_n13705_, new_n13701_ );
and  ( new_n13707_, new_n13705_, new_n13701_ );
or   ( new_n13708_, new_n897_, new_n8995_ );
or   ( new_n13709_, new_n899_, new_n8481_ );
and  ( new_n13710_, new_n13709_, new_n13708_ );
xor  ( new_n13711_, new_n13710_, new_n748_ );
or   ( new_n13712_, new_n13711_, new_n13707_ );
and  ( new_n13713_, new_n13712_, new_n13706_ );
or   ( new_n13714_, new_n13713_, new_n13697_ );
and  ( new_n13715_, new_n13714_, new_n13696_ );
or   ( new_n13716_, new_n7184_, new_n1523_ );
or   ( new_n13717_, new_n7186_, new_n1525_ );
and  ( new_n13718_, new_n13717_, new_n13716_ );
xor  ( new_n13719_, new_n13718_, new_n6638_ );
or   ( new_n13720_, new_n6645_, new_n1899_ );
or   ( new_n13721_, new_n6647_, new_n1754_ );
and  ( new_n13722_, new_n13721_, new_n13720_ );
xor  ( new_n13723_, new_n13722_, new_n6166_ );
or   ( new_n13724_, new_n13723_, new_n13719_ );
and  ( new_n13725_, new_n13723_, new_n13719_ );
or   ( new_n13726_, new_n6173_, new_n2178_ );
or   ( new_n13727_, new_n6175_, new_n2057_ );
and  ( new_n13728_, new_n13727_, new_n13726_ );
xor  ( new_n13729_, new_n13728_, new_n5597_ );
or   ( new_n13730_, new_n13729_, new_n13725_ );
and  ( new_n13731_, new_n13730_, new_n13724_ );
or   ( new_n13732_, new_n8874_, new_n886_ );
or   ( new_n13733_, new_n8876_, new_n805_ );
and  ( new_n13734_, new_n13733_, new_n13732_ );
xor  ( new_n13735_, new_n13734_, new_n8257_ );
or   ( new_n13736_, new_n8264_, new_n1168_ );
or   ( new_n13737_, new_n8266_, new_n986_ );
and  ( new_n13738_, new_n13737_, new_n13736_ );
xor  ( new_n13739_, new_n13738_, new_n7725_ );
or   ( new_n13740_, new_n13739_, new_n13735_ );
and  ( new_n13741_, new_n13739_, new_n13735_ );
or   ( new_n13742_, new_n7732_, new_n1318_ );
or   ( new_n13743_, new_n7734_, new_n1213_ );
and  ( new_n13744_, new_n13743_, new_n13742_ );
xor  ( new_n13745_, new_n13744_, new_n7177_ );
or   ( new_n13746_, new_n13745_, new_n13741_ );
and  ( new_n13747_, new_n13746_, new_n13740_ );
or   ( new_n13748_, new_n13747_, new_n13731_ );
and  ( new_n13749_, new_n13747_, new_n13731_ );
or   ( new_n13750_, new_n10059_, new_n509_ );
or   ( new_n13751_, new_n10061_, new_n443_ );
and  ( new_n13752_, new_n13751_, new_n13750_ );
xor  ( new_n13753_, new_n13752_, new_n9421_ );
and  ( new_n13754_, RIbb2d888_64, RIbb2d360_75 );
or   ( new_n13755_, RIbb2d888_64, new_n419_ );
and  ( new_n13756_, new_n13755_, RIbb2d900_63 );
or   ( new_n13757_, new_n13756_, new_n13754_ );
or   ( new_n13758_, new_n10770_, new_n348_ );
and  ( new_n13759_, new_n13758_, new_n13757_ );
nor  ( new_n13760_, new_n13759_, new_n13753_ );
and  ( new_n13761_, new_n13759_, new_n13753_ );
or   ( new_n13762_, new_n9422_, new_n775_ );
or   ( new_n13763_, new_n9424_, new_n515_ );
and  ( new_n13764_, new_n13763_, new_n13762_ );
xor  ( new_n13765_, new_n13764_, new_n8873_ );
nor  ( new_n13766_, new_n13765_, new_n13761_ );
nor  ( new_n13767_, new_n13766_, new_n13760_ );
or   ( new_n13768_, new_n13767_, new_n13749_ );
and  ( new_n13769_, new_n13768_, new_n13748_ );
or   ( new_n13770_, new_n13769_, new_n13715_ );
or   ( new_n13771_, new_n4302_, new_n3696_ );
or   ( new_n13772_, new_n4304_, new_n3306_ );
and  ( new_n13773_, new_n13772_, new_n13771_ );
xor  ( new_n13774_, new_n13773_, new_n3895_ );
or   ( new_n13775_, new_n3896_, new_n3820_ );
or   ( new_n13776_, new_n3898_, new_n3694_ );
and  ( new_n13777_, new_n13776_, new_n13775_ );
xor  ( new_n13778_, new_n13777_, new_n3460_ );
or   ( new_n13779_, new_n13778_, new_n13774_ );
and  ( new_n13780_, new_n13778_, new_n13774_ );
or   ( new_n13781_, new_n3461_, new_n4267_ );
or   ( new_n13782_, new_n3463_, new_n4069_ );
and  ( new_n13783_, new_n13782_, new_n13781_ );
xor  ( new_n13784_, new_n13783_, new_n3116_ );
or   ( new_n13785_, new_n13784_, new_n13780_ );
and  ( new_n13786_, new_n13785_, new_n13779_ );
or   ( new_n13787_, new_n3117_, new_n4995_ );
or   ( new_n13788_, new_n3119_, new_n4603_ );
and  ( new_n13789_, new_n13788_, new_n13787_ );
xor  ( new_n13790_, new_n13789_, new_n2800_ );
or   ( new_n13791_, new_n2807_, new_n5171_ );
or   ( new_n13792_, new_n2809_, new_n4859_ );
and  ( new_n13793_, new_n13792_, new_n13791_ );
xor  ( new_n13794_, new_n13793_, new_n2424_ );
or   ( new_n13795_, new_n13794_, new_n13790_ );
and  ( new_n13796_, new_n13794_, new_n13790_ );
or   ( new_n13797_, new_n2425_, new_n5570_ );
or   ( new_n13798_, new_n2427_, new_n5428_ );
and  ( new_n13799_, new_n13798_, new_n13797_ );
xor  ( new_n13800_, new_n13799_, new_n2121_ );
or   ( new_n13801_, new_n13800_, new_n13796_ );
and  ( new_n13802_, new_n13801_, new_n13795_ );
nor  ( new_n13803_, new_n13802_, new_n13786_ );
and  ( new_n13804_, new_n13802_, new_n13786_ );
or   ( new_n13805_, new_n5604_, new_n2475_ );
or   ( new_n13806_, new_n5606_, new_n2291_ );
and  ( new_n13807_, new_n13806_, new_n13805_ );
xor  ( new_n13808_, new_n13807_, new_n5206_ );
or   ( new_n13809_, new_n5207_, new_n2751_ );
or   ( new_n13810_, new_n5209_, new_n2646_ );
and  ( new_n13811_, new_n13810_, new_n13809_ );
xor  ( new_n13812_, new_n13811_, new_n4708_ );
nor  ( new_n13813_, new_n13812_, new_n13808_ );
and  ( new_n13814_, new_n13812_, new_n13808_ );
or   ( new_n13815_, new_n4709_, new_n3178_ );
or   ( new_n13816_, new_n4711_, new_n2981_ );
and  ( new_n13817_, new_n13816_, new_n13815_ );
xor  ( new_n13818_, new_n13817_, new_n4295_ );
nor  ( new_n13819_, new_n13818_, new_n13814_ );
nor  ( new_n13820_, new_n13819_, new_n13813_ );
nor  ( new_n13821_, new_n13820_, new_n13804_ );
nor  ( new_n13822_, new_n13821_, new_n13803_ );
and  ( new_n13823_, new_n13769_, new_n13715_ );
or   ( new_n13824_, new_n13823_, new_n13822_ );
and  ( new_n13825_, new_n13824_, new_n13770_ );
and  ( new_n13826_, new_n13825_, new_n13663_ );
nor  ( new_n13827_, new_n13825_, new_n13663_ );
xnor ( new_n13828_, new_n13524_, new_n13520_ );
xor  ( new_n13829_, new_n13828_, new_n13530_ );
xnor ( new_n13830_, new_n13405_, new_n13401_ );
xor  ( new_n13831_, new_n13830_, new_n13411_ );
nor  ( new_n13832_, new_n13831_, new_n13829_ );
nand ( new_n13833_, new_n13831_, new_n13829_ );
xor  ( new_n13834_, new_n13439_, new_n13435_ );
xor  ( new_n13835_, new_n13834_, new_n13445_ );
and  ( new_n13836_, new_n13835_, new_n13833_ );
or   ( new_n13837_, new_n13836_, new_n13832_ );
or   ( new_n13838_, new_n409_, new_n10541_ );
or   ( new_n13839_, new_n411_, new_n10220_ );
and  ( new_n13840_, new_n13839_, new_n13838_ );
xor  ( new_n13841_, new_n13840_, new_n328_ );
and  ( new_n13842_, new_n334_, RIbb31578_128 );
or   ( new_n13843_, new_n13842_, new_n331_ );
nor  ( new_n13844_, RIbb2f1d8_10, RIbb2f160_11 );
or   ( new_n13845_, new_n13844_, new_n332_ );
or   ( new_n13846_, new_n13845_, new_n10841_ );
and  ( new_n13847_, new_n13846_, new_n13843_ );
or   ( new_n13848_, new_n13847_, new_n13841_ );
nand ( new_n13849_, new_n13847_, new_n13841_ );
xor  ( new_n13850_, new_n13421_, new_n13417_ );
xnor ( new_n13851_, new_n13850_, new_n13427_ );
nand ( new_n13852_, new_n13851_, new_n13849_ );
and  ( new_n13853_, new_n13852_, new_n13848_ );
and  ( new_n13854_, new_n13853_, new_n13837_ );
nor  ( new_n13855_, new_n13853_, new_n13837_ );
xnor ( new_n13856_, new_n13457_, new_n13453_ );
xor  ( new_n13857_, new_n13856_, new_n13463_ );
xnor ( new_n13858_, new_n13508_, new_n13504_ );
xor  ( new_n13859_, new_n13858_, new_n13514_ );
nor  ( new_n13860_, new_n13859_, new_n13857_ );
and  ( new_n13861_, new_n13859_, new_n13857_ );
xor  ( new_n13862_, new_n13542_, new_n13538_ );
xnor ( new_n13863_, new_n13862_, new_n13548_ );
nor  ( new_n13864_, new_n13863_, new_n13861_ );
nor  ( new_n13865_, new_n13864_, new_n13860_ );
nor  ( new_n13866_, new_n13865_, new_n13855_ );
nor  ( new_n13867_, new_n13866_, new_n13854_ );
nor  ( new_n13868_, new_n13867_, new_n13827_ );
nor  ( new_n13869_, new_n13868_, new_n13826_ );
or   ( new_n13870_, new_n13869_, new_n13653_ );
and  ( new_n13871_, new_n13870_, new_n13652_ );
or   ( new_n13872_, new_n13871_, new_n13623_ );
and  ( new_n13873_, new_n13872_, new_n13622_ );
xor  ( new_n13874_, new_n13354_, new_n13344_ );
xor  ( new_n13875_, new_n13874_, new_n13597_ );
or   ( new_n13876_, new_n13875_, new_n13873_ );
and  ( new_n13877_, new_n13875_, new_n13873_ );
xor  ( new_n13878_, new_n13334_, new_n13332_ );
xor  ( new_n13879_, new_n13878_, new_n13338_ );
or   ( new_n13880_, new_n13879_, new_n13877_ );
and  ( new_n13881_, new_n13880_, new_n13876_ );
or   ( new_n13882_, new_n13881_, new_n13609_ );
and  ( new_n13883_, new_n13881_, new_n13609_ );
xor  ( new_n13884_, new_n13068_, new_n13058_ );
xor  ( new_n13885_, new_n13884_, new_n13314_ );
or   ( new_n13886_, new_n13885_, new_n13883_ );
and  ( new_n13887_, new_n13886_, new_n13882_ );
nor  ( new_n13888_, new_n13887_, new_n13607_ );
xor  ( new_n13889_, new_n13875_, new_n13873_ );
xor  ( new_n13890_, new_n13889_, new_n13879_ );
xnor ( new_n13891_, new_n13825_, new_n13663_ );
xor  ( new_n13892_, new_n13891_, new_n13867_ );
xnor ( new_n13893_, new_n13635_, new_n13625_ );
xor  ( new_n13894_, new_n13893_, new_n13639_ );
nor  ( new_n13895_, new_n13894_, new_n13892_ );
nand ( new_n13896_, new_n13894_, new_n13892_ );
xor  ( new_n13897_, new_n13645_, new_n13643_ );
xor  ( new_n13898_, new_n13897_, new_n13649_ );
and  ( new_n13899_, new_n13898_, new_n13896_ );
or   ( new_n13900_, new_n13899_, new_n13895_ );
xor  ( new_n13901_, new_n13615_, new_n13613_ );
xor  ( new_n13902_, new_n13901_, new_n13619_ );
nor  ( new_n13903_, new_n13902_, new_n13900_ );
and  ( new_n13904_, new_n13902_, new_n13900_ );
xnor ( new_n13905_, new_n13747_, new_n13731_ );
xor  ( new_n13906_, new_n13905_, new_n13767_ );
xnor ( new_n13907_, new_n13802_, new_n13786_ );
xor  ( new_n13908_, new_n13907_, new_n13820_ );
or   ( new_n13909_, new_n13908_, new_n13906_ );
xor  ( new_n13910_, new_n13695_, new_n13679_ );
xor  ( new_n13911_, new_n13910_, new_n13713_ );
xor  ( new_n13912_, new_n13831_, new_n13829_ );
xor  ( new_n13913_, new_n13912_, new_n13835_ );
nand ( new_n13914_, new_n13913_, new_n13911_ );
nor  ( new_n13915_, new_n13913_, new_n13911_ );
xor  ( new_n13916_, new_n13847_, new_n13841_ );
xor  ( new_n13917_, new_n13916_, new_n13851_ );
or   ( new_n13918_, new_n13917_, new_n13915_ );
and  ( new_n13919_, new_n13918_, new_n13914_ );
or   ( new_n13920_, new_n13919_, new_n13909_ );
and  ( new_n13921_, new_n13919_, new_n13909_ );
xnor ( new_n13922_, new_n13495_, new_n13479_ );
xor  ( new_n13923_, new_n13922_, new_n13465_ );
or   ( new_n13924_, new_n13923_, new_n13921_ );
and  ( new_n13925_, new_n13924_, new_n13920_ );
xnor ( new_n13926_, new_n13853_, new_n13837_ );
xor  ( new_n13927_, new_n13926_, new_n13865_ );
xnor ( new_n13928_, new_n13629_, new_n13627_ );
xor  ( new_n13929_, new_n13928_, new_n13633_ );
nand ( new_n13930_, new_n13929_, new_n13927_ );
nor  ( new_n13931_, new_n13929_, new_n13927_ );
xor  ( new_n13932_, new_n13657_, new_n13655_ );
xnor ( new_n13933_, new_n13932_, new_n13661_ );
or   ( new_n13934_, new_n13933_, new_n13931_ );
and  ( new_n13935_, new_n13934_, new_n13930_ );
nor  ( new_n13936_, new_n13935_, new_n13925_ );
and  ( new_n13937_, new_n13935_, new_n13925_ );
xnor ( new_n13938_, new_n13487_, new_n13483_ );
xor  ( new_n13939_, new_n13938_, new_n13493_ );
xor  ( new_n13940_, new_n13475_, new_n13469_ );
xor  ( new_n13941_, new_n13940_, new_n332_ );
nor  ( new_n13942_, new_n13941_, new_n13939_ );
nand ( new_n13943_, new_n13941_, new_n13939_ );
xor  ( new_n13944_, new_n13859_, new_n13857_ );
xnor ( new_n13945_, new_n13944_, new_n13863_ );
and  ( new_n13946_, new_n13945_, new_n13943_ );
or   ( new_n13947_, new_n13946_, new_n13942_ );
or   ( new_n13948_, new_n6173_, new_n2291_ );
or   ( new_n13949_, new_n6175_, new_n2178_ );
and  ( new_n13950_, new_n13949_, new_n13948_ );
xor  ( new_n13951_, new_n13950_, new_n5597_ );
or   ( new_n13952_, new_n5604_, new_n2646_ );
or   ( new_n13953_, new_n5606_, new_n2475_ );
and  ( new_n13954_, new_n13953_, new_n13952_ );
xor  ( new_n13955_, new_n13954_, new_n5206_ );
or   ( new_n13956_, new_n13955_, new_n13951_ );
and  ( new_n13957_, new_n13955_, new_n13951_ );
or   ( new_n13958_, new_n5207_, new_n2981_ );
or   ( new_n13959_, new_n5209_, new_n2751_ );
and  ( new_n13960_, new_n13959_, new_n13958_ );
xor  ( new_n13961_, new_n13960_, new_n4708_ );
or   ( new_n13962_, new_n13961_, new_n13957_ );
and  ( new_n13963_, new_n13962_, new_n13956_ );
or   ( new_n13964_, new_n3461_, new_n4603_ );
or   ( new_n13965_, new_n3463_, new_n4267_ );
and  ( new_n13966_, new_n13965_, new_n13964_ );
xor  ( new_n13967_, new_n13966_, new_n3116_ );
or   ( new_n13968_, new_n3117_, new_n4859_ );
or   ( new_n13969_, new_n3119_, new_n4995_ );
and  ( new_n13970_, new_n13969_, new_n13968_ );
xor  ( new_n13971_, new_n13970_, new_n2800_ );
or   ( new_n13972_, new_n13971_, new_n13967_ );
and  ( new_n13973_, new_n13971_, new_n13967_ );
or   ( new_n13974_, new_n2807_, new_n5428_ );
or   ( new_n13975_, new_n2809_, new_n5171_ );
and  ( new_n13976_, new_n13975_, new_n13974_ );
xor  ( new_n13977_, new_n13976_, new_n2424_ );
or   ( new_n13978_, new_n13977_, new_n13973_ );
and  ( new_n13979_, new_n13978_, new_n13972_ );
or   ( new_n13980_, new_n13979_, new_n13963_ );
and  ( new_n13981_, new_n13979_, new_n13963_ );
or   ( new_n13982_, new_n4709_, new_n3306_ );
or   ( new_n13983_, new_n4711_, new_n3178_ );
and  ( new_n13984_, new_n13983_, new_n13982_ );
xor  ( new_n13985_, new_n13984_, new_n4295_ );
or   ( new_n13986_, new_n4302_, new_n3694_ );
or   ( new_n13987_, new_n4304_, new_n3696_ );
and  ( new_n13988_, new_n13987_, new_n13986_ );
xor  ( new_n13989_, new_n13988_, new_n3895_ );
or   ( new_n13990_, new_n13989_, new_n13985_ );
and  ( new_n13991_, new_n13989_, new_n13985_ );
or   ( new_n13992_, new_n3896_, new_n4069_ );
or   ( new_n13993_, new_n3898_, new_n3820_ );
and  ( new_n13994_, new_n13993_, new_n13992_ );
xor  ( new_n13995_, new_n13994_, new_n3460_ );
or   ( new_n13996_, new_n13995_, new_n13991_ );
and  ( new_n13997_, new_n13996_, new_n13990_ );
or   ( new_n13998_, new_n13997_, new_n13981_ );
and  ( new_n13999_, new_n13998_, new_n13980_ );
or   ( new_n14000_, new_n9422_, new_n805_ );
or   ( new_n14001_, new_n9424_, new_n775_ );
and  ( new_n14002_, new_n14001_, new_n14000_ );
xor  ( new_n14003_, new_n14002_, new_n8873_ );
or   ( new_n14004_, new_n8874_, new_n986_ );
or   ( new_n14005_, new_n8876_, new_n886_ );
and  ( new_n14006_, new_n14005_, new_n14004_ );
xor  ( new_n14007_, new_n14006_, new_n8257_ );
nor  ( new_n14008_, new_n14007_, new_n14003_ );
and  ( new_n14009_, new_n14007_, new_n14003_ );
or   ( new_n14010_, new_n8264_, new_n1213_ );
or   ( new_n14011_, new_n8266_, new_n1168_ );
and  ( new_n14012_, new_n14011_, new_n14010_ );
xor  ( new_n14013_, new_n14012_, new_n7725_ );
nor  ( new_n14014_, new_n14013_, new_n14009_ );
nor  ( new_n14015_, new_n14014_, new_n14008_ );
or   ( new_n14016_, new_n10059_, new_n515_ );
or   ( new_n14017_, new_n10061_, new_n509_ );
and  ( new_n14018_, new_n14017_, new_n14016_ );
xor  ( new_n14019_, new_n14018_, new_n9421_ );
and  ( new_n14020_, RIbb2d888_64, RIbb2d2e8_76 );
or   ( new_n14021_, RIbb2d888_64, new_n443_ );
and  ( new_n14022_, new_n14021_, RIbb2d900_63 );
or   ( new_n14023_, new_n14022_, new_n14020_ );
or   ( new_n14024_, new_n10770_, new_n419_ );
and  ( new_n14025_, new_n14024_, new_n14023_ );
nor  ( new_n14026_, new_n14025_, new_n14019_ );
and  ( new_n14027_, new_n14025_, new_n14019_ );
nor  ( new_n14028_, new_n14027_, new_n327_ );
nor  ( new_n14029_, new_n14028_, new_n14026_ );
or   ( new_n14030_, new_n7732_, new_n1525_ );
or   ( new_n14031_, new_n7734_, new_n1318_ );
and  ( new_n14032_, new_n14031_, new_n14030_ );
xor  ( new_n14033_, new_n14032_, new_n7177_ );
or   ( new_n14034_, new_n7184_, new_n1754_ );
or   ( new_n14035_, new_n7186_, new_n1523_ );
and  ( new_n14036_, new_n14035_, new_n14034_ );
xor  ( new_n14037_, new_n14036_, new_n6638_ );
or   ( new_n14038_, new_n14037_, new_n14033_ );
and  ( new_n14039_, new_n14037_, new_n14033_ );
or   ( new_n14040_, new_n6645_, new_n2057_ );
or   ( new_n14041_, new_n6647_, new_n1899_ );
and  ( new_n14042_, new_n14041_, new_n14040_ );
xor  ( new_n14043_, new_n14042_, new_n6166_ );
or   ( new_n14044_, new_n14043_, new_n14039_ );
and  ( new_n14045_, new_n14044_, new_n14038_ );
and  ( new_n14046_, new_n14045_, new_n14029_ );
or   ( new_n14047_, new_n14046_, new_n14015_ );
or   ( new_n14048_, new_n14045_, new_n14029_ );
and  ( new_n14049_, new_n14048_, new_n14047_ );
or   ( new_n14050_, new_n14049_, new_n13999_ );
or   ( new_n14051_, new_n2425_, new_n5899_ );
or   ( new_n14052_, new_n2427_, new_n5570_ );
and  ( new_n14053_, new_n14052_, new_n14051_ );
xor  ( new_n14054_, new_n14053_, new_n2121_ );
or   ( new_n14055_, new_n2122_, new_n6425_ );
or   ( new_n14056_, new_n2124_, new_n6219_ );
and  ( new_n14057_, new_n14056_, new_n14055_ );
xor  ( new_n14058_, new_n14057_, new_n1843_ );
or   ( new_n14059_, new_n14058_, new_n14054_ );
and  ( new_n14060_, new_n14058_, new_n14054_ );
or   ( new_n14061_, new_n1844_, new_n6943_ );
or   ( new_n14062_, new_n1846_, new_n6589_ );
and  ( new_n14063_, new_n14062_, new_n14061_ );
xor  ( new_n14064_, new_n14063_, new_n1586_ );
or   ( new_n14065_, new_n14064_, new_n14060_ );
and  ( new_n14066_, new_n14065_, new_n14059_ );
or   ( new_n14067_, new_n897_, new_n9099_ );
or   ( new_n14068_, new_n899_, new_n8995_ );
and  ( new_n14069_, new_n14068_, new_n14067_ );
xor  ( new_n14070_, new_n14069_, new_n748_ );
or   ( new_n14071_, new_n755_, new_n9679_ );
or   ( new_n14072_, new_n757_, new_n9681_ );
and  ( new_n14073_, new_n14072_, new_n14071_ );
xor  ( new_n14074_, new_n14073_, new_n523_ );
or   ( new_n14075_, new_n14074_, new_n14070_ );
and  ( new_n14076_, new_n14074_, new_n14070_ );
or   ( new_n14077_, new_n524_, new_n10541_ );
or   ( new_n14078_, new_n526_, new_n10220_ );
and  ( new_n14079_, new_n14078_, new_n14077_ );
xor  ( new_n14080_, new_n14079_, new_n403_ );
or   ( new_n14081_, new_n14080_, new_n14076_ );
and  ( new_n14082_, new_n14081_, new_n14075_ );
nor  ( new_n14083_, new_n14082_, new_n14066_ );
and  ( new_n14084_, new_n14082_, new_n14066_ );
or   ( new_n14085_, new_n1593_, new_n7373_ );
or   ( new_n14086_, new_n1595_, new_n7149_ );
and  ( new_n14087_, new_n14086_, new_n14085_ );
xor  ( new_n14088_, new_n14087_, new_n1358_ );
or   ( new_n14089_, new_n1364_, new_n8115_ );
or   ( new_n14090_, new_n1366_, new_n8117_ );
and  ( new_n14091_, new_n14090_, new_n14089_ );
xor  ( new_n14092_, new_n14091_, new_n1129_ );
nor  ( new_n14093_, new_n14092_, new_n14088_ );
and  ( new_n14094_, new_n14092_, new_n14088_ );
or   ( new_n14095_, new_n1135_, new_n8481_ );
or   ( new_n14096_, new_n1137_, new_n8352_ );
and  ( new_n14097_, new_n14096_, new_n14095_ );
xor  ( new_n14098_, new_n14097_, new_n896_ );
nor  ( new_n14099_, new_n14098_, new_n14094_ );
nor  ( new_n14100_, new_n14099_, new_n14093_ );
nor  ( new_n14101_, new_n14100_, new_n14084_ );
nor  ( new_n14102_, new_n14101_, new_n14083_ );
and  ( new_n14103_, new_n14049_, new_n13999_ );
or   ( new_n14104_, new_n14103_, new_n14102_ );
and  ( new_n14105_, new_n14104_, new_n14050_ );
and  ( new_n14106_, new_n14105_, new_n13947_ );
nor  ( new_n14107_, new_n14105_, new_n13947_ );
xnor ( new_n14108_, new_n13687_, new_n13683_ );
xor  ( new_n14109_, new_n14108_, new_n13693_ );
xnor ( new_n14110_, new_n13671_, new_n13667_ );
xor  ( new_n14111_, new_n14110_, new_n13677_ );
or   ( new_n14112_, new_n14111_, new_n14109_ );
and  ( new_n14113_, new_n14111_, new_n14109_ );
xor  ( new_n14114_, new_n13705_, new_n13701_ );
xnor ( new_n14115_, new_n14114_, new_n13711_ );
or   ( new_n14116_, new_n14115_, new_n14113_ );
and  ( new_n14117_, new_n14116_, new_n14112_ );
xnor ( new_n14118_, new_n13739_, new_n13735_ );
xor  ( new_n14119_, new_n14118_, new_n13745_ );
xnor ( new_n14120_, new_n13723_, new_n13719_ );
xor  ( new_n14121_, new_n14120_, new_n13729_ );
or   ( new_n14122_, new_n14121_, new_n14119_ );
and  ( new_n14123_, new_n14121_, new_n14119_ );
xor  ( new_n14124_, new_n13759_, new_n13753_ );
xnor ( new_n14125_, new_n14124_, new_n13765_ );
or   ( new_n14126_, new_n14125_, new_n14123_ );
and  ( new_n14127_, new_n14126_, new_n14122_ );
nor  ( new_n14128_, new_n14127_, new_n14117_ );
and  ( new_n14129_, new_n14127_, new_n14117_ );
xnor ( new_n14130_, new_n13794_, new_n13790_ );
xor  ( new_n14131_, new_n14130_, new_n13800_ );
xnor ( new_n14132_, new_n13778_, new_n13774_ );
xor  ( new_n14133_, new_n14132_, new_n13784_ );
nor  ( new_n14134_, new_n14133_, new_n14131_ );
and  ( new_n14135_, new_n14133_, new_n14131_ );
xor  ( new_n14136_, new_n13812_, new_n13808_ );
xnor ( new_n14137_, new_n14136_, new_n13818_ );
nor  ( new_n14138_, new_n14137_, new_n14135_ );
nor  ( new_n14139_, new_n14138_, new_n14134_ );
nor  ( new_n14140_, new_n14139_, new_n14129_ );
nor  ( new_n14141_, new_n14140_, new_n14128_ );
nor  ( new_n14142_, new_n14141_, new_n14107_ );
nor  ( new_n14143_, new_n14142_, new_n14106_ );
nor  ( new_n14144_, new_n14143_, new_n13937_ );
nor  ( new_n14145_, new_n14144_, new_n13936_ );
nor  ( new_n14146_, new_n14145_, new_n13904_ );
or   ( new_n14147_, new_n14146_, new_n13903_ );
xnor ( new_n14148_, new_n13385_, new_n13375_ );
xor  ( new_n14149_, new_n14148_, new_n13595_ );
nand ( new_n14150_, new_n14149_, new_n14147_ );
nor  ( new_n14151_, new_n14149_, new_n14147_ );
xor  ( new_n14152_, new_n13621_, new_n13611_ );
xor  ( new_n14153_, new_n14152_, new_n13871_ );
or   ( new_n14154_, new_n14153_, new_n14151_ );
and  ( new_n14155_, new_n14154_, new_n14150_ );
nor  ( new_n14156_, new_n14155_, new_n13890_ );
xnor ( new_n14157_, new_n13881_, new_n13609_ );
xor  ( new_n14158_, new_n14157_, new_n13885_ );
and  ( new_n14159_, new_n14158_, new_n14156_ );
xor  ( new_n14160_, new_n14149_, new_n14147_ );
xor  ( new_n14161_, new_n14160_, new_n14153_ );
xor  ( new_n14162_, new_n13908_, new_n13906_ );
xnor ( new_n14163_, new_n13913_, new_n13911_ );
xor  ( new_n14164_, new_n14163_, new_n13917_ );
and  ( new_n14165_, new_n14164_, new_n14162_ );
nor  ( new_n14166_, new_n14164_, new_n14162_ );
xor  ( new_n14167_, new_n13979_, new_n13963_ );
xor  ( new_n14168_, new_n14167_, new_n13997_ );
xor  ( new_n14169_, new_n14045_, new_n14029_ );
xor  ( new_n14170_, new_n14169_, new_n14015_ );
and  ( new_n14171_, new_n14170_, new_n14168_ );
nor  ( new_n14172_, new_n14170_, new_n14168_ );
xor  ( new_n14173_, new_n14082_, new_n14066_ );
xnor ( new_n14174_, new_n14173_, new_n14100_ );
nor  ( new_n14175_, new_n14174_, new_n14172_ );
nor  ( new_n14176_, new_n14175_, new_n14171_ );
nor  ( new_n14177_, new_n14176_, new_n14166_ );
nor  ( new_n14178_, new_n14177_, new_n14165_ );
xnor ( new_n14179_, new_n14133_, new_n14131_ );
xor  ( new_n14180_, new_n14179_, new_n14137_ );
xnor ( new_n14181_, new_n14111_, new_n14109_ );
xor  ( new_n14182_, new_n14181_, new_n14115_ );
nor  ( new_n14183_, new_n14182_, new_n14180_ );
and  ( new_n14184_, new_n14182_, new_n14180_ );
xor  ( new_n14185_, new_n14121_, new_n14119_ );
xnor ( new_n14186_, new_n14185_, new_n14125_ );
nor  ( new_n14187_, new_n14186_, new_n14184_ );
nor  ( new_n14188_, new_n14187_, new_n14183_ );
or   ( new_n14189_, new_n5604_, new_n2751_ );
or   ( new_n14190_, new_n5606_, new_n2646_ );
and  ( new_n14191_, new_n14190_, new_n14189_ );
xor  ( new_n14192_, new_n14191_, new_n5206_ );
or   ( new_n14193_, new_n5207_, new_n3178_ );
or   ( new_n14194_, new_n5209_, new_n2981_ );
and  ( new_n14195_, new_n14194_, new_n14193_ );
xor  ( new_n14196_, new_n14195_, new_n4708_ );
or   ( new_n14197_, new_n14196_, new_n14192_ );
and  ( new_n14198_, new_n14196_, new_n14192_ );
or   ( new_n14199_, new_n4709_, new_n3696_ );
or   ( new_n14200_, new_n4711_, new_n3306_ );
and  ( new_n14201_, new_n14200_, new_n14199_ );
xor  ( new_n14202_, new_n14201_, new_n4295_ );
or   ( new_n14203_, new_n14202_, new_n14198_ );
and  ( new_n14204_, new_n14203_, new_n14197_ );
or   ( new_n14205_, new_n4302_, new_n3820_ );
or   ( new_n14206_, new_n4304_, new_n3694_ );
and  ( new_n14207_, new_n14206_, new_n14205_ );
xor  ( new_n14208_, new_n14207_, new_n3895_ );
or   ( new_n14209_, new_n3896_, new_n4267_ );
or   ( new_n14210_, new_n3898_, new_n4069_ );
and  ( new_n14211_, new_n14210_, new_n14209_ );
xor  ( new_n14212_, new_n14211_, new_n3460_ );
or   ( new_n14213_, new_n14212_, new_n14208_ );
and  ( new_n14214_, new_n14212_, new_n14208_ );
or   ( new_n14215_, new_n3461_, new_n4995_ );
or   ( new_n14216_, new_n3463_, new_n4603_ );
and  ( new_n14217_, new_n14216_, new_n14215_ );
xor  ( new_n14218_, new_n14217_, new_n3116_ );
or   ( new_n14219_, new_n14218_, new_n14214_ );
and  ( new_n14220_, new_n14219_, new_n14213_ );
or   ( new_n14221_, new_n14220_, new_n14204_ );
and  ( new_n14222_, new_n14220_, new_n14204_ );
or   ( new_n14223_, new_n3117_, new_n5171_ );
or   ( new_n14224_, new_n3119_, new_n4859_ );
and  ( new_n14225_, new_n14224_, new_n14223_ );
xor  ( new_n14226_, new_n14225_, new_n2800_ );
or   ( new_n14227_, new_n2807_, new_n5570_ );
or   ( new_n14228_, new_n2809_, new_n5428_ );
and  ( new_n14229_, new_n14228_, new_n14227_ );
xor  ( new_n14230_, new_n14229_, new_n2424_ );
or   ( new_n14231_, new_n14230_, new_n14226_ );
and  ( new_n14232_, new_n14230_, new_n14226_ );
or   ( new_n14233_, new_n2425_, new_n6219_ );
or   ( new_n14234_, new_n2427_, new_n5899_ );
and  ( new_n14235_, new_n14234_, new_n14233_ );
xor  ( new_n14236_, new_n14235_, new_n2121_ );
or   ( new_n14237_, new_n14236_, new_n14232_ );
and  ( new_n14238_, new_n14237_, new_n14231_ );
or   ( new_n14239_, new_n14238_, new_n14222_ );
and  ( new_n14240_, new_n14239_, new_n14221_ );
or   ( new_n14241_, new_n1364_, new_n8352_ );
or   ( new_n14242_, new_n1366_, new_n8115_ );
and  ( new_n14243_, new_n14242_, new_n14241_ );
xor  ( new_n14244_, new_n14243_, new_n1129_ );
or   ( new_n14245_, new_n1135_, new_n8995_ );
or   ( new_n14246_, new_n1137_, new_n8481_ );
and  ( new_n14247_, new_n14246_, new_n14245_ );
xor  ( new_n14248_, new_n14247_, new_n896_ );
nor  ( new_n14249_, new_n14248_, new_n14244_ );
and  ( new_n14250_, new_n14248_, new_n14244_ );
or   ( new_n14251_, new_n897_, new_n9681_ );
or   ( new_n14252_, new_n899_, new_n9099_ );
and  ( new_n14253_, new_n14252_, new_n14251_ );
xor  ( new_n14254_, new_n14253_, new_n748_ );
nor  ( new_n14255_, new_n14254_, new_n14250_ );
nor  ( new_n14256_, new_n14255_, new_n14249_ );
or   ( new_n14257_, new_n755_, new_n10220_ );
or   ( new_n14258_, new_n757_, new_n9679_ );
and  ( new_n14259_, new_n14258_, new_n14257_ );
xor  ( new_n14260_, new_n14259_, new_n523_ );
or   ( new_n14261_, new_n524_, new_n10841_ );
or   ( new_n14262_, new_n526_, new_n10541_ );
and  ( new_n14263_, new_n14262_, new_n14261_ );
xor  ( new_n14264_, new_n14263_, new_n403_ );
and  ( new_n14265_, new_n14264_, new_n14260_ );
or   ( new_n14266_, new_n2122_, new_n6589_ );
or   ( new_n14267_, new_n2124_, new_n6425_ );
and  ( new_n14268_, new_n14267_, new_n14266_ );
xor  ( new_n14269_, new_n14268_, new_n1843_ );
or   ( new_n14270_, new_n1844_, new_n7149_ );
or   ( new_n14271_, new_n1846_, new_n6943_ );
and  ( new_n14272_, new_n14271_, new_n14270_ );
xor  ( new_n14273_, new_n14272_, new_n1586_ );
or   ( new_n14274_, new_n14273_, new_n14269_ );
and  ( new_n14275_, new_n14273_, new_n14269_ );
or   ( new_n14276_, new_n1593_, new_n8117_ );
or   ( new_n14277_, new_n1595_, new_n7373_ );
and  ( new_n14278_, new_n14277_, new_n14276_ );
xor  ( new_n14279_, new_n14278_, new_n1358_ );
or   ( new_n14280_, new_n14279_, new_n14275_ );
and  ( new_n14281_, new_n14280_, new_n14274_ );
and  ( new_n14282_, new_n14281_, new_n14265_ );
or   ( new_n14283_, new_n14282_, new_n14256_ );
or   ( new_n14284_, new_n14281_, new_n14265_ );
and  ( new_n14285_, new_n14284_, new_n14283_ );
nor  ( new_n14286_, new_n14285_, new_n14240_ );
or   ( new_n14287_, new_n10059_, new_n775_ );
or   ( new_n14288_, new_n10061_, new_n515_ );
and  ( new_n14289_, new_n14288_, new_n14287_ );
xor  ( new_n14290_, new_n14289_, new_n9421_ );
and  ( new_n14291_, RIbb2d888_64, RIbb2d270_77 );
or   ( new_n14292_, RIbb2d888_64, new_n509_ );
and  ( new_n14293_, new_n14292_, RIbb2d900_63 );
or   ( new_n14294_, new_n14293_, new_n14291_ );
or   ( new_n14295_, new_n10770_, new_n443_ );
and  ( new_n14296_, new_n14295_, new_n14294_ );
or   ( new_n14297_, new_n14296_, new_n14290_ );
and  ( new_n14298_, new_n14296_, new_n14290_ );
or   ( new_n14299_, new_n9422_, new_n886_ );
or   ( new_n14300_, new_n9424_, new_n805_ );
and  ( new_n14301_, new_n14300_, new_n14299_ );
xor  ( new_n14302_, new_n14301_, new_n8873_ );
or   ( new_n14303_, new_n14302_, new_n14298_ );
and  ( new_n14304_, new_n14303_, new_n14297_ );
or   ( new_n14305_, new_n7184_, new_n1899_ );
or   ( new_n14306_, new_n7186_, new_n1754_ );
and  ( new_n14307_, new_n14306_, new_n14305_ );
xor  ( new_n14308_, new_n14307_, new_n6638_ );
or   ( new_n14309_, new_n6645_, new_n2178_ );
or   ( new_n14310_, new_n6647_, new_n2057_ );
and  ( new_n14311_, new_n14310_, new_n14309_ );
xor  ( new_n14312_, new_n14311_, new_n6166_ );
or   ( new_n14313_, new_n14312_, new_n14308_ );
and  ( new_n14314_, new_n14312_, new_n14308_ );
or   ( new_n14315_, new_n6173_, new_n2475_ );
or   ( new_n14316_, new_n6175_, new_n2291_ );
and  ( new_n14317_, new_n14316_, new_n14315_ );
xor  ( new_n14318_, new_n14317_, new_n5597_ );
or   ( new_n14319_, new_n14318_, new_n14314_ );
and  ( new_n14320_, new_n14319_, new_n14313_ );
nor  ( new_n14321_, new_n14320_, new_n14304_ );
and  ( new_n14322_, new_n14320_, new_n14304_ );
or   ( new_n14323_, new_n8874_, new_n1168_ );
or   ( new_n14324_, new_n8876_, new_n986_ );
and  ( new_n14325_, new_n14324_, new_n14323_ );
xor  ( new_n14326_, new_n14325_, new_n8257_ );
or   ( new_n14327_, new_n8264_, new_n1318_ );
or   ( new_n14328_, new_n8266_, new_n1213_ );
and  ( new_n14329_, new_n14328_, new_n14327_ );
xor  ( new_n14330_, new_n14329_, new_n7725_ );
nor  ( new_n14331_, new_n14330_, new_n14326_ );
and  ( new_n14332_, new_n14330_, new_n14326_ );
or   ( new_n14333_, new_n7732_, new_n1523_ );
or   ( new_n14334_, new_n7734_, new_n1525_ );
and  ( new_n14335_, new_n14334_, new_n14333_ );
xor  ( new_n14336_, new_n14335_, new_n7177_ );
nor  ( new_n14337_, new_n14336_, new_n14332_ );
nor  ( new_n14338_, new_n14337_, new_n14331_ );
nor  ( new_n14339_, new_n14338_, new_n14322_ );
nor  ( new_n14340_, new_n14339_, new_n14321_ );
and  ( new_n14341_, new_n14285_, new_n14240_ );
nor  ( new_n14342_, new_n14341_, new_n14340_ );
nor  ( new_n14343_, new_n14342_, new_n14286_ );
and  ( new_n14344_, new_n14343_, new_n14188_ );
nor  ( new_n14345_, new_n14343_, new_n14188_ );
and  ( new_n14346_, new_n371_, RIbb31578_128 );
or   ( new_n14347_, new_n14346_, new_n328_ );
nand ( new_n14348_, new_n14346_, new_n325_ );
and  ( new_n14349_, new_n14348_, new_n14347_ );
xnor ( new_n14350_, new_n14092_, new_n14088_ );
xor  ( new_n14351_, new_n14350_, new_n14098_ );
or   ( new_n14352_, new_n14351_, new_n14349_ );
and  ( new_n14353_, new_n14351_, new_n14349_ );
xor  ( new_n14354_, new_n14074_, new_n14070_ );
xnor ( new_n14355_, new_n14354_, new_n14080_ );
or   ( new_n14356_, new_n14355_, new_n14353_ );
and  ( new_n14357_, new_n14356_, new_n14352_ );
xnor ( new_n14358_, new_n14007_, new_n14003_ );
xor  ( new_n14359_, new_n14358_, new_n14013_ );
xnor ( new_n14360_, new_n14037_, new_n14033_ );
xor  ( new_n14361_, new_n14360_, new_n14043_ );
or   ( new_n14362_, new_n14361_, new_n14359_ );
and  ( new_n14363_, new_n14361_, new_n14359_ );
xor  ( new_n14364_, new_n13955_, new_n13951_ );
xnor ( new_n14365_, new_n14364_, new_n13961_ );
or   ( new_n14366_, new_n14365_, new_n14363_ );
and  ( new_n14367_, new_n14366_, new_n14362_ );
nor  ( new_n14368_, new_n14367_, new_n14357_ );
and  ( new_n14369_, new_n14367_, new_n14357_ );
xnor ( new_n14370_, new_n14058_, new_n14054_ );
xor  ( new_n14371_, new_n14370_, new_n14064_ );
xnor ( new_n14372_, new_n13971_, new_n13967_ );
xor  ( new_n14373_, new_n14372_, new_n13977_ );
nor  ( new_n14374_, new_n14373_, new_n14371_ );
and  ( new_n14375_, new_n14373_, new_n14371_ );
xor  ( new_n14376_, new_n13989_, new_n13985_ );
xnor ( new_n14377_, new_n14376_, new_n13995_ );
nor  ( new_n14378_, new_n14377_, new_n14375_ );
nor  ( new_n14379_, new_n14378_, new_n14374_ );
nor  ( new_n14380_, new_n14379_, new_n14369_ );
nor  ( new_n14381_, new_n14380_, new_n14368_ );
nor  ( new_n14382_, new_n14381_, new_n14345_ );
nor  ( new_n14383_, new_n14382_, new_n14344_ );
and  ( new_n14384_, new_n14383_, new_n14178_ );
not  ( new_n14385_, new_n14384_ );
xor  ( new_n14386_, new_n14127_, new_n14117_ );
xor  ( new_n14387_, new_n14386_, new_n14139_ );
xnor ( new_n14388_, new_n14049_, new_n13999_ );
xor  ( new_n14389_, new_n14388_, new_n14102_ );
nor  ( new_n14390_, new_n14389_, new_n14387_ );
and  ( new_n14391_, new_n14389_, new_n14387_ );
xor  ( new_n14392_, new_n13941_, new_n13939_ );
xnor ( new_n14393_, new_n14392_, new_n13945_ );
nor  ( new_n14394_, new_n14393_, new_n14391_ );
nor  ( new_n14395_, new_n14394_, new_n14390_ );
not  ( new_n14396_, new_n14395_ );
and  ( new_n14397_, new_n14396_, new_n14385_ );
nor  ( new_n14398_, new_n14383_, new_n14178_ );
nor  ( new_n14399_, new_n14398_, new_n14397_ );
xor  ( new_n14400_, new_n13894_, new_n13892_ );
xor  ( new_n14401_, new_n14400_, new_n13898_ );
and  ( new_n14402_, new_n14401_, new_n14399_ );
xnor ( new_n14403_, new_n13769_, new_n13715_ );
xor  ( new_n14404_, new_n14403_, new_n13822_ );
xor  ( new_n14405_, new_n13919_, new_n13909_ );
xor  ( new_n14406_, new_n14405_, new_n13923_ );
nor  ( new_n14407_, new_n14406_, new_n14404_ );
and  ( new_n14408_, new_n14406_, new_n14404_ );
xor  ( new_n14409_, new_n13929_, new_n13927_ );
xnor ( new_n14410_, new_n14409_, new_n13933_ );
not  ( new_n14411_, new_n14410_ );
nor  ( new_n14412_, new_n14411_, new_n14408_ );
nor  ( new_n14413_, new_n14412_, new_n14407_ );
nor  ( new_n14414_, new_n14413_, new_n14402_ );
nor  ( new_n14415_, new_n14401_, new_n14399_ );
or   ( new_n14416_, new_n14415_, new_n14414_ );
xnor ( new_n14417_, new_n13651_, new_n13641_ );
xor  ( new_n14418_, new_n14417_, new_n13869_ );
nand ( new_n14419_, new_n14418_, new_n14416_ );
nor  ( new_n14420_, new_n14418_, new_n14416_ );
xor  ( new_n14421_, new_n13902_, new_n13900_ );
xor  ( new_n14422_, new_n14421_, new_n14145_ );
or   ( new_n14423_, new_n14422_, new_n14420_ );
and  ( new_n14424_, new_n14423_, new_n14419_ );
nor  ( new_n14425_, new_n14424_, new_n14161_ );
xor  ( new_n14426_, new_n14155_, new_n13890_ );
and  ( new_n14427_, new_n14426_, new_n14425_ );
xor  ( new_n14428_, new_n14383_, new_n14178_ );
nor  ( new_n14429_, new_n14428_, new_n14396_ );
not  ( new_n14430_, new_n14398_ );
and  ( new_n14431_, new_n14430_, new_n14397_ );
nor  ( new_n14432_, new_n14431_, new_n14429_ );
xor  ( new_n14433_, new_n14406_, new_n14404_ );
xor  ( new_n14434_, new_n14433_, new_n14410_ );
nand ( new_n14435_, new_n14434_, new_n14432_ );
xnor ( new_n14436_, new_n14343_, new_n14188_ );
xor  ( new_n14437_, new_n14436_, new_n14381_ );
xnor ( new_n14438_, new_n14389_, new_n14387_ );
xor  ( new_n14439_, new_n14438_, new_n14393_ );
nor  ( new_n14440_, new_n14439_, new_n14437_ );
nand ( new_n14441_, new_n14439_, new_n14437_ );
xor  ( new_n14442_, new_n14164_, new_n14162_ );
xor  ( new_n14443_, new_n14442_, new_n14176_ );
and  ( new_n14444_, new_n14443_, new_n14441_ );
or   ( new_n14445_, new_n14444_, new_n14440_ );
xor  ( new_n14446_, new_n14105_, new_n13947_ );
xor  ( new_n14447_, new_n14446_, new_n14141_ );
or   ( new_n14448_, new_n14447_, new_n14445_ );
and  ( new_n14449_, new_n14447_, new_n14445_ );
xor  ( new_n14450_, new_n14285_, new_n14240_ );
xnor ( new_n14451_, new_n14450_, new_n14340_ );
not  ( new_n14452_, new_n14451_ );
xnor ( new_n14453_, new_n14367_, new_n14357_ );
xor  ( new_n14454_, new_n14453_, new_n14379_ );
and  ( new_n14455_, new_n14454_, new_n14452_ );
xnor ( new_n14456_, new_n14212_, new_n14208_ );
xor  ( new_n14457_, new_n14456_, new_n14218_ );
xnor ( new_n14458_, new_n14196_, new_n14192_ );
xor  ( new_n14459_, new_n14458_, new_n14202_ );
or   ( new_n14460_, new_n14459_, new_n14457_ );
and  ( new_n14461_, new_n14459_, new_n14457_ );
xor  ( new_n14462_, new_n14230_, new_n14226_ );
xnor ( new_n14463_, new_n14462_, new_n14236_ );
or   ( new_n14464_, new_n14463_, new_n14461_ );
and  ( new_n14465_, new_n14464_, new_n14460_ );
xnor ( new_n14466_, new_n14248_, new_n14244_ );
xor  ( new_n14467_, new_n14466_, new_n14254_ );
xnor ( new_n14468_, new_n14273_, new_n14269_ );
xor  ( new_n14469_, new_n14468_, new_n14279_ );
or   ( new_n14470_, new_n14469_, new_n14467_ );
nand ( new_n14471_, new_n14469_, new_n14467_ );
xor  ( new_n14472_, new_n14264_, new_n14260_ );
nand ( new_n14473_, new_n14472_, new_n14471_ );
and  ( new_n14474_, new_n14473_, new_n14470_ );
nor  ( new_n14475_, new_n14474_, new_n14465_ );
nand ( new_n14476_, new_n14474_, new_n14465_ );
xnor ( new_n14477_, new_n14312_, new_n14308_ );
xor  ( new_n14478_, new_n14477_, new_n14318_ );
xnor ( new_n14479_, new_n14296_, new_n14290_ );
xor  ( new_n14480_, new_n14479_, new_n14302_ );
nor  ( new_n14481_, new_n14480_, new_n14478_ );
nand ( new_n14482_, new_n14480_, new_n14478_ );
xor  ( new_n14483_, new_n14330_, new_n14326_ );
xor  ( new_n14484_, new_n14483_, new_n14336_ );
and  ( new_n14485_, new_n14484_, new_n14482_ );
or   ( new_n14486_, new_n14485_, new_n14481_ );
and  ( new_n14487_, new_n14486_, new_n14476_ );
or   ( new_n14488_, new_n14487_, new_n14475_ );
or   ( new_n14489_, new_n6173_, new_n2646_ );
or   ( new_n14490_, new_n6175_, new_n2475_ );
and  ( new_n14491_, new_n14490_, new_n14489_ );
xor  ( new_n14492_, new_n14491_, new_n5597_ );
or   ( new_n14493_, new_n5604_, new_n2981_ );
or   ( new_n14494_, new_n5606_, new_n2751_ );
and  ( new_n14495_, new_n14494_, new_n14493_ );
xor  ( new_n14496_, new_n14495_, new_n5206_ );
or   ( new_n14497_, new_n14496_, new_n14492_ );
and  ( new_n14498_, new_n14496_, new_n14492_ );
or   ( new_n14499_, new_n5207_, new_n3306_ );
or   ( new_n14500_, new_n5209_, new_n3178_ );
and  ( new_n14501_, new_n14500_, new_n14499_ );
xor  ( new_n14502_, new_n14501_, new_n4708_ );
or   ( new_n14503_, new_n14502_, new_n14498_ );
and  ( new_n14504_, new_n14503_, new_n14497_ );
or   ( new_n14505_, new_n4709_, new_n3694_ );
or   ( new_n14506_, new_n4711_, new_n3696_ );
and  ( new_n14507_, new_n14506_, new_n14505_ );
xor  ( new_n14508_, new_n14507_, new_n4295_ );
or   ( new_n14509_, new_n4302_, new_n4069_ );
or   ( new_n14510_, new_n4304_, new_n3820_ );
and  ( new_n14511_, new_n14510_, new_n14509_ );
xor  ( new_n14512_, new_n14511_, new_n3895_ );
or   ( new_n14513_, new_n14512_, new_n14508_ );
and  ( new_n14514_, new_n14512_, new_n14508_ );
or   ( new_n14515_, new_n3896_, new_n4603_ );
or   ( new_n14516_, new_n3898_, new_n4267_ );
and  ( new_n14517_, new_n14516_, new_n14515_ );
xor  ( new_n14518_, new_n14517_, new_n3460_ );
or   ( new_n14519_, new_n14518_, new_n14514_ );
and  ( new_n14520_, new_n14519_, new_n14513_ );
or   ( new_n14521_, new_n14520_, new_n14504_ );
and  ( new_n14522_, new_n14520_, new_n14504_ );
or   ( new_n14523_, new_n3461_, new_n4859_ );
or   ( new_n14524_, new_n3463_, new_n4995_ );
and  ( new_n14525_, new_n14524_, new_n14523_ );
xor  ( new_n14526_, new_n14525_, new_n3116_ );
or   ( new_n14527_, new_n3117_, new_n5428_ );
or   ( new_n14528_, new_n3119_, new_n5171_ );
and  ( new_n14529_, new_n14528_, new_n14527_ );
xor  ( new_n14530_, new_n14529_, new_n2800_ );
or   ( new_n14531_, new_n14530_, new_n14526_ );
and  ( new_n14532_, new_n14530_, new_n14526_ );
or   ( new_n14533_, new_n2807_, new_n5899_ );
or   ( new_n14534_, new_n2809_, new_n5570_ );
and  ( new_n14535_, new_n14534_, new_n14533_ );
xor  ( new_n14536_, new_n14535_, new_n2424_ );
or   ( new_n14537_, new_n14536_, new_n14532_ );
and  ( new_n14538_, new_n14537_, new_n14531_ );
or   ( new_n14539_, new_n14538_, new_n14522_ );
and  ( new_n14540_, new_n14539_, new_n14521_ );
or   ( new_n14541_, new_n7732_, new_n1754_ );
or   ( new_n14542_, new_n7734_, new_n1523_ );
and  ( new_n14543_, new_n14542_, new_n14541_ );
xor  ( new_n14544_, new_n14543_, new_n7177_ );
or   ( new_n14545_, new_n7184_, new_n2057_ );
or   ( new_n14546_, new_n7186_, new_n1899_ );
and  ( new_n14547_, new_n14546_, new_n14545_ );
xor  ( new_n14548_, new_n14547_, new_n6638_ );
nor  ( new_n14549_, new_n14548_, new_n14544_ );
and  ( new_n14550_, new_n14548_, new_n14544_ );
or   ( new_n14551_, new_n6645_, new_n2291_ );
or   ( new_n14552_, new_n6647_, new_n2178_ );
and  ( new_n14553_, new_n14552_, new_n14551_ );
xor  ( new_n14554_, new_n14553_, new_n6166_ );
nor  ( new_n14555_, new_n14554_, new_n14550_ );
nor  ( new_n14556_, new_n14555_, new_n14549_ );
or   ( new_n14557_, new_n10059_, new_n805_ );
or   ( new_n14558_, new_n10061_, new_n775_ );
and  ( new_n14559_, new_n14558_, new_n14557_ );
xor  ( new_n14560_, new_n14559_, new_n9421_ );
and  ( new_n14561_, RIbb2d888_64, RIbb2d1f8_78 );
or   ( new_n14562_, RIbb2d888_64, new_n515_ );
and  ( new_n14563_, new_n14562_, RIbb2d900_63 );
or   ( new_n14564_, new_n14563_, new_n14561_ );
or   ( new_n14565_, new_n10770_, new_n509_ );
and  ( new_n14566_, new_n14565_, new_n14564_ );
nor  ( new_n14567_, new_n14566_, new_n14560_ );
and  ( new_n14568_, new_n14566_, new_n14560_ );
nor  ( new_n14569_, new_n14568_, new_n402_ );
nor  ( new_n14570_, new_n14569_, new_n14567_ );
or   ( new_n14571_, new_n9422_, new_n986_ );
or   ( new_n14572_, new_n9424_, new_n886_ );
and  ( new_n14573_, new_n14572_, new_n14571_ );
xor  ( new_n14574_, new_n14573_, new_n8873_ );
or   ( new_n14575_, new_n8874_, new_n1213_ );
or   ( new_n14576_, new_n8876_, new_n1168_ );
and  ( new_n14577_, new_n14576_, new_n14575_ );
xor  ( new_n14578_, new_n14577_, new_n8257_ );
or   ( new_n14579_, new_n14578_, new_n14574_ );
and  ( new_n14580_, new_n14578_, new_n14574_ );
or   ( new_n14581_, new_n8264_, new_n1525_ );
or   ( new_n14582_, new_n8266_, new_n1318_ );
and  ( new_n14583_, new_n14582_, new_n14581_ );
xor  ( new_n14584_, new_n14583_, new_n7725_ );
or   ( new_n14585_, new_n14584_, new_n14580_ );
and  ( new_n14586_, new_n14585_, new_n14579_ );
and  ( new_n14587_, new_n14586_, new_n14570_ );
or   ( new_n14588_, new_n14587_, new_n14556_ );
or   ( new_n14589_, new_n14586_, new_n14570_ );
and  ( new_n14590_, new_n14589_, new_n14588_ );
or   ( new_n14591_, new_n14590_, new_n14540_ );
and  ( new_n14592_, new_n14590_, new_n14540_ );
or   ( new_n14593_, new_n1593_, new_n8115_ );
or   ( new_n14594_, new_n1595_, new_n8117_ );
and  ( new_n14595_, new_n14594_, new_n14593_ );
xor  ( new_n14596_, new_n14595_, new_n1358_ );
or   ( new_n14597_, new_n1364_, new_n8481_ );
or   ( new_n14598_, new_n1366_, new_n8352_ );
and  ( new_n14599_, new_n14598_, new_n14597_ );
xor  ( new_n14600_, new_n14599_, new_n1129_ );
nor  ( new_n14601_, new_n14600_, new_n14596_ );
and  ( new_n14602_, new_n14600_, new_n14596_ );
or   ( new_n14603_, new_n1135_, new_n9099_ );
or   ( new_n14604_, new_n1137_, new_n8995_ );
and  ( new_n14605_, new_n14604_, new_n14603_ );
xor  ( new_n14606_, new_n14605_, new_n896_ );
nor  ( new_n14607_, new_n14606_, new_n14602_ );
nor  ( new_n14608_, new_n14607_, new_n14601_ );
or   ( new_n14609_, new_n2425_, new_n6425_ );
or   ( new_n14610_, new_n2427_, new_n6219_ );
and  ( new_n14611_, new_n14610_, new_n14609_ );
xor  ( new_n14612_, new_n14611_, new_n2121_ );
or   ( new_n14613_, new_n2122_, new_n6943_ );
or   ( new_n14614_, new_n2124_, new_n6589_ );
and  ( new_n14615_, new_n14614_, new_n14613_ );
xor  ( new_n14616_, new_n14615_, new_n1843_ );
or   ( new_n14617_, new_n14616_, new_n14612_ );
and  ( new_n14618_, new_n14616_, new_n14612_ );
or   ( new_n14619_, new_n1844_, new_n7373_ );
or   ( new_n14620_, new_n1846_, new_n7149_ );
and  ( new_n14621_, new_n14620_, new_n14619_ );
xor  ( new_n14622_, new_n14621_, new_n1586_ );
or   ( new_n14623_, new_n14622_, new_n14618_ );
and  ( new_n14624_, new_n14623_, new_n14617_ );
and  ( new_n14625_, new_n14624_, new_n14608_ );
or   ( new_n14626_, new_n14624_, new_n14608_ );
or   ( new_n14627_, new_n897_, new_n9679_ );
or   ( new_n14628_, new_n899_, new_n9681_ );
and  ( new_n14629_, new_n14628_, new_n14627_ );
xor  ( new_n14630_, new_n14629_, new_n748_ );
or   ( new_n14631_, new_n755_, new_n10541_ );
or   ( new_n14632_, new_n757_, new_n10220_ );
and  ( new_n14633_, new_n14632_, new_n14631_ );
xor  ( new_n14634_, new_n14633_, new_n523_ );
and  ( new_n14635_, new_n14634_, new_n14630_ );
or   ( new_n14636_, new_n14634_, new_n14630_ );
and  ( new_n14637_, new_n454_, RIbb31578_128 );
nor  ( new_n14638_, new_n14637_, new_n403_ );
and  ( new_n14639_, new_n14637_, new_n400_ );
or   ( new_n14640_, new_n14639_, new_n14638_ );
and  ( new_n14641_, new_n14640_, new_n14636_ );
or   ( new_n14642_, new_n14641_, new_n14635_ );
and  ( new_n14643_, new_n14642_, new_n14626_ );
or   ( new_n14644_, new_n14643_, new_n14625_ );
or   ( new_n14645_, new_n14644_, new_n14592_ );
and  ( new_n14646_, new_n14645_, new_n14591_ );
or   ( new_n14647_, new_n14646_, new_n14488_ );
and  ( new_n14648_, new_n14646_, new_n14488_ );
xor  ( new_n14649_, new_n14025_, new_n14019_ );
xor  ( new_n14650_, new_n14649_, new_n327_ );
xnor ( new_n14651_, new_n14361_, new_n14359_ );
xor  ( new_n14652_, new_n14651_, new_n14365_ );
and  ( new_n14653_, new_n14652_, new_n14650_ );
or   ( new_n14654_, new_n14652_, new_n14650_ );
xor  ( new_n14655_, new_n14373_, new_n14371_ );
xnor ( new_n14656_, new_n14655_, new_n14377_ );
and  ( new_n14657_, new_n14656_, new_n14654_ );
or   ( new_n14658_, new_n14657_, new_n14653_ );
or   ( new_n14659_, new_n14658_, new_n14648_ );
and  ( new_n14660_, new_n14659_, new_n14647_ );
and  ( new_n14661_, new_n14660_, new_n14455_ );
nor  ( new_n14662_, new_n14660_, new_n14455_ );
xor  ( new_n14663_, new_n14182_, new_n14180_ );
xor  ( new_n14664_, new_n14663_, new_n14186_ );
xnor ( new_n14665_, new_n14170_, new_n14168_ );
xor  ( new_n14666_, new_n14665_, new_n14174_ );
and  ( new_n14667_, new_n14666_, new_n14664_ );
nor  ( new_n14668_, new_n14666_, new_n14664_ );
xor  ( new_n14669_, new_n14220_, new_n14204_ );
xor  ( new_n14670_, new_n14669_, new_n14238_ );
xor  ( new_n14671_, new_n14281_, new_n14265_ );
xor  ( new_n14672_, new_n14671_, new_n14256_ );
and  ( new_n14673_, new_n14672_, new_n14670_ );
nor  ( new_n14674_, new_n14672_, new_n14670_ );
xor  ( new_n14675_, new_n14351_, new_n14349_ );
xnor ( new_n14676_, new_n14675_, new_n14355_ );
not  ( new_n14677_, new_n14676_ );
nor  ( new_n14678_, new_n14677_, new_n14674_ );
nor  ( new_n14679_, new_n14678_, new_n14673_ );
nor  ( new_n14680_, new_n14679_, new_n14668_ );
nor  ( new_n14681_, new_n14680_, new_n14667_ );
nor  ( new_n14682_, new_n14681_, new_n14662_ );
nor  ( new_n14683_, new_n14682_, new_n14661_ );
or   ( new_n14684_, new_n14683_, new_n14449_ );
and  ( new_n14685_, new_n14684_, new_n14448_ );
nor  ( new_n14686_, new_n14685_, new_n14435_ );
nand ( new_n14687_, new_n14685_, new_n14435_ );
xor  ( new_n14688_, new_n13935_, new_n13925_ );
xnor ( new_n14689_, new_n14688_, new_n14143_ );
and  ( new_n14690_, new_n14689_, new_n14687_ );
or   ( new_n14691_, new_n14690_, new_n14686_ );
xnor ( new_n14692_, new_n14418_, new_n14416_ );
xor  ( new_n14693_, new_n14692_, new_n14422_ );
and  ( new_n14694_, new_n14693_, new_n14691_ );
xor  ( new_n14695_, new_n14424_, new_n14161_ );
and  ( new_n14696_, new_n14695_, new_n14694_ );
xor  ( new_n14697_, new_n14685_, new_n14435_ );
xnor ( new_n14698_, new_n14697_, new_n14689_ );
xor  ( new_n14699_, new_n14401_, new_n14399_ );
xor  ( new_n14700_, new_n14699_, new_n14413_ );
nor  ( new_n14701_, new_n14700_, new_n14698_ );
xor  ( new_n14702_, new_n14693_, new_n14691_ );
and  ( new_n14703_, new_n14702_, new_n14701_ );
xnor ( new_n14704_, new_n14700_, new_n14698_ );
xor  ( new_n14705_, new_n14520_, new_n14504_ );
xor  ( new_n14706_, new_n14705_, new_n14538_ );
xor  ( new_n14707_, new_n14586_, new_n14570_ );
xor  ( new_n14708_, new_n14707_, new_n14556_ );
nor  ( new_n14709_, new_n14708_, new_n14706_ );
nand ( new_n14710_, new_n14708_, new_n14706_ );
xnor ( new_n14711_, new_n14624_, new_n14608_ );
xor  ( new_n14712_, new_n14711_, new_n14642_ );
and  ( new_n14713_, new_n14712_, new_n14710_ );
or   ( new_n14714_, new_n14713_, new_n14709_ );
xnor ( new_n14715_, new_n14320_, new_n14304_ );
xor  ( new_n14716_, new_n14715_, new_n14338_ );
nor  ( new_n14717_, new_n14716_, new_n14714_ );
and  ( new_n14718_, new_n14716_, new_n14714_ );
xor  ( new_n14719_, new_n14672_, new_n14670_ );
xor  ( new_n14720_, new_n14719_, new_n14676_ );
not  ( new_n14721_, new_n14720_ );
nor  ( new_n14722_, new_n14721_, new_n14718_ );
nor  ( new_n14723_, new_n14722_, new_n14717_ );
xor  ( new_n14724_, new_n14480_, new_n14478_ );
xor  ( new_n14725_, new_n14724_, new_n14484_ );
xnor ( new_n14726_, new_n14459_, new_n14457_ );
xor  ( new_n14727_, new_n14726_, new_n14463_ );
or   ( new_n14728_, new_n14727_, new_n14725_ );
and  ( new_n14729_, new_n14727_, new_n14725_ );
xor  ( new_n14730_, new_n14469_, new_n14467_ );
xor  ( new_n14731_, new_n14730_, new_n14472_ );
or   ( new_n14732_, new_n14731_, new_n14729_ );
and  ( new_n14733_, new_n14732_, new_n14728_ );
or   ( new_n14734_, new_n10059_, new_n886_ );
or   ( new_n14735_, new_n10061_, new_n805_ );
and  ( new_n14736_, new_n14735_, new_n14734_ );
xor  ( new_n14737_, new_n14736_, new_n9421_ );
and  ( new_n14738_, RIbb2d888_64, RIbb2d180_79 );
or   ( new_n14739_, RIbb2d888_64, new_n775_ );
and  ( new_n14740_, new_n14739_, RIbb2d900_63 );
or   ( new_n14741_, new_n14740_, new_n14738_ );
or   ( new_n14742_, new_n10770_, new_n515_ );
and  ( new_n14743_, new_n14742_, new_n14741_ );
or   ( new_n14744_, new_n14743_, new_n14737_ );
and  ( new_n14745_, new_n14743_, new_n14737_ );
or   ( new_n14746_, new_n9422_, new_n1168_ );
or   ( new_n14747_, new_n9424_, new_n986_ );
and  ( new_n14748_, new_n14747_, new_n14746_ );
xor  ( new_n14749_, new_n14748_, new_n8873_ );
or   ( new_n14750_, new_n14749_, new_n14745_ );
and  ( new_n14751_, new_n14750_, new_n14744_ );
or   ( new_n14752_, new_n7184_, new_n2178_ );
or   ( new_n14753_, new_n7186_, new_n2057_ );
and  ( new_n14754_, new_n14753_, new_n14752_ );
xor  ( new_n14755_, new_n14754_, new_n6638_ );
or   ( new_n14756_, new_n6645_, new_n2475_ );
or   ( new_n14757_, new_n6647_, new_n2291_ );
and  ( new_n14758_, new_n14757_, new_n14756_ );
xor  ( new_n14759_, new_n14758_, new_n6166_ );
or   ( new_n14760_, new_n14759_, new_n14755_ );
and  ( new_n14761_, new_n14759_, new_n14755_ );
or   ( new_n14762_, new_n6173_, new_n2751_ );
or   ( new_n14763_, new_n6175_, new_n2646_ );
and  ( new_n14764_, new_n14763_, new_n14762_ );
xor  ( new_n14765_, new_n14764_, new_n5597_ );
or   ( new_n14766_, new_n14765_, new_n14761_ );
and  ( new_n14767_, new_n14766_, new_n14760_ );
or   ( new_n14768_, new_n14767_, new_n14751_ );
and  ( new_n14769_, new_n14767_, new_n14751_ );
or   ( new_n14770_, new_n8874_, new_n1318_ );
or   ( new_n14771_, new_n8876_, new_n1213_ );
and  ( new_n14772_, new_n14771_, new_n14770_ );
xor  ( new_n14773_, new_n14772_, new_n8257_ );
or   ( new_n14774_, new_n8264_, new_n1523_ );
or   ( new_n14775_, new_n8266_, new_n1525_ );
and  ( new_n14776_, new_n14775_, new_n14774_ );
xor  ( new_n14777_, new_n14776_, new_n7725_ );
nor  ( new_n14778_, new_n14777_, new_n14773_ );
and  ( new_n14779_, new_n14777_, new_n14773_ );
or   ( new_n14780_, new_n7732_, new_n1899_ );
or   ( new_n14781_, new_n7734_, new_n1754_ );
and  ( new_n14782_, new_n14781_, new_n14780_ );
xor  ( new_n14783_, new_n14782_, new_n7177_ );
nor  ( new_n14784_, new_n14783_, new_n14779_ );
nor  ( new_n14785_, new_n14784_, new_n14778_ );
or   ( new_n14786_, new_n14785_, new_n14769_ );
and  ( new_n14787_, new_n14786_, new_n14768_ );
xor  ( new_n14788_, new_n14634_, new_n14630_ );
xor  ( new_n14789_, new_n14788_, new_n14640_ );
or   ( new_n14790_, new_n1364_, new_n8995_ );
or   ( new_n14791_, new_n1366_, new_n8481_ );
and  ( new_n14792_, new_n14791_, new_n14790_ );
xor  ( new_n14793_, new_n14792_, new_n1129_ );
or   ( new_n14794_, new_n1135_, new_n9681_ );
or   ( new_n14795_, new_n1137_, new_n9099_ );
and  ( new_n14796_, new_n14795_, new_n14794_ );
xor  ( new_n14797_, new_n14796_, new_n896_ );
or   ( new_n14798_, new_n14797_, new_n14793_ );
and  ( new_n14799_, new_n14797_, new_n14793_ );
or   ( new_n14800_, new_n897_, new_n10220_ );
or   ( new_n14801_, new_n899_, new_n9679_ );
and  ( new_n14802_, new_n14801_, new_n14800_ );
xor  ( new_n14803_, new_n14802_, new_n748_ );
or   ( new_n14804_, new_n14803_, new_n14799_ );
and  ( new_n14805_, new_n14804_, new_n14798_ );
or   ( new_n14806_, new_n14805_, new_n14789_ );
and  ( new_n14807_, new_n14805_, new_n14789_ );
or   ( new_n14808_, new_n2122_, new_n7149_ );
or   ( new_n14809_, new_n2124_, new_n6943_ );
and  ( new_n14810_, new_n14809_, new_n14808_ );
xor  ( new_n14811_, new_n14810_, new_n1843_ );
or   ( new_n14812_, new_n1844_, new_n8117_ );
or   ( new_n14813_, new_n1846_, new_n7373_ );
and  ( new_n14814_, new_n14813_, new_n14812_ );
xor  ( new_n14815_, new_n14814_, new_n1586_ );
nor  ( new_n14816_, new_n14815_, new_n14811_ );
and  ( new_n14817_, new_n14815_, new_n14811_ );
or   ( new_n14818_, new_n1593_, new_n8352_ );
or   ( new_n14819_, new_n1595_, new_n8115_ );
and  ( new_n14820_, new_n14819_, new_n14818_ );
xor  ( new_n14821_, new_n14820_, new_n1358_ );
nor  ( new_n14822_, new_n14821_, new_n14817_ );
nor  ( new_n14823_, new_n14822_, new_n14816_ );
or   ( new_n14824_, new_n14823_, new_n14807_ );
and  ( new_n14825_, new_n14824_, new_n14806_ );
or   ( new_n14826_, new_n14825_, new_n14787_ );
and  ( new_n14827_, new_n14825_, new_n14787_ );
or   ( new_n14828_, new_n5604_, new_n3178_ );
or   ( new_n14829_, new_n5606_, new_n2981_ );
and  ( new_n14830_, new_n14829_, new_n14828_ );
xor  ( new_n14831_, new_n14830_, new_n5206_ );
or   ( new_n14832_, new_n5207_, new_n3696_ );
or   ( new_n14833_, new_n5209_, new_n3306_ );
and  ( new_n14834_, new_n14833_, new_n14832_ );
xor  ( new_n14835_, new_n14834_, new_n4708_ );
or   ( new_n14836_, new_n14835_, new_n14831_ );
and  ( new_n14837_, new_n14835_, new_n14831_ );
or   ( new_n14838_, new_n4709_, new_n3820_ );
or   ( new_n14839_, new_n4711_, new_n3694_ );
and  ( new_n14840_, new_n14839_, new_n14838_ );
xor  ( new_n14841_, new_n14840_, new_n4295_ );
or   ( new_n14842_, new_n14841_, new_n14837_ );
and  ( new_n14843_, new_n14842_, new_n14836_ );
or   ( new_n14844_, new_n4302_, new_n4267_ );
or   ( new_n14845_, new_n4304_, new_n4069_ );
and  ( new_n14846_, new_n14845_, new_n14844_ );
xor  ( new_n14847_, new_n14846_, new_n3895_ );
or   ( new_n14848_, new_n3896_, new_n4995_ );
or   ( new_n14849_, new_n3898_, new_n4603_ );
and  ( new_n14850_, new_n14849_, new_n14848_ );
xor  ( new_n14851_, new_n14850_, new_n3460_ );
or   ( new_n14852_, new_n14851_, new_n14847_ );
and  ( new_n14853_, new_n14851_, new_n14847_ );
or   ( new_n14854_, new_n3461_, new_n5171_ );
or   ( new_n14855_, new_n3463_, new_n4859_ );
and  ( new_n14856_, new_n14855_, new_n14854_ );
xor  ( new_n14857_, new_n14856_, new_n3116_ );
or   ( new_n14858_, new_n14857_, new_n14853_ );
and  ( new_n14859_, new_n14858_, new_n14852_ );
nor  ( new_n14860_, new_n14859_, new_n14843_ );
and  ( new_n14861_, new_n14859_, new_n14843_ );
or   ( new_n14862_, new_n3117_, new_n5570_ );
or   ( new_n14863_, new_n3119_, new_n5428_ );
and  ( new_n14864_, new_n14863_, new_n14862_ );
xor  ( new_n14865_, new_n14864_, new_n2800_ );
or   ( new_n14866_, new_n2807_, new_n6219_ );
or   ( new_n14867_, new_n2809_, new_n5899_ );
and  ( new_n14868_, new_n14867_, new_n14866_ );
xor  ( new_n14869_, new_n14868_, new_n2424_ );
nor  ( new_n14870_, new_n14869_, new_n14865_ );
and  ( new_n14871_, new_n14869_, new_n14865_ );
or   ( new_n14872_, new_n2425_, new_n6589_ );
or   ( new_n14873_, new_n2427_, new_n6425_ );
and  ( new_n14874_, new_n14873_, new_n14872_ );
xor  ( new_n14875_, new_n14874_, new_n2121_ );
nor  ( new_n14876_, new_n14875_, new_n14871_ );
nor  ( new_n14877_, new_n14876_, new_n14870_ );
nor  ( new_n14878_, new_n14877_, new_n14861_ );
nor  ( new_n14879_, new_n14878_, new_n14860_ );
or   ( new_n14880_, new_n14879_, new_n14827_ );
and  ( new_n14881_, new_n14880_, new_n14826_ );
and  ( new_n14882_, new_n14881_, new_n14733_ );
nor  ( new_n14883_, new_n14881_, new_n14733_ );
xor  ( new_n14884_, new_n14578_, new_n14574_ );
xnor ( new_n14885_, new_n14884_, new_n14584_ );
xor  ( new_n14886_, new_n14566_, new_n14560_ );
xor  ( new_n14887_, new_n14886_, new_n403_ );
or   ( new_n14888_, new_n14887_, new_n14885_ );
xnor ( new_n14889_, new_n14616_, new_n14612_ );
xor  ( new_n14890_, new_n14889_, new_n14622_ );
xnor ( new_n14891_, new_n14530_, new_n14526_ );
xor  ( new_n14892_, new_n14891_, new_n14536_ );
or   ( new_n14893_, new_n14892_, new_n14890_ );
and  ( new_n14894_, new_n14892_, new_n14890_ );
xor  ( new_n14895_, new_n14600_, new_n14596_ );
xnor ( new_n14896_, new_n14895_, new_n14606_ );
or   ( new_n14897_, new_n14896_, new_n14894_ );
and  ( new_n14898_, new_n14897_, new_n14893_ );
nor  ( new_n14899_, new_n14898_, new_n14888_ );
and  ( new_n14900_, new_n14898_, new_n14888_ );
xnor ( new_n14901_, new_n14512_, new_n14508_ );
xor  ( new_n14902_, new_n14901_, new_n14518_ );
xnor ( new_n14903_, new_n14496_, new_n14492_ );
xor  ( new_n14904_, new_n14903_, new_n14502_ );
nor  ( new_n14905_, new_n14904_, new_n14902_ );
and  ( new_n14906_, new_n14904_, new_n14902_ );
xor  ( new_n14907_, new_n14548_, new_n14544_ );
xnor ( new_n14908_, new_n14907_, new_n14554_ );
nor  ( new_n14909_, new_n14908_, new_n14906_ );
nor  ( new_n14910_, new_n14909_, new_n14905_ );
nor  ( new_n14911_, new_n14910_, new_n14900_ );
nor  ( new_n14912_, new_n14911_, new_n14899_ );
nor  ( new_n14913_, new_n14912_, new_n14883_ );
nor  ( new_n14914_, new_n14913_, new_n14882_ );
and  ( new_n14915_, new_n14914_, new_n14723_ );
xor  ( new_n14916_, new_n14590_, new_n14540_ );
xor  ( new_n14917_, new_n14916_, new_n14644_ );
xor  ( new_n14918_, new_n14474_, new_n14465_ );
xor  ( new_n14919_, new_n14918_, new_n14486_ );
and  ( new_n14920_, new_n14919_, new_n14917_ );
nor  ( new_n14921_, new_n14919_, new_n14917_ );
xor  ( new_n14922_, new_n14652_, new_n14650_ );
xnor ( new_n14923_, new_n14922_, new_n14656_ );
nor  ( new_n14924_, new_n14923_, new_n14921_ );
nor  ( new_n14925_, new_n14924_, new_n14920_ );
nor  ( new_n14926_, new_n14925_, new_n14915_ );
nor  ( new_n14927_, new_n14914_, new_n14723_ );
nor  ( new_n14928_, new_n14927_, new_n14926_ );
xor  ( new_n14929_, new_n14439_, new_n14437_ );
xor  ( new_n14930_, new_n14929_, new_n14443_ );
and  ( new_n14931_, new_n14930_, new_n14928_ );
xor  ( new_n14932_, new_n14646_, new_n14488_ );
xor  ( new_n14933_, new_n14932_, new_n14658_ );
xnor ( new_n14934_, new_n14666_, new_n14664_ );
xor  ( new_n14935_, new_n14934_, new_n14679_ );
and  ( new_n14936_, new_n14935_, new_n14933_ );
nor  ( new_n14937_, new_n14935_, new_n14933_ );
xor  ( new_n14938_, new_n14454_, new_n14452_ );
not  ( new_n14939_, new_n14938_ );
nor  ( new_n14940_, new_n14939_, new_n14937_ );
nor  ( new_n14941_, new_n14940_, new_n14936_ );
nor  ( new_n14942_, new_n14941_, new_n14931_ );
nor  ( new_n14943_, new_n14930_, new_n14928_ );
or   ( new_n14944_, new_n14943_, new_n14942_ );
xnor ( new_n14945_, new_n14447_, new_n14445_ );
xor  ( new_n14946_, new_n14945_, new_n14683_ );
nand ( new_n14947_, new_n14946_, new_n14944_ );
nor  ( new_n14948_, new_n14946_, new_n14944_ );
xnor ( new_n14949_, new_n14434_, new_n14432_ );
or   ( new_n14950_, new_n14949_, new_n14948_ );
and  ( new_n14951_, new_n14950_, new_n14947_ );
nor  ( new_n14952_, new_n14951_, new_n14704_ );
xor  ( new_n14953_, new_n14946_, new_n14944_ );
xor  ( new_n14954_, new_n14953_, new_n14949_ );
xnor ( new_n14955_, new_n14914_, new_n14723_ );
nand ( new_n14956_, new_n14955_, new_n14925_ );
or   ( new_n14957_, new_n14925_, new_n14915_ );
or   ( new_n14958_, new_n14927_, new_n14957_ );
and  ( new_n14959_, new_n14958_, new_n14956_ );
xor  ( new_n14960_, new_n14919_, new_n14917_ );
xor  ( new_n14961_, new_n14960_, new_n14923_ );
xnor ( new_n14962_, new_n14892_, new_n14890_ );
xor  ( new_n14963_, new_n14962_, new_n14896_ );
xnor ( new_n14964_, new_n14904_, new_n14902_ );
xor  ( new_n14965_, new_n14964_, new_n14908_ );
or   ( new_n14966_, new_n14965_, new_n14963_ );
and  ( new_n14967_, new_n14965_, new_n14963_ );
xor  ( new_n14968_, new_n14887_, new_n14885_ );
or   ( new_n14969_, new_n14968_, new_n14967_ );
and  ( new_n14970_, new_n14969_, new_n14966_ );
or   ( new_n14971_, new_n6173_, new_n2981_ );
or   ( new_n14972_, new_n6175_, new_n2751_ );
and  ( new_n14973_, new_n14972_, new_n14971_ );
xor  ( new_n14974_, new_n14973_, new_n5597_ );
or   ( new_n14975_, new_n5604_, new_n3306_ );
or   ( new_n14976_, new_n5606_, new_n3178_ );
and  ( new_n14977_, new_n14976_, new_n14975_ );
xor  ( new_n14978_, new_n14977_, new_n5206_ );
or   ( new_n14979_, new_n14978_, new_n14974_ );
and  ( new_n14980_, new_n14978_, new_n14974_ );
or   ( new_n14981_, new_n5207_, new_n3694_ );
or   ( new_n14982_, new_n5209_, new_n3696_ );
and  ( new_n14983_, new_n14982_, new_n14981_ );
xor  ( new_n14984_, new_n14983_, new_n4708_ );
or   ( new_n14985_, new_n14984_, new_n14980_ );
and  ( new_n14986_, new_n14985_, new_n14979_ );
or   ( new_n14987_, new_n4709_, new_n4069_ );
or   ( new_n14988_, new_n4711_, new_n3820_ );
and  ( new_n14989_, new_n14988_, new_n14987_ );
xor  ( new_n14990_, new_n14989_, new_n4295_ );
or   ( new_n14991_, new_n4302_, new_n4603_ );
or   ( new_n14992_, new_n4304_, new_n4267_ );
and  ( new_n14993_, new_n14992_, new_n14991_ );
xor  ( new_n14994_, new_n14993_, new_n3895_ );
or   ( new_n14995_, new_n14994_, new_n14990_ );
and  ( new_n14996_, new_n14994_, new_n14990_ );
or   ( new_n14997_, new_n3896_, new_n4859_ );
or   ( new_n14998_, new_n3898_, new_n4995_ );
and  ( new_n14999_, new_n14998_, new_n14997_ );
xor  ( new_n15000_, new_n14999_, new_n3460_ );
or   ( new_n15001_, new_n15000_, new_n14996_ );
and  ( new_n15002_, new_n15001_, new_n14995_ );
or   ( new_n15003_, new_n15002_, new_n14986_ );
and  ( new_n15004_, new_n15002_, new_n14986_ );
or   ( new_n15005_, new_n3461_, new_n5428_ );
or   ( new_n15006_, new_n3463_, new_n5171_ );
and  ( new_n15007_, new_n15006_, new_n15005_ );
xor  ( new_n15008_, new_n15007_, new_n3116_ );
or   ( new_n15009_, new_n3117_, new_n5899_ );
or   ( new_n15010_, new_n3119_, new_n5570_ );
and  ( new_n15011_, new_n15010_, new_n15009_ );
xor  ( new_n15012_, new_n15011_, new_n2800_ );
nor  ( new_n15013_, new_n15012_, new_n15008_ );
and  ( new_n15014_, new_n15012_, new_n15008_ );
or   ( new_n15015_, new_n2807_, new_n6425_ );
or   ( new_n15016_, new_n2809_, new_n6219_ );
and  ( new_n15017_, new_n15016_, new_n15015_ );
xor  ( new_n15018_, new_n15017_, new_n2424_ );
nor  ( new_n15019_, new_n15018_, new_n15014_ );
nor  ( new_n15020_, new_n15019_, new_n15013_ );
or   ( new_n15021_, new_n15020_, new_n15004_ );
and  ( new_n15022_, new_n15021_, new_n15003_ );
or   ( new_n15023_, new_n755_, new_n10841_ );
or   ( new_n15024_, new_n757_, new_n10541_ );
and  ( new_n15025_, new_n15024_, new_n15023_ );
xor  ( new_n15026_, new_n15025_, new_n523_ );
or   ( new_n15027_, new_n2425_, new_n6943_ );
or   ( new_n15028_, new_n2427_, new_n6589_ );
and  ( new_n15029_, new_n15028_, new_n15027_ );
xor  ( new_n15030_, new_n15029_, new_n2121_ );
or   ( new_n15031_, new_n2122_, new_n7373_ );
or   ( new_n15032_, new_n2124_, new_n7149_ );
and  ( new_n15033_, new_n15032_, new_n15031_ );
xor  ( new_n15034_, new_n15033_, new_n1843_ );
or   ( new_n15035_, new_n15034_, new_n15030_ );
and  ( new_n15036_, new_n15034_, new_n15030_ );
or   ( new_n15037_, new_n1844_, new_n8115_ );
or   ( new_n15038_, new_n1846_, new_n8117_ );
and  ( new_n15039_, new_n15038_, new_n15037_ );
xor  ( new_n15040_, new_n15039_, new_n1586_ );
or   ( new_n15041_, new_n15040_, new_n15036_ );
and  ( new_n15042_, new_n15041_, new_n15035_ );
or   ( new_n15043_, new_n15042_, new_n15026_ );
and  ( new_n15044_, new_n15042_, new_n15026_ );
or   ( new_n15045_, new_n1593_, new_n8481_ );
or   ( new_n15046_, new_n1595_, new_n8352_ );
and  ( new_n15047_, new_n15046_, new_n15045_ );
xor  ( new_n15048_, new_n15047_, new_n1358_ );
or   ( new_n15049_, new_n1364_, new_n9099_ );
or   ( new_n15050_, new_n1366_, new_n8995_ );
and  ( new_n15051_, new_n15050_, new_n15049_ );
xor  ( new_n15052_, new_n15051_, new_n1129_ );
nor  ( new_n15053_, new_n15052_, new_n15048_ );
and  ( new_n15054_, new_n15052_, new_n15048_ );
or   ( new_n15055_, new_n1135_, new_n9679_ );
or   ( new_n15056_, new_n1137_, new_n9681_ );
and  ( new_n15057_, new_n15056_, new_n15055_ );
xor  ( new_n15058_, new_n15057_, new_n896_ );
nor  ( new_n15059_, new_n15058_, new_n15054_ );
nor  ( new_n15060_, new_n15059_, new_n15053_ );
or   ( new_n15061_, new_n15060_, new_n15044_ );
and  ( new_n15062_, new_n15061_, new_n15043_ );
or   ( new_n15063_, new_n15062_, new_n15022_ );
and  ( new_n15064_, new_n15062_, new_n15022_ );
or   ( new_n15065_, new_n7732_, new_n2057_ );
or   ( new_n15066_, new_n7734_, new_n1899_ );
and  ( new_n15067_, new_n15066_, new_n15065_ );
xor  ( new_n15068_, new_n15067_, new_n7177_ );
or   ( new_n15069_, new_n7184_, new_n2291_ );
or   ( new_n15070_, new_n7186_, new_n2178_ );
and  ( new_n15071_, new_n15070_, new_n15069_ );
xor  ( new_n15072_, new_n15071_, new_n6638_ );
nor  ( new_n15073_, new_n15072_, new_n15068_ );
and  ( new_n15074_, new_n15072_, new_n15068_ );
or   ( new_n15075_, new_n6645_, new_n2646_ );
or   ( new_n15076_, new_n6647_, new_n2475_ );
and  ( new_n15077_, new_n15076_, new_n15075_ );
xor  ( new_n15078_, new_n15077_, new_n6166_ );
nor  ( new_n15079_, new_n15078_, new_n15074_ );
nor  ( new_n15080_, new_n15079_, new_n15073_ );
or   ( new_n15081_, new_n10059_, new_n986_ );
or   ( new_n15082_, new_n10061_, new_n886_ );
and  ( new_n15083_, new_n15082_, new_n15081_ );
xor  ( new_n15084_, new_n15083_, new_n9421_ );
and  ( new_n15085_, RIbb2d888_64, RIbb2d108_80 );
or   ( new_n15086_, RIbb2d888_64, new_n805_ );
and  ( new_n15087_, new_n15086_, RIbb2d900_63 );
or   ( new_n15088_, new_n15087_, new_n15085_ );
or   ( new_n15089_, new_n10770_, new_n775_ );
and  ( new_n15090_, new_n15089_, new_n15088_ );
nor  ( new_n15091_, new_n15090_, new_n15084_ );
and  ( new_n15092_, new_n15090_, new_n15084_ );
nor  ( new_n15093_, new_n15092_, new_n522_ );
nor  ( new_n15094_, new_n15093_, new_n15091_ );
or   ( new_n15095_, new_n9422_, new_n1213_ );
or   ( new_n15096_, new_n9424_, new_n1168_ );
and  ( new_n15097_, new_n15096_, new_n15095_ );
xor  ( new_n15098_, new_n15097_, new_n8873_ );
or   ( new_n15099_, new_n8874_, new_n1525_ );
or   ( new_n15100_, new_n8876_, new_n1318_ );
and  ( new_n15101_, new_n15100_, new_n15099_ );
xor  ( new_n15102_, new_n15101_, new_n8257_ );
nor  ( new_n15103_, new_n15102_, new_n15098_ );
and  ( new_n15104_, new_n15102_, new_n15098_ );
or   ( new_n15105_, new_n8264_, new_n1754_ );
or   ( new_n15106_, new_n8266_, new_n1523_ );
and  ( new_n15107_, new_n15106_, new_n15105_ );
xor  ( new_n15108_, new_n15107_, new_n7725_ );
nor  ( new_n15109_, new_n15108_, new_n15104_ );
nor  ( new_n15110_, new_n15109_, new_n15103_ );
and  ( new_n15111_, new_n15110_, new_n15094_ );
nor  ( new_n15112_, new_n15111_, new_n15080_ );
nor  ( new_n15113_, new_n15110_, new_n15094_ );
nor  ( new_n15114_, new_n15113_, new_n15112_ );
or   ( new_n15115_, new_n15114_, new_n15064_ );
and  ( new_n15116_, new_n15115_, new_n15063_ );
nand ( new_n15117_, new_n15116_, new_n14970_ );
nor  ( new_n15118_, new_n15116_, new_n14970_ );
xor  ( new_n15119_, new_n14743_, new_n14737_ );
xnor ( new_n15120_, new_n15119_, new_n14749_ );
xnor ( new_n15121_, new_n14777_, new_n14773_ );
xor  ( new_n15122_, new_n15121_, new_n14783_ );
or   ( new_n15123_, new_n15122_, new_n15120_ );
xnor ( new_n15124_, new_n14797_, new_n14793_ );
xor  ( new_n15125_, new_n15124_, new_n14803_ );
xnor ( new_n15126_, new_n14869_, new_n14865_ );
xor  ( new_n15127_, new_n15126_, new_n14875_ );
or   ( new_n15128_, new_n15127_, new_n15125_ );
and  ( new_n15129_, new_n15127_, new_n15125_ );
xor  ( new_n15130_, new_n14815_, new_n14811_ );
xnor ( new_n15131_, new_n15130_, new_n14821_ );
or   ( new_n15132_, new_n15131_, new_n15129_ );
and  ( new_n15133_, new_n15132_, new_n15128_ );
or   ( new_n15134_, new_n15133_, new_n15123_ );
and  ( new_n15135_, new_n15133_, new_n15123_ );
xnor ( new_n15136_, new_n14851_, new_n14847_ );
xor  ( new_n15137_, new_n15136_, new_n14857_ );
xnor ( new_n15138_, new_n14835_, new_n14831_ );
xor  ( new_n15139_, new_n15138_, new_n14841_ );
nor  ( new_n15140_, new_n15139_, new_n15137_ );
and  ( new_n15141_, new_n15139_, new_n15137_ );
xor  ( new_n15142_, new_n14759_, new_n14755_ );
xnor ( new_n15143_, new_n15142_, new_n14765_ );
nor  ( new_n15144_, new_n15143_, new_n15141_ );
nor  ( new_n15145_, new_n15144_, new_n15140_ );
or   ( new_n15146_, new_n15145_, new_n15135_ );
and  ( new_n15147_, new_n15146_, new_n15134_ );
or   ( new_n15148_, new_n15147_, new_n15118_ );
and  ( new_n15149_, new_n15148_, new_n15117_ );
nand ( new_n15150_, new_n15149_, new_n14961_ );
or   ( new_n15151_, new_n15149_, new_n14961_ );
xnor ( new_n15152_, new_n14727_, new_n14725_ );
xor  ( new_n15153_, new_n15152_, new_n14731_ );
xor  ( new_n15154_, new_n14708_, new_n14706_ );
xor  ( new_n15155_, new_n15154_, new_n14712_ );
nor  ( new_n15156_, new_n15155_, new_n15153_ );
and  ( new_n15157_, new_n15155_, new_n15153_ );
xnor ( new_n15158_, new_n14767_, new_n14751_ );
xor  ( new_n15159_, new_n15158_, new_n14785_ );
xnor ( new_n15160_, new_n14859_, new_n14843_ );
xor  ( new_n15161_, new_n15160_, new_n14877_ );
nor  ( new_n15162_, new_n15161_, new_n15159_ );
and  ( new_n15163_, new_n15161_, new_n15159_ );
xor  ( new_n15164_, new_n14805_, new_n14789_ );
xnor ( new_n15165_, new_n15164_, new_n14823_ );
nor  ( new_n15166_, new_n15165_, new_n15163_ );
nor  ( new_n15167_, new_n15166_, new_n15162_ );
nor  ( new_n15168_, new_n15167_, new_n15157_ );
nor  ( new_n15169_, new_n15168_, new_n15156_ );
nand ( new_n15170_, new_n15169_, new_n15151_ );
and  ( new_n15171_, new_n15170_, new_n15150_ );
and  ( new_n15172_, new_n15171_, new_n14959_ );
or   ( new_n15173_, new_n15171_, new_n14959_ );
xor  ( new_n15174_, new_n14935_, new_n14933_ );
xor  ( new_n15175_, new_n15174_, new_n14938_ );
and  ( new_n15176_, new_n15175_, new_n15173_ );
or   ( new_n15177_, new_n15176_, new_n15172_ );
xnor ( new_n15178_, new_n14660_, new_n14455_ );
xor  ( new_n15179_, new_n15178_, new_n14681_ );
nand ( new_n15180_, new_n15179_, new_n15177_ );
nor  ( new_n15181_, new_n15179_, new_n15177_ );
xor  ( new_n15182_, new_n14930_, new_n14928_ );
xor  ( new_n15183_, new_n15182_, new_n14941_ );
or   ( new_n15184_, new_n15183_, new_n15181_ );
and  ( new_n15185_, new_n15184_, new_n15180_ );
nor  ( new_n15186_, new_n15185_, new_n14954_ );
xor  ( new_n15187_, new_n15179_, new_n15177_ );
xor  ( new_n15188_, new_n15187_, new_n15183_ );
xor  ( new_n15189_, new_n14881_, new_n14733_ );
xnor ( new_n15190_, new_n15189_, new_n14912_ );
xor  ( new_n15191_, new_n15149_, new_n14961_ );
xnor ( new_n15192_, new_n15191_, new_n15169_ );
nand ( new_n15193_, new_n15192_, new_n15190_ );
xor  ( new_n15194_, new_n14716_, new_n14714_ );
xor  ( new_n15195_, new_n15194_, new_n14721_ );
xor  ( new_n15196_, new_n15116_, new_n14970_ );
xor  ( new_n15197_, new_n15196_, new_n15147_ );
xnor ( new_n15198_, new_n14825_, new_n14787_ );
xor  ( new_n15199_, new_n15198_, new_n14879_ );
or   ( new_n15200_, new_n15199_, new_n15197_ );
and  ( new_n15201_, new_n15199_, new_n15197_ );
xor  ( new_n15202_, new_n15155_, new_n15153_ );
xor  ( new_n15203_, new_n15202_, new_n15167_ );
or   ( new_n15204_, new_n15203_, new_n15201_ );
and  ( new_n15205_, new_n15204_, new_n15200_ );
or   ( new_n15206_, new_n15205_, new_n15195_ );
and  ( new_n15207_, new_n15205_, new_n15195_ );
xnor ( new_n15208_, new_n15002_, new_n14986_ );
xor  ( new_n15209_, new_n15208_, new_n15020_ );
xnor ( new_n15210_, new_n15042_, new_n15026_ );
xor  ( new_n15211_, new_n15210_, new_n15060_ );
nor  ( new_n15212_, new_n15211_, new_n15209_ );
nand ( new_n15213_, new_n15211_, new_n15209_ );
xnor ( new_n15214_, new_n15110_, new_n15094_ );
xnor ( new_n15215_, new_n15214_, new_n15080_ );
and  ( new_n15216_, new_n15215_, new_n15213_ );
or   ( new_n15217_, new_n15216_, new_n15212_ );
xnor ( new_n15218_, new_n15161_, new_n15159_ );
xor  ( new_n15219_, new_n15218_, new_n15165_ );
and  ( new_n15220_, new_n15219_, new_n15217_ );
nor  ( new_n15221_, new_n15219_, new_n15217_ );
xor  ( new_n15222_, new_n14965_, new_n14963_ );
xnor ( new_n15223_, new_n15222_, new_n14968_ );
nor  ( new_n15224_, new_n15223_, new_n15221_ );
or   ( new_n15225_, new_n15224_, new_n15220_ );
xnor ( new_n15226_, new_n14898_, new_n14888_ );
xor  ( new_n15227_, new_n15226_, new_n14910_ );
and  ( new_n15228_, new_n15227_, new_n15225_ );
nor  ( new_n15229_, new_n15227_, new_n15225_ );
not  ( new_n15230_, new_n15229_ );
and  ( new_n15231_, new_n660_, RIbb31578_128 );
or   ( new_n15232_, new_n15231_, new_n523_ );
nand ( new_n15233_, new_n15231_, new_n520_ );
and  ( new_n15234_, new_n15233_, new_n15232_ );
xnor ( new_n15235_, new_n15052_, new_n15048_ );
xor  ( new_n15236_, new_n15235_, new_n15058_ );
or   ( new_n15237_, new_n15236_, new_n15234_ );
and  ( new_n15238_, new_n15236_, new_n15234_ );
xor  ( new_n15239_, new_n15034_, new_n15030_ );
xnor ( new_n15240_, new_n15239_, new_n15040_ );
or   ( new_n15241_, new_n15240_, new_n15238_ );
and  ( new_n15242_, new_n15241_, new_n15237_ );
xnor ( new_n15243_, new_n15072_, new_n15068_ );
xor  ( new_n15244_, new_n15243_, new_n15078_ );
xnor ( new_n15245_, new_n15102_, new_n15098_ );
xor  ( new_n15246_, new_n15245_, new_n15108_ );
or   ( new_n15247_, new_n15246_, new_n15244_ );
and  ( new_n15248_, new_n15246_, new_n15244_ );
xor  ( new_n15249_, new_n15090_, new_n15084_ );
xor  ( new_n15250_, new_n15249_, new_n523_ );
or   ( new_n15251_, new_n15250_, new_n15248_ );
and  ( new_n15252_, new_n15251_, new_n15247_ );
nor  ( new_n15253_, new_n15252_, new_n15242_ );
and  ( new_n15254_, new_n15252_, new_n15242_ );
xnor ( new_n15255_, new_n14994_, new_n14990_ );
xor  ( new_n15256_, new_n15255_, new_n15000_ );
xnor ( new_n15257_, new_n14978_, new_n14974_ );
xor  ( new_n15258_, new_n15257_, new_n14984_ );
nor  ( new_n15259_, new_n15258_, new_n15256_ );
and  ( new_n15260_, new_n15258_, new_n15256_ );
xor  ( new_n15261_, new_n15012_, new_n15008_ );
xnor ( new_n15262_, new_n15261_, new_n15018_ );
nor  ( new_n15263_, new_n15262_, new_n15260_ );
nor  ( new_n15264_, new_n15263_, new_n15259_ );
nor  ( new_n15265_, new_n15264_, new_n15254_ );
or   ( new_n15266_, new_n15265_, new_n15253_ );
or   ( new_n15267_, new_n3117_, new_n6219_ );
or   ( new_n15268_, new_n3119_, new_n5899_ );
and  ( new_n15269_, new_n15268_, new_n15267_ );
xor  ( new_n15270_, new_n15269_, new_n2800_ );
or   ( new_n15271_, new_n2807_, new_n6589_ );
or   ( new_n15272_, new_n2809_, new_n6425_ );
and  ( new_n15273_, new_n15272_, new_n15271_ );
xor  ( new_n15274_, new_n15273_, new_n2424_ );
or   ( new_n15275_, new_n15274_, new_n15270_ );
and  ( new_n15276_, new_n15274_, new_n15270_ );
or   ( new_n15277_, new_n2425_, new_n7149_ );
or   ( new_n15278_, new_n2427_, new_n6943_ );
and  ( new_n15279_, new_n15278_, new_n15277_ );
xor  ( new_n15280_, new_n15279_, new_n2121_ );
or   ( new_n15281_, new_n15280_, new_n15276_ );
and  ( new_n15282_, new_n15281_, new_n15275_ );
or   ( new_n15283_, new_n4302_, new_n4995_ );
or   ( new_n15284_, new_n4304_, new_n4603_ );
and  ( new_n15285_, new_n15284_, new_n15283_ );
xor  ( new_n15286_, new_n15285_, new_n3895_ );
or   ( new_n15287_, new_n3896_, new_n5171_ );
or   ( new_n15288_, new_n3898_, new_n4859_ );
and  ( new_n15289_, new_n15288_, new_n15287_ );
xor  ( new_n15290_, new_n15289_, new_n3460_ );
or   ( new_n15291_, new_n15290_, new_n15286_ );
and  ( new_n15292_, new_n15290_, new_n15286_ );
or   ( new_n15293_, new_n3461_, new_n5570_ );
or   ( new_n15294_, new_n3463_, new_n5428_ );
and  ( new_n15295_, new_n15294_, new_n15293_ );
xor  ( new_n15296_, new_n15295_, new_n3116_ );
or   ( new_n15297_, new_n15296_, new_n15292_ );
and  ( new_n15298_, new_n15297_, new_n15291_ );
or   ( new_n15299_, new_n15298_, new_n15282_ );
and  ( new_n15300_, new_n15298_, new_n15282_ );
or   ( new_n15301_, new_n5604_, new_n3696_ );
or   ( new_n15302_, new_n5606_, new_n3306_ );
and  ( new_n15303_, new_n15302_, new_n15301_ );
xor  ( new_n15304_, new_n15303_, new_n5206_ );
or   ( new_n15305_, new_n5207_, new_n3820_ );
or   ( new_n15306_, new_n5209_, new_n3694_ );
and  ( new_n15307_, new_n15306_, new_n15305_ );
xor  ( new_n15308_, new_n15307_, new_n4708_ );
nor  ( new_n15309_, new_n15308_, new_n15304_ );
and  ( new_n15310_, new_n15308_, new_n15304_ );
or   ( new_n15311_, new_n4709_, new_n4267_ );
or   ( new_n15312_, new_n4711_, new_n4069_ );
and  ( new_n15313_, new_n15312_, new_n15311_ );
xor  ( new_n15314_, new_n15313_, new_n4295_ );
nor  ( new_n15315_, new_n15314_, new_n15310_ );
nor  ( new_n15316_, new_n15315_, new_n15309_ );
or   ( new_n15317_, new_n15316_, new_n15300_ );
and  ( new_n15318_, new_n15317_, new_n15299_ );
or   ( new_n15319_, new_n897_, new_n10541_ );
or   ( new_n15320_, new_n899_, new_n10220_ );
and  ( new_n15321_, new_n15320_, new_n15319_ );
xor  ( new_n15322_, new_n15321_, new_n748_ );
or   ( new_n15323_, new_n2122_, new_n8117_ );
or   ( new_n15324_, new_n2124_, new_n7373_ );
and  ( new_n15325_, new_n15324_, new_n15323_ );
xor  ( new_n15326_, new_n15325_, new_n1843_ );
or   ( new_n15327_, new_n1844_, new_n8352_ );
or   ( new_n15328_, new_n1846_, new_n8115_ );
and  ( new_n15329_, new_n15328_, new_n15327_ );
xor  ( new_n15330_, new_n15329_, new_n1586_ );
or   ( new_n15331_, new_n15330_, new_n15326_ );
and  ( new_n15332_, new_n15330_, new_n15326_ );
or   ( new_n15333_, new_n1593_, new_n8995_ );
or   ( new_n15334_, new_n1595_, new_n8481_ );
and  ( new_n15335_, new_n15334_, new_n15333_ );
xor  ( new_n15336_, new_n15335_, new_n1358_ );
or   ( new_n15337_, new_n15336_, new_n15332_ );
and  ( new_n15338_, new_n15337_, new_n15331_ );
or   ( new_n15339_, new_n15338_, new_n15322_ );
and  ( new_n15340_, new_n15338_, new_n15322_ );
or   ( new_n15341_, new_n1364_, new_n9681_ );
or   ( new_n15342_, new_n1366_, new_n9099_ );
and  ( new_n15343_, new_n15342_, new_n15341_ );
xor  ( new_n15344_, new_n15343_, new_n1129_ );
or   ( new_n15345_, new_n1135_, new_n10220_ );
or   ( new_n15346_, new_n1137_, new_n9679_ );
and  ( new_n15347_, new_n15346_, new_n15345_ );
xor  ( new_n15348_, new_n15347_, new_n896_ );
nor  ( new_n15349_, new_n15348_, new_n15344_ );
and  ( new_n15350_, new_n15348_, new_n15344_ );
or   ( new_n15351_, new_n897_, new_n10841_ );
or   ( new_n15352_, new_n899_, new_n10541_ );
and  ( new_n15353_, new_n15352_, new_n15351_ );
xor  ( new_n15354_, new_n15353_, new_n748_ );
nor  ( new_n15355_, new_n15354_, new_n15350_ );
nor  ( new_n15356_, new_n15355_, new_n15349_ );
or   ( new_n15357_, new_n15356_, new_n15340_ );
and  ( new_n15358_, new_n15357_, new_n15339_ );
or   ( new_n15359_, new_n15358_, new_n15318_ );
and  ( new_n15360_, new_n15358_, new_n15318_ );
or   ( new_n15361_, new_n8874_, new_n1523_ );
or   ( new_n15362_, new_n8876_, new_n1525_ );
and  ( new_n15363_, new_n15362_, new_n15361_ );
xor  ( new_n15364_, new_n15363_, new_n8257_ );
or   ( new_n15365_, new_n8264_, new_n1899_ );
or   ( new_n15366_, new_n8266_, new_n1754_ );
and  ( new_n15367_, new_n15366_, new_n15365_ );
xor  ( new_n15368_, new_n15367_, new_n7725_ );
or   ( new_n15369_, new_n15368_, new_n15364_ );
and  ( new_n15370_, new_n15368_, new_n15364_ );
or   ( new_n15371_, new_n7732_, new_n2178_ );
or   ( new_n15372_, new_n7734_, new_n2057_ );
and  ( new_n15373_, new_n15372_, new_n15371_ );
xor  ( new_n15374_, new_n15373_, new_n7177_ );
or   ( new_n15375_, new_n15374_, new_n15370_ );
and  ( new_n15376_, new_n15375_, new_n15369_ );
or   ( new_n15377_, new_n10059_, new_n1168_ );
or   ( new_n15378_, new_n10061_, new_n986_ );
and  ( new_n15379_, new_n15378_, new_n15377_ );
xor  ( new_n15380_, new_n15379_, new_n9421_ );
and  ( new_n15381_, RIbb2d888_64, RIbb2d090_81 );
or   ( new_n15382_, RIbb2d888_64, new_n886_ );
and  ( new_n15383_, new_n15382_, RIbb2d900_63 );
or   ( new_n15384_, new_n15383_, new_n15381_ );
or   ( new_n15385_, new_n10770_, new_n805_ );
and  ( new_n15386_, new_n15385_, new_n15384_ );
or   ( new_n15387_, new_n15386_, new_n15380_ );
and  ( new_n15388_, new_n15386_, new_n15380_ );
or   ( new_n15389_, new_n9422_, new_n1318_ );
or   ( new_n15390_, new_n9424_, new_n1213_ );
and  ( new_n15391_, new_n15390_, new_n15389_ );
xor  ( new_n15392_, new_n15391_, new_n8873_ );
or   ( new_n15393_, new_n15392_, new_n15388_ );
and  ( new_n15394_, new_n15393_, new_n15387_ );
nor  ( new_n15395_, new_n15394_, new_n15376_ );
and  ( new_n15396_, new_n15394_, new_n15376_ );
or   ( new_n15397_, new_n7184_, new_n2475_ );
or   ( new_n15398_, new_n7186_, new_n2291_ );
and  ( new_n15399_, new_n15398_, new_n15397_ );
xor  ( new_n15400_, new_n15399_, new_n6638_ );
or   ( new_n15401_, new_n6645_, new_n2751_ );
or   ( new_n15402_, new_n6647_, new_n2646_ );
and  ( new_n15403_, new_n15402_, new_n15401_ );
xor  ( new_n15404_, new_n15403_, new_n6166_ );
nor  ( new_n15405_, new_n15404_, new_n15400_ );
and  ( new_n15406_, new_n15404_, new_n15400_ );
or   ( new_n15407_, new_n6173_, new_n3178_ );
or   ( new_n15408_, new_n6175_, new_n2981_ );
and  ( new_n15409_, new_n15408_, new_n15407_ );
xor  ( new_n15410_, new_n15409_, new_n5597_ );
nor  ( new_n15411_, new_n15410_, new_n15406_ );
nor  ( new_n15412_, new_n15411_, new_n15405_ );
nor  ( new_n15413_, new_n15412_, new_n15396_ );
nor  ( new_n15414_, new_n15413_, new_n15395_ );
or   ( new_n15415_, new_n15414_, new_n15360_ );
and  ( new_n15416_, new_n15415_, new_n15359_ );
nor  ( new_n15417_, new_n15416_, new_n15266_ );
and  ( new_n15418_, new_n15416_, new_n15266_ );
xnor ( new_n15419_, new_n15127_, new_n15125_ );
xor  ( new_n15420_, new_n15419_, new_n15131_ );
xnor ( new_n15421_, new_n15139_, new_n15137_ );
xor  ( new_n15422_, new_n15421_, new_n15143_ );
nor  ( new_n15423_, new_n15422_, new_n15420_ );
and  ( new_n15424_, new_n15422_, new_n15420_ );
xor  ( new_n15425_, new_n15122_, new_n15120_ );
nor  ( new_n15426_, new_n15425_, new_n15424_ );
nor  ( new_n15427_, new_n15426_, new_n15423_ );
nor  ( new_n15428_, new_n15427_, new_n15418_ );
nor  ( new_n15429_, new_n15428_, new_n15417_ );
and  ( new_n15430_, new_n15429_, new_n15230_ );
nor  ( new_n15431_, new_n15430_, new_n15228_ );
or   ( new_n15432_, new_n15431_, new_n15207_ );
and  ( new_n15433_, new_n15432_, new_n15206_ );
or   ( new_n15434_, new_n15433_, new_n15193_ );
and  ( new_n15435_, new_n15433_, new_n15193_ );
xnor ( new_n15436_, new_n15171_, new_n14959_ );
xor  ( new_n15437_, new_n15436_, new_n15175_ );
or   ( new_n15438_, new_n15437_, new_n15435_ );
and  ( new_n15439_, new_n15438_, new_n15434_ );
nor  ( new_n15440_, new_n15439_, new_n15188_ );
xor  ( new_n15441_, new_n15433_, new_n15193_ );
xor  ( new_n15442_, new_n15441_, new_n15437_ );
xor  ( new_n15443_, new_n15199_, new_n15197_ );
xor  ( new_n15444_, new_n15443_, new_n15203_ );
xnor ( new_n15445_, new_n15416_, new_n15266_ );
xor  ( new_n15446_, new_n15445_, new_n15427_ );
xnor ( new_n15447_, new_n15062_, new_n15022_ );
xor  ( new_n15448_, new_n15447_, new_n15114_ );
or   ( new_n15449_, new_n15448_, new_n15446_ );
and  ( new_n15450_, new_n15448_, new_n15446_ );
xor  ( new_n15451_, new_n15219_, new_n15217_ );
xor  ( new_n15452_, new_n15451_, new_n15223_ );
or   ( new_n15453_, new_n15452_, new_n15450_ );
and  ( new_n15454_, new_n15453_, new_n15449_ );
nor  ( new_n15455_, new_n15454_, new_n15444_ );
and  ( new_n15456_, new_n15454_, new_n15444_ );
xor  ( new_n15457_, new_n15252_, new_n15242_ );
xor  ( new_n15458_, new_n15457_, new_n15264_ );
xnor ( new_n15459_, new_n15211_, new_n15209_ );
xor  ( new_n15460_, new_n15459_, new_n15215_ );
nor  ( new_n15461_, new_n15460_, new_n15458_ );
and  ( new_n15462_, new_n15460_, new_n15458_ );
xor  ( new_n15463_, new_n15422_, new_n15420_ );
xnor ( new_n15464_, new_n15463_, new_n15425_ );
nor  ( new_n15465_, new_n15464_, new_n15462_ );
or   ( new_n15466_, new_n15465_, new_n15461_ );
xnor ( new_n15467_, new_n15133_, new_n15123_ );
xor  ( new_n15468_, new_n15467_, new_n15145_ );
and  ( new_n15469_, new_n15468_, new_n15466_ );
nor  ( new_n15470_, new_n15468_, new_n15466_ );
xor  ( new_n15471_, new_n15258_, new_n15256_ );
xor  ( new_n15472_, new_n15471_, new_n15262_ );
xnor ( new_n15473_, new_n15338_, new_n15322_ );
xor  ( new_n15474_, new_n15473_, new_n15356_ );
or   ( new_n15475_, new_n15474_, new_n15472_ );
nand ( new_n15476_, new_n15474_, new_n15472_ );
xor  ( new_n15477_, new_n15236_, new_n15234_ );
xnor ( new_n15478_, new_n15477_, new_n15240_ );
nand ( new_n15479_, new_n15478_, new_n15476_ );
and  ( new_n15480_, new_n15479_, new_n15475_ );
xor  ( new_n15481_, new_n15246_, new_n15244_ );
xor  ( new_n15482_, new_n15481_, new_n15250_ );
xnor ( new_n15483_, new_n15368_, new_n15364_ );
xor  ( new_n15484_, new_n15483_, new_n15374_ );
xnor ( new_n15485_, new_n15308_, new_n15304_ );
xor  ( new_n15486_, new_n15485_, new_n15314_ );
or   ( new_n15487_, new_n15486_, new_n15484_ );
and  ( new_n15488_, new_n15486_, new_n15484_ );
xor  ( new_n15489_, new_n15404_, new_n15400_ );
xnor ( new_n15490_, new_n15489_, new_n15410_ );
or   ( new_n15491_, new_n15490_, new_n15488_ );
and  ( new_n15492_, new_n15491_, new_n15487_ );
or   ( new_n15493_, new_n15492_, new_n15482_ );
and  ( new_n15494_, new_n15492_, new_n15482_ );
xnor ( new_n15495_, new_n15330_, new_n15326_ );
xor  ( new_n15496_, new_n15495_, new_n15336_ );
xnor ( new_n15497_, new_n15290_, new_n15286_ );
xor  ( new_n15498_, new_n15497_, new_n15296_ );
nor  ( new_n15499_, new_n15498_, new_n15496_ );
and  ( new_n15500_, new_n15498_, new_n15496_ );
xor  ( new_n15501_, new_n15274_, new_n15270_ );
xnor ( new_n15502_, new_n15501_, new_n15280_ );
nor  ( new_n15503_, new_n15502_, new_n15500_ );
nor  ( new_n15504_, new_n15503_, new_n15499_ );
or   ( new_n15505_, new_n15504_, new_n15494_ );
and  ( new_n15506_, new_n15505_, new_n15493_ );
nor  ( new_n15507_, new_n15506_, new_n15480_ );
and  ( new_n15508_, new_n15506_, new_n15480_ );
or   ( new_n15509_, new_n4709_, new_n4603_ );
or   ( new_n15510_, new_n4711_, new_n4267_ );
and  ( new_n15511_, new_n15510_, new_n15509_ );
xor  ( new_n15512_, new_n15511_, new_n4295_ );
or   ( new_n15513_, new_n4302_, new_n4859_ );
or   ( new_n15514_, new_n4304_, new_n4995_ );
and  ( new_n15515_, new_n15514_, new_n15513_ );
xor  ( new_n15516_, new_n15515_, new_n3895_ );
or   ( new_n15517_, new_n15516_, new_n15512_ );
and  ( new_n15518_, new_n15516_, new_n15512_ );
or   ( new_n15519_, new_n3896_, new_n5428_ );
or   ( new_n15520_, new_n3898_, new_n5171_ );
and  ( new_n15521_, new_n15520_, new_n15519_ );
xor  ( new_n15522_, new_n15521_, new_n3460_ );
or   ( new_n15523_, new_n15522_, new_n15518_ );
and  ( new_n15524_, new_n15523_, new_n15517_ );
or   ( new_n15525_, new_n3461_, new_n5899_ );
or   ( new_n15526_, new_n3463_, new_n5570_ );
and  ( new_n15527_, new_n15526_, new_n15525_ );
xor  ( new_n15528_, new_n15527_, new_n3116_ );
or   ( new_n15529_, new_n3117_, new_n6425_ );
or   ( new_n15530_, new_n3119_, new_n6219_ );
and  ( new_n15531_, new_n15530_, new_n15529_ );
xor  ( new_n15532_, new_n15531_, new_n2800_ );
or   ( new_n15533_, new_n15532_, new_n15528_ );
and  ( new_n15534_, new_n15532_, new_n15528_ );
or   ( new_n15535_, new_n2807_, new_n6943_ );
or   ( new_n15536_, new_n2809_, new_n6589_ );
and  ( new_n15537_, new_n15536_, new_n15535_ );
xor  ( new_n15538_, new_n15537_, new_n2424_ );
or   ( new_n15539_, new_n15538_, new_n15534_ );
and  ( new_n15540_, new_n15539_, new_n15533_ );
or   ( new_n15541_, new_n15540_, new_n15524_ );
and  ( new_n15542_, new_n15540_, new_n15524_ );
or   ( new_n15543_, new_n6173_, new_n3306_ );
or   ( new_n15544_, new_n6175_, new_n3178_ );
and  ( new_n15545_, new_n15544_, new_n15543_ );
xor  ( new_n15546_, new_n15545_, new_n5597_ );
or   ( new_n15547_, new_n5604_, new_n3694_ );
or   ( new_n15548_, new_n5606_, new_n3696_ );
and  ( new_n15549_, new_n15548_, new_n15547_ );
xor  ( new_n15550_, new_n15549_, new_n5206_ );
or   ( new_n15551_, new_n15550_, new_n15546_ );
and  ( new_n15552_, new_n15550_, new_n15546_ );
or   ( new_n15553_, new_n5207_, new_n4069_ );
or   ( new_n15554_, new_n5209_, new_n3820_ );
and  ( new_n15555_, new_n15554_, new_n15553_ );
xor  ( new_n15556_, new_n15555_, new_n4708_ );
or   ( new_n15557_, new_n15556_, new_n15552_ );
and  ( new_n15558_, new_n15557_, new_n15551_ );
or   ( new_n15559_, new_n15558_, new_n15542_ );
and  ( new_n15560_, new_n15559_, new_n15541_ );
xor  ( new_n15561_, new_n15348_, new_n15344_ );
xor  ( new_n15562_, new_n15561_, new_n15354_ );
or   ( new_n15563_, new_n2425_, new_n7373_ );
or   ( new_n15564_, new_n2427_, new_n7149_ );
and  ( new_n15565_, new_n15564_, new_n15563_ );
xor  ( new_n15566_, new_n15565_, new_n2121_ );
or   ( new_n15567_, new_n2122_, new_n8115_ );
or   ( new_n15568_, new_n2124_, new_n8117_ );
and  ( new_n15569_, new_n15568_, new_n15567_ );
xor  ( new_n15570_, new_n15569_, new_n1843_ );
or   ( new_n15571_, new_n15570_, new_n15566_ );
and  ( new_n15572_, new_n15570_, new_n15566_ );
or   ( new_n15573_, new_n1844_, new_n8481_ );
or   ( new_n15574_, new_n1846_, new_n8352_ );
and  ( new_n15575_, new_n15574_, new_n15573_ );
xor  ( new_n15576_, new_n15575_, new_n1586_ );
or   ( new_n15577_, new_n15576_, new_n15572_ );
and  ( new_n15578_, new_n15577_, new_n15571_ );
or   ( new_n15579_, new_n15578_, new_n15562_ );
and  ( new_n15580_, new_n15578_, new_n15562_ );
or   ( new_n15581_, new_n1593_, new_n9099_ );
or   ( new_n15582_, new_n1595_, new_n8995_ );
and  ( new_n15583_, new_n15582_, new_n15581_ );
xor  ( new_n15584_, new_n15583_, new_n1358_ );
or   ( new_n15585_, new_n1364_, new_n9679_ );
or   ( new_n15586_, new_n1366_, new_n9681_ );
and  ( new_n15587_, new_n15586_, new_n15585_ );
xor  ( new_n15588_, new_n15587_, new_n1129_ );
nor  ( new_n15589_, new_n15588_, new_n15584_ );
and  ( new_n15590_, new_n15588_, new_n15584_ );
or   ( new_n15591_, new_n1135_, new_n10541_ );
or   ( new_n15592_, new_n1137_, new_n10220_ );
and  ( new_n15593_, new_n15592_, new_n15591_ );
xor  ( new_n15594_, new_n15593_, new_n896_ );
nor  ( new_n15595_, new_n15594_, new_n15590_ );
nor  ( new_n15596_, new_n15595_, new_n15589_ );
or   ( new_n15597_, new_n15596_, new_n15580_ );
and  ( new_n15598_, new_n15597_, new_n15579_ );
nor  ( new_n15599_, new_n15598_, new_n15560_ );
and  ( new_n15600_, new_n15598_, new_n15560_ );
or   ( new_n15601_, new_n9422_, new_n1525_ );
or   ( new_n15602_, new_n9424_, new_n1318_ );
and  ( new_n15603_, new_n15602_, new_n15601_ );
xor  ( new_n15604_, new_n15603_, new_n8873_ );
or   ( new_n15605_, new_n8874_, new_n1754_ );
or   ( new_n15606_, new_n8876_, new_n1523_ );
and  ( new_n15607_, new_n15606_, new_n15605_ );
xor  ( new_n15608_, new_n15607_, new_n8257_ );
nor  ( new_n15609_, new_n15608_, new_n15604_ );
and  ( new_n15610_, new_n15608_, new_n15604_ );
or   ( new_n15611_, new_n8264_, new_n2057_ );
or   ( new_n15612_, new_n8266_, new_n1899_ );
and  ( new_n15613_, new_n15612_, new_n15611_ );
xor  ( new_n15614_, new_n15613_, new_n7725_ );
nor  ( new_n15615_, new_n15614_, new_n15610_ );
nor  ( new_n15616_, new_n15615_, new_n15609_ );
or   ( new_n15617_, new_n10059_, new_n1213_ );
or   ( new_n15618_, new_n10061_, new_n1168_ );
and  ( new_n15619_, new_n15618_, new_n15617_ );
xor  ( new_n15620_, new_n15619_, new_n9421_ );
and  ( new_n15621_, RIbb2d888_64, RIbb2d018_82 );
or   ( new_n15622_, RIbb2d888_64, new_n986_ );
and  ( new_n15623_, new_n15622_, RIbb2d900_63 );
or   ( new_n15624_, new_n15623_, new_n15621_ );
or   ( new_n15625_, new_n10770_, new_n886_ );
and  ( new_n15626_, new_n15625_, new_n15624_ );
nor  ( new_n15627_, new_n15626_, new_n15620_ );
and  ( new_n15628_, new_n15626_, new_n15620_ );
nor  ( new_n15629_, new_n15628_, new_n747_ );
nor  ( new_n15630_, new_n15629_, new_n15627_ );
or   ( new_n15631_, new_n7732_, new_n2291_ );
or   ( new_n15632_, new_n7734_, new_n2178_ );
and  ( new_n15633_, new_n15632_, new_n15631_ );
xor  ( new_n15634_, new_n15633_, new_n7177_ );
or   ( new_n15635_, new_n7184_, new_n2646_ );
or   ( new_n15636_, new_n7186_, new_n2475_ );
and  ( new_n15637_, new_n15636_, new_n15635_ );
xor  ( new_n15638_, new_n15637_, new_n6638_ );
nor  ( new_n15639_, new_n15638_, new_n15634_ );
and  ( new_n15640_, new_n15638_, new_n15634_ );
or   ( new_n15641_, new_n6645_, new_n2981_ );
or   ( new_n15642_, new_n6647_, new_n2751_ );
and  ( new_n15643_, new_n15642_, new_n15641_ );
xor  ( new_n15644_, new_n15643_, new_n6166_ );
nor  ( new_n15645_, new_n15644_, new_n15640_ );
nor  ( new_n15646_, new_n15645_, new_n15639_ );
and  ( new_n15647_, new_n15646_, new_n15630_ );
nor  ( new_n15648_, new_n15647_, new_n15616_ );
nor  ( new_n15649_, new_n15646_, new_n15630_ );
nor  ( new_n15650_, new_n15649_, new_n15648_ );
nor  ( new_n15651_, new_n15650_, new_n15600_ );
nor  ( new_n15652_, new_n15651_, new_n15599_ );
not  ( new_n15653_, new_n15652_ );
nor  ( new_n15654_, new_n15653_, new_n15508_ );
nor  ( new_n15655_, new_n15654_, new_n15507_ );
nor  ( new_n15656_, new_n15655_, new_n15470_ );
nor  ( new_n15657_, new_n15656_, new_n15469_ );
nor  ( new_n15658_, new_n15657_, new_n15456_ );
or   ( new_n15659_, new_n15658_, new_n15455_ );
xnor ( new_n15660_, new_n15205_, new_n15195_ );
xor  ( new_n15661_, new_n15660_, new_n15431_ );
nand ( new_n15662_, new_n15661_, new_n15659_ );
nor  ( new_n15663_, new_n15661_, new_n15659_ );
xnor ( new_n15664_, new_n15192_, new_n15190_ );
or   ( new_n15665_, new_n15664_, new_n15663_ );
and  ( new_n15666_, new_n15665_, new_n15662_ );
nor  ( new_n15667_, new_n15666_, new_n15442_ );
xor  ( new_n15668_, new_n15661_, new_n15659_ );
xor  ( new_n15669_, new_n15668_, new_n15664_ );
xor  ( new_n15670_, new_n15448_, new_n15446_ );
xor  ( new_n15671_, new_n15670_, new_n15452_ );
xnor ( new_n15672_, new_n15358_, new_n15318_ );
xor  ( new_n15673_, new_n15672_, new_n15414_ );
xor  ( new_n15674_, new_n15506_, new_n15480_ );
xor  ( new_n15675_, new_n15674_, new_n15653_ );
or   ( new_n15676_, new_n15675_, new_n15673_ );
and  ( new_n15677_, new_n15675_, new_n15673_ );
xor  ( new_n15678_, new_n15460_, new_n15458_ );
xor  ( new_n15679_, new_n15678_, new_n15464_ );
or   ( new_n15680_, new_n15679_, new_n15677_ );
and  ( new_n15681_, new_n15680_, new_n15676_ );
nor  ( new_n15682_, new_n15681_, new_n15671_ );
nand ( new_n15683_, new_n15681_, new_n15671_ );
xor  ( new_n15684_, new_n15492_, new_n15482_ );
xnor ( new_n15685_, new_n15684_, new_n15504_ );
not  ( new_n15686_, new_n15685_ );
xnor ( new_n15687_, new_n15598_, new_n15560_ );
xor  ( new_n15688_, new_n15687_, new_n15650_ );
or   ( new_n15689_, new_n15688_, new_n15686_ );
xnor ( new_n15690_, new_n15386_, new_n15380_ );
xor  ( new_n15691_, new_n15690_, new_n15392_ );
xnor ( new_n15692_, new_n15608_, new_n15604_ );
xor  ( new_n15693_, new_n15692_, new_n15614_ );
xnor ( new_n15694_, new_n15550_, new_n15546_ );
xor  ( new_n15695_, new_n15694_, new_n15556_ );
or   ( new_n15696_, new_n15695_, new_n15693_ );
and  ( new_n15697_, new_n15695_, new_n15693_ );
xor  ( new_n15698_, new_n15638_, new_n15634_ );
xnor ( new_n15699_, new_n15698_, new_n15644_ );
or   ( new_n15700_, new_n15699_, new_n15697_ );
and  ( new_n15701_, new_n15700_, new_n15696_ );
nor  ( new_n15702_, new_n15701_, new_n15691_ );
and  ( new_n15703_, new_n15701_, new_n15691_ );
xnor ( new_n15704_, new_n15532_, new_n15528_ );
xor  ( new_n15705_, new_n15704_, new_n15538_ );
xnor ( new_n15706_, new_n15570_, new_n15566_ );
xor  ( new_n15707_, new_n15706_, new_n15576_ );
nor  ( new_n15708_, new_n15707_, new_n15705_ );
and  ( new_n15709_, new_n15707_, new_n15705_ );
xor  ( new_n15710_, new_n15516_, new_n15512_ );
xnor ( new_n15711_, new_n15710_, new_n15522_ );
nor  ( new_n15712_, new_n15711_, new_n15709_ );
nor  ( new_n15713_, new_n15712_, new_n15708_ );
nor  ( new_n15714_, new_n15713_, new_n15703_ );
nor  ( new_n15715_, new_n15714_, new_n15702_ );
or   ( new_n15716_, new_n7184_, new_n2751_ );
or   ( new_n15717_, new_n7186_, new_n2646_ );
and  ( new_n15718_, new_n15717_, new_n15716_ );
xor  ( new_n15719_, new_n15718_, new_n6638_ );
or   ( new_n15720_, new_n6645_, new_n3178_ );
or   ( new_n15721_, new_n6647_, new_n2981_ );
and  ( new_n15722_, new_n15721_, new_n15720_ );
xor  ( new_n15723_, new_n15722_, new_n6166_ );
or   ( new_n15724_, new_n15723_, new_n15719_ );
and  ( new_n15725_, new_n15723_, new_n15719_ );
or   ( new_n15726_, new_n6173_, new_n3696_ );
or   ( new_n15727_, new_n6175_, new_n3306_ );
and  ( new_n15728_, new_n15727_, new_n15726_ );
xor  ( new_n15729_, new_n15728_, new_n5597_ );
or   ( new_n15730_, new_n15729_, new_n15725_ );
and  ( new_n15731_, new_n15730_, new_n15724_ );
or   ( new_n15732_, new_n8874_, new_n1899_ );
or   ( new_n15733_, new_n8876_, new_n1754_ );
and  ( new_n15734_, new_n15733_, new_n15732_ );
xor  ( new_n15735_, new_n15734_, new_n8257_ );
or   ( new_n15736_, new_n8264_, new_n2178_ );
or   ( new_n15737_, new_n8266_, new_n2057_ );
and  ( new_n15738_, new_n15737_, new_n15736_ );
xor  ( new_n15739_, new_n15738_, new_n7725_ );
or   ( new_n15740_, new_n15739_, new_n15735_ );
and  ( new_n15741_, new_n15739_, new_n15735_ );
or   ( new_n15742_, new_n7732_, new_n2475_ );
or   ( new_n15743_, new_n7734_, new_n2291_ );
and  ( new_n15744_, new_n15743_, new_n15742_ );
xor  ( new_n15745_, new_n15744_, new_n7177_ );
or   ( new_n15746_, new_n15745_, new_n15741_ );
and  ( new_n15747_, new_n15746_, new_n15740_ );
nor  ( new_n15748_, new_n15747_, new_n15731_ );
and  ( new_n15749_, new_n15747_, new_n15731_ );
or   ( new_n15750_, new_n10059_, new_n1318_ );
or   ( new_n15751_, new_n10061_, new_n1213_ );
and  ( new_n15752_, new_n15751_, new_n15750_ );
xor  ( new_n15753_, new_n15752_, new_n9421_ );
and  ( new_n15754_, RIbb2d888_64, RIbb2cfa0_83 );
or   ( new_n15755_, RIbb2d888_64, new_n1168_ );
and  ( new_n15756_, new_n15755_, RIbb2d900_63 );
or   ( new_n15757_, new_n15756_, new_n15754_ );
or   ( new_n15758_, new_n10770_, new_n986_ );
and  ( new_n15759_, new_n15758_, new_n15757_ );
nor  ( new_n15760_, new_n15759_, new_n15753_ );
and  ( new_n15761_, new_n15759_, new_n15753_ );
or   ( new_n15762_, new_n9422_, new_n1523_ );
or   ( new_n15763_, new_n9424_, new_n1525_ );
and  ( new_n15764_, new_n15763_, new_n15762_ );
xor  ( new_n15765_, new_n15764_, new_n8873_ );
nor  ( new_n15766_, new_n15765_, new_n15761_ );
nor  ( new_n15767_, new_n15766_, new_n15760_ );
nor  ( new_n15768_, new_n15767_, new_n15749_ );
nor  ( new_n15769_, new_n15768_, new_n15748_ );
or   ( new_n15770_, new_n4302_, new_n5171_ );
or   ( new_n15771_, new_n4304_, new_n4859_ );
and  ( new_n15772_, new_n15771_, new_n15770_ );
xor  ( new_n15773_, new_n15772_, new_n3895_ );
or   ( new_n15774_, new_n3896_, new_n5570_ );
or   ( new_n15775_, new_n3898_, new_n5428_ );
and  ( new_n15776_, new_n15775_, new_n15774_ );
xor  ( new_n15777_, new_n15776_, new_n3460_ );
or   ( new_n15778_, new_n15777_, new_n15773_ );
and  ( new_n15779_, new_n15777_, new_n15773_ );
or   ( new_n15780_, new_n3461_, new_n6219_ );
or   ( new_n15781_, new_n3463_, new_n5899_ );
and  ( new_n15782_, new_n15781_, new_n15780_ );
xor  ( new_n15783_, new_n15782_, new_n3116_ );
or   ( new_n15784_, new_n15783_, new_n15779_ );
and  ( new_n15785_, new_n15784_, new_n15778_ );
or   ( new_n15786_, new_n5604_, new_n3820_ );
or   ( new_n15787_, new_n5606_, new_n3694_ );
and  ( new_n15788_, new_n15787_, new_n15786_ );
xor  ( new_n15789_, new_n15788_, new_n5206_ );
or   ( new_n15790_, new_n5207_, new_n4267_ );
or   ( new_n15791_, new_n5209_, new_n4069_ );
and  ( new_n15792_, new_n15791_, new_n15790_ );
xor  ( new_n15793_, new_n15792_, new_n4708_ );
or   ( new_n15794_, new_n15793_, new_n15789_ );
and  ( new_n15795_, new_n15793_, new_n15789_ );
or   ( new_n15796_, new_n4709_, new_n4995_ );
or   ( new_n15797_, new_n4711_, new_n4603_ );
and  ( new_n15798_, new_n15797_, new_n15796_ );
xor  ( new_n15799_, new_n15798_, new_n4295_ );
or   ( new_n15800_, new_n15799_, new_n15795_ );
and  ( new_n15801_, new_n15800_, new_n15794_ );
nor  ( new_n15802_, new_n15801_, new_n15785_ );
and  ( new_n15803_, new_n15801_, new_n15785_ );
or   ( new_n15804_, new_n3117_, new_n6589_ );
or   ( new_n15805_, new_n3119_, new_n6425_ );
and  ( new_n15806_, new_n15805_, new_n15804_ );
xor  ( new_n15807_, new_n15806_, new_n2800_ );
or   ( new_n15808_, new_n2807_, new_n7149_ );
or   ( new_n15809_, new_n2809_, new_n6943_ );
and  ( new_n15810_, new_n15809_, new_n15808_ );
xor  ( new_n15811_, new_n15810_, new_n2424_ );
nor  ( new_n15812_, new_n15811_, new_n15807_ );
and  ( new_n15813_, new_n15811_, new_n15807_ );
or   ( new_n15814_, new_n2425_, new_n8117_ );
or   ( new_n15815_, new_n2427_, new_n7373_ );
and  ( new_n15816_, new_n15815_, new_n15814_ );
xor  ( new_n15817_, new_n15816_, new_n2121_ );
nor  ( new_n15818_, new_n15817_, new_n15813_ );
nor  ( new_n15819_, new_n15818_, new_n15812_ );
nor  ( new_n15820_, new_n15819_, new_n15803_ );
nor  ( new_n15821_, new_n15820_, new_n15802_ );
and  ( new_n15822_, new_n15821_, new_n15769_ );
nor  ( new_n15823_, new_n15821_, new_n15769_ );
and  ( new_n15824_, new_n820_, RIbb31578_128 );
or   ( new_n15825_, new_n15824_, new_n748_ );
nand ( new_n15826_, new_n15824_, new_n745_ );
and  ( new_n15827_, new_n15826_, new_n15825_ );
xnor ( new_n15828_, new_n15588_, new_n15584_ );
xor  ( new_n15829_, new_n15828_, new_n15594_ );
nor  ( new_n15830_, new_n15829_, new_n15827_ );
and  ( new_n15831_, new_n15829_, new_n15827_ );
not  ( new_n15832_, new_n15831_ );
or   ( new_n15833_, new_n2122_, new_n8352_ );
or   ( new_n15834_, new_n2124_, new_n8115_ );
and  ( new_n15835_, new_n15834_, new_n15833_ );
xor  ( new_n15836_, new_n15835_, new_n1843_ );
or   ( new_n15837_, new_n1844_, new_n8995_ );
or   ( new_n15838_, new_n1846_, new_n8481_ );
and  ( new_n15839_, new_n15838_, new_n15837_ );
xor  ( new_n15840_, new_n15839_, new_n1586_ );
nor  ( new_n15841_, new_n15840_, new_n15836_ );
and  ( new_n15842_, new_n15840_, new_n15836_ );
or   ( new_n15843_, new_n1593_, new_n9681_ );
or   ( new_n15844_, new_n1595_, new_n9099_ );
and  ( new_n15845_, new_n15844_, new_n15843_ );
xor  ( new_n15846_, new_n15845_, new_n1358_ );
nor  ( new_n15847_, new_n15846_, new_n15842_ );
nor  ( new_n15848_, new_n15847_, new_n15841_ );
and  ( new_n15849_, new_n15848_, new_n15832_ );
nor  ( new_n15850_, new_n15849_, new_n15830_ );
nor  ( new_n15851_, new_n15850_, new_n15823_ );
nor  ( new_n15852_, new_n15851_, new_n15822_ );
and  ( new_n15853_, new_n15852_, new_n15715_ );
xnor ( new_n15854_, new_n15498_, new_n15496_ );
xor  ( new_n15855_, new_n15854_, new_n15502_ );
xnor ( new_n15856_, new_n15486_, new_n15484_ );
xor  ( new_n15857_, new_n15856_, new_n15490_ );
and  ( new_n15858_, new_n15857_, new_n15855_ );
nor  ( new_n15859_, new_n15857_, new_n15855_ );
xor  ( new_n15860_, new_n15578_, new_n15562_ );
xnor ( new_n15861_, new_n15860_, new_n15596_ );
nor  ( new_n15862_, new_n15861_, new_n15859_ );
nor  ( new_n15863_, new_n15862_, new_n15858_ );
nor  ( new_n15864_, new_n15863_, new_n15853_ );
nor  ( new_n15865_, new_n15852_, new_n15715_ );
nor  ( new_n15866_, new_n15865_, new_n15864_ );
nor  ( new_n15867_, new_n15866_, new_n15689_ );
and  ( new_n15868_, new_n15866_, new_n15689_ );
xnor ( new_n15869_, new_n15394_, new_n15376_ );
xor  ( new_n15870_, new_n15869_, new_n15412_ );
xnor ( new_n15871_, new_n15298_, new_n15282_ );
xor  ( new_n15872_, new_n15871_, new_n15316_ );
nor  ( new_n15873_, new_n15872_, new_n15870_ );
and  ( new_n15874_, new_n15872_, new_n15870_ );
xor  ( new_n15875_, new_n15474_, new_n15472_ );
xor  ( new_n15876_, new_n15875_, new_n15478_ );
not  ( new_n15877_, new_n15876_ );
nor  ( new_n15878_, new_n15877_, new_n15874_ );
nor  ( new_n15879_, new_n15878_, new_n15873_ );
nor  ( new_n15880_, new_n15879_, new_n15868_ );
nor  ( new_n15881_, new_n15880_, new_n15867_ );
not  ( new_n15882_, new_n15881_ );
and  ( new_n15883_, new_n15882_, new_n15683_ );
or   ( new_n15884_, new_n15883_, new_n15682_ );
xor  ( new_n15885_, new_n15227_, new_n15225_ );
xor  ( new_n15886_, new_n15885_, new_n15429_ );
nand ( new_n15887_, new_n15886_, new_n15884_ );
nor  ( new_n15888_, new_n15886_, new_n15884_ );
xor  ( new_n15889_, new_n15454_, new_n15444_ );
xor  ( new_n15890_, new_n15889_, new_n15657_ );
or   ( new_n15891_, new_n15890_, new_n15888_ );
and  ( new_n15892_, new_n15891_, new_n15887_ );
nor  ( new_n15893_, new_n15892_, new_n15669_ );
xor  ( new_n15894_, new_n15886_, new_n15884_ );
xor  ( new_n15895_, new_n15894_, new_n15890_ );
xor  ( new_n15896_, new_n15675_, new_n15673_ );
xor  ( new_n15897_, new_n15896_, new_n15679_ );
xnor ( new_n15898_, new_n15852_, new_n15715_ );
and  ( new_n15899_, new_n15898_, new_n15863_ );
not  ( new_n15900_, new_n15865_ );
and  ( new_n15901_, new_n15900_, new_n15864_ );
or   ( new_n15902_, new_n15901_, new_n15899_ );
xor  ( new_n15903_, new_n15872_, new_n15870_ );
xor  ( new_n15904_, new_n15903_, new_n15877_ );
or   ( new_n15905_, new_n15904_, new_n15902_ );
nand ( new_n15906_, new_n15904_, new_n15902_ );
xor  ( new_n15907_, new_n15688_, new_n15686_ );
nand ( new_n15908_, new_n15907_, new_n15906_ );
and  ( new_n15909_, new_n15908_, new_n15905_ );
nor  ( new_n15910_, new_n15909_, new_n15897_ );
nand ( new_n15911_, new_n15909_, new_n15897_ );
xnor ( new_n15912_, new_n15821_, new_n15769_ );
xor  ( new_n15913_, new_n15912_, new_n15850_ );
xnor ( new_n15914_, new_n15701_, new_n15691_ );
xor  ( new_n15915_, new_n15914_, new_n15713_ );
nand ( new_n15916_, new_n15915_, new_n15913_ );
or   ( new_n15917_, new_n10059_, new_n1525_ );
or   ( new_n15918_, new_n10061_, new_n1318_ );
and  ( new_n15919_, new_n15918_, new_n15917_ );
xor  ( new_n15920_, new_n15919_, new_n9421_ );
and  ( new_n15921_, RIbb2d888_64, RIbb2cf28_84 );
or   ( new_n15922_, RIbb2d888_64, new_n1213_ );
and  ( new_n15923_, new_n15922_, RIbb2d900_63 );
or   ( new_n15924_, new_n15923_, new_n15921_ );
or   ( new_n15925_, new_n10770_, new_n1168_ );
and  ( new_n15926_, new_n15925_, new_n15924_ );
or   ( new_n15927_, new_n15926_, new_n15920_ );
and  ( new_n15928_, new_n15926_, new_n15920_ );
or   ( new_n15929_, new_n15928_, new_n895_ );
and  ( new_n15930_, new_n15929_, new_n15927_ );
or   ( new_n15931_, new_n7732_, new_n2646_ );
or   ( new_n15932_, new_n7734_, new_n2475_ );
and  ( new_n15933_, new_n15932_, new_n15931_ );
xor  ( new_n15934_, new_n15933_, new_n7177_ );
or   ( new_n15935_, new_n7184_, new_n2981_ );
or   ( new_n15936_, new_n7186_, new_n2751_ );
and  ( new_n15937_, new_n15936_, new_n15935_ );
xor  ( new_n15938_, new_n15937_, new_n6638_ );
or   ( new_n15939_, new_n15938_, new_n15934_ );
and  ( new_n15940_, new_n15938_, new_n15934_ );
or   ( new_n15941_, new_n6645_, new_n3306_ );
or   ( new_n15942_, new_n6647_, new_n3178_ );
and  ( new_n15943_, new_n15942_, new_n15941_ );
xor  ( new_n15944_, new_n15943_, new_n6166_ );
or   ( new_n15945_, new_n15944_, new_n15940_ );
and  ( new_n15946_, new_n15945_, new_n15939_ );
or   ( new_n15947_, new_n15946_, new_n15930_ );
and  ( new_n15948_, new_n15946_, new_n15930_ );
or   ( new_n15949_, new_n9422_, new_n1754_ );
or   ( new_n15950_, new_n9424_, new_n1523_ );
and  ( new_n15951_, new_n15950_, new_n15949_ );
xor  ( new_n15952_, new_n15951_, new_n8873_ );
or   ( new_n15953_, new_n8874_, new_n2057_ );
or   ( new_n15954_, new_n8876_, new_n1899_ );
and  ( new_n15955_, new_n15954_, new_n15953_ );
xor  ( new_n15956_, new_n15955_, new_n8257_ );
nor  ( new_n15957_, new_n15956_, new_n15952_ );
and  ( new_n15958_, new_n15956_, new_n15952_ );
or   ( new_n15959_, new_n8264_, new_n2291_ );
or   ( new_n15960_, new_n8266_, new_n2178_ );
and  ( new_n15961_, new_n15960_, new_n15959_ );
xor  ( new_n15962_, new_n15961_, new_n7725_ );
nor  ( new_n15963_, new_n15962_, new_n15958_ );
nor  ( new_n15964_, new_n15963_, new_n15957_ );
or   ( new_n15965_, new_n15964_, new_n15948_ );
and  ( new_n15966_, new_n15965_, new_n15947_ );
or   ( new_n15967_, new_n1364_, new_n10220_ );
or   ( new_n15968_, new_n1366_, new_n9679_ );
and  ( new_n15969_, new_n15968_, new_n15967_ );
xor  ( new_n15970_, new_n15969_, new_n1128_ );
or   ( new_n15971_, new_n1593_, new_n9679_ );
or   ( new_n15972_, new_n1595_, new_n9681_ );
and  ( new_n15973_, new_n15972_, new_n15971_ );
xor  ( new_n15974_, new_n15973_, new_n1358_ );
or   ( new_n15975_, new_n1364_, new_n10541_ );
or   ( new_n15976_, new_n1366_, new_n10220_ );
and  ( new_n15977_, new_n15976_, new_n15975_ );
xor  ( new_n15978_, new_n15977_, new_n1129_ );
nand ( new_n15979_, new_n15978_, new_n15974_ );
nor  ( new_n15980_, new_n15978_, new_n15974_ );
and  ( new_n15981_, new_n1040_, RIbb31578_128 );
nor  ( new_n15982_, new_n15981_, new_n896_ );
and  ( new_n15983_, new_n15981_, new_n893_ );
nor  ( new_n15984_, new_n15983_, new_n15982_ );
or   ( new_n15985_, new_n15984_, new_n15980_ );
and  ( new_n15986_, new_n15985_, new_n15979_ );
nand ( new_n15987_, new_n15986_, new_n15970_ );
nor  ( new_n15988_, new_n15986_, new_n15970_ );
or   ( new_n15989_, new_n2425_, new_n8115_ );
or   ( new_n15990_, new_n2427_, new_n8117_ );
and  ( new_n15991_, new_n15990_, new_n15989_ );
xor  ( new_n15992_, new_n15991_, new_n2121_ );
or   ( new_n15993_, new_n2122_, new_n8481_ );
or   ( new_n15994_, new_n2124_, new_n8352_ );
and  ( new_n15995_, new_n15994_, new_n15993_ );
xor  ( new_n15996_, new_n15995_, new_n1843_ );
nor  ( new_n15997_, new_n15996_, new_n15992_ );
and  ( new_n15998_, new_n15996_, new_n15992_ );
or   ( new_n15999_, new_n1844_, new_n9099_ );
or   ( new_n16000_, new_n1846_, new_n8995_ );
and  ( new_n16001_, new_n16000_, new_n15999_ );
xor  ( new_n16002_, new_n16001_, new_n1586_ );
nor  ( new_n16003_, new_n16002_, new_n15998_ );
nor  ( new_n16004_, new_n16003_, new_n15997_ );
or   ( new_n16005_, new_n16004_, new_n15988_ );
and  ( new_n16006_, new_n16005_, new_n15987_ );
nor  ( new_n16007_, new_n16006_, new_n15966_ );
nand ( new_n16008_, new_n16006_, new_n15966_ );
or   ( new_n16009_, new_n4709_, new_n4859_ );
or   ( new_n16010_, new_n4711_, new_n4995_ );
and  ( new_n16011_, new_n16010_, new_n16009_ );
xor  ( new_n16012_, new_n16011_, new_n4295_ );
or   ( new_n16013_, new_n4302_, new_n5428_ );
or   ( new_n16014_, new_n4304_, new_n5171_ );
and  ( new_n16015_, new_n16014_, new_n16013_ );
xor  ( new_n16016_, new_n16015_, new_n3895_ );
or   ( new_n16017_, new_n16016_, new_n16012_ );
and  ( new_n16018_, new_n16016_, new_n16012_ );
or   ( new_n16019_, new_n3896_, new_n5899_ );
or   ( new_n16020_, new_n3898_, new_n5570_ );
and  ( new_n16021_, new_n16020_, new_n16019_ );
xor  ( new_n16022_, new_n16021_, new_n3460_ );
or   ( new_n16023_, new_n16022_, new_n16018_ );
and  ( new_n16024_, new_n16023_, new_n16017_ );
or   ( new_n16025_, new_n6173_, new_n3694_ );
or   ( new_n16026_, new_n6175_, new_n3696_ );
and  ( new_n16027_, new_n16026_, new_n16025_ );
xor  ( new_n16028_, new_n16027_, new_n5597_ );
or   ( new_n16029_, new_n5604_, new_n4069_ );
or   ( new_n16030_, new_n5606_, new_n3820_ );
and  ( new_n16031_, new_n16030_, new_n16029_ );
xor  ( new_n16032_, new_n16031_, new_n5206_ );
or   ( new_n16033_, new_n16032_, new_n16028_ );
and  ( new_n16034_, new_n16032_, new_n16028_ );
or   ( new_n16035_, new_n5207_, new_n4603_ );
or   ( new_n16036_, new_n5209_, new_n4267_ );
and  ( new_n16037_, new_n16036_, new_n16035_ );
xor  ( new_n16038_, new_n16037_, new_n4708_ );
or   ( new_n16039_, new_n16038_, new_n16034_ );
and  ( new_n16040_, new_n16039_, new_n16033_ );
nor  ( new_n16041_, new_n16040_, new_n16024_ );
nand ( new_n16042_, new_n16040_, new_n16024_ );
or   ( new_n16043_, new_n3461_, new_n6425_ );
or   ( new_n16044_, new_n3463_, new_n6219_ );
and  ( new_n16045_, new_n16044_, new_n16043_ );
xor  ( new_n16046_, new_n16045_, new_n3116_ );
or   ( new_n16047_, new_n3117_, new_n6943_ );
or   ( new_n16048_, new_n3119_, new_n6589_ );
and  ( new_n16049_, new_n16048_, new_n16047_ );
xor  ( new_n16050_, new_n16049_, new_n2800_ );
nor  ( new_n16051_, new_n16050_, new_n16046_ );
and  ( new_n16052_, new_n16050_, new_n16046_ );
or   ( new_n16053_, new_n2807_, new_n7373_ );
or   ( new_n16054_, new_n2809_, new_n7149_ );
and  ( new_n16055_, new_n16054_, new_n16053_ );
xor  ( new_n16056_, new_n16055_, new_n2424_ );
nor  ( new_n16057_, new_n16056_, new_n16052_ );
or   ( new_n16058_, new_n16057_, new_n16051_ );
and  ( new_n16059_, new_n16058_, new_n16042_ );
or   ( new_n16060_, new_n16059_, new_n16041_ );
and  ( new_n16061_, new_n16060_, new_n16008_ );
or   ( new_n16062_, new_n16061_, new_n16007_ );
or   ( new_n16063_, new_n1135_, new_n10841_ );
or   ( new_n16064_, new_n1137_, new_n10541_ );
and  ( new_n16065_, new_n16064_, new_n16063_ );
xor  ( new_n16066_, new_n16065_, new_n895_ );
xnor ( new_n16067_, new_n15811_, new_n15807_ );
xor  ( new_n16068_, new_n16067_, new_n15817_ );
and  ( new_n16069_, new_n16068_, new_n16066_ );
or   ( new_n16070_, new_n16068_, new_n16066_ );
xnor ( new_n16071_, new_n15840_, new_n15836_ );
xor  ( new_n16072_, new_n16071_, new_n15846_ );
and  ( new_n16073_, new_n16072_, new_n16070_ );
or   ( new_n16074_, new_n16073_, new_n16069_ );
xnor ( new_n16075_, new_n15793_, new_n15789_ );
xor  ( new_n16076_, new_n16075_, new_n15799_ );
xnor ( new_n16077_, new_n15777_, new_n15773_ );
xor  ( new_n16078_, new_n16077_, new_n15783_ );
or   ( new_n16079_, new_n16078_, new_n16076_ );
and  ( new_n16080_, new_n16078_, new_n16076_ );
xor  ( new_n16081_, new_n15723_, new_n15719_ );
xnor ( new_n16082_, new_n16081_, new_n15729_ );
or   ( new_n16083_, new_n16082_, new_n16080_ );
and  ( new_n16084_, new_n16083_, new_n16079_ );
or   ( new_n16085_, new_n16084_, new_n16074_ );
and  ( new_n16086_, new_n16084_, new_n16074_ );
xor  ( new_n16087_, new_n15626_, new_n15620_ );
xor  ( new_n16088_, new_n16087_, new_n748_ );
or   ( new_n16089_, new_n16088_, new_n16086_ );
and  ( new_n16090_, new_n16089_, new_n16085_ );
or   ( new_n16091_, new_n16090_, new_n16062_ );
and  ( new_n16092_, new_n16090_, new_n16062_ );
xor  ( new_n16093_, new_n15829_, new_n15827_ );
xor  ( new_n16094_, new_n16093_, new_n15848_ );
xnor ( new_n16095_, new_n15695_, new_n15693_ );
xor  ( new_n16096_, new_n16095_, new_n15699_ );
nor  ( new_n16097_, new_n16096_, new_n16094_ );
nand ( new_n16098_, new_n16096_, new_n16094_ );
xor  ( new_n16099_, new_n15707_, new_n15705_ );
xnor ( new_n16100_, new_n16099_, new_n15711_ );
not  ( new_n16101_, new_n16100_ );
and  ( new_n16102_, new_n16101_, new_n16098_ );
or   ( new_n16103_, new_n16102_, new_n16097_ );
or   ( new_n16104_, new_n16103_, new_n16092_ );
and  ( new_n16105_, new_n16104_, new_n16091_ );
nor  ( new_n16106_, new_n16105_, new_n15916_ );
and  ( new_n16107_, new_n16105_, new_n15916_ );
xor  ( new_n16108_, new_n15540_, new_n15524_ );
xor  ( new_n16109_, new_n16108_, new_n15558_ );
xor  ( new_n16110_, new_n15646_, new_n15630_ );
xor  ( new_n16111_, new_n16110_, new_n15616_ );
and  ( new_n16112_, new_n16111_, new_n16109_ );
nor  ( new_n16113_, new_n16111_, new_n16109_ );
xor  ( new_n16114_, new_n15857_, new_n15855_ );
xnor ( new_n16115_, new_n16114_, new_n15861_ );
not  ( new_n16116_, new_n16115_ );
nor  ( new_n16117_, new_n16116_, new_n16113_ );
nor  ( new_n16118_, new_n16117_, new_n16112_ );
nor  ( new_n16119_, new_n16118_, new_n16107_ );
nor  ( new_n16120_, new_n16119_, new_n16106_ );
not  ( new_n16121_, new_n16120_ );
and  ( new_n16122_, new_n16121_, new_n15911_ );
or   ( new_n16123_, new_n16122_, new_n15910_ );
xnor ( new_n16124_, new_n15468_, new_n15466_ );
xor  ( new_n16125_, new_n16124_, new_n15655_ );
nand ( new_n16126_, new_n16125_, new_n16123_ );
or   ( new_n16127_, new_n16125_, new_n16123_ );
xor  ( new_n16128_, new_n15681_, new_n15671_ );
xor  ( new_n16129_, new_n16128_, new_n15882_ );
nand ( new_n16130_, new_n16129_, new_n16127_ );
and  ( new_n16131_, new_n16130_, new_n16126_ );
nor  ( new_n16132_, new_n16131_, new_n15895_ );
xor  ( new_n16133_, new_n15904_, new_n15902_ );
xor  ( new_n16134_, new_n16133_, new_n15907_ );
xnor ( new_n16135_, new_n15801_, new_n15785_ );
xor  ( new_n16136_, new_n16135_, new_n15819_ );
xnor ( new_n16137_, new_n15946_, new_n15930_ );
xor  ( new_n16138_, new_n16137_, new_n15964_ );
xor  ( new_n16139_, new_n16040_, new_n16024_ );
xor  ( new_n16140_, new_n16139_, new_n16058_ );
or   ( new_n16141_, new_n16140_, new_n16138_ );
and  ( new_n16142_, new_n16140_, new_n16138_ );
xor  ( new_n16143_, new_n15986_, new_n15970_ );
xnor ( new_n16144_, new_n16143_, new_n16004_ );
or   ( new_n16145_, new_n16144_, new_n16142_ );
and  ( new_n16146_, new_n16145_, new_n16141_ );
nor  ( new_n16147_, new_n16146_, new_n16136_ );
and  ( new_n16148_, new_n16146_, new_n16136_ );
xor  ( new_n16149_, new_n15747_, new_n15731_ );
xnor ( new_n16150_, new_n16149_, new_n15767_ );
nor  ( new_n16151_, new_n16150_, new_n16148_ );
or   ( new_n16152_, new_n16151_, new_n16147_ );
xnor ( new_n16153_, new_n15739_, new_n15735_ );
xor  ( new_n16154_, new_n16153_, new_n15745_ );
xor  ( new_n16155_, new_n15926_, new_n15920_ );
xor  ( new_n16156_, new_n16155_, new_n896_ );
xnor ( new_n16157_, new_n15938_, new_n15934_ );
xor  ( new_n16158_, new_n16157_, new_n15944_ );
or   ( new_n16159_, new_n16158_, new_n16156_ );
and  ( new_n16160_, new_n16158_, new_n16156_ );
xnor ( new_n16161_, new_n15956_, new_n15952_ );
xor  ( new_n16162_, new_n16161_, new_n15962_ );
or   ( new_n16163_, new_n16162_, new_n16160_ );
and  ( new_n16164_, new_n16163_, new_n16159_ );
nor  ( new_n16165_, new_n16164_, new_n16154_ );
nand ( new_n16166_, new_n16164_, new_n16154_ );
xnor ( new_n16167_, new_n16032_, new_n16028_ );
xor  ( new_n16168_, new_n16167_, new_n16038_ );
xnor ( new_n16169_, new_n16016_, new_n16012_ );
xor  ( new_n16170_, new_n16169_, new_n16022_ );
nor  ( new_n16171_, new_n16170_, new_n16168_ );
nand ( new_n16172_, new_n16170_, new_n16168_ );
xor  ( new_n16173_, new_n16050_, new_n16046_ );
xor  ( new_n16174_, new_n16173_, new_n16056_ );
and  ( new_n16175_, new_n16174_, new_n16172_ );
or   ( new_n16176_, new_n16175_, new_n16171_ );
and  ( new_n16177_, new_n16176_, new_n16166_ );
or   ( new_n16178_, new_n16177_, new_n16165_ );
or   ( new_n16179_, new_n8874_, new_n2178_ );
or   ( new_n16180_, new_n8876_, new_n2057_ );
and  ( new_n16181_, new_n16180_, new_n16179_ );
xor  ( new_n16182_, new_n16181_, new_n8257_ );
or   ( new_n16183_, new_n8264_, new_n2475_ );
or   ( new_n16184_, new_n8266_, new_n2291_ );
and  ( new_n16185_, new_n16184_, new_n16183_ );
xor  ( new_n16186_, new_n16185_, new_n7725_ );
or   ( new_n16187_, new_n16186_, new_n16182_ );
and  ( new_n16188_, new_n16186_, new_n16182_ );
or   ( new_n16189_, new_n7732_, new_n2751_ );
or   ( new_n16190_, new_n7734_, new_n2646_ );
and  ( new_n16191_, new_n16190_, new_n16189_ );
xor  ( new_n16192_, new_n16191_, new_n7177_ );
or   ( new_n16193_, new_n16192_, new_n16188_ );
and  ( new_n16194_, new_n16193_, new_n16187_ );
or   ( new_n16195_, new_n10059_, new_n1523_ );
or   ( new_n16196_, new_n10061_, new_n1525_ );
and  ( new_n16197_, new_n16196_, new_n16195_ );
xor  ( new_n16198_, new_n16197_, new_n9421_ );
and  ( new_n16199_, RIbb2d888_64, RIbb2ceb0_85 );
or   ( new_n16200_, RIbb2d888_64, new_n1318_ );
and  ( new_n16201_, new_n16200_, RIbb2d900_63 );
or   ( new_n16202_, new_n16201_, new_n16199_ );
or   ( new_n16203_, new_n10770_, new_n1213_ );
and  ( new_n16204_, new_n16203_, new_n16202_ );
or   ( new_n16205_, new_n16204_, new_n16198_ );
and  ( new_n16206_, new_n16204_, new_n16198_ );
or   ( new_n16207_, new_n9422_, new_n1899_ );
or   ( new_n16208_, new_n9424_, new_n1754_ );
and  ( new_n16209_, new_n16208_, new_n16207_ );
xor  ( new_n16210_, new_n16209_, new_n8873_ );
or   ( new_n16211_, new_n16210_, new_n16206_ );
and  ( new_n16212_, new_n16211_, new_n16205_ );
or   ( new_n16213_, new_n16212_, new_n16194_ );
and  ( new_n16214_, new_n16212_, new_n16194_ );
or   ( new_n16215_, new_n7184_, new_n3178_ );
or   ( new_n16216_, new_n7186_, new_n2981_ );
and  ( new_n16217_, new_n16216_, new_n16215_ );
xor  ( new_n16218_, new_n16217_, new_n6638_ );
or   ( new_n16219_, new_n6645_, new_n3696_ );
or   ( new_n16220_, new_n6647_, new_n3306_ );
and  ( new_n16221_, new_n16220_, new_n16219_ );
xor  ( new_n16222_, new_n16221_, new_n6166_ );
or   ( new_n16223_, new_n16222_, new_n16218_ );
and  ( new_n16224_, new_n16222_, new_n16218_ );
or   ( new_n16225_, new_n6173_, new_n3820_ );
or   ( new_n16226_, new_n6175_, new_n3694_ );
and  ( new_n16227_, new_n16226_, new_n16225_ );
xor  ( new_n16228_, new_n16227_, new_n5597_ );
or   ( new_n16229_, new_n16228_, new_n16224_ );
and  ( new_n16230_, new_n16229_, new_n16223_ );
or   ( new_n16231_, new_n16230_, new_n16214_ );
and  ( new_n16232_, new_n16231_, new_n16213_ );
xor  ( new_n16233_, new_n15996_, new_n15992_ );
xor  ( new_n16234_, new_n16233_, new_n16002_ );
or   ( new_n16235_, new_n2122_, new_n8995_ );
or   ( new_n16236_, new_n2124_, new_n8481_ );
and  ( new_n16237_, new_n16236_, new_n16235_ );
xor  ( new_n16238_, new_n16237_, new_n1843_ );
or   ( new_n16239_, new_n1844_, new_n9681_ );
or   ( new_n16240_, new_n1846_, new_n9099_ );
and  ( new_n16241_, new_n16240_, new_n16239_ );
xor  ( new_n16242_, new_n16241_, new_n1586_ );
or   ( new_n16243_, new_n16242_, new_n16238_ );
and  ( new_n16244_, new_n16242_, new_n16238_ );
or   ( new_n16245_, new_n1593_, new_n10220_ );
or   ( new_n16246_, new_n1595_, new_n9679_ );
and  ( new_n16247_, new_n16246_, new_n16245_ );
xor  ( new_n16248_, new_n16247_, new_n1358_ );
or   ( new_n16249_, new_n16248_, new_n16244_ );
and  ( new_n16250_, new_n16249_, new_n16243_ );
or   ( new_n16251_, new_n16250_, new_n16234_ );
and  ( new_n16252_, new_n16250_, new_n16234_ );
xor  ( new_n16253_, new_n15978_, new_n15974_ );
xnor ( new_n16254_, new_n16253_, new_n15984_ );
or   ( new_n16255_, new_n16254_, new_n16252_ );
and  ( new_n16256_, new_n16255_, new_n16251_ );
or   ( new_n16257_, new_n16256_, new_n16232_ );
and  ( new_n16258_, new_n16256_, new_n16232_ );
or   ( new_n16259_, new_n3117_, new_n7149_ );
or   ( new_n16260_, new_n3119_, new_n6943_ );
and  ( new_n16261_, new_n16260_, new_n16259_ );
xor  ( new_n16262_, new_n16261_, new_n2800_ );
or   ( new_n16263_, new_n2807_, new_n8117_ );
or   ( new_n16264_, new_n2809_, new_n7373_ );
and  ( new_n16265_, new_n16264_, new_n16263_ );
xor  ( new_n16266_, new_n16265_, new_n2424_ );
or   ( new_n16267_, new_n16266_, new_n16262_ );
and  ( new_n16268_, new_n16266_, new_n16262_ );
or   ( new_n16269_, new_n2425_, new_n8352_ );
or   ( new_n16270_, new_n2427_, new_n8115_ );
and  ( new_n16271_, new_n16270_, new_n16269_ );
xor  ( new_n16272_, new_n16271_, new_n2121_ );
or   ( new_n16273_, new_n16272_, new_n16268_ );
and  ( new_n16274_, new_n16273_, new_n16267_ );
or   ( new_n16275_, new_n4302_, new_n5570_ );
or   ( new_n16276_, new_n4304_, new_n5428_ );
and  ( new_n16277_, new_n16276_, new_n16275_ );
xor  ( new_n16278_, new_n16277_, new_n3895_ );
or   ( new_n16279_, new_n3896_, new_n6219_ );
or   ( new_n16280_, new_n3898_, new_n5899_ );
and  ( new_n16281_, new_n16280_, new_n16279_ );
xor  ( new_n16282_, new_n16281_, new_n3460_ );
or   ( new_n16283_, new_n16282_, new_n16278_ );
and  ( new_n16284_, new_n16282_, new_n16278_ );
or   ( new_n16285_, new_n3461_, new_n6589_ );
or   ( new_n16286_, new_n3463_, new_n6425_ );
and  ( new_n16287_, new_n16286_, new_n16285_ );
xor  ( new_n16288_, new_n16287_, new_n3116_ );
or   ( new_n16289_, new_n16288_, new_n16284_ );
and  ( new_n16290_, new_n16289_, new_n16283_ );
nor  ( new_n16291_, new_n16290_, new_n16274_ );
and  ( new_n16292_, new_n16290_, new_n16274_ );
or   ( new_n16293_, new_n5604_, new_n4267_ );
or   ( new_n16294_, new_n5606_, new_n4069_ );
and  ( new_n16295_, new_n16294_, new_n16293_ );
xor  ( new_n16296_, new_n16295_, new_n5206_ );
or   ( new_n16297_, new_n5207_, new_n4995_ );
or   ( new_n16298_, new_n5209_, new_n4603_ );
and  ( new_n16299_, new_n16298_, new_n16297_ );
xor  ( new_n16300_, new_n16299_, new_n4708_ );
nor  ( new_n16301_, new_n16300_, new_n16296_ );
and  ( new_n16302_, new_n16300_, new_n16296_ );
or   ( new_n16303_, new_n4709_, new_n5171_ );
or   ( new_n16304_, new_n4711_, new_n4859_ );
and  ( new_n16305_, new_n16304_, new_n16303_ );
xor  ( new_n16306_, new_n16305_, new_n4295_ );
nor  ( new_n16307_, new_n16306_, new_n16302_ );
nor  ( new_n16308_, new_n16307_, new_n16301_ );
nor  ( new_n16309_, new_n16308_, new_n16292_ );
nor  ( new_n16310_, new_n16309_, new_n16291_ );
or   ( new_n16311_, new_n16310_, new_n16258_ );
and  ( new_n16312_, new_n16311_, new_n16257_ );
or   ( new_n16313_, new_n16312_, new_n16178_ );
nand ( new_n16314_, new_n16312_, new_n16178_ );
xnor ( new_n16315_, new_n15759_, new_n15753_ );
xor  ( new_n16316_, new_n16315_, new_n15765_ );
xor  ( new_n16317_, new_n16068_, new_n16066_ );
xor  ( new_n16318_, new_n16317_, new_n16072_ );
nor  ( new_n16319_, new_n16318_, new_n16316_ );
and  ( new_n16320_, new_n16318_, new_n16316_ );
xor  ( new_n16321_, new_n16078_, new_n16076_ );
xnor ( new_n16322_, new_n16321_, new_n16082_ );
not  ( new_n16323_, new_n16322_ );
nor  ( new_n16324_, new_n16323_, new_n16320_ );
nor  ( new_n16325_, new_n16324_, new_n16319_ );
nand ( new_n16326_, new_n16325_, new_n16314_ );
and  ( new_n16327_, new_n16326_, new_n16313_ );
or   ( new_n16328_, new_n16327_, new_n16152_ );
nand ( new_n16329_, new_n16327_, new_n16152_ );
xor  ( new_n16330_, new_n16084_, new_n16074_ );
xor  ( new_n16331_, new_n16330_, new_n16088_ );
xor  ( new_n16332_, new_n16006_, new_n15966_ );
xor  ( new_n16333_, new_n16332_, new_n16060_ );
nor  ( new_n16334_, new_n16333_, new_n16331_ );
and  ( new_n16335_, new_n16333_, new_n16331_ );
xor  ( new_n16336_, new_n16096_, new_n16094_ );
xor  ( new_n16337_, new_n16336_, new_n16101_ );
nor  ( new_n16338_, new_n16337_, new_n16335_ );
nor  ( new_n16339_, new_n16338_, new_n16334_ );
nand ( new_n16340_, new_n16339_, new_n16329_ );
and  ( new_n16341_, new_n16340_, new_n16328_ );
or   ( new_n16342_, new_n16341_, new_n16134_ );
nand ( new_n16343_, new_n16341_, new_n16134_ );
xor  ( new_n16344_, new_n16090_, new_n16062_ );
xor  ( new_n16345_, new_n16344_, new_n16103_ );
xor  ( new_n16346_, new_n16111_, new_n16109_ );
xor  ( new_n16347_, new_n16346_, new_n16116_ );
nor  ( new_n16348_, new_n16347_, new_n16345_ );
and  ( new_n16349_, new_n16347_, new_n16345_ );
xor  ( new_n16350_, new_n15915_, new_n15913_ );
not  ( new_n16351_, new_n16350_ );
nor  ( new_n16352_, new_n16351_, new_n16349_ );
nor  ( new_n16353_, new_n16352_, new_n16348_ );
nand ( new_n16354_, new_n16353_, new_n16343_ );
and  ( new_n16355_, new_n16354_, new_n16342_ );
xnor ( new_n16356_, new_n15866_, new_n15689_ );
xor  ( new_n16357_, new_n16356_, new_n15879_ );
or   ( new_n16358_, new_n16357_, new_n16355_ );
and  ( new_n16359_, new_n16357_, new_n16355_ );
xor  ( new_n16360_, new_n15909_, new_n15897_ );
xor  ( new_n16361_, new_n16360_, new_n16121_ );
or   ( new_n16362_, new_n16361_, new_n16359_ );
and  ( new_n16363_, new_n16362_, new_n16358_ );
xor  ( new_n16364_, new_n16125_, new_n16123_ );
xor  ( new_n16365_, new_n16364_, new_n16129_ );
and  ( new_n16366_, new_n16365_, new_n16363_ );
xnor ( new_n16367_, new_n16357_, new_n16355_ );
xor  ( new_n16368_, new_n16367_, new_n16361_ );
xnor ( new_n16369_, new_n16333_, new_n16331_ );
xor  ( new_n16370_, new_n16369_, new_n16337_ );
or   ( new_n16371_, new_n6173_, new_n4069_ );
or   ( new_n16372_, new_n6175_, new_n3820_ );
and  ( new_n16373_, new_n16372_, new_n16371_ );
xor  ( new_n16374_, new_n16373_, new_n5597_ );
or   ( new_n16375_, new_n5604_, new_n4603_ );
or   ( new_n16376_, new_n5606_, new_n4267_ );
and  ( new_n16377_, new_n16376_, new_n16375_ );
xor  ( new_n16378_, new_n16377_, new_n5206_ );
or   ( new_n16379_, new_n16378_, new_n16374_ );
and  ( new_n16380_, new_n16378_, new_n16374_ );
or   ( new_n16381_, new_n5207_, new_n4859_ );
or   ( new_n16382_, new_n5209_, new_n4995_ );
and  ( new_n16383_, new_n16382_, new_n16381_ );
xor  ( new_n16384_, new_n16383_, new_n4708_ );
or   ( new_n16385_, new_n16384_, new_n16380_ );
and  ( new_n16386_, new_n16385_, new_n16379_ );
or   ( new_n16387_, new_n3461_, new_n6943_ );
or   ( new_n16388_, new_n3463_, new_n6589_ );
and  ( new_n16389_, new_n16388_, new_n16387_ );
xor  ( new_n16390_, new_n16389_, new_n3116_ );
or   ( new_n16391_, new_n3117_, new_n7373_ );
or   ( new_n16392_, new_n3119_, new_n7149_ );
and  ( new_n16393_, new_n16392_, new_n16391_ );
xor  ( new_n16394_, new_n16393_, new_n2800_ );
or   ( new_n16395_, new_n16394_, new_n16390_ );
and  ( new_n16396_, new_n16394_, new_n16390_ );
or   ( new_n16397_, new_n2807_, new_n8115_ );
or   ( new_n16398_, new_n2809_, new_n8117_ );
and  ( new_n16399_, new_n16398_, new_n16397_ );
xor  ( new_n16400_, new_n16399_, new_n2424_ );
or   ( new_n16401_, new_n16400_, new_n16396_ );
and  ( new_n16402_, new_n16401_, new_n16395_ );
or   ( new_n16403_, new_n16402_, new_n16386_ );
and  ( new_n16404_, new_n16402_, new_n16386_ );
or   ( new_n16405_, new_n4709_, new_n5428_ );
or   ( new_n16406_, new_n4711_, new_n5171_ );
and  ( new_n16407_, new_n16406_, new_n16405_ );
xor  ( new_n16408_, new_n16407_, new_n4295_ );
or   ( new_n16409_, new_n4302_, new_n5899_ );
or   ( new_n16410_, new_n4304_, new_n5570_ );
and  ( new_n16411_, new_n16410_, new_n16409_ );
xor  ( new_n16412_, new_n16411_, new_n3895_ );
nor  ( new_n16413_, new_n16412_, new_n16408_ );
and  ( new_n16414_, new_n16412_, new_n16408_ );
or   ( new_n16415_, new_n3896_, new_n6425_ );
or   ( new_n16416_, new_n3898_, new_n6219_ );
and  ( new_n16417_, new_n16416_, new_n16415_ );
xor  ( new_n16418_, new_n16417_, new_n3460_ );
nor  ( new_n16419_, new_n16418_, new_n16414_ );
nor  ( new_n16420_, new_n16419_, new_n16413_ );
or   ( new_n16421_, new_n16420_, new_n16404_ );
and  ( new_n16422_, new_n16421_, new_n16403_ );
or   ( new_n16423_, new_n1593_, new_n10541_ );
or   ( new_n16424_, new_n1595_, new_n10220_ );
and  ( new_n16425_, new_n16424_, new_n16423_ );
xor  ( new_n16426_, new_n16425_, new_n1358_ );
not  ( new_n16427_, new_n16426_ );
and  ( new_n16428_, new_n1251_, RIbb31578_128 );
or   ( new_n16429_, new_n16428_, new_n1129_ );
nand ( new_n16430_, new_n16428_, new_n1126_ );
and  ( new_n16431_, new_n16430_, new_n16429_ );
nor  ( new_n16432_, new_n16431_, new_n16427_ );
or   ( new_n16433_, new_n1364_, new_n10841_ );
or   ( new_n16434_, new_n1366_, new_n10541_ );
and  ( new_n16435_, new_n16434_, new_n16433_ );
xor  ( new_n16436_, new_n16435_, new_n1129_ );
or   ( new_n16437_, new_n16436_, new_n16432_ );
and  ( new_n16438_, new_n16436_, new_n16432_ );
or   ( new_n16439_, new_n2425_, new_n8481_ );
or   ( new_n16440_, new_n2427_, new_n8352_ );
and  ( new_n16441_, new_n16440_, new_n16439_ );
xor  ( new_n16442_, new_n16441_, new_n2121_ );
or   ( new_n16443_, new_n2122_, new_n9099_ );
or   ( new_n16444_, new_n2124_, new_n8995_ );
and  ( new_n16445_, new_n16444_, new_n16443_ );
xor  ( new_n16446_, new_n16445_, new_n1843_ );
nor  ( new_n16447_, new_n16446_, new_n16442_ );
and  ( new_n16448_, new_n16446_, new_n16442_ );
or   ( new_n16449_, new_n1844_, new_n9679_ );
or   ( new_n16450_, new_n1846_, new_n9681_ );
and  ( new_n16451_, new_n16450_, new_n16449_ );
xor  ( new_n16452_, new_n16451_, new_n1586_ );
nor  ( new_n16453_, new_n16452_, new_n16448_ );
nor  ( new_n16454_, new_n16453_, new_n16447_ );
or   ( new_n16455_, new_n16454_, new_n16438_ );
and  ( new_n16456_, new_n16455_, new_n16437_ );
nor  ( new_n16457_, new_n16456_, new_n16422_ );
nand ( new_n16458_, new_n16456_, new_n16422_ );
or   ( new_n16459_, new_n10059_, new_n1754_ );
or   ( new_n16460_, new_n10061_, new_n1523_ );
and  ( new_n16461_, new_n16460_, new_n16459_ );
xor  ( new_n16462_, new_n16461_, new_n9421_ );
and  ( new_n16463_, RIbb2d888_64, RIbb2ce38_86 );
or   ( new_n16464_, RIbb2d888_64, new_n1525_ );
and  ( new_n16465_, new_n16464_, RIbb2d900_63 );
or   ( new_n16466_, new_n16465_, new_n16463_ );
or   ( new_n16467_, new_n10770_, new_n1318_ );
and  ( new_n16468_, new_n16467_, new_n16466_ );
or   ( new_n16469_, new_n16468_, new_n16462_ );
and  ( new_n16470_, new_n16468_, new_n16462_ );
or   ( new_n16471_, new_n16470_, new_n1128_ );
and  ( new_n16472_, new_n16471_, new_n16469_ );
or   ( new_n16473_, new_n7732_, new_n2981_ );
or   ( new_n16474_, new_n7734_, new_n2751_ );
and  ( new_n16475_, new_n16474_, new_n16473_ );
xor  ( new_n16476_, new_n16475_, new_n7177_ );
or   ( new_n16477_, new_n7184_, new_n3306_ );
or   ( new_n16478_, new_n7186_, new_n3178_ );
and  ( new_n16479_, new_n16478_, new_n16477_ );
xor  ( new_n16480_, new_n16479_, new_n6638_ );
or   ( new_n16481_, new_n16480_, new_n16476_ );
and  ( new_n16482_, new_n16480_, new_n16476_ );
or   ( new_n16483_, new_n6645_, new_n3694_ );
or   ( new_n16484_, new_n6647_, new_n3696_ );
and  ( new_n16485_, new_n16484_, new_n16483_ );
xor  ( new_n16486_, new_n16485_, new_n6166_ );
or   ( new_n16487_, new_n16486_, new_n16482_ );
and  ( new_n16488_, new_n16487_, new_n16481_ );
nor  ( new_n16489_, new_n16488_, new_n16472_ );
and  ( new_n16490_, new_n16488_, new_n16472_ );
or   ( new_n16491_, new_n9422_, new_n2057_ );
or   ( new_n16492_, new_n9424_, new_n1899_ );
and  ( new_n16493_, new_n16492_, new_n16491_ );
xor  ( new_n16494_, new_n16493_, new_n8873_ );
or   ( new_n16495_, new_n8874_, new_n2291_ );
or   ( new_n16496_, new_n8876_, new_n2178_ );
and  ( new_n16497_, new_n16496_, new_n16495_ );
xor  ( new_n16498_, new_n16497_, new_n8257_ );
nor  ( new_n16499_, new_n16498_, new_n16494_ );
and  ( new_n16500_, new_n16498_, new_n16494_ );
or   ( new_n16501_, new_n8264_, new_n2646_ );
or   ( new_n16502_, new_n8266_, new_n2475_ );
and  ( new_n16503_, new_n16502_, new_n16501_ );
xor  ( new_n16504_, new_n16503_, new_n7725_ );
nor  ( new_n16505_, new_n16504_, new_n16500_ );
nor  ( new_n16506_, new_n16505_, new_n16499_ );
nor  ( new_n16507_, new_n16506_, new_n16490_ );
nor  ( new_n16508_, new_n16507_, new_n16489_ );
not  ( new_n16509_, new_n16508_ );
and  ( new_n16510_, new_n16509_, new_n16458_ );
or   ( new_n16511_, new_n16510_, new_n16457_ );
xor  ( new_n16512_, new_n16158_, new_n16156_ );
xor  ( new_n16513_, new_n16512_, new_n16162_ );
xnor ( new_n16514_, new_n16282_, new_n16278_ );
xor  ( new_n16515_, new_n16514_, new_n16288_ );
xnor ( new_n16516_, new_n16242_, new_n16238_ );
xor  ( new_n16517_, new_n16516_, new_n16248_ );
or   ( new_n16518_, new_n16517_, new_n16515_ );
and  ( new_n16519_, new_n16517_, new_n16515_ );
xnor ( new_n16520_, new_n16266_, new_n16262_ );
xor  ( new_n16521_, new_n16520_, new_n16272_ );
or   ( new_n16522_, new_n16521_, new_n16519_ );
and  ( new_n16523_, new_n16522_, new_n16518_ );
or   ( new_n16524_, new_n16523_, new_n16513_ );
and  ( new_n16525_, new_n16523_, new_n16513_ );
xnor ( new_n16526_, new_n16186_, new_n16182_ );
xor  ( new_n16527_, new_n16526_, new_n16192_ );
xnor ( new_n16528_, new_n16300_, new_n16296_ );
xor  ( new_n16529_, new_n16528_, new_n16306_ );
nor  ( new_n16530_, new_n16529_, new_n16527_ );
and  ( new_n16531_, new_n16529_, new_n16527_ );
xor  ( new_n16532_, new_n16222_, new_n16218_ );
xnor ( new_n16533_, new_n16532_, new_n16228_ );
nor  ( new_n16534_, new_n16533_, new_n16531_ );
nor  ( new_n16535_, new_n16534_, new_n16530_ );
or   ( new_n16536_, new_n16535_, new_n16525_ );
and  ( new_n16537_, new_n16536_, new_n16524_ );
nand ( new_n16538_, new_n16537_, new_n16511_ );
or   ( new_n16539_, new_n16537_, new_n16511_ );
xor  ( new_n16540_, new_n16290_, new_n16274_ );
xor  ( new_n16541_, new_n16540_, new_n16308_ );
xor  ( new_n16542_, new_n16170_, new_n16168_ );
xor  ( new_n16543_, new_n16542_, new_n16174_ );
and  ( new_n16544_, new_n16543_, new_n16541_ );
nor  ( new_n16545_, new_n16543_, new_n16541_ );
xor  ( new_n16546_, new_n16250_, new_n16234_ );
xnor ( new_n16547_, new_n16546_, new_n16254_ );
nor  ( new_n16548_, new_n16547_, new_n16545_ );
nor  ( new_n16549_, new_n16548_, new_n16544_ );
nand ( new_n16550_, new_n16549_, new_n16539_ );
and  ( new_n16551_, new_n16550_, new_n16538_ );
nor  ( new_n16552_, new_n16551_, new_n16370_ );
nand ( new_n16553_, new_n16551_, new_n16370_ );
xnor ( new_n16554_, new_n16140_, new_n16138_ );
xor  ( new_n16555_, new_n16554_, new_n16144_ );
xor  ( new_n16556_, new_n16164_, new_n16154_ );
xor  ( new_n16557_, new_n16556_, new_n16176_ );
nand ( new_n16558_, new_n16557_, new_n16555_ );
nor  ( new_n16559_, new_n16557_, new_n16555_ );
xor  ( new_n16560_, new_n16318_, new_n16316_ );
xor  ( new_n16561_, new_n16560_, new_n16323_ );
or   ( new_n16562_, new_n16561_, new_n16559_ );
and  ( new_n16563_, new_n16562_, new_n16558_ );
and  ( new_n16564_, new_n16563_, new_n16553_ );
or   ( new_n16565_, new_n16564_, new_n16552_ );
xor  ( new_n16566_, new_n16327_, new_n16152_ );
xor  ( new_n16567_, new_n16566_, new_n16339_ );
nor  ( new_n16568_, new_n16567_, new_n16565_ );
and  ( new_n16569_, new_n16567_, new_n16565_ );
xor  ( new_n16570_, new_n16347_, new_n16345_ );
xor  ( new_n16571_, new_n16570_, new_n16351_ );
nor  ( new_n16572_, new_n16571_, new_n16569_ );
or   ( new_n16573_, new_n16572_, new_n16568_ );
xnor ( new_n16574_, new_n16105_, new_n15916_ );
xor  ( new_n16575_, new_n16574_, new_n16118_ );
nand ( new_n16576_, new_n16575_, new_n16573_ );
nor  ( new_n16577_, new_n16575_, new_n16573_ );
xor  ( new_n16578_, new_n16341_, new_n16134_ );
xor  ( new_n16579_, new_n16578_, new_n16353_ );
or   ( new_n16580_, new_n16579_, new_n16577_ );
and  ( new_n16581_, new_n16580_, new_n16576_ );
nor  ( new_n16582_, new_n16581_, new_n16368_ );
xor  ( new_n16583_, new_n16575_, new_n16573_ );
xor  ( new_n16584_, new_n16583_, new_n16579_ );
xor  ( new_n16585_, new_n16312_, new_n16178_ );
xor  ( new_n16586_, new_n16585_, new_n16325_ );
xor  ( new_n16587_, new_n16551_, new_n16370_ );
xor  ( new_n16588_, new_n16587_, new_n16563_ );
or   ( new_n16589_, new_n16588_, new_n16586_ );
xor  ( new_n16590_, new_n16537_, new_n16511_ );
xor  ( new_n16591_, new_n16590_, new_n16549_ );
xnor ( new_n16592_, new_n16557_, new_n16555_ );
xnor ( new_n16593_, new_n16592_, new_n16561_ );
or   ( new_n16594_, new_n16593_, new_n16591_ );
xor  ( new_n16595_, new_n16212_, new_n16194_ );
xor  ( new_n16596_, new_n16595_, new_n16230_ );
xnor ( new_n16597_, new_n16523_, new_n16513_ );
xor  ( new_n16598_, new_n16597_, new_n16535_ );
nand ( new_n16599_, new_n16598_, new_n16596_ );
nor  ( new_n16600_, new_n16598_, new_n16596_ );
xor  ( new_n16601_, new_n16543_, new_n16541_ );
xor  ( new_n16602_, new_n16601_, new_n16547_ );
or   ( new_n16603_, new_n16602_, new_n16600_ );
and  ( new_n16604_, new_n16603_, new_n16599_ );
xnor ( new_n16605_, new_n16256_, new_n16232_ );
xor  ( new_n16606_, new_n16605_, new_n16310_ );
or   ( new_n16607_, new_n16606_, new_n16604_ );
and  ( new_n16608_, new_n16606_, new_n16604_ );
xnor ( new_n16609_, new_n16204_, new_n16198_ );
xor  ( new_n16610_, new_n16609_, new_n16210_ );
xnor ( new_n16611_, new_n16394_, new_n16390_ );
xor  ( new_n16612_, new_n16611_, new_n16400_ );
xnor ( new_n16613_, new_n16378_, new_n16374_ );
xor  ( new_n16614_, new_n16613_, new_n16384_ );
or   ( new_n16615_, new_n16614_, new_n16612_ );
and  ( new_n16616_, new_n16614_, new_n16612_ );
xor  ( new_n16617_, new_n16412_, new_n16408_ );
xnor ( new_n16618_, new_n16617_, new_n16418_ );
or   ( new_n16619_, new_n16618_, new_n16616_ );
and  ( new_n16620_, new_n16619_, new_n16615_ );
nor  ( new_n16621_, new_n16620_, new_n16610_ );
and  ( new_n16622_, new_n16620_, new_n16610_ );
xor  ( new_n16623_, new_n16468_, new_n16462_ );
xor  ( new_n16624_, new_n16623_, new_n1129_ );
xnor ( new_n16625_, new_n16480_, new_n16476_ );
xor  ( new_n16626_, new_n16625_, new_n16486_ );
nor  ( new_n16627_, new_n16626_, new_n16624_ );
and  ( new_n16628_, new_n16626_, new_n16624_ );
xor  ( new_n16629_, new_n16498_, new_n16494_ );
xnor ( new_n16630_, new_n16629_, new_n16504_ );
nor  ( new_n16631_, new_n16630_, new_n16628_ );
nor  ( new_n16632_, new_n16631_, new_n16627_ );
nor  ( new_n16633_, new_n16632_, new_n16622_ );
or   ( new_n16634_, new_n16633_, new_n16621_ );
xor  ( new_n16635_, new_n16517_, new_n16515_ );
xor  ( new_n16636_, new_n16635_, new_n16521_ );
xnor ( new_n16637_, new_n16436_, new_n16432_ );
xor  ( new_n16638_, new_n16637_, new_n16454_ );
nand ( new_n16639_, new_n16638_, new_n16636_ );
nor  ( new_n16640_, new_n16638_, new_n16636_ );
xor  ( new_n16641_, new_n16529_, new_n16527_ );
xnor ( new_n16642_, new_n16641_, new_n16533_ );
or   ( new_n16643_, new_n16642_, new_n16640_ );
and  ( new_n16644_, new_n16643_, new_n16639_ );
nor  ( new_n16645_, new_n16644_, new_n16634_ );
nand ( new_n16646_, new_n16644_, new_n16634_ );
or   ( new_n16647_, new_n3117_, new_n8117_ );
or   ( new_n16648_, new_n3119_, new_n7373_ );
and  ( new_n16649_, new_n16648_, new_n16647_ );
xor  ( new_n16650_, new_n16649_, new_n2800_ );
or   ( new_n16651_, new_n2807_, new_n8352_ );
or   ( new_n16652_, new_n2809_, new_n8115_ );
and  ( new_n16653_, new_n16652_, new_n16651_ );
xor  ( new_n16654_, new_n16653_, new_n2424_ );
or   ( new_n16655_, new_n16654_, new_n16650_ );
and  ( new_n16656_, new_n16654_, new_n16650_ );
or   ( new_n16657_, new_n2425_, new_n8995_ );
or   ( new_n16658_, new_n2427_, new_n8481_ );
and  ( new_n16659_, new_n16658_, new_n16657_ );
xor  ( new_n16660_, new_n16659_, new_n2121_ );
or   ( new_n16661_, new_n16660_, new_n16656_ );
and  ( new_n16662_, new_n16661_, new_n16655_ );
or   ( new_n16663_, new_n4302_, new_n6219_ );
or   ( new_n16664_, new_n4304_, new_n5899_ );
and  ( new_n16665_, new_n16664_, new_n16663_ );
xor  ( new_n16666_, new_n16665_, new_n3895_ );
or   ( new_n16667_, new_n3896_, new_n6589_ );
or   ( new_n16668_, new_n3898_, new_n6425_ );
and  ( new_n16669_, new_n16668_, new_n16667_ );
xor  ( new_n16670_, new_n16669_, new_n3460_ );
or   ( new_n16671_, new_n16670_, new_n16666_ );
and  ( new_n16672_, new_n16670_, new_n16666_ );
or   ( new_n16673_, new_n3461_, new_n7149_ );
or   ( new_n16674_, new_n3463_, new_n6943_ );
and  ( new_n16675_, new_n16674_, new_n16673_ );
xor  ( new_n16676_, new_n16675_, new_n3116_ );
or   ( new_n16677_, new_n16676_, new_n16672_ );
and  ( new_n16678_, new_n16677_, new_n16671_ );
or   ( new_n16679_, new_n16678_, new_n16662_ );
and  ( new_n16680_, new_n16678_, new_n16662_ );
or   ( new_n16681_, new_n5604_, new_n4995_ );
or   ( new_n16682_, new_n5606_, new_n4603_ );
and  ( new_n16683_, new_n16682_, new_n16681_ );
xor  ( new_n16684_, new_n16683_, new_n5206_ );
or   ( new_n16685_, new_n5207_, new_n5171_ );
or   ( new_n16686_, new_n5209_, new_n4859_ );
and  ( new_n16687_, new_n16686_, new_n16685_ );
xor  ( new_n16688_, new_n16687_, new_n4708_ );
or   ( new_n16689_, new_n16688_, new_n16684_ );
and  ( new_n16690_, new_n16688_, new_n16684_ );
or   ( new_n16691_, new_n4709_, new_n5570_ );
or   ( new_n16692_, new_n4711_, new_n5428_ );
and  ( new_n16693_, new_n16692_, new_n16691_ );
xor  ( new_n16694_, new_n16693_, new_n4295_ );
or   ( new_n16695_, new_n16694_, new_n16690_ );
and  ( new_n16696_, new_n16695_, new_n16689_ );
or   ( new_n16697_, new_n16696_, new_n16680_ );
and  ( new_n16698_, new_n16697_, new_n16679_ );
xor  ( new_n16699_, new_n16446_, new_n16442_ );
xor  ( new_n16700_, new_n16699_, new_n16452_ );
or   ( new_n16701_, new_n2122_, new_n9681_ );
or   ( new_n16702_, new_n2124_, new_n9099_ );
and  ( new_n16703_, new_n16702_, new_n16701_ );
xor  ( new_n16704_, new_n16703_, new_n1843_ );
or   ( new_n16705_, new_n1844_, new_n10220_ );
or   ( new_n16706_, new_n1846_, new_n9679_ );
and  ( new_n16707_, new_n16706_, new_n16705_ );
xor  ( new_n16708_, new_n16707_, new_n1586_ );
or   ( new_n16709_, new_n16708_, new_n16704_ );
and  ( new_n16710_, new_n16708_, new_n16704_ );
or   ( new_n16711_, new_n1593_, new_n10841_ );
or   ( new_n16712_, new_n1595_, new_n10541_ );
and  ( new_n16713_, new_n16712_, new_n16711_ );
xor  ( new_n16714_, new_n16713_, new_n1358_ );
or   ( new_n16715_, new_n16714_, new_n16710_ );
and  ( new_n16716_, new_n16715_, new_n16709_ );
or   ( new_n16717_, new_n16716_, new_n16700_ );
and  ( new_n16718_, new_n16716_, new_n16700_ );
xor  ( new_n16719_, new_n16431_, new_n16427_ );
or   ( new_n16720_, new_n16719_, new_n16718_ );
and  ( new_n16721_, new_n16720_, new_n16717_ );
nor  ( new_n16722_, new_n16721_, new_n16698_ );
nand ( new_n16723_, new_n16721_, new_n16698_ );
or   ( new_n16724_, new_n8874_, new_n2475_ );
or   ( new_n16725_, new_n8876_, new_n2291_ );
and  ( new_n16726_, new_n16725_, new_n16724_ );
xor  ( new_n16727_, new_n16726_, new_n8257_ );
or   ( new_n16728_, new_n8264_, new_n2751_ );
or   ( new_n16729_, new_n8266_, new_n2646_ );
and  ( new_n16730_, new_n16729_, new_n16728_ );
xor  ( new_n16731_, new_n16730_, new_n7725_ );
or   ( new_n16732_, new_n16731_, new_n16727_ );
and  ( new_n16733_, new_n16731_, new_n16727_ );
or   ( new_n16734_, new_n7732_, new_n3178_ );
or   ( new_n16735_, new_n7734_, new_n2981_ );
and  ( new_n16736_, new_n16735_, new_n16734_ );
xor  ( new_n16737_, new_n16736_, new_n7177_ );
or   ( new_n16738_, new_n16737_, new_n16733_ );
and  ( new_n16739_, new_n16738_, new_n16732_ );
or   ( new_n16740_, new_n7184_, new_n3696_ );
or   ( new_n16741_, new_n7186_, new_n3306_ );
and  ( new_n16742_, new_n16741_, new_n16740_ );
xor  ( new_n16743_, new_n16742_, new_n6638_ );
or   ( new_n16744_, new_n6645_, new_n3820_ );
or   ( new_n16745_, new_n6647_, new_n3694_ );
and  ( new_n16746_, new_n16745_, new_n16744_ );
xor  ( new_n16747_, new_n16746_, new_n6166_ );
or   ( new_n16748_, new_n16747_, new_n16743_ );
and  ( new_n16749_, new_n16747_, new_n16743_ );
or   ( new_n16750_, new_n6173_, new_n4267_ );
or   ( new_n16751_, new_n6175_, new_n4069_ );
and  ( new_n16752_, new_n16751_, new_n16750_ );
xor  ( new_n16753_, new_n16752_, new_n5597_ );
or   ( new_n16754_, new_n16753_, new_n16749_ );
and  ( new_n16755_, new_n16754_, new_n16748_ );
nor  ( new_n16756_, new_n16755_, new_n16739_ );
nand ( new_n16757_, new_n16755_, new_n16739_ );
or   ( new_n16758_, new_n10059_, new_n1899_ );
or   ( new_n16759_, new_n10061_, new_n1754_ );
and  ( new_n16760_, new_n16759_, new_n16758_ );
xor  ( new_n16761_, new_n16760_, new_n9421_ );
and  ( new_n16762_, RIbb2d888_64, RIbb2cdc0_87 );
or   ( new_n16763_, RIbb2d888_64, new_n1523_ );
and  ( new_n16764_, new_n16763_, RIbb2d900_63 );
or   ( new_n16765_, new_n16764_, new_n16762_ );
or   ( new_n16766_, new_n10770_, new_n1525_ );
and  ( new_n16767_, new_n16766_, new_n16765_ );
nor  ( new_n16768_, new_n16767_, new_n16761_ );
nand ( new_n16769_, new_n16767_, new_n16761_ );
or   ( new_n16770_, new_n9422_, new_n2178_ );
or   ( new_n16771_, new_n9424_, new_n2057_ );
and  ( new_n16772_, new_n16771_, new_n16770_ );
xor  ( new_n16773_, new_n16772_, new_n8872_ );
and  ( new_n16774_, new_n16773_, new_n16769_ );
or   ( new_n16775_, new_n16774_, new_n16768_ );
and  ( new_n16776_, new_n16775_, new_n16757_ );
or   ( new_n16777_, new_n16776_, new_n16756_ );
and  ( new_n16778_, new_n16777_, new_n16723_ );
or   ( new_n16779_, new_n16778_, new_n16722_ );
and  ( new_n16780_, new_n16779_, new_n16646_ );
or   ( new_n16781_, new_n16780_, new_n16645_ );
or   ( new_n16782_, new_n16781_, new_n16608_ );
and  ( new_n16783_, new_n16782_, new_n16607_ );
or   ( new_n16784_, new_n16783_, new_n16594_ );
and  ( new_n16785_, new_n16783_, new_n16594_ );
xor  ( new_n16786_, new_n16146_, new_n16136_ );
xor  ( new_n16787_, new_n16786_, new_n16150_ );
or   ( new_n16788_, new_n16787_, new_n16785_ );
and  ( new_n16789_, new_n16788_, new_n16784_ );
or   ( new_n16790_, new_n16789_, new_n16589_ );
and  ( new_n16791_, new_n16789_, new_n16589_ );
xor  ( new_n16792_, new_n16567_, new_n16565_ );
xor  ( new_n16793_, new_n16792_, new_n16571_ );
or   ( new_n16794_, new_n16793_, new_n16791_ );
and  ( new_n16795_, new_n16794_, new_n16790_ );
nor  ( new_n16796_, new_n16795_, new_n16584_ );
xor  ( new_n16797_, new_n16789_, new_n16589_ );
xor  ( new_n16798_, new_n16797_, new_n16793_ );
xor  ( new_n16799_, new_n16783_, new_n16594_ );
xor  ( new_n16800_, new_n16799_, new_n16787_ );
xnor ( new_n16801_, new_n16402_, new_n16386_ );
xor  ( new_n16802_, new_n16801_, new_n16420_ );
xnor ( new_n16803_, new_n16488_, new_n16472_ );
xor  ( new_n16804_, new_n16803_, new_n16506_ );
nor  ( new_n16805_, new_n16804_, new_n16802_ );
and  ( new_n16806_, new_n16804_, new_n16802_ );
xor  ( new_n16807_, new_n16638_, new_n16636_ );
xnor ( new_n16808_, new_n16807_, new_n16642_ );
nor  ( new_n16809_, new_n16808_, new_n16806_ );
or   ( new_n16810_, new_n16809_, new_n16805_ );
xor  ( new_n16811_, new_n16708_, new_n16704_ );
xor  ( new_n16812_, new_n16811_, new_n16714_ );
or   ( new_n16813_, new_n2425_, new_n9099_ );
or   ( new_n16814_, new_n2427_, new_n8995_ );
and  ( new_n16815_, new_n16814_, new_n16813_ );
xor  ( new_n16816_, new_n16815_, new_n2121_ );
or   ( new_n16817_, new_n2122_, new_n9679_ );
or   ( new_n16818_, new_n2124_, new_n9681_ );
and  ( new_n16819_, new_n16818_, new_n16817_ );
xor  ( new_n16820_, new_n16819_, new_n1843_ );
or   ( new_n16821_, new_n16820_, new_n16816_ );
and  ( new_n16822_, new_n16820_, new_n16816_ );
or   ( new_n16823_, new_n1844_, new_n10541_ );
or   ( new_n16824_, new_n1846_, new_n10220_ );
and  ( new_n16825_, new_n16824_, new_n16823_ );
xor  ( new_n16826_, new_n16825_, new_n1586_ );
or   ( new_n16827_, new_n16826_, new_n16822_ );
and  ( new_n16828_, new_n16827_, new_n16821_ );
or   ( new_n16829_, new_n16828_, new_n16812_ );
nand ( new_n16830_, new_n16828_, new_n16812_ );
xor  ( new_n16831_, new_n16654_, new_n16650_ );
xnor ( new_n16832_, new_n16831_, new_n16660_ );
nand ( new_n16833_, new_n16832_, new_n16830_ );
and  ( new_n16834_, new_n16833_, new_n16829_ );
or   ( new_n16835_, new_n7732_, new_n3306_ );
or   ( new_n16836_, new_n7734_, new_n3178_ );
and  ( new_n16837_, new_n16836_, new_n16835_ );
xor  ( new_n16838_, new_n16837_, new_n7177_ );
or   ( new_n16839_, new_n7184_, new_n3694_ );
or   ( new_n16840_, new_n7186_, new_n3696_ );
and  ( new_n16841_, new_n16840_, new_n16839_ );
xor  ( new_n16842_, new_n16841_, new_n6638_ );
or   ( new_n16843_, new_n16842_, new_n16838_ );
and  ( new_n16844_, new_n16842_, new_n16838_ );
or   ( new_n16845_, new_n6645_, new_n4069_ );
or   ( new_n16846_, new_n6647_, new_n3820_ );
and  ( new_n16847_, new_n16846_, new_n16845_ );
xor  ( new_n16848_, new_n16847_, new_n6166_ );
or   ( new_n16849_, new_n16848_, new_n16844_ );
and  ( new_n16850_, new_n16849_, new_n16843_ );
or   ( new_n16851_, new_n10059_, new_n2057_ );
or   ( new_n16852_, new_n10061_, new_n1899_ );
and  ( new_n16853_, new_n16852_, new_n16851_ );
xor  ( new_n16854_, new_n16853_, new_n9421_ );
and  ( new_n16855_, RIbb2d888_64, RIbb2cd48_88 );
or   ( new_n16856_, RIbb2d888_64, new_n1754_ );
and  ( new_n16857_, new_n16856_, RIbb2d900_63 );
or   ( new_n16858_, new_n16857_, new_n16855_ );
or   ( new_n16859_, new_n10770_, new_n1523_ );
and  ( new_n16860_, new_n16859_, new_n16858_ );
nor  ( new_n16861_, new_n16860_, new_n16854_ );
and  ( new_n16862_, new_n16860_, new_n16854_ );
nor  ( new_n16863_, new_n16862_, new_n1357_ );
nor  ( new_n16864_, new_n16863_, new_n16861_ );
or   ( new_n16865_, new_n9422_, new_n2291_ );
or   ( new_n16866_, new_n9424_, new_n2178_ );
and  ( new_n16867_, new_n16866_, new_n16865_ );
xor  ( new_n16868_, new_n16867_, new_n8873_ );
or   ( new_n16869_, new_n8874_, new_n2646_ );
or   ( new_n16870_, new_n8876_, new_n2475_ );
and  ( new_n16871_, new_n16870_, new_n16869_ );
xor  ( new_n16872_, new_n16871_, new_n8257_ );
or   ( new_n16873_, new_n16872_, new_n16868_ );
and  ( new_n16874_, new_n16872_, new_n16868_ );
or   ( new_n16875_, new_n8264_, new_n2981_ );
or   ( new_n16876_, new_n8266_, new_n2751_ );
and  ( new_n16877_, new_n16876_, new_n16875_ );
xor  ( new_n16878_, new_n16877_, new_n7725_ );
or   ( new_n16879_, new_n16878_, new_n16874_ );
and  ( new_n16880_, new_n16879_, new_n16873_ );
and  ( new_n16881_, new_n16880_, new_n16864_ );
or   ( new_n16882_, new_n16881_, new_n16850_ );
or   ( new_n16883_, new_n16880_, new_n16864_ );
and  ( new_n16884_, new_n16883_, new_n16882_ );
nor  ( new_n16885_, new_n16884_, new_n16834_ );
nand ( new_n16886_, new_n16884_, new_n16834_ );
or   ( new_n16887_, new_n6173_, new_n4603_ );
or   ( new_n16888_, new_n6175_, new_n4267_ );
and  ( new_n16889_, new_n16888_, new_n16887_ );
xor  ( new_n16890_, new_n16889_, new_n5597_ );
or   ( new_n16891_, new_n5604_, new_n4859_ );
or   ( new_n16892_, new_n5606_, new_n4995_ );
and  ( new_n16893_, new_n16892_, new_n16891_ );
xor  ( new_n16894_, new_n16893_, new_n5206_ );
or   ( new_n16895_, new_n16894_, new_n16890_ );
and  ( new_n16896_, new_n16894_, new_n16890_ );
or   ( new_n16897_, new_n5207_, new_n5428_ );
or   ( new_n16898_, new_n5209_, new_n5171_ );
and  ( new_n16899_, new_n16898_, new_n16897_ );
xor  ( new_n16900_, new_n16899_, new_n4708_ );
or   ( new_n16901_, new_n16900_, new_n16896_ );
and  ( new_n16902_, new_n16901_, new_n16895_ );
or   ( new_n16903_, new_n3461_, new_n7373_ );
or   ( new_n16904_, new_n3463_, new_n7149_ );
and  ( new_n16905_, new_n16904_, new_n16903_ );
xor  ( new_n16906_, new_n16905_, new_n3116_ );
or   ( new_n16907_, new_n3117_, new_n8115_ );
or   ( new_n16908_, new_n3119_, new_n8117_ );
and  ( new_n16909_, new_n16908_, new_n16907_ );
xor  ( new_n16910_, new_n16909_, new_n2800_ );
or   ( new_n16911_, new_n16910_, new_n16906_ );
and  ( new_n16912_, new_n16910_, new_n16906_ );
or   ( new_n16913_, new_n2807_, new_n8481_ );
or   ( new_n16914_, new_n2809_, new_n8352_ );
and  ( new_n16915_, new_n16914_, new_n16913_ );
xor  ( new_n16916_, new_n16915_, new_n2424_ );
or   ( new_n16917_, new_n16916_, new_n16912_ );
and  ( new_n16918_, new_n16917_, new_n16911_ );
nor  ( new_n16919_, new_n16918_, new_n16902_ );
and  ( new_n16920_, new_n16918_, new_n16902_ );
or   ( new_n16921_, new_n4709_, new_n5899_ );
or   ( new_n16922_, new_n4711_, new_n5570_ );
and  ( new_n16923_, new_n16922_, new_n16921_ );
xor  ( new_n16924_, new_n16923_, new_n4295_ );
or   ( new_n16925_, new_n4302_, new_n6425_ );
or   ( new_n16926_, new_n4304_, new_n6219_ );
and  ( new_n16927_, new_n16926_, new_n16925_ );
xor  ( new_n16928_, new_n16927_, new_n3895_ );
nor  ( new_n16929_, new_n16928_, new_n16924_ );
and  ( new_n16930_, new_n16928_, new_n16924_ );
or   ( new_n16931_, new_n3896_, new_n6943_ );
or   ( new_n16932_, new_n3898_, new_n6589_ );
and  ( new_n16933_, new_n16932_, new_n16931_ );
xor  ( new_n16934_, new_n16933_, new_n3460_ );
nor  ( new_n16935_, new_n16934_, new_n16930_ );
nor  ( new_n16936_, new_n16935_, new_n16929_ );
nor  ( new_n16937_, new_n16936_, new_n16920_ );
nor  ( new_n16938_, new_n16937_, new_n16919_ );
not  ( new_n16939_, new_n16938_ );
and  ( new_n16940_, new_n16939_, new_n16886_ );
or   ( new_n16941_, new_n16940_, new_n16885_ );
xor  ( new_n16942_, new_n16731_, new_n16727_ );
xnor ( new_n16943_, new_n16942_, new_n16737_ );
xor  ( new_n16944_, new_n16767_, new_n16761_ );
xor  ( new_n16945_, new_n16944_, new_n16773_ );
or   ( new_n16946_, new_n16945_, new_n16943_ );
xnor ( new_n16947_, new_n16670_, new_n16666_ );
xor  ( new_n16948_, new_n16947_, new_n16676_ );
xnor ( new_n16949_, new_n16747_, new_n16743_ );
xor  ( new_n16950_, new_n16949_, new_n16753_ );
or   ( new_n16951_, new_n16950_, new_n16948_ );
and  ( new_n16952_, new_n16950_, new_n16948_ );
xnor ( new_n16953_, new_n16688_, new_n16684_ );
xor  ( new_n16954_, new_n16953_, new_n16694_ );
or   ( new_n16955_, new_n16954_, new_n16952_ );
and  ( new_n16956_, new_n16955_, new_n16951_ );
or   ( new_n16957_, new_n16956_, new_n16946_ );
and  ( new_n16958_, new_n16956_, new_n16946_ );
xor  ( new_n16959_, new_n16626_, new_n16624_ );
xor  ( new_n16960_, new_n16959_, new_n16630_ );
or   ( new_n16961_, new_n16960_, new_n16958_ );
and  ( new_n16962_, new_n16961_, new_n16957_ );
nand ( new_n16963_, new_n16962_, new_n16941_ );
or   ( new_n16964_, new_n16962_, new_n16941_ );
xor  ( new_n16965_, new_n16678_, new_n16662_ );
xor  ( new_n16966_, new_n16965_, new_n16696_ );
xnor ( new_n16967_, new_n16614_, new_n16612_ );
xor  ( new_n16968_, new_n16967_, new_n16618_ );
and  ( new_n16969_, new_n16968_, new_n16966_ );
nor  ( new_n16970_, new_n16968_, new_n16966_ );
xor  ( new_n16971_, new_n16716_, new_n16700_ );
xnor ( new_n16972_, new_n16971_, new_n16719_ );
nor  ( new_n16973_, new_n16972_, new_n16970_ );
nor  ( new_n16974_, new_n16973_, new_n16969_ );
nand ( new_n16975_, new_n16974_, new_n16964_ );
and  ( new_n16976_, new_n16975_, new_n16963_ );
nor  ( new_n16977_, new_n16976_, new_n16810_ );
nand ( new_n16978_, new_n16976_, new_n16810_ );
xor  ( new_n16979_, new_n16456_, new_n16422_ );
xor  ( new_n16980_, new_n16979_, new_n16509_ );
and  ( new_n16981_, new_n16980_, new_n16978_ );
or   ( new_n16982_, new_n16981_, new_n16977_ );
xor  ( new_n16983_, new_n16606_, new_n16604_ );
xor  ( new_n16984_, new_n16983_, new_n16781_ );
or   ( new_n16985_, new_n16984_, new_n16982_ );
and  ( new_n16986_, new_n16984_, new_n16982_ );
xnor ( new_n16987_, new_n16593_, new_n16591_ );
or   ( new_n16988_, new_n16987_, new_n16986_ );
and  ( new_n16989_, new_n16988_, new_n16985_ );
or   ( new_n16990_, new_n16989_, new_n16800_ );
and  ( new_n16991_, new_n16989_, new_n16800_ );
xnor ( new_n16992_, new_n16588_, new_n16586_ );
or   ( new_n16993_, new_n16992_, new_n16991_ );
and  ( new_n16994_, new_n16993_, new_n16990_ );
nor  ( new_n16995_, new_n16994_, new_n16798_ );
xor  ( new_n16996_, new_n16989_, new_n16800_ );
xor  ( new_n16997_, new_n16996_, new_n16992_ );
xor  ( new_n16998_, new_n16976_, new_n16810_ );
xor  ( new_n16999_, new_n16998_, new_n16980_ );
xor  ( new_n17000_, new_n16644_, new_n16634_ );
xor  ( new_n17001_, new_n17000_, new_n16779_ );
or   ( new_n17002_, new_n17001_, new_n16999_ );
xor  ( new_n17003_, new_n16598_, new_n16596_ );
xor  ( new_n17004_, new_n17003_, new_n16602_ );
xor  ( new_n17005_, new_n16620_, new_n16610_ );
xor  ( new_n17006_, new_n17005_, new_n16632_ );
and  ( new_n17007_, new_n1474_, RIbb31578_128 );
or   ( new_n17008_, new_n17007_, new_n1358_ );
nand ( new_n17009_, new_n17007_, new_n1355_ );
and  ( new_n17010_, new_n17009_, new_n17008_ );
xnor ( new_n17011_, new_n16820_, new_n16816_ );
xor  ( new_n17012_, new_n17011_, new_n16826_ );
nor  ( new_n17013_, new_n17012_, new_n17010_ );
nand ( new_n17014_, new_n17012_, new_n17010_ );
xor  ( new_n17015_, new_n16910_, new_n16906_ );
xnor ( new_n17016_, new_n17015_, new_n16916_ );
not  ( new_n17017_, new_n17016_ );
and  ( new_n17018_, new_n17017_, new_n17014_ );
or   ( new_n17019_, new_n17018_, new_n17013_ );
or   ( new_n17020_, new_n8874_, new_n2751_ );
or   ( new_n17021_, new_n8876_, new_n2646_ );
and  ( new_n17022_, new_n17021_, new_n17020_ );
xor  ( new_n17023_, new_n17022_, new_n8257_ );
or   ( new_n17024_, new_n8264_, new_n3178_ );
or   ( new_n17025_, new_n8266_, new_n2981_ );
and  ( new_n17026_, new_n17025_, new_n17024_ );
xor  ( new_n17027_, new_n17026_, new_n7725_ );
or   ( new_n17028_, new_n17027_, new_n17023_ );
and  ( new_n17029_, new_n17027_, new_n17023_ );
or   ( new_n17030_, new_n7732_, new_n3696_ );
or   ( new_n17031_, new_n7734_, new_n3306_ );
and  ( new_n17032_, new_n17031_, new_n17030_ );
xor  ( new_n17033_, new_n17032_, new_n7177_ );
or   ( new_n17034_, new_n17033_, new_n17029_ );
and  ( new_n17035_, new_n17034_, new_n17028_ );
or   ( new_n17036_, new_n10059_, new_n2178_ );
or   ( new_n17037_, new_n10061_, new_n2057_ );
and  ( new_n17038_, new_n17037_, new_n17036_ );
xor  ( new_n17039_, new_n17038_, new_n9421_ );
and  ( new_n17040_, RIbb2d888_64, RIbb2ccd0_89 );
or   ( new_n17041_, RIbb2d888_64, new_n1899_ );
and  ( new_n17042_, new_n17041_, RIbb2d900_63 );
or   ( new_n17043_, new_n17042_, new_n17040_ );
or   ( new_n17044_, new_n10770_, new_n1754_ );
and  ( new_n17045_, new_n17044_, new_n17043_ );
or   ( new_n17046_, new_n17045_, new_n17039_ );
and  ( new_n17047_, new_n17045_, new_n17039_ );
or   ( new_n17048_, new_n9422_, new_n2475_ );
or   ( new_n17049_, new_n9424_, new_n2291_ );
and  ( new_n17050_, new_n17049_, new_n17048_ );
xor  ( new_n17051_, new_n17050_, new_n8873_ );
or   ( new_n17052_, new_n17051_, new_n17047_ );
and  ( new_n17053_, new_n17052_, new_n17046_ );
or   ( new_n17054_, new_n17053_, new_n17035_ );
and  ( new_n17055_, new_n17053_, new_n17035_ );
or   ( new_n17056_, new_n7184_, new_n3820_ );
or   ( new_n17057_, new_n7186_, new_n3694_ );
and  ( new_n17058_, new_n17057_, new_n17056_ );
xor  ( new_n17059_, new_n17058_, new_n6638_ );
or   ( new_n17060_, new_n6645_, new_n4267_ );
or   ( new_n17061_, new_n6647_, new_n4069_ );
and  ( new_n17062_, new_n17061_, new_n17060_ );
xor  ( new_n17063_, new_n17062_, new_n6166_ );
nor  ( new_n17064_, new_n17063_, new_n17059_ );
and  ( new_n17065_, new_n17063_, new_n17059_ );
or   ( new_n17066_, new_n6173_, new_n4995_ );
or   ( new_n17067_, new_n6175_, new_n4603_ );
and  ( new_n17068_, new_n17067_, new_n17066_ );
xor  ( new_n17069_, new_n17068_, new_n5597_ );
nor  ( new_n17070_, new_n17069_, new_n17065_ );
nor  ( new_n17071_, new_n17070_, new_n17064_ );
or   ( new_n17072_, new_n17071_, new_n17055_ );
and  ( new_n17073_, new_n17072_, new_n17054_ );
nor  ( new_n17074_, new_n17073_, new_n17019_ );
nand ( new_n17075_, new_n17073_, new_n17019_ );
or   ( new_n17076_, new_n5604_, new_n5171_ );
or   ( new_n17077_, new_n5606_, new_n4859_ );
and  ( new_n17078_, new_n17077_, new_n17076_ );
xor  ( new_n17079_, new_n17078_, new_n5206_ );
or   ( new_n17080_, new_n5207_, new_n5570_ );
or   ( new_n17081_, new_n5209_, new_n5428_ );
and  ( new_n17082_, new_n17081_, new_n17080_ );
xor  ( new_n17083_, new_n17082_, new_n4708_ );
or   ( new_n17084_, new_n17083_, new_n17079_ );
and  ( new_n17085_, new_n17083_, new_n17079_ );
or   ( new_n17086_, new_n4709_, new_n6219_ );
or   ( new_n17087_, new_n4711_, new_n5899_ );
and  ( new_n17088_, new_n17087_, new_n17086_ );
xor  ( new_n17089_, new_n17088_, new_n4295_ );
or   ( new_n17090_, new_n17089_, new_n17085_ );
and  ( new_n17091_, new_n17090_, new_n17084_ );
or   ( new_n17092_, new_n4302_, new_n6589_ );
or   ( new_n17093_, new_n4304_, new_n6425_ );
and  ( new_n17094_, new_n17093_, new_n17092_ );
xor  ( new_n17095_, new_n17094_, new_n3895_ );
or   ( new_n17096_, new_n3896_, new_n7149_ );
or   ( new_n17097_, new_n3898_, new_n6943_ );
and  ( new_n17098_, new_n17097_, new_n17096_ );
xor  ( new_n17099_, new_n17098_, new_n3460_ );
or   ( new_n17100_, new_n17099_, new_n17095_ );
and  ( new_n17101_, new_n17099_, new_n17095_ );
or   ( new_n17102_, new_n3461_, new_n8117_ );
or   ( new_n17103_, new_n3463_, new_n7373_ );
and  ( new_n17104_, new_n17103_, new_n17102_ );
xor  ( new_n17105_, new_n17104_, new_n3116_ );
or   ( new_n17106_, new_n17105_, new_n17101_ );
and  ( new_n17107_, new_n17106_, new_n17100_ );
nor  ( new_n17108_, new_n17107_, new_n17091_ );
nand ( new_n17109_, new_n17107_, new_n17091_ );
or   ( new_n17110_, new_n3117_, new_n8352_ );
or   ( new_n17111_, new_n3119_, new_n8115_ );
and  ( new_n17112_, new_n17111_, new_n17110_ );
xor  ( new_n17113_, new_n17112_, new_n2800_ );
or   ( new_n17114_, new_n2807_, new_n8995_ );
or   ( new_n17115_, new_n2809_, new_n8481_ );
and  ( new_n17116_, new_n17115_, new_n17114_ );
xor  ( new_n17117_, new_n17116_, new_n2424_ );
nor  ( new_n17118_, new_n17117_, new_n17113_ );
nand ( new_n17119_, new_n17117_, new_n17113_ );
or   ( new_n17120_, new_n2425_, new_n9681_ );
or   ( new_n17121_, new_n2427_, new_n9099_ );
and  ( new_n17122_, new_n17121_, new_n17120_ );
xor  ( new_n17123_, new_n17122_, new_n2121_ );
not  ( new_n17124_, new_n17123_ );
and  ( new_n17125_, new_n17124_, new_n17119_ );
or   ( new_n17126_, new_n17125_, new_n17118_ );
and  ( new_n17127_, new_n17126_, new_n17109_ );
or   ( new_n17128_, new_n17127_, new_n17108_ );
and  ( new_n17129_, new_n17128_, new_n17075_ );
or   ( new_n17130_, new_n17129_, new_n17074_ );
xnor ( new_n17131_, new_n16880_, new_n16864_ );
xor  ( new_n17132_, new_n17131_, new_n16850_ );
xnor ( new_n17133_, new_n16918_, new_n16902_ );
xor  ( new_n17134_, new_n17133_, new_n16936_ );
or   ( new_n17135_, new_n17134_, new_n17132_ );
and  ( new_n17136_, new_n17134_, new_n17132_ );
xor  ( new_n17137_, new_n16828_, new_n16812_ );
xor  ( new_n17138_, new_n17137_, new_n16832_ );
or   ( new_n17139_, new_n17138_, new_n17136_ );
and  ( new_n17140_, new_n17139_, new_n17135_ );
and  ( new_n17141_, new_n17140_, new_n17130_ );
or   ( new_n17142_, new_n17140_, new_n17130_ );
xor  ( new_n17143_, new_n16950_, new_n16948_ );
xor  ( new_n17144_, new_n17143_, new_n16954_ );
xnor ( new_n17145_, new_n16842_, new_n16838_ );
xor  ( new_n17146_, new_n17145_, new_n16848_ );
xnor ( new_n17147_, new_n16894_, new_n16890_ );
xor  ( new_n17148_, new_n17147_, new_n16900_ );
or   ( new_n17149_, new_n17148_, new_n17146_ );
and  ( new_n17150_, new_n17148_, new_n17146_ );
xor  ( new_n17151_, new_n16928_, new_n16924_ );
xnor ( new_n17152_, new_n17151_, new_n16934_ );
or   ( new_n17153_, new_n17152_, new_n17150_ );
and  ( new_n17154_, new_n17153_, new_n17149_ );
nor  ( new_n17155_, new_n17154_, new_n17144_ );
and  ( new_n17156_, new_n17154_, new_n17144_ );
xor  ( new_n17157_, new_n16945_, new_n16943_ );
not  ( new_n17158_, new_n17157_ );
nor  ( new_n17159_, new_n17158_, new_n17156_ );
nor  ( new_n17160_, new_n17159_, new_n17155_ );
and  ( new_n17161_, new_n17160_, new_n17142_ );
or   ( new_n17162_, new_n17161_, new_n17141_ );
or   ( new_n17163_, new_n17162_, new_n17006_ );
and  ( new_n17164_, new_n17162_, new_n17006_ );
xor  ( new_n17165_, new_n16755_, new_n16739_ );
xor  ( new_n17166_, new_n17165_, new_n16775_ );
xor  ( new_n17167_, new_n16956_, new_n16946_ );
xor  ( new_n17168_, new_n17167_, new_n16960_ );
or   ( new_n17169_, new_n17168_, new_n17166_ );
and  ( new_n17170_, new_n17168_, new_n17166_ );
xor  ( new_n17171_, new_n16968_, new_n16966_ );
xor  ( new_n17172_, new_n17171_, new_n16972_ );
or   ( new_n17173_, new_n17172_, new_n17170_ );
and  ( new_n17174_, new_n17173_, new_n17169_ );
or   ( new_n17175_, new_n17174_, new_n17164_ );
and  ( new_n17176_, new_n17175_, new_n17163_ );
and  ( new_n17177_, new_n17176_, new_n17004_ );
xor  ( new_n17178_, new_n16962_, new_n16941_ );
xor  ( new_n17179_, new_n17178_, new_n16974_ );
xor  ( new_n17180_, new_n16721_, new_n16698_ );
xor  ( new_n17181_, new_n17180_, new_n16777_ );
or   ( new_n17182_, new_n17181_, new_n17179_ );
and  ( new_n17183_, new_n17181_, new_n17179_ );
xor  ( new_n17184_, new_n16804_, new_n16802_ );
xor  ( new_n17185_, new_n17184_, new_n16808_ );
or   ( new_n17186_, new_n17185_, new_n17183_ );
and  ( new_n17187_, new_n17186_, new_n17182_ );
or   ( new_n17188_, new_n17187_, new_n17177_ );
or   ( new_n17189_, new_n17176_, new_n17004_ );
and  ( new_n17190_, new_n17189_, new_n17188_ );
or   ( new_n17191_, new_n17190_, new_n17002_ );
and  ( new_n17192_, new_n17190_, new_n17002_ );
xor  ( new_n17193_, new_n16984_, new_n16982_ );
xor  ( new_n17194_, new_n17193_, new_n16987_ );
or   ( new_n17195_, new_n17194_, new_n17192_ );
and  ( new_n17196_, new_n17195_, new_n17191_ );
nor  ( new_n17197_, new_n17196_, new_n16997_ );
xor  ( new_n17198_, new_n17190_, new_n17002_ );
xor  ( new_n17199_, new_n17198_, new_n17194_ );
xor  ( new_n17200_, new_n17176_, new_n17004_ );
xor  ( new_n17201_, new_n17200_, new_n17187_ );
xor  ( new_n17202_, new_n17140_, new_n17130_ );
xor  ( new_n17203_, new_n17202_, new_n17160_ );
xor  ( new_n17204_, new_n17168_, new_n17166_ );
xor  ( new_n17205_, new_n17204_, new_n17172_ );
or   ( new_n17206_, new_n17205_, new_n17203_ );
xnor ( new_n17207_, new_n16872_, new_n16868_ );
xor  ( new_n17208_, new_n17207_, new_n16878_ );
xnor ( new_n17209_, new_n17099_, new_n17095_ );
xor  ( new_n17210_, new_n17209_, new_n17105_ );
xnor ( new_n17211_, new_n17083_, new_n17079_ );
xor  ( new_n17212_, new_n17211_, new_n17089_ );
or   ( new_n17213_, new_n17212_, new_n17210_ );
and  ( new_n17214_, new_n17212_, new_n17210_ );
xor  ( new_n17215_, new_n17117_, new_n17113_ );
xor  ( new_n17216_, new_n17215_, new_n17124_ );
or   ( new_n17217_, new_n17216_, new_n17214_ );
and  ( new_n17218_, new_n17217_, new_n17213_ );
nor  ( new_n17219_, new_n17218_, new_n17208_ );
and  ( new_n17220_, new_n17218_, new_n17208_ );
xnor ( new_n17221_, new_n17045_, new_n17039_ );
xor  ( new_n17222_, new_n17221_, new_n17051_ );
xnor ( new_n17223_, new_n17027_, new_n17023_ );
xor  ( new_n17224_, new_n17223_, new_n17033_ );
nor  ( new_n17225_, new_n17224_, new_n17222_ );
and  ( new_n17226_, new_n17224_, new_n17222_ );
xor  ( new_n17227_, new_n17063_, new_n17059_ );
xnor ( new_n17228_, new_n17227_, new_n17069_ );
nor  ( new_n17229_, new_n17228_, new_n17226_ );
nor  ( new_n17230_, new_n17229_, new_n17225_ );
nor  ( new_n17231_, new_n17230_, new_n17220_ );
nor  ( new_n17232_, new_n17231_, new_n17219_ );
or   ( new_n17233_, new_n3461_, new_n8115_ );
or   ( new_n17234_, new_n3463_, new_n8117_ );
and  ( new_n17235_, new_n17234_, new_n17233_ );
xor  ( new_n17236_, new_n17235_, new_n3116_ );
or   ( new_n17237_, new_n3117_, new_n8481_ );
or   ( new_n17238_, new_n3119_, new_n8352_ );
and  ( new_n17239_, new_n17238_, new_n17237_ );
xor  ( new_n17240_, new_n17239_, new_n2800_ );
or   ( new_n17241_, new_n17240_, new_n17236_ );
and  ( new_n17242_, new_n17240_, new_n17236_ );
or   ( new_n17243_, new_n2807_, new_n9099_ );
or   ( new_n17244_, new_n2809_, new_n8995_ );
and  ( new_n17245_, new_n17244_, new_n17243_ );
xor  ( new_n17246_, new_n17245_, new_n2424_ );
or   ( new_n17247_, new_n17246_, new_n17242_ );
and  ( new_n17248_, new_n17247_, new_n17241_ );
or   ( new_n17249_, new_n6173_, new_n4859_ );
or   ( new_n17250_, new_n6175_, new_n4995_ );
and  ( new_n17251_, new_n17250_, new_n17249_ );
xor  ( new_n17252_, new_n17251_, new_n5597_ );
or   ( new_n17253_, new_n5604_, new_n5428_ );
or   ( new_n17254_, new_n5606_, new_n5171_ );
and  ( new_n17255_, new_n17254_, new_n17253_ );
xor  ( new_n17256_, new_n17255_, new_n5206_ );
or   ( new_n17257_, new_n17256_, new_n17252_ );
and  ( new_n17258_, new_n17256_, new_n17252_ );
or   ( new_n17259_, new_n5207_, new_n5899_ );
or   ( new_n17260_, new_n5209_, new_n5570_ );
and  ( new_n17261_, new_n17260_, new_n17259_ );
xor  ( new_n17262_, new_n17261_, new_n4708_ );
or   ( new_n17263_, new_n17262_, new_n17258_ );
and  ( new_n17264_, new_n17263_, new_n17257_ );
nor  ( new_n17265_, new_n17264_, new_n17248_ );
and  ( new_n17266_, new_n17264_, new_n17248_ );
or   ( new_n17267_, new_n4709_, new_n6425_ );
or   ( new_n17268_, new_n4711_, new_n6219_ );
and  ( new_n17269_, new_n17268_, new_n17267_ );
xor  ( new_n17270_, new_n17269_, new_n4295_ );
or   ( new_n17271_, new_n4302_, new_n6943_ );
or   ( new_n17272_, new_n4304_, new_n6589_ );
and  ( new_n17273_, new_n17272_, new_n17271_ );
xor  ( new_n17274_, new_n17273_, new_n3895_ );
nor  ( new_n17275_, new_n17274_, new_n17270_ );
and  ( new_n17276_, new_n17274_, new_n17270_ );
or   ( new_n17277_, new_n3896_, new_n7373_ );
or   ( new_n17278_, new_n3898_, new_n7149_ );
and  ( new_n17279_, new_n17278_, new_n17277_ );
xor  ( new_n17280_, new_n17279_, new_n3460_ );
nor  ( new_n17281_, new_n17280_, new_n17276_ );
nor  ( new_n17282_, new_n17281_, new_n17275_ );
nor  ( new_n17283_, new_n17282_, new_n17266_ );
nor  ( new_n17284_, new_n17283_, new_n17265_ );
or   ( new_n17285_, new_n10059_, new_n2291_ );
or   ( new_n17286_, new_n10061_, new_n2178_ );
and  ( new_n17287_, new_n17286_, new_n17285_ );
xor  ( new_n17288_, new_n17287_, new_n9421_ );
and  ( new_n17289_, RIbb2d888_64, RIbb2cc58_90 );
or   ( new_n17290_, RIbb2d888_64, new_n2057_ );
and  ( new_n17291_, new_n17290_, RIbb2d900_63 );
or   ( new_n17292_, new_n17291_, new_n17289_ );
or   ( new_n17293_, new_n10770_, new_n1899_ );
and  ( new_n17294_, new_n17293_, new_n17292_ );
or   ( new_n17295_, new_n17294_, new_n17288_ );
and  ( new_n17296_, new_n17294_, new_n17288_ );
or   ( new_n17297_, new_n17296_, new_n1585_ );
and  ( new_n17298_, new_n17297_, new_n17295_ );
or   ( new_n17299_, new_n7732_, new_n3694_ );
or   ( new_n17300_, new_n7734_, new_n3696_ );
and  ( new_n17301_, new_n17300_, new_n17299_ );
xor  ( new_n17302_, new_n17301_, new_n7177_ );
or   ( new_n17303_, new_n7184_, new_n4069_ );
or   ( new_n17304_, new_n7186_, new_n3820_ );
and  ( new_n17305_, new_n17304_, new_n17303_ );
xor  ( new_n17306_, new_n17305_, new_n6638_ );
or   ( new_n17307_, new_n17306_, new_n17302_ );
and  ( new_n17308_, new_n17306_, new_n17302_ );
or   ( new_n17309_, new_n6645_, new_n4603_ );
or   ( new_n17310_, new_n6647_, new_n4267_ );
and  ( new_n17311_, new_n17310_, new_n17309_ );
xor  ( new_n17312_, new_n17311_, new_n6166_ );
or   ( new_n17313_, new_n17312_, new_n17308_ );
and  ( new_n17314_, new_n17313_, new_n17307_ );
nor  ( new_n17315_, new_n17314_, new_n17298_ );
and  ( new_n17316_, new_n17314_, new_n17298_ );
or   ( new_n17317_, new_n9422_, new_n2646_ );
or   ( new_n17318_, new_n9424_, new_n2475_ );
and  ( new_n17319_, new_n17318_, new_n17317_ );
xor  ( new_n17320_, new_n17319_, new_n8873_ );
or   ( new_n17321_, new_n8874_, new_n2981_ );
or   ( new_n17322_, new_n8876_, new_n2751_ );
and  ( new_n17323_, new_n17322_, new_n17321_ );
xor  ( new_n17324_, new_n17323_, new_n8257_ );
nor  ( new_n17325_, new_n17324_, new_n17320_ );
and  ( new_n17326_, new_n17324_, new_n17320_ );
or   ( new_n17327_, new_n8264_, new_n3306_ );
or   ( new_n17328_, new_n8266_, new_n3178_ );
and  ( new_n17329_, new_n17328_, new_n17327_ );
xor  ( new_n17330_, new_n17329_, new_n7725_ );
nor  ( new_n17331_, new_n17330_, new_n17326_ );
nor  ( new_n17332_, new_n17331_, new_n17325_ );
nor  ( new_n17333_, new_n17332_, new_n17316_ );
nor  ( new_n17334_, new_n17333_, new_n17315_ );
and  ( new_n17335_, new_n17334_, new_n17284_ );
nor  ( new_n17336_, new_n17334_, new_n17284_ );
or   ( new_n17337_, new_n2122_, new_n10220_ );
or   ( new_n17338_, new_n2124_, new_n9679_ );
and  ( new_n17339_, new_n17338_, new_n17337_ );
xor  ( new_n17340_, new_n17339_, new_n1842_ );
or   ( new_n17341_, new_n2425_, new_n9679_ );
or   ( new_n17342_, new_n2427_, new_n9681_ );
and  ( new_n17343_, new_n17342_, new_n17341_ );
xor  ( new_n17344_, new_n17343_, new_n2121_ );
or   ( new_n17345_, new_n2122_, new_n10541_ );
or   ( new_n17346_, new_n2124_, new_n10220_ );
and  ( new_n17347_, new_n17346_, new_n17345_ );
xor  ( new_n17348_, new_n17347_, new_n1843_ );
nand ( new_n17349_, new_n17348_, new_n17344_ );
nor  ( new_n17350_, new_n17348_, new_n17344_ );
and  ( new_n17351_, new_n1739_, RIbb31578_128 );
or   ( new_n17352_, new_n17351_, new_n1586_ );
nand ( new_n17353_, new_n17351_, new_n1583_ );
and  ( new_n17354_, new_n17353_, new_n17352_ );
or   ( new_n17355_, new_n17354_, new_n17350_ );
and  ( new_n17356_, new_n17355_, new_n17349_ );
nor  ( new_n17357_, new_n17356_, new_n17340_ );
and  ( new_n17358_, new_n17356_, new_n17340_ );
not  ( new_n17359_, new_n17358_ );
or   ( new_n17360_, new_n1844_, new_n10841_ );
or   ( new_n17361_, new_n1846_, new_n10541_ );
and  ( new_n17362_, new_n17361_, new_n17360_ );
xor  ( new_n17363_, new_n17362_, new_n1586_ );
and  ( new_n17364_, new_n17363_, new_n17359_ );
nor  ( new_n17365_, new_n17364_, new_n17357_ );
nor  ( new_n17366_, new_n17365_, new_n17336_ );
nor  ( new_n17367_, new_n17366_, new_n17335_ );
and  ( new_n17368_, new_n17367_, new_n17232_ );
not  ( new_n17369_, new_n17368_ );
xor  ( new_n17370_, new_n16860_, new_n16854_ );
xor  ( new_n17371_, new_n17370_, new_n1357_ );
xnor ( new_n17372_, new_n17148_, new_n17146_ );
xor  ( new_n17373_, new_n17372_, new_n17152_ );
and  ( new_n17374_, new_n17373_, new_n17371_ );
nor  ( new_n17375_, new_n17373_, new_n17371_ );
xor  ( new_n17376_, new_n17012_, new_n17010_ );
xor  ( new_n17377_, new_n17376_, new_n17017_ );
not  ( new_n17378_, new_n17377_ );
nor  ( new_n17379_, new_n17378_, new_n17375_ );
nor  ( new_n17380_, new_n17379_, new_n17374_ );
not  ( new_n17381_, new_n17380_ );
and  ( new_n17382_, new_n17381_, new_n17369_ );
nor  ( new_n17383_, new_n17367_, new_n17232_ );
nor  ( new_n17384_, new_n17383_, new_n17382_ );
xor  ( new_n17385_, new_n17134_, new_n17132_ );
xor  ( new_n17386_, new_n17385_, new_n17138_ );
xor  ( new_n17387_, new_n17073_, new_n17019_ );
xor  ( new_n17388_, new_n17387_, new_n17128_ );
or   ( new_n17389_, new_n17388_, new_n17386_ );
nand ( new_n17390_, new_n17388_, new_n17386_ );
xor  ( new_n17391_, new_n17154_, new_n17144_ );
xor  ( new_n17392_, new_n17391_, new_n17157_ );
nand ( new_n17393_, new_n17392_, new_n17390_ );
and  ( new_n17394_, new_n17393_, new_n17389_ );
and  ( new_n17395_, new_n17394_, new_n17384_ );
xor  ( new_n17396_, new_n16884_, new_n16834_ );
xor  ( new_n17397_, new_n17396_, new_n16939_ );
or   ( new_n17398_, new_n17397_, new_n17395_ );
or   ( new_n17399_, new_n17394_, new_n17384_ );
and  ( new_n17400_, new_n17399_, new_n17398_ );
or   ( new_n17401_, new_n17400_, new_n17206_ );
and  ( new_n17402_, new_n17400_, new_n17206_ );
xor  ( new_n17403_, new_n17181_, new_n17179_ );
xor  ( new_n17404_, new_n17403_, new_n17185_ );
or   ( new_n17405_, new_n17404_, new_n17402_ );
and  ( new_n17406_, new_n17405_, new_n17401_ );
or   ( new_n17407_, new_n17406_, new_n17201_ );
and  ( new_n17408_, new_n17406_, new_n17201_ );
xnor ( new_n17409_, new_n17001_, new_n16999_ );
or   ( new_n17410_, new_n17409_, new_n17408_ );
and  ( new_n17411_, new_n17410_, new_n17407_ );
nor  ( new_n17412_, new_n17411_, new_n17199_ );
xor  ( new_n17413_, new_n17406_, new_n17201_ );
xor  ( new_n17414_, new_n17413_, new_n17409_ );
xor  ( new_n17415_, new_n17174_, new_n17006_ );
xor  ( new_n17416_, new_n17415_, new_n17162_ );
xor  ( new_n17417_, new_n17314_, new_n17298_ );
xor  ( new_n17418_, new_n17417_, new_n17332_ );
xor  ( new_n17419_, new_n17356_, new_n17340_ );
xor  ( new_n17420_, new_n17419_, new_n17363_ );
and  ( new_n17421_, new_n17420_, new_n17418_ );
nor  ( new_n17422_, new_n17420_, new_n17418_ );
xor  ( new_n17423_, new_n17264_, new_n17248_ );
xnor ( new_n17424_, new_n17423_, new_n17282_ );
nor  ( new_n17425_, new_n17424_, new_n17422_ );
nor  ( new_n17426_, new_n17425_, new_n17421_ );
or   ( new_n17427_, new_n8874_, new_n3178_ );
or   ( new_n17428_, new_n8876_, new_n2981_ );
and  ( new_n17429_, new_n17428_, new_n17427_ );
xor  ( new_n17430_, new_n17429_, new_n8257_ );
or   ( new_n17431_, new_n8264_, new_n3696_ );
or   ( new_n17432_, new_n8266_, new_n3306_ );
and  ( new_n17433_, new_n17432_, new_n17431_ );
xor  ( new_n17434_, new_n17433_, new_n7725_ );
or   ( new_n17435_, new_n17434_, new_n17430_ );
and  ( new_n17436_, new_n17434_, new_n17430_ );
or   ( new_n17437_, new_n7732_, new_n3820_ );
or   ( new_n17438_, new_n7734_, new_n3694_ );
and  ( new_n17439_, new_n17438_, new_n17437_ );
xor  ( new_n17440_, new_n17439_, new_n7177_ );
or   ( new_n17441_, new_n17440_, new_n17436_ );
and  ( new_n17442_, new_n17441_, new_n17435_ );
or   ( new_n17443_, new_n7184_, new_n4267_ );
or   ( new_n17444_, new_n7186_, new_n4069_ );
and  ( new_n17445_, new_n17444_, new_n17443_ );
xor  ( new_n17446_, new_n17445_, new_n6638_ );
or   ( new_n17447_, new_n6645_, new_n4995_ );
or   ( new_n17448_, new_n6647_, new_n4603_ );
and  ( new_n17449_, new_n17448_, new_n17447_ );
xor  ( new_n17450_, new_n17449_, new_n6166_ );
or   ( new_n17451_, new_n17450_, new_n17446_ );
and  ( new_n17452_, new_n17450_, new_n17446_ );
or   ( new_n17453_, new_n6173_, new_n5171_ );
or   ( new_n17454_, new_n6175_, new_n4859_ );
and  ( new_n17455_, new_n17454_, new_n17453_ );
xor  ( new_n17456_, new_n17455_, new_n5597_ );
or   ( new_n17457_, new_n17456_, new_n17452_ );
and  ( new_n17458_, new_n17457_, new_n17451_ );
nor  ( new_n17459_, new_n17458_, new_n17442_ );
and  ( new_n17460_, new_n17458_, new_n17442_ );
or   ( new_n17461_, new_n10059_, new_n2475_ );
or   ( new_n17462_, new_n10061_, new_n2291_ );
and  ( new_n17463_, new_n17462_, new_n17461_ );
xor  ( new_n17464_, new_n17463_, new_n9421_ );
and  ( new_n17465_, RIbb2d888_64, RIbb2cbe0_91 );
or   ( new_n17466_, RIbb2d888_64, new_n2178_ );
and  ( new_n17467_, new_n17466_, RIbb2d900_63 );
or   ( new_n17468_, new_n17467_, new_n17465_ );
or   ( new_n17469_, new_n10770_, new_n2057_ );
and  ( new_n17470_, new_n17469_, new_n17468_ );
nor  ( new_n17471_, new_n17470_, new_n17464_ );
and  ( new_n17472_, new_n17470_, new_n17464_ );
or   ( new_n17473_, new_n9422_, new_n2751_ );
or   ( new_n17474_, new_n9424_, new_n2646_ );
and  ( new_n17475_, new_n17474_, new_n17473_ );
xor  ( new_n17476_, new_n17475_, new_n8873_ );
nor  ( new_n17477_, new_n17476_, new_n17472_ );
nor  ( new_n17478_, new_n17477_, new_n17471_ );
nor  ( new_n17479_, new_n17478_, new_n17460_ );
nor  ( new_n17480_, new_n17479_, new_n17459_ );
or   ( new_n17481_, new_n5604_, new_n5570_ );
or   ( new_n17482_, new_n5606_, new_n5428_ );
and  ( new_n17483_, new_n17482_, new_n17481_ );
xor  ( new_n17484_, new_n17483_, new_n5206_ );
or   ( new_n17485_, new_n5207_, new_n6219_ );
or   ( new_n17486_, new_n5209_, new_n5899_ );
and  ( new_n17487_, new_n17486_, new_n17485_ );
xor  ( new_n17488_, new_n17487_, new_n4708_ );
or   ( new_n17489_, new_n17488_, new_n17484_ );
and  ( new_n17490_, new_n17488_, new_n17484_ );
or   ( new_n17491_, new_n4709_, new_n6589_ );
or   ( new_n17492_, new_n4711_, new_n6425_ );
and  ( new_n17493_, new_n17492_, new_n17491_ );
xor  ( new_n17494_, new_n17493_, new_n4295_ );
or   ( new_n17495_, new_n17494_, new_n17490_ );
and  ( new_n17496_, new_n17495_, new_n17489_ );
or   ( new_n17497_, new_n3117_, new_n8995_ );
or   ( new_n17498_, new_n3119_, new_n8481_ );
and  ( new_n17499_, new_n17498_, new_n17497_ );
xor  ( new_n17500_, new_n17499_, new_n2800_ );
or   ( new_n17501_, new_n2807_, new_n9681_ );
or   ( new_n17502_, new_n2809_, new_n9099_ );
and  ( new_n17503_, new_n17502_, new_n17501_ );
xor  ( new_n17504_, new_n17503_, new_n2424_ );
or   ( new_n17505_, new_n17504_, new_n17500_ );
and  ( new_n17506_, new_n17504_, new_n17500_ );
or   ( new_n17507_, new_n2425_, new_n10220_ );
or   ( new_n17508_, new_n2427_, new_n9679_ );
and  ( new_n17509_, new_n17508_, new_n17507_ );
xor  ( new_n17510_, new_n17509_, new_n2121_ );
or   ( new_n17511_, new_n17510_, new_n17506_ );
and  ( new_n17512_, new_n17511_, new_n17505_ );
nor  ( new_n17513_, new_n17512_, new_n17496_ );
and  ( new_n17514_, new_n17512_, new_n17496_ );
or   ( new_n17515_, new_n4302_, new_n7149_ );
or   ( new_n17516_, new_n4304_, new_n6943_ );
and  ( new_n17517_, new_n17516_, new_n17515_ );
xor  ( new_n17518_, new_n17517_, new_n3895_ );
or   ( new_n17519_, new_n3896_, new_n8117_ );
or   ( new_n17520_, new_n3898_, new_n7373_ );
and  ( new_n17521_, new_n17520_, new_n17519_ );
xor  ( new_n17522_, new_n17521_, new_n3460_ );
nor  ( new_n17523_, new_n17522_, new_n17518_ );
and  ( new_n17524_, new_n17522_, new_n17518_ );
or   ( new_n17525_, new_n3461_, new_n8352_ );
or   ( new_n17526_, new_n3463_, new_n8115_ );
and  ( new_n17527_, new_n17526_, new_n17525_ );
xor  ( new_n17528_, new_n17527_, new_n3116_ );
nor  ( new_n17529_, new_n17528_, new_n17524_ );
nor  ( new_n17530_, new_n17529_, new_n17523_ );
nor  ( new_n17531_, new_n17530_, new_n17514_ );
nor  ( new_n17532_, new_n17531_, new_n17513_ );
and  ( new_n17533_, new_n17532_, new_n17480_ );
nor  ( new_n17534_, new_n17532_, new_n17480_ );
xor  ( new_n17535_, new_n17348_, new_n17344_ );
xor  ( new_n17536_, new_n17535_, new_n17354_ );
xnor ( new_n17537_, new_n17240_, new_n17236_ );
xor  ( new_n17538_, new_n17537_, new_n17246_ );
nor  ( new_n17539_, new_n17538_, new_n17536_ );
and  ( new_n17540_, new_n17538_, new_n17536_ );
xor  ( new_n17541_, new_n17274_, new_n17270_ );
xnor ( new_n17542_, new_n17541_, new_n17280_ );
nor  ( new_n17543_, new_n17542_, new_n17540_ );
nor  ( new_n17544_, new_n17543_, new_n17539_ );
nor  ( new_n17545_, new_n17544_, new_n17534_ );
nor  ( new_n17546_, new_n17545_, new_n17533_ );
and  ( new_n17547_, new_n17546_, new_n17426_ );
not  ( new_n17548_, new_n17547_ );
xor  ( new_n17549_, new_n17224_, new_n17222_ );
xor  ( new_n17550_, new_n17549_, new_n17228_ );
xnor ( new_n17551_, new_n17256_, new_n17252_ );
xor  ( new_n17552_, new_n17551_, new_n17262_ );
xnor ( new_n17553_, new_n17306_, new_n17302_ );
xor  ( new_n17554_, new_n17553_, new_n17312_ );
or   ( new_n17555_, new_n17554_, new_n17552_ );
and  ( new_n17556_, new_n17554_, new_n17552_ );
xnor ( new_n17557_, new_n17324_, new_n17320_ );
xor  ( new_n17558_, new_n17557_, new_n17330_ );
or   ( new_n17559_, new_n17558_, new_n17556_ );
and  ( new_n17560_, new_n17559_, new_n17555_ );
nor  ( new_n17561_, new_n17560_, new_n17550_ );
and  ( new_n17562_, new_n17560_, new_n17550_ );
xor  ( new_n17563_, new_n17212_, new_n17210_ );
xnor ( new_n17564_, new_n17563_, new_n17216_ );
not  ( new_n17565_, new_n17564_ );
nor  ( new_n17566_, new_n17565_, new_n17562_ );
nor  ( new_n17567_, new_n17566_, new_n17561_ );
not  ( new_n17568_, new_n17567_ );
and  ( new_n17569_, new_n17568_, new_n17548_ );
nor  ( new_n17570_, new_n17546_, new_n17426_ );
or   ( new_n17571_, new_n17570_, new_n17569_ );
xor  ( new_n17572_, new_n17388_, new_n17386_ );
xor  ( new_n17573_, new_n17572_, new_n17392_ );
or   ( new_n17574_, new_n17573_, new_n17571_ );
nand ( new_n17575_, new_n17573_, new_n17571_ );
xnor ( new_n17576_, new_n17053_, new_n17035_ );
xor  ( new_n17577_, new_n17576_, new_n17071_ );
xor  ( new_n17578_, new_n17107_, new_n17091_ );
xor  ( new_n17579_, new_n17578_, new_n17126_ );
nor  ( new_n17580_, new_n17579_, new_n17577_ );
and  ( new_n17581_, new_n17579_, new_n17577_ );
xor  ( new_n17582_, new_n17373_, new_n17371_ );
xor  ( new_n17583_, new_n17582_, new_n17377_ );
not  ( new_n17584_, new_n17583_ );
nor  ( new_n17585_, new_n17584_, new_n17581_ );
nor  ( new_n17586_, new_n17585_, new_n17580_ );
nand ( new_n17587_, new_n17586_, new_n17575_ );
and  ( new_n17588_, new_n17587_, new_n17574_ );
xnor ( new_n17589_, new_n17394_, new_n17384_ );
xor  ( new_n17590_, new_n17589_, new_n17397_ );
nand ( new_n17591_, new_n17590_, new_n17588_ );
nor  ( new_n17592_, new_n17590_, new_n17588_ );
xnor ( new_n17593_, new_n17205_, new_n17203_ );
or   ( new_n17594_, new_n17593_, new_n17592_ );
and  ( new_n17595_, new_n17594_, new_n17591_ );
or   ( new_n17596_, new_n17595_, new_n17416_ );
and  ( new_n17597_, new_n17595_, new_n17416_ );
xor  ( new_n17598_, new_n17400_, new_n17206_ );
xor  ( new_n17599_, new_n17598_, new_n17404_ );
or   ( new_n17600_, new_n17599_, new_n17597_ );
and  ( new_n17601_, new_n17600_, new_n17596_ );
nor  ( new_n17602_, new_n17601_, new_n17414_ );
xor  ( new_n17603_, new_n17546_, new_n17426_ );
or   ( new_n17604_, new_n17603_, new_n17568_ );
not  ( new_n17605_, new_n17569_ );
or   ( new_n17606_, new_n17570_, new_n17605_ );
and  ( new_n17607_, new_n17606_, new_n17604_ );
xnor ( new_n17608_, new_n17334_, new_n17284_ );
xor  ( new_n17609_, new_n17608_, new_n17365_ );
nand ( new_n17610_, new_n17609_, new_n17607_ );
nor  ( new_n17611_, new_n17609_, new_n17607_ );
xor  ( new_n17612_, new_n17579_, new_n17577_ );
xor  ( new_n17613_, new_n17612_, new_n17584_ );
or   ( new_n17614_, new_n17613_, new_n17611_ );
and  ( new_n17615_, new_n17614_, new_n17610_ );
or   ( new_n17616_, new_n2122_, new_n10841_ );
or   ( new_n17617_, new_n2124_, new_n10541_ );
and  ( new_n17618_, new_n17617_, new_n17616_ );
xor  ( new_n17619_, new_n17618_, new_n1842_ );
xnor ( new_n17620_, new_n17504_, new_n17500_ );
xor  ( new_n17621_, new_n17620_, new_n17510_ );
nand ( new_n17622_, new_n17621_, new_n17619_ );
or   ( new_n17623_, new_n17621_, new_n17619_ );
xor  ( new_n17624_, new_n17522_, new_n17518_ );
xnor ( new_n17625_, new_n17624_, new_n17528_ );
nand ( new_n17626_, new_n17625_, new_n17623_ );
and  ( new_n17627_, new_n17626_, new_n17622_ );
or   ( new_n17628_, new_n7732_, new_n4069_ );
or   ( new_n17629_, new_n7734_, new_n3820_ );
and  ( new_n17630_, new_n17629_, new_n17628_ );
xor  ( new_n17631_, new_n17630_, new_n7177_ );
or   ( new_n17632_, new_n7184_, new_n4603_ );
or   ( new_n17633_, new_n7186_, new_n4267_ );
and  ( new_n17634_, new_n17633_, new_n17632_ );
xor  ( new_n17635_, new_n17634_, new_n6638_ );
nor  ( new_n17636_, new_n17635_, new_n17631_ );
and  ( new_n17637_, new_n17635_, new_n17631_ );
or   ( new_n17638_, new_n6645_, new_n4859_ );
or   ( new_n17639_, new_n6647_, new_n4995_ );
and  ( new_n17640_, new_n17639_, new_n17638_ );
xor  ( new_n17641_, new_n17640_, new_n6166_ );
nor  ( new_n17642_, new_n17641_, new_n17637_ );
nor  ( new_n17643_, new_n17642_, new_n17636_ );
or   ( new_n17644_, new_n10059_, new_n2646_ );
or   ( new_n17645_, new_n10061_, new_n2475_ );
and  ( new_n17646_, new_n17645_, new_n17644_ );
xor  ( new_n17647_, new_n17646_, new_n9421_ );
and  ( new_n17648_, RIbb2d888_64, RIbb2cb68_92 );
or   ( new_n17649_, RIbb2d888_64, new_n2291_ );
and  ( new_n17650_, new_n17649_, RIbb2d900_63 );
or   ( new_n17651_, new_n17650_, new_n17648_ );
or   ( new_n17652_, new_n10770_, new_n2178_ );
and  ( new_n17653_, new_n17652_, new_n17651_ );
nor  ( new_n17654_, new_n17653_, new_n17647_ );
and  ( new_n17655_, new_n17653_, new_n17647_ );
nor  ( new_n17656_, new_n17655_, new_n1842_ );
nor  ( new_n17657_, new_n17656_, new_n17654_ );
or   ( new_n17658_, new_n9422_, new_n2981_ );
or   ( new_n17659_, new_n9424_, new_n2751_ );
and  ( new_n17660_, new_n17659_, new_n17658_ );
xor  ( new_n17661_, new_n17660_, new_n8873_ );
or   ( new_n17662_, new_n8874_, new_n3306_ );
or   ( new_n17663_, new_n8876_, new_n3178_ );
and  ( new_n17664_, new_n17663_, new_n17662_ );
xor  ( new_n17665_, new_n17664_, new_n8257_ );
or   ( new_n17666_, new_n17665_, new_n17661_ );
and  ( new_n17667_, new_n17665_, new_n17661_ );
or   ( new_n17668_, new_n8264_, new_n3694_ );
or   ( new_n17669_, new_n8266_, new_n3696_ );
and  ( new_n17670_, new_n17669_, new_n17668_ );
xor  ( new_n17671_, new_n17670_, new_n7725_ );
or   ( new_n17672_, new_n17671_, new_n17667_ );
and  ( new_n17673_, new_n17672_, new_n17666_ );
and  ( new_n17674_, new_n17673_, new_n17657_ );
or   ( new_n17675_, new_n17674_, new_n17643_ );
or   ( new_n17676_, new_n17673_, new_n17657_ );
and  ( new_n17677_, new_n17676_, new_n17675_ );
nor  ( new_n17678_, new_n17677_, new_n17627_ );
nand ( new_n17679_, new_n17677_, new_n17627_ );
or   ( new_n17680_, new_n6173_, new_n5428_ );
or   ( new_n17681_, new_n6175_, new_n5171_ );
and  ( new_n17682_, new_n17681_, new_n17680_ );
xor  ( new_n17683_, new_n17682_, new_n5597_ );
or   ( new_n17684_, new_n5604_, new_n5899_ );
or   ( new_n17685_, new_n5606_, new_n5570_ );
and  ( new_n17686_, new_n17685_, new_n17684_ );
xor  ( new_n17687_, new_n17686_, new_n5206_ );
or   ( new_n17688_, new_n17687_, new_n17683_ );
and  ( new_n17689_, new_n17687_, new_n17683_ );
or   ( new_n17690_, new_n5207_, new_n6425_ );
or   ( new_n17691_, new_n5209_, new_n6219_ );
and  ( new_n17692_, new_n17691_, new_n17690_ );
xor  ( new_n17693_, new_n17692_, new_n4708_ );
or   ( new_n17694_, new_n17693_, new_n17689_ );
and  ( new_n17695_, new_n17694_, new_n17688_ );
or   ( new_n17696_, new_n3461_, new_n8481_ );
or   ( new_n17697_, new_n3463_, new_n8352_ );
and  ( new_n17698_, new_n17697_, new_n17696_ );
xor  ( new_n17699_, new_n17698_, new_n3116_ );
or   ( new_n17700_, new_n3117_, new_n9099_ );
or   ( new_n17701_, new_n3119_, new_n8995_ );
and  ( new_n17702_, new_n17701_, new_n17700_ );
xor  ( new_n17703_, new_n17702_, new_n2800_ );
or   ( new_n17704_, new_n17703_, new_n17699_ );
and  ( new_n17705_, new_n17703_, new_n17699_ );
or   ( new_n17706_, new_n2807_, new_n9679_ );
or   ( new_n17707_, new_n2809_, new_n9681_ );
and  ( new_n17708_, new_n17707_, new_n17706_ );
xor  ( new_n17709_, new_n17708_, new_n2424_ );
or   ( new_n17710_, new_n17709_, new_n17705_ );
and  ( new_n17711_, new_n17710_, new_n17704_ );
nor  ( new_n17712_, new_n17711_, new_n17695_ );
and  ( new_n17713_, new_n17711_, new_n17695_ );
or   ( new_n17714_, new_n4709_, new_n6943_ );
or   ( new_n17715_, new_n4711_, new_n6589_ );
and  ( new_n17716_, new_n17715_, new_n17714_ );
xor  ( new_n17717_, new_n17716_, new_n4295_ );
or   ( new_n17718_, new_n4302_, new_n7373_ );
or   ( new_n17719_, new_n4304_, new_n7149_ );
and  ( new_n17720_, new_n17719_, new_n17718_ );
xor  ( new_n17721_, new_n17720_, new_n3895_ );
nor  ( new_n17722_, new_n17721_, new_n17717_ );
and  ( new_n17723_, new_n17721_, new_n17717_ );
or   ( new_n17724_, new_n3896_, new_n8115_ );
or   ( new_n17725_, new_n3898_, new_n8117_ );
and  ( new_n17726_, new_n17725_, new_n17724_ );
xor  ( new_n17727_, new_n17726_, new_n3460_ );
nor  ( new_n17728_, new_n17727_, new_n17723_ );
nor  ( new_n17729_, new_n17728_, new_n17722_ );
nor  ( new_n17730_, new_n17729_, new_n17713_ );
or   ( new_n17731_, new_n17730_, new_n17712_ );
and  ( new_n17732_, new_n17731_, new_n17679_ );
or   ( new_n17733_, new_n17732_, new_n17678_ );
xor  ( new_n17734_, new_n17294_, new_n17288_ );
xor  ( new_n17735_, new_n17734_, new_n1586_ );
xnor ( new_n17736_, new_n17450_, new_n17446_ );
xor  ( new_n17737_, new_n17736_, new_n17456_ );
xnor ( new_n17738_, new_n17488_, new_n17484_ );
xor  ( new_n17739_, new_n17738_, new_n17494_ );
or   ( new_n17740_, new_n17739_, new_n17737_ );
and  ( new_n17741_, new_n17739_, new_n17737_ );
xor  ( new_n17742_, new_n17434_, new_n17430_ );
xnor ( new_n17743_, new_n17742_, new_n17440_ );
or   ( new_n17744_, new_n17743_, new_n17741_ );
and  ( new_n17745_, new_n17744_, new_n17740_ );
or   ( new_n17746_, new_n17745_, new_n17735_ );
and  ( new_n17747_, new_n17745_, new_n17735_ );
xor  ( new_n17748_, new_n17554_, new_n17552_ );
xor  ( new_n17749_, new_n17748_, new_n17558_ );
or   ( new_n17750_, new_n17749_, new_n17747_ );
and  ( new_n17751_, new_n17750_, new_n17746_ );
and  ( new_n17752_, new_n17751_, new_n17733_ );
or   ( new_n17753_, new_n17751_, new_n17733_ );
xnor ( new_n17754_, new_n17512_, new_n17496_ );
xor  ( new_n17755_, new_n17754_, new_n17530_ );
xnor ( new_n17756_, new_n17458_, new_n17442_ );
xor  ( new_n17757_, new_n17756_, new_n17478_ );
or   ( new_n17758_, new_n17757_, new_n17755_ );
and  ( new_n17759_, new_n17757_, new_n17755_ );
xor  ( new_n17760_, new_n17538_, new_n17536_ );
xnor ( new_n17761_, new_n17760_, new_n17542_ );
not  ( new_n17762_, new_n17761_ );
or   ( new_n17763_, new_n17762_, new_n17759_ );
and  ( new_n17764_, new_n17763_, new_n17758_ );
and  ( new_n17765_, new_n17764_, new_n17753_ );
or   ( new_n17766_, new_n17765_, new_n17752_ );
xnor ( new_n17767_, new_n17532_, new_n17480_ );
xor  ( new_n17768_, new_n17767_, new_n17544_ );
xnor ( new_n17769_, new_n17420_, new_n17418_ );
xor  ( new_n17770_, new_n17769_, new_n17424_ );
nand ( new_n17771_, new_n17770_, new_n17768_ );
nor  ( new_n17772_, new_n17770_, new_n17768_ );
xor  ( new_n17773_, new_n17560_, new_n17550_ );
xor  ( new_n17774_, new_n17773_, new_n17565_ );
or   ( new_n17775_, new_n17774_, new_n17772_ );
and  ( new_n17776_, new_n17775_, new_n17771_ );
or   ( new_n17777_, new_n17776_, new_n17766_ );
and  ( new_n17778_, new_n17776_, new_n17766_ );
xor  ( new_n17779_, new_n17218_, new_n17208_ );
xor  ( new_n17780_, new_n17779_, new_n17230_ );
or   ( new_n17781_, new_n17780_, new_n17778_ );
and  ( new_n17782_, new_n17781_, new_n17777_ );
nor  ( new_n17783_, new_n17782_, new_n17615_ );
and  ( new_n17784_, new_n17782_, new_n17615_ );
xor  ( new_n17785_, new_n17367_, new_n17232_ );
nor  ( new_n17786_, new_n17785_, new_n17381_ );
not  ( new_n17787_, new_n17383_ );
and  ( new_n17788_, new_n17787_, new_n17382_ );
nor  ( new_n17789_, new_n17788_, new_n17786_ );
not  ( new_n17790_, new_n17789_ );
nor  ( new_n17791_, new_n17790_, new_n17784_ );
nor  ( new_n17792_, new_n17791_, new_n17783_ );
xor  ( new_n17793_, new_n17590_, new_n17588_ );
xor  ( new_n17794_, new_n17793_, new_n17593_ );
or   ( new_n17795_, new_n17794_, new_n17792_ );
xor  ( new_n17796_, new_n17595_, new_n17416_ );
xor  ( new_n17797_, new_n17796_, new_n17599_ );
nor  ( new_n17798_, new_n17797_, new_n17795_ );
xnor ( new_n17799_, new_n17794_, new_n17792_ );
xor  ( new_n17800_, new_n17782_, new_n17615_ );
xor  ( new_n17801_, new_n17800_, new_n17790_ );
xnor ( new_n17802_, new_n17770_, new_n17768_ );
xor  ( new_n17803_, new_n17802_, new_n17774_ );
or   ( new_n17804_, new_n8874_, new_n3696_ );
or   ( new_n17805_, new_n8876_, new_n3306_ );
and  ( new_n17806_, new_n17805_, new_n17804_ );
xor  ( new_n17807_, new_n17806_, new_n8257_ );
or   ( new_n17808_, new_n8264_, new_n3820_ );
or   ( new_n17809_, new_n8266_, new_n3694_ );
and  ( new_n17810_, new_n17809_, new_n17808_ );
xor  ( new_n17811_, new_n17810_, new_n7725_ );
or   ( new_n17812_, new_n17811_, new_n17807_ );
and  ( new_n17813_, new_n17811_, new_n17807_ );
or   ( new_n17814_, new_n7732_, new_n4267_ );
or   ( new_n17815_, new_n7734_, new_n4069_ );
and  ( new_n17816_, new_n17815_, new_n17814_ );
xor  ( new_n17817_, new_n17816_, new_n7177_ );
or   ( new_n17818_, new_n17817_, new_n17813_ );
and  ( new_n17819_, new_n17818_, new_n17812_ );
or   ( new_n17820_, new_n10059_, new_n2751_ );
or   ( new_n17821_, new_n10061_, new_n2646_ );
and  ( new_n17822_, new_n17821_, new_n17820_ );
xor  ( new_n17823_, new_n17822_, new_n9421_ );
and  ( new_n17824_, RIbb2d888_64, RIbb2caf0_93 );
or   ( new_n17825_, RIbb2d888_64, new_n2475_ );
and  ( new_n17826_, new_n17825_, RIbb2d900_63 );
or   ( new_n17827_, new_n17826_, new_n17824_ );
or   ( new_n17828_, new_n10770_, new_n2291_ );
and  ( new_n17829_, new_n17828_, new_n17827_ );
or   ( new_n17830_, new_n17829_, new_n17823_ );
and  ( new_n17831_, new_n17829_, new_n17823_ );
or   ( new_n17832_, new_n9422_, new_n3178_ );
or   ( new_n17833_, new_n9424_, new_n2981_ );
and  ( new_n17834_, new_n17833_, new_n17832_ );
xor  ( new_n17835_, new_n17834_, new_n8873_ );
or   ( new_n17836_, new_n17835_, new_n17831_ );
and  ( new_n17837_, new_n17836_, new_n17830_ );
or   ( new_n17838_, new_n17837_, new_n17819_ );
and  ( new_n17839_, new_n17837_, new_n17819_ );
or   ( new_n17840_, new_n7184_, new_n4995_ );
or   ( new_n17841_, new_n7186_, new_n4603_ );
and  ( new_n17842_, new_n17841_, new_n17840_ );
xor  ( new_n17843_, new_n17842_, new_n6638_ );
or   ( new_n17844_, new_n6645_, new_n5171_ );
or   ( new_n17845_, new_n6647_, new_n4859_ );
and  ( new_n17846_, new_n17845_, new_n17844_ );
xor  ( new_n17847_, new_n17846_, new_n6166_ );
nor  ( new_n17848_, new_n17847_, new_n17843_ );
and  ( new_n17849_, new_n17847_, new_n17843_ );
or   ( new_n17850_, new_n6173_, new_n5570_ );
or   ( new_n17851_, new_n6175_, new_n5428_ );
and  ( new_n17852_, new_n17851_, new_n17850_ );
xor  ( new_n17853_, new_n17852_, new_n5597_ );
nor  ( new_n17854_, new_n17853_, new_n17849_ );
nor  ( new_n17855_, new_n17854_, new_n17848_ );
or   ( new_n17856_, new_n17855_, new_n17839_ );
and  ( new_n17857_, new_n17856_, new_n17838_ );
or   ( new_n17858_, new_n2425_, new_n10541_ );
or   ( new_n17859_, new_n2427_, new_n10220_ );
and  ( new_n17860_, new_n17859_, new_n17858_ );
xor  ( new_n17861_, new_n17860_, new_n2120_ );
and  ( new_n17862_, new_n2000_, RIbb31578_128 );
or   ( new_n17863_, new_n17862_, new_n1843_ );
nand ( new_n17864_, new_n17862_, new_n1840_ );
and  ( new_n17865_, new_n17864_, new_n17863_ );
nand ( new_n17866_, new_n17865_, new_n17861_ );
or   ( new_n17867_, new_n17865_, new_n17861_ );
xor  ( new_n17868_, new_n17703_, new_n17699_ );
xnor ( new_n17869_, new_n17868_, new_n17709_ );
nand ( new_n17870_, new_n17869_, new_n17867_ );
and  ( new_n17871_, new_n17870_, new_n17866_ );
nor  ( new_n17872_, new_n17871_, new_n17857_ );
nand ( new_n17873_, new_n17871_, new_n17857_ );
or   ( new_n17874_, new_n4302_, new_n8117_ );
or   ( new_n17875_, new_n4304_, new_n7373_ );
and  ( new_n17876_, new_n17875_, new_n17874_ );
xor  ( new_n17877_, new_n17876_, new_n3895_ );
or   ( new_n17878_, new_n3896_, new_n8352_ );
or   ( new_n17879_, new_n3898_, new_n8115_ );
and  ( new_n17880_, new_n17879_, new_n17878_ );
xor  ( new_n17881_, new_n17880_, new_n3460_ );
or   ( new_n17882_, new_n17881_, new_n17877_ );
and  ( new_n17883_, new_n17881_, new_n17877_ );
or   ( new_n17884_, new_n3461_, new_n8995_ );
or   ( new_n17885_, new_n3463_, new_n8481_ );
and  ( new_n17886_, new_n17885_, new_n17884_ );
xor  ( new_n17887_, new_n17886_, new_n3116_ );
or   ( new_n17888_, new_n17887_, new_n17883_ );
and  ( new_n17889_, new_n17888_, new_n17882_ );
or   ( new_n17890_, new_n3117_, new_n9681_ );
or   ( new_n17891_, new_n3119_, new_n9099_ );
and  ( new_n17892_, new_n17891_, new_n17890_ );
xor  ( new_n17893_, new_n17892_, new_n2800_ );
or   ( new_n17894_, new_n2807_, new_n10220_ );
or   ( new_n17895_, new_n2809_, new_n9679_ );
and  ( new_n17896_, new_n17895_, new_n17894_ );
xor  ( new_n17897_, new_n17896_, new_n2424_ );
or   ( new_n17898_, new_n17897_, new_n17893_ );
and  ( new_n17899_, new_n17897_, new_n17893_ );
or   ( new_n17900_, new_n2425_, new_n10841_ );
or   ( new_n17901_, new_n2427_, new_n10541_ );
and  ( new_n17902_, new_n17901_, new_n17900_ );
xor  ( new_n17903_, new_n17902_, new_n2121_ );
or   ( new_n17904_, new_n17903_, new_n17899_ );
and  ( new_n17905_, new_n17904_, new_n17898_ );
nor  ( new_n17906_, new_n17905_, new_n17889_ );
nand ( new_n17907_, new_n17905_, new_n17889_ );
or   ( new_n17908_, new_n5604_, new_n6219_ );
or   ( new_n17909_, new_n5606_, new_n5899_ );
and  ( new_n17910_, new_n17909_, new_n17908_ );
xor  ( new_n17911_, new_n17910_, new_n5206_ );
or   ( new_n17912_, new_n5207_, new_n6589_ );
or   ( new_n17913_, new_n5209_, new_n6425_ );
and  ( new_n17914_, new_n17913_, new_n17912_ );
xor  ( new_n17915_, new_n17914_, new_n4708_ );
nor  ( new_n17916_, new_n17915_, new_n17911_ );
nand ( new_n17917_, new_n17915_, new_n17911_ );
or   ( new_n17918_, new_n4709_, new_n7149_ );
or   ( new_n17919_, new_n4711_, new_n6943_ );
and  ( new_n17920_, new_n17919_, new_n17918_ );
xor  ( new_n17921_, new_n17920_, new_n4295_ );
not  ( new_n17922_, new_n17921_ );
and  ( new_n17923_, new_n17922_, new_n17917_ );
or   ( new_n17924_, new_n17923_, new_n17916_ );
and  ( new_n17925_, new_n17924_, new_n17907_ );
or   ( new_n17926_, new_n17925_, new_n17906_ );
and  ( new_n17927_, new_n17926_, new_n17873_ );
or   ( new_n17928_, new_n17927_, new_n17872_ );
xor  ( new_n17929_, new_n17665_, new_n17661_ );
xnor ( new_n17930_, new_n17929_, new_n17671_ );
xor  ( new_n17931_, new_n17653_, new_n17647_ );
xor  ( new_n17932_, new_n17931_, new_n1843_ );
or   ( new_n17933_, new_n17932_, new_n17930_ );
xnor ( new_n17934_, new_n17635_, new_n17631_ );
xor  ( new_n17935_, new_n17934_, new_n17641_ );
xnor ( new_n17936_, new_n17687_, new_n17683_ );
xor  ( new_n17937_, new_n17936_, new_n17693_ );
or   ( new_n17938_, new_n17937_, new_n17935_ );
and  ( new_n17939_, new_n17937_, new_n17935_ );
xnor ( new_n17940_, new_n17721_, new_n17717_ );
xor  ( new_n17941_, new_n17940_, new_n17727_ );
or   ( new_n17942_, new_n17941_, new_n17939_ );
and  ( new_n17943_, new_n17942_, new_n17938_ );
or   ( new_n17944_, new_n17943_, new_n17933_ );
and  ( new_n17945_, new_n17943_, new_n17933_ );
xor  ( new_n17946_, new_n17470_, new_n17464_ );
xnor ( new_n17947_, new_n17946_, new_n17476_ );
or   ( new_n17948_, new_n17947_, new_n17945_ );
and  ( new_n17949_, new_n17948_, new_n17944_ );
nand ( new_n17950_, new_n17949_, new_n17928_ );
or   ( new_n17951_, new_n17949_, new_n17928_ );
xor  ( new_n17952_, new_n17711_, new_n17695_ );
xor  ( new_n17953_, new_n17952_, new_n17729_ );
xnor ( new_n17954_, new_n17739_, new_n17737_ );
xor  ( new_n17955_, new_n17954_, new_n17743_ );
and  ( new_n17956_, new_n17955_, new_n17953_ );
nor  ( new_n17957_, new_n17955_, new_n17953_ );
xor  ( new_n17958_, new_n17621_, new_n17619_ );
xor  ( new_n17959_, new_n17958_, new_n17625_ );
nor  ( new_n17960_, new_n17959_, new_n17957_ );
nor  ( new_n17961_, new_n17960_, new_n17956_ );
nand ( new_n17962_, new_n17961_, new_n17951_ );
and  ( new_n17963_, new_n17962_, new_n17950_ );
nor  ( new_n17964_, new_n17963_, new_n17803_ );
nand ( new_n17965_, new_n17963_, new_n17803_ );
xor  ( new_n17966_, new_n17745_, new_n17735_ );
xor  ( new_n17967_, new_n17966_, new_n17749_ );
xor  ( new_n17968_, new_n17677_, new_n17627_ );
xor  ( new_n17969_, new_n17968_, new_n17731_ );
nor  ( new_n17970_, new_n17969_, new_n17967_ );
and  ( new_n17971_, new_n17969_, new_n17967_ );
xor  ( new_n17972_, new_n17757_, new_n17755_ );
xor  ( new_n17973_, new_n17972_, new_n17762_ );
nor  ( new_n17974_, new_n17973_, new_n17971_ );
nor  ( new_n17975_, new_n17974_, new_n17970_ );
and  ( new_n17976_, new_n17975_, new_n17965_ );
or   ( new_n17977_, new_n17976_, new_n17964_ );
xor  ( new_n17978_, new_n17776_, new_n17766_ );
xor  ( new_n17979_, new_n17978_, new_n17780_ );
or   ( new_n17980_, new_n17979_, new_n17977_ );
and  ( new_n17981_, new_n17979_, new_n17977_ );
xor  ( new_n17982_, new_n17609_, new_n17607_ );
xor  ( new_n17983_, new_n17982_, new_n17613_ );
or   ( new_n17984_, new_n17983_, new_n17981_ );
and  ( new_n17985_, new_n17984_, new_n17980_ );
or   ( new_n17986_, new_n17985_, new_n17801_ );
and  ( new_n17987_, new_n17985_, new_n17801_ );
xor  ( new_n17988_, new_n17573_, new_n17571_ );
xor  ( new_n17989_, new_n17988_, new_n17586_ );
or   ( new_n17990_, new_n17989_, new_n17987_ );
and  ( new_n17991_, new_n17990_, new_n17986_ );
nor  ( new_n17992_, new_n17991_, new_n17799_ );
xor  ( new_n17993_, new_n17979_, new_n17977_ );
xor  ( new_n17994_, new_n17993_, new_n17983_ );
xor  ( new_n17995_, new_n17751_, new_n17733_ );
xor  ( new_n17996_, new_n17995_, new_n17764_ );
xnor ( new_n17997_, new_n17837_, new_n17819_ );
xor  ( new_n17998_, new_n17997_, new_n17855_ );
xor  ( new_n17999_, new_n17905_, new_n17889_ );
xor  ( new_n18000_, new_n17999_, new_n17924_ );
nor  ( new_n18001_, new_n18000_, new_n17998_ );
and  ( new_n18002_, new_n18000_, new_n17998_ );
xor  ( new_n18003_, new_n17865_, new_n17861_ );
xor  ( new_n18004_, new_n18003_, new_n17869_ );
nor  ( new_n18005_, new_n18004_, new_n18002_ );
nor  ( new_n18006_, new_n18005_, new_n18001_ );
or   ( new_n18007_, new_n4709_, new_n7373_ );
or   ( new_n18008_, new_n4711_, new_n7149_ );
and  ( new_n18009_, new_n18008_, new_n18007_ );
xor  ( new_n18010_, new_n18009_, new_n4295_ );
or   ( new_n18011_, new_n4302_, new_n8115_ );
or   ( new_n18012_, new_n4304_, new_n8117_ );
and  ( new_n18013_, new_n18012_, new_n18011_ );
xor  ( new_n18014_, new_n18013_, new_n3895_ );
or   ( new_n18015_, new_n18014_, new_n18010_ );
and  ( new_n18016_, new_n18014_, new_n18010_ );
or   ( new_n18017_, new_n3896_, new_n8481_ );
or   ( new_n18018_, new_n3898_, new_n8352_ );
and  ( new_n18019_, new_n18018_, new_n18017_ );
xor  ( new_n18020_, new_n18019_, new_n3460_ );
or   ( new_n18021_, new_n18020_, new_n18016_ );
and  ( new_n18022_, new_n18021_, new_n18015_ );
or   ( new_n18023_, new_n6173_, new_n5899_ );
or   ( new_n18024_, new_n6175_, new_n5570_ );
and  ( new_n18025_, new_n18024_, new_n18023_ );
xor  ( new_n18026_, new_n18025_, new_n5597_ );
or   ( new_n18027_, new_n5604_, new_n6425_ );
or   ( new_n18028_, new_n5606_, new_n6219_ );
and  ( new_n18029_, new_n18028_, new_n18027_ );
xor  ( new_n18030_, new_n18029_, new_n5206_ );
or   ( new_n18031_, new_n18030_, new_n18026_ );
and  ( new_n18032_, new_n18030_, new_n18026_ );
or   ( new_n18033_, new_n5207_, new_n6943_ );
or   ( new_n18034_, new_n5209_, new_n6589_ );
and  ( new_n18035_, new_n18034_, new_n18033_ );
xor  ( new_n18036_, new_n18035_, new_n4708_ );
or   ( new_n18037_, new_n18036_, new_n18032_ );
and  ( new_n18038_, new_n18037_, new_n18031_ );
nor  ( new_n18039_, new_n18038_, new_n18022_ );
and  ( new_n18040_, new_n18038_, new_n18022_ );
or   ( new_n18041_, new_n3461_, new_n9099_ );
or   ( new_n18042_, new_n3463_, new_n8995_ );
and  ( new_n18043_, new_n18042_, new_n18041_ );
xor  ( new_n18044_, new_n18043_, new_n3116_ );
or   ( new_n18045_, new_n3117_, new_n9679_ );
or   ( new_n18046_, new_n3119_, new_n9681_ );
and  ( new_n18047_, new_n18046_, new_n18045_ );
xor  ( new_n18048_, new_n18047_, new_n2800_ );
nor  ( new_n18049_, new_n18048_, new_n18044_ );
and  ( new_n18050_, new_n18048_, new_n18044_ );
or   ( new_n18051_, new_n2807_, new_n10541_ );
or   ( new_n18052_, new_n2809_, new_n10220_ );
and  ( new_n18053_, new_n18052_, new_n18051_ );
xor  ( new_n18054_, new_n18053_, new_n2424_ );
nor  ( new_n18055_, new_n18054_, new_n18050_ );
nor  ( new_n18056_, new_n18055_, new_n18049_ );
nor  ( new_n18057_, new_n18056_, new_n18040_ );
nor  ( new_n18058_, new_n18057_, new_n18039_ );
or   ( new_n18059_, new_n10059_, new_n2981_ );
or   ( new_n18060_, new_n10061_, new_n2751_ );
and  ( new_n18061_, new_n18060_, new_n18059_ );
xor  ( new_n18062_, new_n18061_, new_n9421_ );
and  ( new_n18063_, RIbb2d888_64, RIbb2ca78_94 );
or   ( new_n18064_, RIbb2d888_64, new_n2646_ );
and  ( new_n18065_, new_n18064_, RIbb2d900_63 );
or   ( new_n18066_, new_n18065_, new_n18063_ );
or   ( new_n18067_, new_n10770_, new_n2475_ );
and  ( new_n18068_, new_n18067_, new_n18066_ );
or   ( new_n18069_, new_n18068_, new_n18062_ );
and  ( new_n18070_, new_n18068_, new_n18062_ );
or   ( new_n18071_, new_n18070_, new_n2120_ );
and  ( new_n18072_, new_n18071_, new_n18069_ );
or   ( new_n18073_, new_n9422_, new_n3306_ );
or   ( new_n18074_, new_n9424_, new_n3178_ );
and  ( new_n18075_, new_n18074_, new_n18073_ );
xor  ( new_n18076_, new_n18075_, new_n8873_ );
or   ( new_n18077_, new_n8874_, new_n3694_ );
or   ( new_n18078_, new_n8876_, new_n3696_ );
and  ( new_n18079_, new_n18078_, new_n18077_ );
xor  ( new_n18080_, new_n18079_, new_n8257_ );
or   ( new_n18081_, new_n18080_, new_n18076_ );
and  ( new_n18082_, new_n18080_, new_n18076_ );
or   ( new_n18083_, new_n8264_, new_n4069_ );
or   ( new_n18084_, new_n8266_, new_n3820_ );
and  ( new_n18085_, new_n18084_, new_n18083_ );
xor  ( new_n18086_, new_n18085_, new_n7725_ );
or   ( new_n18087_, new_n18086_, new_n18082_ );
and  ( new_n18088_, new_n18087_, new_n18081_ );
nor  ( new_n18089_, new_n18088_, new_n18072_ );
and  ( new_n18090_, new_n18088_, new_n18072_ );
or   ( new_n18091_, new_n7732_, new_n4603_ );
or   ( new_n18092_, new_n7734_, new_n4267_ );
and  ( new_n18093_, new_n18092_, new_n18091_ );
xor  ( new_n18094_, new_n18093_, new_n7177_ );
or   ( new_n18095_, new_n7184_, new_n4859_ );
or   ( new_n18096_, new_n7186_, new_n4995_ );
and  ( new_n18097_, new_n18096_, new_n18095_ );
xor  ( new_n18098_, new_n18097_, new_n6638_ );
nor  ( new_n18099_, new_n18098_, new_n18094_ );
and  ( new_n18100_, new_n18098_, new_n18094_ );
or   ( new_n18101_, new_n6645_, new_n5428_ );
or   ( new_n18102_, new_n6647_, new_n5171_ );
and  ( new_n18103_, new_n18102_, new_n18101_ );
xor  ( new_n18104_, new_n18103_, new_n6166_ );
nor  ( new_n18105_, new_n18104_, new_n18100_ );
nor  ( new_n18106_, new_n18105_, new_n18099_ );
nor  ( new_n18107_, new_n18106_, new_n18090_ );
nor  ( new_n18108_, new_n18107_, new_n18089_ );
and  ( new_n18109_, new_n18108_, new_n18058_ );
nor  ( new_n18110_, new_n18108_, new_n18058_ );
xnor ( new_n18111_, new_n17897_, new_n17893_ );
xor  ( new_n18112_, new_n18111_, new_n17903_ );
xnor ( new_n18113_, new_n17881_, new_n17877_ );
xor  ( new_n18114_, new_n18113_, new_n17887_ );
nor  ( new_n18115_, new_n18114_, new_n18112_ );
and  ( new_n18116_, new_n18114_, new_n18112_ );
xor  ( new_n18117_, new_n17915_, new_n17911_ );
xor  ( new_n18118_, new_n18117_, new_n17922_ );
nor  ( new_n18119_, new_n18118_, new_n18116_ );
nor  ( new_n18120_, new_n18119_, new_n18115_ );
nor  ( new_n18121_, new_n18120_, new_n18110_ );
nor  ( new_n18122_, new_n18121_, new_n18109_ );
and  ( new_n18123_, new_n18122_, new_n18006_ );
xor  ( new_n18124_, new_n17937_, new_n17935_ );
xor  ( new_n18125_, new_n18124_, new_n17941_ );
xnor ( new_n18126_, new_n17829_, new_n17823_ );
xor  ( new_n18127_, new_n18126_, new_n17835_ );
xnor ( new_n18128_, new_n17811_, new_n17807_ );
xor  ( new_n18129_, new_n18128_, new_n17817_ );
or   ( new_n18130_, new_n18129_, new_n18127_ );
and  ( new_n18131_, new_n18129_, new_n18127_ );
xor  ( new_n18132_, new_n17847_, new_n17843_ );
xnor ( new_n18133_, new_n18132_, new_n17853_ );
or   ( new_n18134_, new_n18133_, new_n18131_ );
and  ( new_n18135_, new_n18134_, new_n18130_ );
nor  ( new_n18136_, new_n18135_, new_n18125_ );
and  ( new_n18137_, new_n18135_, new_n18125_ );
xor  ( new_n18138_, new_n17932_, new_n17930_ );
not  ( new_n18139_, new_n18138_ );
nor  ( new_n18140_, new_n18139_, new_n18137_ );
nor  ( new_n18141_, new_n18140_, new_n18136_ );
nor  ( new_n18142_, new_n18141_, new_n18123_ );
nor  ( new_n18143_, new_n18122_, new_n18006_ );
or   ( new_n18144_, new_n18143_, new_n18142_ );
xor  ( new_n18145_, new_n17673_, new_n17657_ );
xor  ( new_n18146_, new_n18145_, new_n17643_ );
xnor ( new_n18147_, new_n17943_, new_n17933_ );
xor  ( new_n18148_, new_n18147_, new_n17947_ );
or   ( new_n18149_, new_n18148_, new_n18146_ );
and  ( new_n18150_, new_n18148_, new_n18146_ );
xor  ( new_n18151_, new_n17955_, new_n17953_ );
xnor ( new_n18152_, new_n18151_, new_n17959_ );
or   ( new_n18153_, new_n18152_, new_n18150_ );
and  ( new_n18154_, new_n18153_, new_n18149_ );
nand ( new_n18155_, new_n18154_, new_n18144_ );
nor  ( new_n18156_, new_n18154_, new_n18144_ );
xor  ( new_n18157_, new_n17969_, new_n17967_ );
xor  ( new_n18158_, new_n18157_, new_n17973_ );
or   ( new_n18159_, new_n18158_, new_n18156_ );
and  ( new_n18160_, new_n18159_, new_n18155_ );
or   ( new_n18161_, new_n18160_, new_n17996_ );
and  ( new_n18162_, new_n18160_, new_n17996_ );
xor  ( new_n18163_, new_n17963_, new_n17803_ );
xor  ( new_n18164_, new_n18163_, new_n17975_ );
or   ( new_n18165_, new_n18164_, new_n18162_ );
and  ( new_n18166_, new_n18165_, new_n18161_ );
nor  ( new_n18167_, new_n18166_, new_n17994_ );
xnor ( new_n18168_, new_n17985_, new_n17801_ );
xor  ( new_n18169_, new_n18168_, new_n17989_ );
and  ( new_n18170_, new_n18169_, new_n18167_ );
not  ( new_n18171_, new_n18141_ );
xor  ( new_n18172_, new_n18122_, new_n18006_ );
nor  ( new_n18173_, new_n18172_, new_n18171_ );
not  ( new_n18174_, new_n18143_ );
and  ( new_n18175_, new_n18174_, new_n18142_ );
nor  ( new_n18176_, new_n18175_, new_n18173_ );
not  ( new_n18177_, new_n18176_ );
xnor ( new_n18178_, new_n18148_, new_n18146_ );
xor  ( new_n18179_, new_n18178_, new_n18152_ );
or   ( new_n18180_, new_n18179_, new_n18177_ );
xnor ( new_n18181_, new_n18108_, new_n18058_ );
xor  ( new_n18182_, new_n18181_, new_n18120_ );
xnor ( new_n18183_, new_n18000_, new_n17998_ );
xor  ( new_n18184_, new_n18183_, new_n18004_ );
nand ( new_n18185_, new_n18184_, new_n18182_ );
or   ( new_n18186_, new_n18184_, new_n18182_ );
xor  ( new_n18187_, new_n18135_, new_n18125_ );
xor  ( new_n18188_, new_n18187_, new_n18138_ );
nand ( new_n18189_, new_n18188_, new_n18186_ );
and  ( new_n18190_, new_n18189_, new_n18185_ );
xor  ( new_n18191_, new_n17871_, new_n17857_ );
xor  ( new_n18192_, new_n18191_, new_n17926_ );
or   ( new_n18193_, new_n18192_, new_n18190_ );
and  ( new_n18194_, new_n18192_, new_n18190_ );
xor  ( new_n18195_, new_n18088_, new_n18072_ );
xnor ( new_n18196_, new_n18195_, new_n18106_ );
xnor ( new_n18197_, new_n18038_, new_n18022_ );
xor  ( new_n18198_, new_n18197_, new_n18056_ );
nor  ( new_n18199_, new_n18198_, new_n18196_ );
and  ( new_n18200_, new_n2242_, RIbb31578_128 );
or   ( new_n18201_, new_n18200_, new_n2121_ );
nand ( new_n18202_, new_n18200_, new_n2118_ );
and  ( new_n18203_, new_n18202_, new_n18201_ );
xnor ( new_n18204_, new_n18048_, new_n18044_ );
xor  ( new_n18205_, new_n18204_, new_n18054_ );
nor  ( new_n18206_, new_n18205_, new_n18203_ );
nand ( new_n18207_, new_n18205_, new_n18203_ );
xor  ( new_n18208_, new_n18014_, new_n18010_ );
xnor ( new_n18209_, new_n18208_, new_n18020_ );
not  ( new_n18210_, new_n18209_ );
and  ( new_n18211_, new_n18210_, new_n18207_ );
or   ( new_n18212_, new_n18211_, new_n18206_ );
or   ( new_n18213_, new_n10059_, new_n3178_ );
or   ( new_n18214_, new_n10061_, new_n2981_ );
and  ( new_n18215_, new_n18214_, new_n18213_ );
xor  ( new_n18216_, new_n18215_, new_n9421_ );
and  ( new_n18217_, RIbb2d888_64, RIbb2ca00_95 );
or   ( new_n18218_, RIbb2d888_64, new_n2751_ );
and  ( new_n18219_, new_n18218_, RIbb2d900_63 );
or   ( new_n18220_, new_n18219_, new_n18217_ );
or   ( new_n18221_, new_n10770_, new_n2646_ );
and  ( new_n18222_, new_n18221_, new_n18220_ );
or   ( new_n18223_, new_n18222_, new_n18216_ );
and  ( new_n18224_, new_n18222_, new_n18216_ );
or   ( new_n18225_, new_n9422_, new_n3696_ );
or   ( new_n18226_, new_n9424_, new_n3306_ );
and  ( new_n18227_, new_n18226_, new_n18225_ );
xor  ( new_n18228_, new_n18227_, new_n8873_ );
or   ( new_n18229_, new_n18228_, new_n18224_ );
and  ( new_n18230_, new_n18229_, new_n18223_ );
or   ( new_n18231_, new_n7184_, new_n5171_ );
or   ( new_n18232_, new_n7186_, new_n4859_ );
and  ( new_n18233_, new_n18232_, new_n18231_ );
xor  ( new_n18234_, new_n18233_, new_n6638_ );
or   ( new_n18235_, new_n6645_, new_n5570_ );
or   ( new_n18236_, new_n6647_, new_n5428_ );
and  ( new_n18237_, new_n18236_, new_n18235_ );
xor  ( new_n18238_, new_n18237_, new_n6166_ );
or   ( new_n18239_, new_n18238_, new_n18234_ );
and  ( new_n18240_, new_n18238_, new_n18234_ );
or   ( new_n18241_, new_n6173_, new_n6219_ );
or   ( new_n18242_, new_n6175_, new_n5899_ );
and  ( new_n18243_, new_n18242_, new_n18241_ );
xor  ( new_n18244_, new_n18243_, new_n5597_ );
or   ( new_n18245_, new_n18244_, new_n18240_ );
and  ( new_n18246_, new_n18245_, new_n18239_ );
or   ( new_n18247_, new_n18246_, new_n18230_ );
and  ( new_n18248_, new_n18246_, new_n18230_ );
or   ( new_n18249_, new_n8874_, new_n3820_ );
or   ( new_n18250_, new_n8876_, new_n3694_ );
and  ( new_n18251_, new_n18250_, new_n18249_ );
xor  ( new_n18252_, new_n18251_, new_n8257_ );
or   ( new_n18253_, new_n8264_, new_n4267_ );
or   ( new_n18254_, new_n8266_, new_n4069_ );
and  ( new_n18255_, new_n18254_, new_n18253_ );
xor  ( new_n18256_, new_n18255_, new_n7725_ );
or   ( new_n18257_, new_n18256_, new_n18252_ );
and  ( new_n18258_, new_n18256_, new_n18252_ );
or   ( new_n18259_, new_n7732_, new_n4995_ );
or   ( new_n18260_, new_n7734_, new_n4603_ );
and  ( new_n18261_, new_n18260_, new_n18259_ );
xor  ( new_n18262_, new_n18261_, new_n7177_ );
or   ( new_n18263_, new_n18262_, new_n18258_ );
and  ( new_n18264_, new_n18263_, new_n18257_ );
or   ( new_n18265_, new_n18264_, new_n18248_ );
and  ( new_n18266_, new_n18265_, new_n18247_ );
or   ( new_n18267_, new_n18266_, new_n18212_ );
and  ( new_n18268_, new_n18266_, new_n18212_ );
or   ( new_n18269_, new_n4302_, new_n8352_ );
or   ( new_n18270_, new_n4304_, new_n8115_ );
and  ( new_n18271_, new_n18270_, new_n18269_ );
xor  ( new_n18272_, new_n18271_, new_n3895_ );
or   ( new_n18273_, new_n3896_, new_n8995_ );
or   ( new_n18274_, new_n3898_, new_n8481_ );
and  ( new_n18275_, new_n18274_, new_n18273_ );
xor  ( new_n18276_, new_n18275_, new_n3460_ );
nor  ( new_n18277_, new_n18276_, new_n18272_ );
and  ( new_n18278_, new_n18276_, new_n18272_ );
or   ( new_n18279_, new_n3461_, new_n9681_ );
or   ( new_n18280_, new_n3463_, new_n9099_ );
and  ( new_n18281_, new_n18280_, new_n18279_ );
xor  ( new_n18282_, new_n18281_, new_n3116_ );
nor  ( new_n18283_, new_n18282_, new_n18278_ );
nor  ( new_n18284_, new_n18283_, new_n18277_ );
or   ( new_n18285_, new_n3117_, new_n10220_ );
or   ( new_n18286_, new_n3119_, new_n9679_ );
and  ( new_n18287_, new_n18286_, new_n18285_ );
xor  ( new_n18288_, new_n18287_, new_n2800_ );
or   ( new_n18289_, new_n2807_, new_n10841_ );
or   ( new_n18290_, new_n2809_, new_n10541_ );
and  ( new_n18291_, new_n18290_, new_n18289_ );
xor  ( new_n18292_, new_n18291_, new_n2424_ );
and  ( new_n18293_, new_n18292_, new_n18288_ );
or   ( new_n18294_, new_n5604_, new_n6589_ );
or   ( new_n18295_, new_n5606_, new_n6425_ );
and  ( new_n18296_, new_n18295_, new_n18294_ );
xor  ( new_n18297_, new_n18296_, new_n5206_ );
or   ( new_n18298_, new_n5207_, new_n7149_ );
or   ( new_n18299_, new_n5209_, new_n6943_ );
and  ( new_n18300_, new_n18299_, new_n18298_ );
xor  ( new_n18301_, new_n18300_, new_n4708_ );
nor  ( new_n18302_, new_n18301_, new_n18297_ );
and  ( new_n18303_, new_n18301_, new_n18297_ );
or   ( new_n18304_, new_n4709_, new_n8117_ );
or   ( new_n18305_, new_n4711_, new_n7373_ );
and  ( new_n18306_, new_n18305_, new_n18304_ );
xor  ( new_n18307_, new_n18306_, new_n4295_ );
nor  ( new_n18308_, new_n18307_, new_n18303_ );
nor  ( new_n18309_, new_n18308_, new_n18302_ );
and  ( new_n18310_, new_n18309_, new_n18293_ );
nor  ( new_n18311_, new_n18310_, new_n18284_ );
nor  ( new_n18312_, new_n18309_, new_n18293_ );
nor  ( new_n18313_, new_n18312_, new_n18311_ );
or   ( new_n18314_, new_n18313_, new_n18268_ );
and  ( new_n18315_, new_n18314_, new_n18267_ );
and  ( new_n18316_, new_n18315_, new_n18199_ );
nor  ( new_n18317_, new_n18315_, new_n18199_ );
xor  ( new_n18318_, new_n18114_, new_n18112_ );
xor  ( new_n18319_, new_n18318_, new_n18118_ );
xnor ( new_n18320_, new_n18080_, new_n18076_ );
xor  ( new_n18321_, new_n18320_, new_n18086_ );
xnor ( new_n18322_, new_n18030_, new_n18026_ );
xor  ( new_n18323_, new_n18322_, new_n18036_ );
or   ( new_n18324_, new_n18323_, new_n18321_ );
and  ( new_n18325_, new_n18323_, new_n18321_ );
xor  ( new_n18326_, new_n18098_, new_n18094_ );
xnor ( new_n18327_, new_n18326_, new_n18104_ );
or   ( new_n18328_, new_n18327_, new_n18325_ );
and  ( new_n18329_, new_n18328_, new_n18324_ );
nor  ( new_n18330_, new_n18329_, new_n18319_ );
and  ( new_n18331_, new_n18329_, new_n18319_ );
xor  ( new_n18332_, new_n18129_, new_n18127_ );
xnor ( new_n18333_, new_n18332_, new_n18133_ );
not  ( new_n18334_, new_n18333_ );
nor  ( new_n18335_, new_n18334_, new_n18331_ );
nor  ( new_n18336_, new_n18335_, new_n18330_ );
nor  ( new_n18337_, new_n18336_, new_n18317_ );
nor  ( new_n18338_, new_n18337_, new_n18316_ );
or   ( new_n18339_, new_n18338_, new_n18194_ );
and  ( new_n18340_, new_n18339_, new_n18193_ );
nor  ( new_n18341_, new_n18340_, new_n18180_ );
and  ( new_n18342_, new_n18340_, new_n18180_ );
xor  ( new_n18343_, new_n17949_, new_n17928_ );
xor  ( new_n18344_, new_n18343_, new_n17961_ );
nor  ( new_n18345_, new_n18344_, new_n18342_ );
or   ( new_n18346_, new_n18345_, new_n18341_ );
xnor ( new_n18347_, new_n18160_, new_n17996_ );
xor  ( new_n18348_, new_n18347_, new_n18164_ );
and  ( new_n18349_, new_n18348_, new_n18346_ );
xor  ( new_n18350_, new_n18166_, new_n17994_ );
and  ( new_n18351_, new_n18350_, new_n18349_ );
xor  ( new_n18352_, new_n18340_, new_n18180_ );
xor  ( new_n18353_, new_n18352_, new_n18344_ );
xor  ( new_n18354_, new_n18154_, new_n18144_ );
xor  ( new_n18355_, new_n18354_, new_n18158_ );
nor  ( new_n18356_, new_n18355_, new_n18353_ );
xor  ( new_n18357_, new_n18348_, new_n18346_ );
and  ( new_n18358_, new_n18357_, new_n18356_ );
xor  ( new_n18359_, new_n18355_, new_n18353_ );
xor  ( new_n18360_, new_n18068_, new_n18062_ );
xor  ( new_n18361_, new_n18360_, new_n2121_ );
xnor ( new_n18362_, new_n18238_, new_n18234_ );
xor  ( new_n18363_, new_n18362_, new_n18244_ );
xnor ( new_n18364_, new_n18222_, new_n18216_ );
xor  ( new_n18365_, new_n18364_, new_n18228_ );
or   ( new_n18366_, new_n18365_, new_n18363_ );
and  ( new_n18367_, new_n18365_, new_n18363_ );
xor  ( new_n18368_, new_n18256_, new_n18252_ );
xnor ( new_n18369_, new_n18368_, new_n18262_ );
or   ( new_n18370_, new_n18369_, new_n18367_ );
and  ( new_n18371_, new_n18370_, new_n18366_ );
nor  ( new_n18372_, new_n18371_, new_n18361_ );
and  ( new_n18373_, new_n18371_, new_n18361_ );
xor  ( new_n18374_, new_n18323_, new_n18321_ );
xnor ( new_n18375_, new_n18374_, new_n18327_ );
not  ( new_n18376_, new_n18375_ );
nor  ( new_n18377_, new_n18376_, new_n18373_ );
nor  ( new_n18378_, new_n18377_, new_n18372_ );
or   ( new_n18379_, new_n7732_, new_n4859_ );
or   ( new_n18380_, new_n7734_, new_n4995_ );
and  ( new_n18381_, new_n18380_, new_n18379_ );
xor  ( new_n18382_, new_n18381_, new_n7177_ );
or   ( new_n18383_, new_n7184_, new_n5428_ );
or   ( new_n18384_, new_n7186_, new_n5171_ );
and  ( new_n18385_, new_n18384_, new_n18383_ );
xor  ( new_n18386_, new_n18385_, new_n6638_ );
nor  ( new_n18387_, new_n18386_, new_n18382_ );
nand ( new_n18388_, new_n18386_, new_n18382_ );
or   ( new_n18389_, new_n6645_, new_n5899_ );
or   ( new_n18390_, new_n6647_, new_n5570_ );
and  ( new_n18391_, new_n18390_, new_n18389_ );
xor  ( new_n18392_, new_n18391_, new_n6165_ );
and  ( new_n18393_, new_n18392_, new_n18388_ );
or   ( new_n18394_, new_n18393_, new_n18387_ );
or   ( new_n18395_, new_n10059_, new_n3306_ );
or   ( new_n18396_, new_n10061_, new_n3178_ );
and  ( new_n18397_, new_n18396_, new_n18395_ );
xor  ( new_n18398_, new_n18397_, new_n9421_ );
and  ( new_n18399_, RIbb2d888_64, RIbb2c988_96 );
or   ( new_n18400_, RIbb2d888_64, new_n2981_ );
and  ( new_n18401_, new_n18400_, RIbb2d900_63 );
or   ( new_n18402_, new_n18401_, new_n18399_ );
or   ( new_n18403_, new_n10770_, new_n2751_ );
and  ( new_n18404_, new_n18403_, new_n18402_ );
nor  ( new_n18405_, new_n18404_, new_n18398_ );
nand ( new_n18406_, new_n18404_, new_n18398_ );
and  ( new_n18407_, new_n18406_, new_n2424_ );
or   ( new_n18408_, new_n18407_, new_n18405_ );
or   ( new_n18409_, new_n9422_, new_n3694_ );
or   ( new_n18410_, new_n9424_, new_n3696_ );
and  ( new_n18411_, new_n18410_, new_n18409_ );
xor  ( new_n18412_, new_n18411_, new_n8873_ );
or   ( new_n18413_, new_n8874_, new_n4069_ );
or   ( new_n18414_, new_n8876_, new_n3820_ );
and  ( new_n18415_, new_n18414_, new_n18413_ );
xor  ( new_n18416_, new_n18415_, new_n8257_ );
nor  ( new_n18417_, new_n18416_, new_n18412_ );
and  ( new_n18418_, new_n18416_, new_n18412_ );
or   ( new_n18419_, new_n8264_, new_n4603_ );
or   ( new_n18420_, new_n8266_, new_n4267_ );
and  ( new_n18421_, new_n18420_, new_n18419_ );
xor  ( new_n18422_, new_n18421_, new_n7725_ );
nor  ( new_n18423_, new_n18422_, new_n18418_ );
nor  ( new_n18424_, new_n18423_, new_n18417_ );
not  ( new_n18425_, new_n18424_ );
or   ( new_n18426_, new_n18425_, new_n18408_ );
and  ( new_n18427_, new_n18426_, new_n18394_ );
and  ( new_n18428_, new_n18425_, new_n18408_ );
or   ( new_n18429_, new_n18428_, new_n18427_ );
or   ( new_n18430_, new_n6173_, new_n6425_ );
or   ( new_n18431_, new_n6175_, new_n6219_ );
and  ( new_n18432_, new_n18431_, new_n18430_ );
xor  ( new_n18433_, new_n18432_, new_n5597_ );
or   ( new_n18434_, new_n5604_, new_n6943_ );
or   ( new_n18435_, new_n5606_, new_n6589_ );
and  ( new_n18436_, new_n18435_, new_n18434_ );
xor  ( new_n18437_, new_n18436_, new_n5206_ );
nor  ( new_n18438_, new_n18437_, new_n18433_ );
nand ( new_n18439_, new_n18437_, new_n18433_ );
or   ( new_n18440_, new_n5207_, new_n7373_ );
or   ( new_n18441_, new_n5209_, new_n7149_ );
and  ( new_n18442_, new_n18441_, new_n18440_ );
xor  ( new_n18443_, new_n18442_, new_n4708_ );
not  ( new_n18444_, new_n18443_ );
and  ( new_n18445_, new_n18444_, new_n18439_ );
or   ( new_n18446_, new_n18445_, new_n18438_ );
or   ( new_n18447_, new_n4709_, new_n8115_ );
or   ( new_n18448_, new_n4711_, new_n8117_ );
and  ( new_n18449_, new_n18448_, new_n18447_ );
xor  ( new_n18450_, new_n18449_, new_n4295_ );
or   ( new_n18451_, new_n4302_, new_n8481_ );
or   ( new_n18452_, new_n4304_, new_n8352_ );
and  ( new_n18453_, new_n18452_, new_n18451_ );
xor  ( new_n18454_, new_n18453_, new_n3895_ );
nor  ( new_n18455_, new_n18454_, new_n18450_ );
and  ( new_n18456_, new_n18454_, new_n18450_ );
or   ( new_n18457_, new_n3896_, new_n9099_ );
or   ( new_n18458_, new_n3898_, new_n8995_ );
and  ( new_n18459_, new_n18458_, new_n18457_ );
xor  ( new_n18460_, new_n18459_, new_n3460_ );
nor  ( new_n18461_, new_n18460_, new_n18456_ );
nor  ( new_n18462_, new_n18461_, new_n18455_ );
not  ( new_n18463_, new_n18462_ );
or   ( new_n18464_, new_n18463_, new_n18446_ );
and  ( new_n18465_, new_n18463_, new_n18446_ );
or   ( new_n18466_, new_n3461_, new_n9679_ );
or   ( new_n18467_, new_n3463_, new_n9681_ );
and  ( new_n18468_, new_n18467_, new_n18466_ );
xor  ( new_n18469_, new_n18468_, new_n3116_ );
or   ( new_n18470_, new_n3117_, new_n10541_ );
or   ( new_n18471_, new_n3119_, new_n10220_ );
and  ( new_n18472_, new_n18471_, new_n18470_ );
xor  ( new_n18473_, new_n18472_, new_n2800_ );
nand ( new_n18474_, new_n18473_, new_n18469_ );
nor  ( new_n18475_, new_n18473_, new_n18469_ );
and  ( new_n18476_, new_n2613_, RIbb31578_128 );
nor  ( new_n18477_, new_n18476_, new_n2424_ );
and  ( new_n18478_, new_n18476_, new_n2421_ );
nor  ( new_n18479_, new_n18478_, new_n18477_ );
or   ( new_n18480_, new_n18479_, new_n18475_ );
and  ( new_n18481_, new_n18480_, new_n18474_ );
or   ( new_n18482_, new_n18481_, new_n18465_ );
and  ( new_n18483_, new_n18482_, new_n18464_ );
nor  ( new_n18484_, new_n18483_, new_n18429_ );
and  ( new_n18485_, new_n18483_, new_n18429_ );
xnor ( new_n18486_, new_n18276_, new_n18272_ );
xor  ( new_n18487_, new_n18486_, new_n18282_ );
xnor ( new_n18488_, new_n18301_, new_n18297_ );
xor  ( new_n18489_, new_n18488_, new_n18307_ );
nor  ( new_n18490_, new_n18489_, new_n18487_ );
and  ( new_n18491_, new_n18489_, new_n18487_ );
xor  ( new_n18492_, new_n18292_, new_n18288_ );
not  ( new_n18493_, new_n18492_ );
nor  ( new_n18494_, new_n18493_, new_n18491_ );
nor  ( new_n18495_, new_n18494_, new_n18490_ );
nor  ( new_n18496_, new_n18495_, new_n18485_ );
nor  ( new_n18497_, new_n18496_, new_n18484_ );
and  ( new_n18498_, new_n18497_, new_n18378_ );
xor  ( new_n18499_, new_n18246_, new_n18230_ );
xor  ( new_n18500_, new_n18499_, new_n18264_ );
xor  ( new_n18501_, new_n18309_, new_n18293_ );
xor  ( new_n18502_, new_n18501_, new_n18284_ );
and  ( new_n18503_, new_n18502_, new_n18500_ );
nor  ( new_n18504_, new_n18502_, new_n18500_ );
not  ( new_n18505_, new_n18504_ );
xor  ( new_n18506_, new_n18205_, new_n18203_ );
xor  ( new_n18507_, new_n18506_, new_n18210_ );
and  ( new_n18508_, new_n18507_, new_n18505_ );
nor  ( new_n18509_, new_n18508_, new_n18503_ );
nor  ( new_n18510_, new_n18509_, new_n18498_ );
nor  ( new_n18511_, new_n18497_, new_n18378_ );
or   ( new_n18512_, new_n18511_, new_n18510_ );
xor  ( new_n18513_, new_n18184_, new_n18182_ );
xor  ( new_n18514_, new_n18513_, new_n18188_ );
or   ( new_n18515_, new_n18514_, new_n18512_ );
nand ( new_n18516_, new_n18514_, new_n18512_ );
xor  ( new_n18517_, new_n18329_, new_n18319_ );
xor  ( new_n18518_, new_n18517_, new_n18334_ );
xnor ( new_n18519_, new_n18266_, new_n18212_ );
xor  ( new_n18520_, new_n18519_, new_n18313_ );
nor  ( new_n18521_, new_n18520_, new_n18518_ );
and  ( new_n18522_, new_n18520_, new_n18518_ );
xor  ( new_n18523_, new_n18198_, new_n18196_ );
not  ( new_n18524_, new_n18523_ );
nor  ( new_n18525_, new_n18524_, new_n18522_ );
nor  ( new_n18526_, new_n18525_, new_n18521_ );
nand ( new_n18527_, new_n18526_, new_n18516_ );
and  ( new_n18528_, new_n18527_, new_n18515_ );
xnor ( new_n18529_, new_n18192_, new_n18190_ );
xor  ( new_n18530_, new_n18529_, new_n18338_ );
or   ( new_n18531_, new_n18530_, new_n18528_ );
and  ( new_n18532_, new_n18530_, new_n18528_ );
xor  ( new_n18533_, new_n18179_, new_n18177_ );
or   ( new_n18534_, new_n18533_, new_n18532_ );
and  ( new_n18535_, new_n18534_, new_n18531_ );
and  ( new_n18536_, new_n18535_, new_n18359_ );
xnor ( new_n18537_, new_n18530_, new_n18528_ );
xor  ( new_n18538_, new_n18537_, new_n18533_ );
xnor ( new_n18539_, new_n18497_, new_n18378_ );
and  ( new_n18540_, new_n18539_, new_n18509_ );
not  ( new_n18541_, new_n18510_ );
nor  ( new_n18542_, new_n18511_, new_n18541_ );
or   ( new_n18543_, new_n18542_, new_n18540_ );
xor  ( new_n18544_, new_n18462_, new_n18446_ );
xor  ( new_n18545_, new_n18544_, new_n18481_ );
xnor ( new_n18546_, new_n18365_, new_n18363_ );
xor  ( new_n18547_, new_n18546_, new_n18369_ );
or   ( new_n18548_, new_n18547_, new_n18545_ );
and  ( new_n18549_, new_n18547_, new_n18545_ );
xor  ( new_n18550_, new_n18489_, new_n18487_ );
xor  ( new_n18551_, new_n18550_, new_n18492_ );
or   ( new_n18552_, new_n18551_, new_n18549_ );
and  ( new_n18553_, new_n18552_, new_n18548_ );
xor  ( new_n18554_, new_n18502_, new_n18500_ );
xor  ( new_n18555_, new_n18554_, new_n18507_ );
nand ( new_n18556_, new_n18555_, new_n18553_ );
nor  ( new_n18557_, new_n18555_, new_n18553_ );
or   ( new_n18558_, new_n10059_, new_n3696_ );
or   ( new_n18559_, new_n10061_, new_n3306_ );
and  ( new_n18560_, new_n18559_, new_n18558_ );
xor  ( new_n18561_, new_n18560_, new_n9421_ );
and  ( new_n18562_, RIbb2d888_64, RIbb2c910_97 );
or   ( new_n18563_, RIbb2d888_64, new_n3178_ );
and  ( new_n18564_, new_n18563_, RIbb2d900_63 );
or   ( new_n18565_, new_n18564_, new_n18562_ );
or   ( new_n18566_, new_n10770_, new_n2981_ );
and  ( new_n18567_, new_n18566_, new_n18565_ );
or   ( new_n18568_, new_n18567_, new_n18561_ );
and  ( new_n18569_, new_n18567_, new_n18561_ );
or   ( new_n18570_, new_n9422_, new_n3820_ );
or   ( new_n18571_, new_n9424_, new_n3694_ );
and  ( new_n18572_, new_n18571_, new_n18570_ );
xor  ( new_n18573_, new_n18572_, new_n8873_ );
or   ( new_n18574_, new_n18573_, new_n18569_ );
and  ( new_n18575_, new_n18574_, new_n18568_ );
or   ( new_n18576_, new_n8874_, new_n4267_ );
or   ( new_n18577_, new_n8876_, new_n4069_ );
and  ( new_n18578_, new_n18577_, new_n18576_ );
xor  ( new_n18579_, new_n18578_, new_n8257_ );
or   ( new_n18580_, new_n8264_, new_n4995_ );
or   ( new_n18581_, new_n8266_, new_n4603_ );
and  ( new_n18582_, new_n18581_, new_n18580_ );
xor  ( new_n18583_, new_n18582_, new_n7725_ );
or   ( new_n18584_, new_n18583_, new_n18579_ );
and  ( new_n18585_, new_n18583_, new_n18579_ );
or   ( new_n18586_, new_n7732_, new_n5171_ );
or   ( new_n18587_, new_n7734_, new_n4859_ );
and  ( new_n18588_, new_n18587_, new_n18586_ );
xor  ( new_n18589_, new_n18588_, new_n7177_ );
or   ( new_n18590_, new_n18589_, new_n18585_ );
and  ( new_n18591_, new_n18590_, new_n18584_ );
or   ( new_n18592_, new_n18591_, new_n18575_ );
and  ( new_n18593_, new_n18591_, new_n18575_ );
or   ( new_n18594_, new_n7184_, new_n5570_ );
or   ( new_n18595_, new_n7186_, new_n5428_ );
and  ( new_n18596_, new_n18595_, new_n18594_ );
xor  ( new_n18597_, new_n18596_, new_n6638_ );
or   ( new_n18598_, new_n6645_, new_n6219_ );
or   ( new_n18599_, new_n6647_, new_n5899_ );
and  ( new_n18600_, new_n18599_, new_n18598_ );
xor  ( new_n18601_, new_n18600_, new_n6166_ );
nor  ( new_n18602_, new_n18601_, new_n18597_ );
and  ( new_n18603_, new_n18601_, new_n18597_ );
or   ( new_n18604_, new_n6173_, new_n6589_ );
or   ( new_n18605_, new_n6175_, new_n6425_ );
and  ( new_n18606_, new_n18605_, new_n18604_ );
xor  ( new_n18607_, new_n18606_, new_n5597_ );
nor  ( new_n18608_, new_n18607_, new_n18603_ );
nor  ( new_n18609_, new_n18608_, new_n18602_ );
or   ( new_n18610_, new_n18609_, new_n18593_ );
and  ( new_n18611_, new_n18610_, new_n18592_ );
xnor ( new_n18612_, new_n18473_, new_n18469_ );
xor  ( new_n18613_, new_n18612_, new_n18479_ );
or   ( new_n18614_, new_n5604_, new_n7149_ );
or   ( new_n18615_, new_n5606_, new_n6943_ );
and  ( new_n18616_, new_n18615_, new_n18614_ );
xor  ( new_n18617_, new_n18616_, new_n5206_ );
or   ( new_n18618_, new_n5207_, new_n8117_ );
or   ( new_n18619_, new_n5209_, new_n7373_ );
and  ( new_n18620_, new_n18619_, new_n18618_ );
xor  ( new_n18621_, new_n18620_, new_n4708_ );
or   ( new_n18622_, new_n18621_, new_n18617_ );
and  ( new_n18623_, new_n18621_, new_n18617_ );
or   ( new_n18624_, new_n4709_, new_n8352_ );
or   ( new_n18625_, new_n4711_, new_n8115_ );
and  ( new_n18626_, new_n18625_, new_n18624_ );
xor  ( new_n18627_, new_n18626_, new_n4295_ );
or   ( new_n18628_, new_n18627_, new_n18623_ );
and  ( new_n18629_, new_n18628_, new_n18622_ );
or   ( new_n18630_, new_n18629_, new_n18613_ );
and  ( new_n18631_, new_n18629_, new_n18613_ );
or   ( new_n18632_, new_n4302_, new_n8995_ );
or   ( new_n18633_, new_n4304_, new_n8481_ );
and  ( new_n18634_, new_n18633_, new_n18632_ );
xor  ( new_n18635_, new_n18634_, new_n3895_ );
or   ( new_n18636_, new_n3896_, new_n9681_ );
or   ( new_n18637_, new_n3898_, new_n9099_ );
and  ( new_n18638_, new_n18637_, new_n18636_ );
xor  ( new_n18639_, new_n18638_, new_n3460_ );
nor  ( new_n18640_, new_n18639_, new_n18635_ );
and  ( new_n18641_, new_n18639_, new_n18635_ );
or   ( new_n18642_, new_n3461_, new_n10220_ );
or   ( new_n18643_, new_n3463_, new_n9679_ );
and  ( new_n18644_, new_n18643_, new_n18642_ );
xor  ( new_n18645_, new_n18644_, new_n3116_ );
nor  ( new_n18646_, new_n18645_, new_n18641_ );
nor  ( new_n18647_, new_n18646_, new_n18640_ );
or   ( new_n18648_, new_n18647_, new_n18631_ );
and  ( new_n18649_, new_n18648_, new_n18630_ );
and  ( new_n18650_, new_n18649_, new_n18611_ );
nor  ( new_n18651_, new_n18649_, new_n18611_ );
xnor ( new_n18652_, new_n18454_, new_n18450_ );
xor  ( new_n18653_, new_n18652_, new_n18460_ );
xor  ( new_n18654_, new_n18386_, new_n18382_ );
xor  ( new_n18655_, new_n18654_, new_n18392_ );
nor  ( new_n18656_, new_n18655_, new_n18653_ );
and  ( new_n18657_, new_n18655_, new_n18653_ );
xor  ( new_n18658_, new_n18437_, new_n18433_ );
xor  ( new_n18659_, new_n18658_, new_n18444_ );
nor  ( new_n18660_, new_n18659_, new_n18657_ );
nor  ( new_n18661_, new_n18660_, new_n18656_ );
nor  ( new_n18662_, new_n18661_, new_n18651_ );
nor  ( new_n18663_, new_n18662_, new_n18650_ );
or   ( new_n18664_, new_n18663_, new_n18557_ );
and  ( new_n18665_, new_n18664_, new_n18556_ );
nor  ( new_n18666_, new_n18665_, new_n18543_ );
and  ( new_n18667_, new_n18665_, new_n18543_ );
xor  ( new_n18668_, new_n18520_, new_n18518_ );
xor  ( new_n18669_, new_n18668_, new_n18524_ );
nor  ( new_n18670_, new_n18669_, new_n18667_ );
or   ( new_n18671_, new_n18670_, new_n18666_ );
xnor ( new_n18672_, new_n18315_, new_n18199_ );
xor  ( new_n18673_, new_n18672_, new_n18336_ );
nand ( new_n18674_, new_n18673_, new_n18671_ );
nor  ( new_n18675_, new_n18673_, new_n18671_ );
xor  ( new_n18676_, new_n18514_, new_n18512_ );
xor  ( new_n18677_, new_n18676_, new_n18526_ );
or   ( new_n18678_, new_n18677_, new_n18675_ );
and  ( new_n18679_, new_n18678_, new_n18674_ );
nor  ( new_n18680_, new_n18679_, new_n18538_ );
xor  ( new_n18681_, new_n18673_, new_n18671_ );
xor  ( new_n18682_, new_n18681_, new_n18677_ );
xor  ( new_n18683_, new_n18483_, new_n18429_ );
xor  ( new_n18684_, new_n18683_, new_n18495_ );
xnor ( new_n18685_, new_n18555_, new_n18553_ );
xnor ( new_n18686_, new_n18685_, new_n18663_ );
or   ( new_n18687_, new_n18686_, new_n18684_ );
xor  ( new_n18688_, new_n18371_, new_n18361_ );
xor  ( new_n18689_, new_n18688_, new_n18376_ );
xor  ( new_n18690_, new_n18424_, new_n18408_ );
xor  ( new_n18691_, new_n18690_, new_n18394_ );
xnor ( new_n18692_, new_n18649_, new_n18611_ );
xor  ( new_n18693_, new_n18692_, new_n18661_ );
nand ( new_n18694_, new_n18693_, new_n18691_ );
nor  ( new_n18695_, new_n18693_, new_n18691_ );
xor  ( new_n18696_, new_n18547_, new_n18545_ );
xnor ( new_n18697_, new_n18696_, new_n18551_ );
or   ( new_n18698_, new_n18697_, new_n18695_ );
and  ( new_n18699_, new_n18698_, new_n18694_ );
or   ( new_n18700_, new_n18699_, new_n18689_ );
and  ( new_n18701_, new_n18699_, new_n18689_ );
xor  ( new_n18702_, new_n18591_, new_n18575_ );
xnor ( new_n18703_, new_n18702_, new_n18609_ );
xnor ( new_n18704_, new_n18629_, new_n18613_ );
xor  ( new_n18705_, new_n18704_, new_n18647_ );
or   ( new_n18706_, new_n18705_, new_n18703_ );
or   ( new_n18707_, new_n3117_, new_n10841_ );
or   ( new_n18708_, new_n3119_, new_n10541_ );
and  ( new_n18709_, new_n18708_, new_n18707_ );
xor  ( new_n18710_, new_n18709_, new_n2800_ );
or   ( new_n18711_, new_n4709_, new_n8481_ );
or   ( new_n18712_, new_n4711_, new_n8352_ );
and  ( new_n18713_, new_n18712_, new_n18711_ );
xor  ( new_n18714_, new_n18713_, new_n4295_ );
or   ( new_n18715_, new_n4302_, new_n9099_ );
or   ( new_n18716_, new_n4304_, new_n8995_ );
and  ( new_n18717_, new_n18716_, new_n18715_ );
xor  ( new_n18718_, new_n18717_, new_n3895_ );
or   ( new_n18719_, new_n18718_, new_n18714_ );
and  ( new_n18720_, new_n18718_, new_n18714_ );
or   ( new_n18721_, new_n3896_, new_n9679_ );
or   ( new_n18722_, new_n3898_, new_n9681_ );
and  ( new_n18723_, new_n18722_, new_n18721_ );
xor  ( new_n18724_, new_n18723_, new_n3460_ );
or   ( new_n18725_, new_n18724_, new_n18720_ );
and  ( new_n18726_, new_n18725_, new_n18719_ );
or   ( new_n18727_, new_n18726_, new_n18710_ );
and  ( new_n18728_, new_n18726_, new_n18710_ );
or   ( new_n18729_, new_n6173_, new_n6943_ );
or   ( new_n18730_, new_n6175_, new_n6589_ );
and  ( new_n18731_, new_n18730_, new_n18729_ );
xor  ( new_n18732_, new_n18731_, new_n5597_ );
or   ( new_n18733_, new_n5604_, new_n7373_ );
or   ( new_n18734_, new_n5606_, new_n7149_ );
and  ( new_n18735_, new_n18734_, new_n18733_ );
xor  ( new_n18736_, new_n18735_, new_n5206_ );
nor  ( new_n18737_, new_n18736_, new_n18732_ );
and  ( new_n18738_, new_n18736_, new_n18732_ );
or   ( new_n18739_, new_n5207_, new_n8115_ );
or   ( new_n18740_, new_n5209_, new_n8117_ );
and  ( new_n18741_, new_n18740_, new_n18739_ );
xor  ( new_n18742_, new_n18741_, new_n4708_ );
nor  ( new_n18743_, new_n18742_, new_n18738_ );
nor  ( new_n18744_, new_n18743_, new_n18737_ );
or   ( new_n18745_, new_n18744_, new_n18728_ );
and  ( new_n18746_, new_n18745_, new_n18727_ );
or   ( new_n18747_, new_n9422_, new_n4069_ );
or   ( new_n18748_, new_n9424_, new_n3820_ );
and  ( new_n18749_, new_n18748_, new_n18747_ );
xor  ( new_n18750_, new_n18749_, new_n8873_ );
or   ( new_n18751_, new_n8874_, new_n4603_ );
or   ( new_n18752_, new_n8876_, new_n4267_ );
and  ( new_n18753_, new_n18752_, new_n18751_ );
xor  ( new_n18754_, new_n18753_, new_n8257_ );
nor  ( new_n18755_, new_n18754_, new_n18750_ );
and  ( new_n18756_, new_n18754_, new_n18750_ );
or   ( new_n18757_, new_n8264_, new_n4859_ );
or   ( new_n18758_, new_n8266_, new_n4995_ );
and  ( new_n18759_, new_n18758_, new_n18757_ );
xor  ( new_n18760_, new_n18759_, new_n7725_ );
nor  ( new_n18761_, new_n18760_, new_n18756_ );
nor  ( new_n18762_, new_n18761_, new_n18755_ );
or   ( new_n18763_, new_n10059_, new_n3694_ );
or   ( new_n18764_, new_n10061_, new_n3696_ );
and  ( new_n18765_, new_n18764_, new_n18763_ );
xor  ( new_n18766_, new_n18765_, new_n9421_ );
and  ( new_n18767_, RIbb2d888_64, RIbb2c898_98 );
or   ( new_n18768_, RIbb2d888_64, new_n3306_ );
and  ( new_n18769_, new_n18768_, RIbb2d900_63 );
or   ( new_n18770_, new_n18769_, new_n18767_ );
or   ( new_n18771_, new_n10770_, new_n3178_ );
and  ( new_n18772_, new_n18771_, new_n18770_ );
nor  ( new_n18773_, new_n18772_, new_n18766_ );
and  ( new_n18774_, new_n18772_, new_n18766_ );
nor  ( new_n18775_, new_n18774_, new_n2799_ );
nor  ( new_n18776_, new_n18775_, new_n18773_ );
or   ( new_n18777_, new_n7732_, new_n5428_ );
or   ( new_n18778_, new_n7734_, new_n5171_ );
and  ( new_n18779_, new_n18778_, new_n18777_ );
xor  ( new_n18780_, new_n18779_, new_n7177_ );
or   ( new_n18781_, new_n7184_, new_n5899_ );
or   ( new_n18782_, new_n7186_, new_n5570_ );
and  ( new_n18783_, new_n18782_, new_n18781_ );
xor  ( new_n18784_, new_n18783_, new_n6638_ );
or   ( new_n18785_, new_n18784_, new_n18780_ );
and  ( new_n18786_, new_n18784_, new_n18780_ );
or   ( new_n18787_, new_n6645_, new_n6425_ );
or   ( new_n18788_, new_n6647_, new_n6219_ );
and  ( new_n18789_, new_n18788_, new_n18787_ );
xor  ( new_n18790_, new_n18789_, new_n6166_ );
or   ( new_n18791_, new_n18790_, new_n18786_ );
and  ( new_n18792_, new_n18791_, new_n18785_ );
and  ( new_n18793_, new_n18792_, new_n18776_ );
or   ( new_n18794_, new_n18793_, new_n18762_ );
or   ( new_n18795_, new_n18792_, new_n18776_ );
and  ( new_n18796_, new_n18795_, new_n18794_ );
nand ( new_n18797_, new_n18796_, new_n18746_ );
nor  ( new_n18798_, new_n18796_, new_n18746_ );
xnor ( new_n18799_, new_n18621_, new_n18617_ );
xor  ( new_n18800_, new_n18799_, new_n18627_ );
xnor ( new_n18801_, new_n18639_, new_n18635_ );
xor  ( new_n18802_, new_n18801_, new_n18645_ );
nor  ( new_n18803_, new_n18802_, new_n18800_ );
and  ( new_n18804_, new_n18802_, new_n18800_ );
xor  ( new_n18805_, new_n18601_, new_n18597_ );
xnor ( new_n18806_, new_n18805_, new_n18607_ );
nor  ( new_n18807_, new_n18806_, new_n18804_ );
nor  ( new_n18808_, new_n18807_, new_n18803_ );
or   ( new_n18809_, new_n18808_, new_n18798_ );
and  ( new_n18810_, new_n18809_, new_n18797_ );
nor  ( new_n18811_, new_n18810_, new_n18706_ );
and  ( new_n18812_, new_n18810_, new_n18706_ );
xor  ( new_n18813_, new_n18404_, new_n18398_ );
xor  ( new_n18814_, new_n18813_, new_n2424_ );
xnor ( new_n18815_, new_n18416_, new_n18412_ );
xor  ( new_n18816_, new_n18815_, new_n18422_ );
nor  ( new_n18817_, new_n18816_, new_n18814_ );
and  ( new_n18818_, new_n18816_, new_n18814_ );
not  ( new_n18819_, new_n18818_ );
xor  ( new_n18820_, new_n18655_, new_n18653_ );
xnor ( new_n18821_, new_n18820_, new_n18659_ );
and  ( new_n18822_, new_n18821_, new_n18819_ );
nor  ( new_n18823_, new_n18822_, new_n18817_ );
nor  ( new_n18824_, new_n18823_, new_n18812_ );
nor  ( new_n18825_, new_n18824_, new_n18811_ );
or   ( new_n18826_, new_n18825_, new_n18701_ );
and  ( new_n18827_, new_n18826_, new_n18700_ );
or   ( new_n18828_, new_n18827_, new_n18687_ );
and  ( new_n18829_, new_n18827_, new_n18687_ );
xor  ( new_n18830_, new_n18665_, new_n18543_ );
xor  ( new_n18831_, new_n18830_, new_n18669_ );
or   ( new_n18832_, new_n18831_, new_n18829_ );
and  ( new_n18833_, new_n18832_, new_n18828_ );
nor  ( new_n18834_, new_n18833_, new_n18682_ );
xnor ( new_n18835_, new_n18693_, new_n18691_ );
xor  ( new_n18836_, new_n18835_, new_n18697_ );
or   ( new_n18837_, new_n8874_, new_n4995_ );
or   ( new_n18838_, new_n8876_, new_n4603_ );
and  ( new_n18839_, new_n18838_, new_n18837_ );
xor  ( new_n18840_, new_n18839_, new_n8257_ );
or   ( new_n18841_, new_n8264_, new_n5171_ );
or   ( new_n18842_, new_n8266_, new_n4859_ );
and  ( new_n18843_, new_n18842_, new_n18841_ );
xor  ( new_n18844_, new_n18843_, new_n7725_ );
or   ( new_n18845_, new_n18844_, new_n18840_ );
and  ( new_n18846_, new_n18844_, new_n18840_ );
or   ( new_n18847_, new_n7732_, new_n5570_ );
or   ( new_n18848_, new_n7734_, new_n5428_ );
and  ( new_n18849_, new_n18848_, new_n18847_ );
xor  ( new_n18850_, new_n18849_, new_n7177_ );
or   ( new_n18851_, new_n18850_, new_n18846_ );
and  ( new_n18852_, new_n18851_, new_n18845_ );
or   ( new_n18853_, new_n7184_, new_n6219_ );
or   ( new_n18854_, new_n7186_, new_n5899_ );
and  ( new_n18855_, new_n18854_, new_n18853_ );
xor  ( new_n18856_, new_n18855_, new_n6638_ );
or   ( new_n18857_, new_n6645_, new_n6589_ );
or   ( new_n18858_, new_n6647_, new_n6425_ );
and  ( new_n18859_, new_n18858_, new_n18857_ );
xor  ( new_n18860_, new_n18859_, new_n6166_ );
or   ( new_n18861_, new_n18860_, new_n18856_ );
and  ( new_n18862_, new_n18860_, new_n18856_ );
or   ( new_n18863_, new_n6173_, new_n7149_ );
or   ( new_n18864_, new_n6175_, new_n6943_ );
and  ( new_n18865_, new_n18864_, new_n18863_ );
xor  ( new_n18866_, new_n18865_, new_n5597_ );
or   ( new_n18867_, new_n18866_, new_n18862_ );
and  ( new_n18868_, new_n18867_, new_n18861_ );
or   ( new_n18869_, new_n18868_, new_n18852_ );
and  ( new_n18870_, new_n18868_, new_n18852_ );
or   ( new_n18871_, new_n10059_, new_n3820_ );
or   ( new_n18872_, new_n10061_, new_n3694_ );
and  ( new_n18873_, new_n18872_, new_n18871_ );
xor  ( new_n18874_, new_n18873_, new_n9421_ );
and  ( new_n18875_, RIbb2d888_64, RIbb2c820_99 );
or   ( new_n18876_, RIbb2d888_64, new_n3696_ );
and  ( new_n18877_, new_n18876_, RIbb2d900_63 );
or   ( new_n18878_, new_n18877_, new_n18875_ );
or   ( new_n18879_, new_n10770_, new_n3306_ );
and  ( new_n18880_, new_n18879_, new_n18878_ );
nor  ( new_n18881_, new_n18880_, new_n18874_ );
and  ( new_n18882_, new_n18880_, new_n18874_ );
or   ( new_n18883_, new_n9422_, new_n4267_ );
or   ( new_n18884_, new_n9424_, new_n4069_ );
and  ( new_n18885_, new_n18884_, new_n18883_ );
xor  ( new_n18886_, new_n18885_, new_n8873_ );
nor  ( new_n18887_, new_n18886_, new_n18882_ );
nor  ( new_n18888_, new_n18887_, new_n18881_ );
or   ( new_n18889_, new_n18888_, new_n18870_ );
and  ( new_n18890_, new_n18889_, new_n18869_ );
or   ( new_n18891_, new_n3461_, new_n10541_ );
or   ( new_n18892_, new_n3463_, new_n10220_ );
and  ( new_n18893_, new_n18892_, new_n18891_ );
xor  ( new_n18894_, new_n18893_, new_n3116_ );
or   ( new_n18895_, new_n4302_, new_n9681_ );
or   ( new_n18896_, new_n4304_, new_n9099_ );
and  ( new_n18897_, new_n18896_, new_n18895_ );
xor  ( new_n18898_, new_n18897_, new_n3895_ );
or   ( new_n18899_, new_n3896_, new_n10220_ );
or   ( new_n18900_, new_n3898_, new_n9679_ );
and  ( new_n18901_, new_n18900_, new_n18899_ );
xor  ( new_n18902_, new_n18901_, new_n3460_ );
or   ( new_n18903_, new_n18902_, new_n18898_ );
and  ( new_n18904_, new_n18902_, new_n18898_ );
or   ( new_n18905_, new_n3461_, new_n10841_ );
or   ( new_n18906_, new_n3463_, new_n10541_ );
and  ( new_n18907_, new_n18906_, new_n18905_ );
xor  ( new_n18908_, new_n18907_, new_n3116_ );
or   ( new_n18909_, new_n18908_, new_n18904_ );
and  ( new_n18910_, new_n18909_, new_n18903_ );
or   ( new_n18911_, new_n18910_, new_n18894_ );
and  ( new_n18912_, new_n18910_, new_n18894_ );
or   ( new_n18913_, new_n5604_, new_n8117_ );
or   ( new_n18914_, new_n5606_, new_n7373_ );
and  ( new_n18915_, new_n18914_, new_n18913_ );
xor  ( new_n18916_, new_n18915_, new_n5206_ );
or   ( new_n18917_, new_n5207_, new_n8352_ );
or   ( new_n18918_, new_n5209_, new_n8115_ );
and  ( new_n18919_, new_n18918_, new_n18917_ );
xor  ( new_n18920_, new_n18919_, new_n4708_ );
nor  ( new_n18921_, new_n18920_, new_n18916_ );
and  ( new_n18922_, new_n18920_, new_n18916_ );
or   ( new_n18923_, new_n4709_, new_n8995_ );
or   ( new_n18924_, new_n4711_, new_n8481_ );
and  ( new_n18925_, new_n18924_, new_n18923_ );
xor  ( new_n18926_, new_n18925_, new_n4295_ );
nor  ( new_n18927_, new_n18926_, new_n18922_ );
nor  ( new_n18928_, new_n18927_, new_n18921_ );
or   ( new_n18929_, new_n18928_, new_n18912_ );
and  ( new_n18930_, new_n18929_, new_n18911_ );
nor  ( new_n18931_, new_n18930_, new_n18890_ );
nand ( new_n18932_, new_n18930_, new_n18890_ );
and  ( new_n18933_, new_n2928_, RIbb31578_128 );
or   ( new_n18934_, new_n18933_, new_n2800_ );
nand ( new_n18935_, new_n18933_, new_n2797_ );
and  ( new_n18936_, new_n18935_, new_n18934_ );
xnor ( new_n18937_, new_n18736_, new_n18732_ );
xor  ( new_n18938_, new_n18937_, new_n18742_ );
nor  ( new_n18939_, new_n18938_, new_n18936_ );
and  ( new_n18940_, new_n18938_, new_n18936_ );
xor  ( new_n18941_, new_n18718_, new_n18714_ );
xnor ( new_n18942_, new_n18941_, new_n18724_ );
nor  ( new_n18943_, new_n18942_, new_n18940_ );
nor  ( new_n18944_, new_n18943_, new_n18939_ );
and  ( new_n18945_, new_n18944_, new_n18932_ );
or   ( new_n18946_, new_n18945_, new_n18931_ );
xor  ( new_n18947_, new_n18802_, new_n18800_ );
xor  ( new_n18948_, new_n18947_, new_n18806_ );
xnor ( new_n18949_, new_n18726_, new_n18710_ );
xor  ( new_n18950_, new_n18949_, new_n18744_ );
or   ( new_n18951_, new_n18950_, new_n18948_ );
and  ( new_n18952_, new_n18950_, new_n18948_ );
xnor ( new_n18953_, new_n18792_, new_n18776_ );
xnor ( new_n18954_, new_n18953_, new_n18762_ );
not  ( new_n18955_, new_n18954_ );
or   ( new_n18956_, new_n18955_, new_n18952_ );
and  ( new_n18957_, new_n18956_, new_n18951_ );
nand ( new_n18958_, new_n18957_, new_n18946_ );
or   ( new_n18959_, new_n18957_, new_n18946_ );
xnor ( new_n18960_, new_n18583_, new_n18579_ );
xor  ( new_n18961_, new_n18960_, new_n18589_ );
xnor ( new_n18962_, new_n18754_, new_n18750_ );
xor  ( new_n18963_, new_n18962_, new_n18760_ );
xnor ( new_n18964_, new_n18784_, new_n18780_ );
xor  ( new_n18965_, new_n18964_, new_n18790_ );
or   ( new_n18966_, new_n18965_, new_n18963_ );
and  ( new_n18967_, new_n18965_, new_n18963_ );
xor  ( new_n18968_, new_n18772_, new_n18766_ );
xor  ( new_n18969_, new_n18968_, new_n2800_ );
or   ( new_n18970_, new_n18969_, new_n18967_ );
and  ( new_n18971_, new_n18970_, new_n18966_ );
nor  ( new_n18972_, new_n18971_, new_n18961_ );
and  ( new_n18973_, new_n18971_, new_n18961_ );
xor  ( new_n18974_, new_n18567_, new_n18561_ );
xnor ( new_n18975_, new_n18974_, new_n18573_ );
nor  ( new_n18976_, new_n18975_, new_n18973_ );
nor  ( new_n18977_, new_n18976_, new_n18972_ );
nand ( new_n18978_, new_n18977_, new_n18959_ );
and  ( new_n18979_, new_n18978_, new_n18958_ );
or   ( new_n18980_, new_n18979_, new_n18836_ );
nand ( new_n18981_, new_n18979_, new_n18836_ );
xor  ( new_n18982_, new_n18816_, new_n18814_ );
xor  ( new_n18983_, new_n18982_, new_n18821_ );
xnor ( new_n18984_, new_n18796_, new_n18746_ );
xor  ( new_n18985_, new_n18984_, new_n18808_ );
and  ( new_n18986_, new_n18985_, new_n18983_ );
nor  ( new_n18987_, new_n18985_, new_n18983_ );
xor  ( new_n18988_, new_n18705_, new_n18703_ );
not  ( new_n18989_, new_n18988_ );
nor  ( new_n18990_, new_n18989_, new_n18987_ );
nor  ( new_n18991_, new_n18990_, new_n18986_ );
nand ( new_n18992_, new_n18991_, new_n18981_ );
and  ( new_n18993_, new_n18992_, new_n18980_ );
xnor ( new_n18994_, new_n18699_, new_n18689_ );
xor  ( new_n18995_, new_n18994_, new_n18825_ );
nor  ( new_n18996_, new_n18995_, new_n18993_ );
nand ( new_n18997_, new_n18995_, new_n18993_ );
xnor ( new_n18998_, new_n18686_, new_n18684_ );
and  ( new_n18999_, new_n18998_, new_n18997_ );
or   ( new_n19000_, new_n18999_, new_n18996_ );
xor  ( new_n19001_, new_n18827_, new_n18687_ );
xor  ( new_n19002_, new_n19001_, new_n18831_ );
nor  ( new_n19003_, new_n19002_, new_n19000_ );
xor  ( new_n19004_, new_n18995_, new_n18993_ );
xor  ( new_n19005_, new_n19004_, new_n18998_ );
xor  ( new_n19006_, new_n18930_, new_n18890_ );
xnor ( new_n19007_, new_n19006_, new_n18944_ );
xnor ( new_n19008_, new_n18971_, new_n18961_ );
xor  ( new_n19009_, new_n19008_, new_n18975_ );
nand ( new_n19010_, new_n19009_, new_n19007_ );
xor  ( new_n19011_, new_n18965_, new_n18963_ );
xor  ( new_n19012_, new_n19011_, new_n18969_ );
xnor ( new_n19013_, new_n18910_, new_n18894_ );
xor  ( new_n19014_, new_n19013_, new_n18928_ );
or   ( new_n19015_, new_n19014_, new_n19012_ );
nand ( new_n19016_, new_n19014_, new_n19012_ );
xor  ( new_n19017_, new_n18938_, new_n18936_ );
xnor ( new_n19018_, new_n19017_, new_n18942_ );
nand ( new_n19019_, new_n19018_, new_n19016_ );
and  ( new_n19020_, new_n19019_, new_n19015_ );
xor  ( new_n19021_, new_n18902_, new_n18898_ );
xor  ( new_n19022_, new_n19021_, new_n18908_ );
or   ( new_n19023_, new_n6173_, new_n7373_ );
or   ( new_n19024_, new_n6175_, new_n7149_ );
and  ( new_n19025_, new_n19024_, new_n19023_ );
xor  ( new_n19026_, new_n19025_, new_n5597_ );
or   ( new_n19027_, new_n5604_, new_n8115_ );
or   ( new_n19028_, new_n5606_, new_n8117_ );
and  ( new_n19029_, new_n19028_, new_n19027_ );
xor  ( new_n19030_, new_n19029_, new_n5206_ );
or   ( new_n19031_, new_n19030_, new_n19026_ );
and  ( new_n19032_, new_n19030_, new_n19026_ );
or   ( new_n19033_, new_n5207_, new_n8481_ );
or   ( new_n19034_, new_n5209_, new_n8352_ );
and  ( new_n19035_, new_n19034_, new_n19033_ );
xor  ( new_n19036_, new_n19035_, new_n4708_ );
or   ( new_n19037_, new_n19036_, new_n19032_ );
and  ( new_n19038_, new_n19037_, new_n19031_ );
or   ( new_n19039_, new_n19038_, new_n19022_ );
and  ( new_n19040_, new_n19038_, new_n19022_ );
or   ( new_n19041_, new_n4709_, new_n9099_ );
or   ( new_n19042_, new_n4711_, new_n8995_ );
and  ( new_n19043_, new_n19042_, new_n19041_ );
xor  ( new_n19044_, new_n19043_, new_n4295_ );
or   ( new_n19045_, new_n4302_, new_n9679_ );
or   ( new_n19046_, new_n4304_, new_n9681_ );
and  ( new_n19047_, new_n19046_, new_n19045_ );
xor  ( new_n19048_, new_n19047_, new_n3895_ );
nor  ( new_n19049_, new_n19048_, new_n19044_ );
and  ( new_n19050_, new_n19048_, new_n19044_ );
or   ( new_n19051_, new_n3896_, new_n10541_ );
or   ( new_n19052_, new_n3898_, new_n10220_ );
and  ( new_n19053_, new_n19052_, new_n19051_ );
xor  ( new_n19054_, new_n19053_, new_n3460_ );
nor  ( new_n19055_, new_n19054_, new_n19050_ );
nor  ( new_n19056_, new_n19055_, new_n19049_ );
or   ( new_n19057_, new_n19056_, new_n19040_ );
and  ( new_n19058_, new_n19057_, new_n19039_ );
or   ( new_n19059_, new_n7732_, new_n5899_ );
or   ( new_n19060_, new_n7734_, new_n5570_ );
and  ( new_n19061_, new_n19060_, new_n19059_ );
xor  ( new_n19062_, new_n19061_, new_n7177_ );
or   ( new_n19063_, new_n7184_, new_n6425_ );
or   ( new_n19064_, new_n7186_, new_n6219_ );
and  ( new_n19065_, new_n19064_, new_n19063_ );
xor  ( new_n19066_, new_n19065_, new_n6638_ );
nor  ( new_n19067_, new_n19066_, new_n19062_ );
and  ( new_n19068_, new_n19066_, new_n19062_ );
or   ( new_n19069_, new_n6645_, new_n6943_ );
or   ( new_n19070_, new_n6647_, new_n6589_ );
and  ( new_n19071_, new_n19070_, new_n19069_ );
xor  ( new_n19072_, new_n19071_, new_n6166_ );
nor  ( new_n19073_, new_n19072_, new_n19068_ );
nor  ( new_n19074_, new_n19073_, new_n19067_ );
or   ( new_n19075_, new_n10059_, new_n4069_ );
or   ( new_n19076_, new_n10061_, new_n3820_ );
and  ( new_n19077_, new_n19076_, new_n19075_ );
xor  ( new_n19078_, new_n19077_, new_n9421_ );
and  ( new_n19079_, RIbb2d888_64, RIbb2c7a8_100 );
or   ( new_n19080_, RIbb2d888_64, new_n3694_ );
and  ( new_n19081_, new_n19080_, RIbb2d900_63 );
or   ( new_n19082_, new_n19081_, new_n19079_ );
or   ( new_n19083_, new_n10770_, new_n3696_ );
and  ( new_n19084_, new_n19083_, new_n19082_ );
nor  ( new_n19085_, new_n19084_, new_n19078_ );
and  ( new_n19086_, new_n19084_, new_n19078_ );
nor  ( new_n19087_, new_n19086_, new_n3115_ );
nor  ( new_n19088_, new_n19087_, new_n19085_ );
or   ( new_n19089_, new_n9422_, new_n4603_ );
or   ( new_n19090_, new_n9424_, new_n4267_ );
and  ( new_n19091_, new_n19090_, new_n19089_ );
xor  ( new_n19092_, new_n19091_, new_n8873_ );
or   ( new_n19093_, new_n8874_, new_n4859_ );
or   ( new_n19094_, new_n8876_, new_n4995_ );
and  ( new_n19095_, new_n19094_, new_n19093_ );
xor  ( new_n19096_, new_n19095_, new_n8257_ );
or   ( new_n19097_, new_n19096_, new_n19092_ );
and  ( new_n19098_, new_n19096_, new_n19092_ );
or   ( new_n19099_, new_n8264_, new_n5428_ );
or   ( new_n19100_, new_n8266_, new_n5171_ );
and  ( new_n19101_, new_n19100_, new_n19099_ );
xor  ( new_n19102_, new_n19101_, new_n7725_ );
or   ( new_n19103_, new_n19102_, new_n19098_ );
and  ( new_n19104_, new_n19103_, new_n19097_ );
and  ( new_n19105_, new_n19104_, new_n19088_ );
or   ( new_n19106_, new_n19105_, new_n19074_ );
or   ( new_n19107_, new_n19104_, new_n19088_ );
and  ( new_n19108_, new_n19107_, new_n19106_ );
nand ( new_n19109_, new_n19108_, new_n19058_ );
nor  ( new_n19110_, new_n19108_, new_n19058_ );
xnor ( new_n19111_, new_n18860_, new_n18856_ );
xor  ( new_n19112_, new_n19111_, new_n18866_ );
xnor ( new_n19113_, new_n18844_, new_n18840_ );
xor  ( new_n19114_, new_n19113_, new_n18850_ );
nor  ( new_n19115_, new_n19114_, new_n19112_ );
and  ( new_n19116_, new_n19114_, new_n19112_ );
xor  ( new_n19117_, new_n18920_, new_n18916_ );
xnor ( new_n19118_, new_n19117_, new_n18926_ );
nor  ( new_n19119_, new_n19118_, new_n19116_ );
nor  ( new_n19120_, new_n19119_, new_n19115_ );
or   ( new_n19121_, new_n19120_, new_n19110_ );
and  ( new_n19122_, new_n19121_, new_n19109_ );
or   ( new_n19123_, new_n19122_, new_n19020_ );
and  ( new_n19124_, new_n19122_, new_n19020_ );
xor  ( new_n19125_, new_n18950_, new_n18948_ );
xor  ( new_n19126_, new_n19125_, new_n18955_ );
or   ( new_n19127_, new_n19126_, new_n19124_ );
and  ( new_n19128_, new_n19127_, new_n19123_ );
nor  ( new_n19129_, new_n19128_, new_n19010_ );
nand ( new_n19130_, new_n19128_, new_n19010_ );
xor  ( new_n19131_, new_n18985_, new_n18983_ );
xor  ( new_n19132_, new_n19131_, new_n18988_ );
and  ( new_n19133_, new_n19132_, new_n19130_ );
or   ( new_n19134_, new_n19133_, new_n19129_ );
xnor ( new_n19135_, new_n18810_, new_n18706_ );
xor  ( new_n19136_, new_n19135_, new_n18823_ );
nand ( new_n19137_, new_n19136_, new_n19134_ );
nor  ( new_n19138_, new_n19136_, new_n19134_ );
xor  ( new_n19139_, new_n18979_, new_n18836_ );
xor  ( new_n19140_, new_n19139_, new_n18991_ );
or   ( new_n19141_, new_n19140_, new_n19138_ );
and  ( new_n19142_, new_n19141_, new_n19137_ );
nor  ( new_n19143_, new_n19142_, new_n19005_ );
xor  ( new_n19144_, new_n19136_, new_n19134_ );
xor  ( new_n19145_, new_n19144_, new_n19140_ );
or   ( new_n19146_, new_n7184_, new_n6589_ );
or   ( new_n19147_, new_n7186_, new_n6425_ );
and  ( new_n19148_, new_n19147_, new_n19146_ );
xor  ( new_n19149_, new_n19148_, new_n6638_ );
or   ( new_n19150_, new_n6645_, new_n7149_ );
or   ( new_n19151_, new_n6647_, new_n6943_ );
and  ( new_n19152_, new_n19151_, new_n19150_ );
xor  ( new_n19153_, new_n19152_, new_n6166_ );
or   ( new_n19154_, new_n19153_, new_n19149_ );
and  ( new_n19155_, new_n19153_, new_n19149_ );
or   ( new_n19156_, new_n6173_, new_n8117_ );
or   ( new_n19157_, new_n6175_, new_n7373_ );
and  ( new_n19158_, new_n19157_, new_n19156_ );
xor  ( new_n19159_, new_n19158_, new_n5597_ );
or   ( new_n19160_, new_n19159_, new_n19155_ );
and  ( new_n19161_, new_n19160_, new_n19154_ );
or   ( new_n19162_, new_n10059_, new_n4267_ );
or   ( new_n19163_, new_n10061_, new_n4069_ );
and  ( new_n19164_, new_n19163_, new_n19162_ );
xor  ( new_n19165_, new_n19164_, new_n9421_ );
and  ( new_n19166_, RIbb2d888_64, RIbb2c730_101 );
or   ( new_n19167_, RIbb2d888_64, new_n3820_ );
and  ( new_n19168_, new_n19167_, RIbb2d900_63 );
or   ( new_n19169_, new_n19168_, new_n19166_ );
or   ( new_n19170_, new_n10770_, new_n3694_ );
and  ( new_n19171_, new_n19170_, new_n19169_ );
or   ( new_n19172_, new_n19171_, new_n19165_ );
and  ( new_n19173_, new_n19171_, new_n19165_ );
or   ( new_n19174_, new_n9422_, new_n4995_ );
or   ( new_n19175_, new_n9424_, new_n4603_ );
and  ( new_n19176_, new_n19175_, new_n19174_ );
xor  ( new_n19177_, new_n19176_, new_n8873_ );
or   ( new_n19178_, new_n19177_, new_n19173_ );
and  ( new_n19179_, new_n19178_, new_n19172_ );
nor  ( new_n19180_, new_n19179_, new_n19161_ );
nand ( new_n19181_, new_n19179_, new_n19161_ );
or   ( new_n19182_, new_n8874_, new_n5171_ );
or   ( new_n19183_, new_n8876_, new_n4859_ );
and  ( new_n19184_, new_n19183_, new_n19182_ );
xor  ( new_n19185_, new_n19184_, new_n8257_ );
or   ( new_n19186_, new_n8264_, new_n5570_ );
or   ( new_n19187_, new_n8266_, new_n5428_ );
and  ( new_n19188_, new_n19187_, new_n19186_ );
xor  ( new_n19189_, new_n19188_, new_n7725_ );
nor  ( new_n19190_, new_n19189_, new_n19185_ );
nand ( new_n19191_, new_n19189_, new_n19185_ );
or   ( new_n19192_, new_n7732_, new_n6219_ );
or   ( new_n19193_, new_n7734_, new_n5899_ );
and  ( new_n19194_, new_n19193_, new_n19192_ );
xor  ( new_n19195_, new_n19194_, new_n7176_ );
and  ( new_n19196_, new_n19195_, new_n19191_ );
or   ( new_n19197_, new_n19196_, new_n19190_ );
and  ( new_n19198_, new_n19197_, new_n19181_ );
or   ( new_n19199_, new_n19198_, new_n19180_ );
and  ( new_n19200_, new_n3291_, RIbb31578_128 );
or   ( new_n19201_, new_n19200_, new_n3116_ );
nand ( new_n19202_, new_n19200_, new_n3113_ );
and  ( new_n19203_, new_n19202_, new_n19201_ );
xnor ( new_n19204_, new_n19048_, new_n19044_ );
xor  ( new_n19205_, new_n19204_, new_n19054_ );
or   ( new_n19206_, new_n19205_, new_n19203_ );
and  ( new_n19207_, new_n19205_, new_n19203_ );
or   ( new_n19208_, new_n5604_, new_n8352_ );
or   ( new_n19209_, new_n5606_, new_n8115_ );
and  ( new_n19210_, new_n19209_, new_n19208_ );
xor  ( new_n19211_, new_n19210_, new_n5206_ );
or   ( new_n19212_, new_n5207_, new_n8995_ );
or   ( new_n19213_, new_n5209_, new_n8481_ );
and  ( new_n19214_, new_n19213_, new_n19212_ );
xor  ( new_n19215_, new_n19214_, new_n4708_ );
nor  ( new_n19216_, new_n19215_, new_n19211_ );
and  ( new_n19217_, new_n19215_, new_n19211_ );
or   ( new_n19218_, new_n4709_, new_n9681_ );
or   ( new_n19219_, new_n4711_, new_n9099_ );
and  ( new_n19220_, new_n19219_, new_n19218_ );
xor  ( new_n19221_, new_n19220_, new_n4295_ );
nor  ( new_n19222_, new_n19221_, new_n19217_ );
nor  ( new_n19223_, new_n19222_, new_n19216_ );
not  ( new_n19224_, new_n19223_ );
or   ( new_n19225_, new_n19224_, new_n19207_ );
and  ( new_n19226_, new_n19225_, new_n19206_ );
and  ( new_n19227_, new_n19226_, new_n19199_ );
xnor ( new_n19228_, new_n19066_, new_n19062_ );
xor  ( new_n19229_, new_n19228_, new_n19072_ );
xnor ( new_n19230_, new_n19096_, new_n19092_ );
xor  ( new_n19231_, new_n19230_, new_n19102_ );
nor  ( new_n19232_, new_n19231_, new_n19229_ );
and  ( new_n19233_, new_n19231_, new_n19229_ );
xor  ( new_n19234_, new_n19030_, new_n19026_ );
xnor ( new_n19235_, new_n19234_, new_n19036_ );
nor  ( new_n19236_, new_n19235_, new_n19233_ );
nor  ( new_n19237_, new_n19236_, new_n19232_ );
or   ( new_n19238_, new_n19237_, new_n19227_ );
or   ( new_n19239_, new_n19226_, new_n19199_ );
and  ( new_n19240_, new_n19239_, new_n19238_ );
xnor ( new_n19241_, new_n18868_, new_n18852_ );
xor  ( new_n19242_, new_n19241_, new_n18888_ );
and  ( new_n19243_, new_n19242_, new_n19240_ );
xor  ( new_n19244_, new_n19114_, new_n19112_ );
xor  ( new_n19245_, new_n19244_, new_n19118_ );
xnor ( new_n19246_, new_n19038_, new_n19022_ );
xor  ( new_n19247_, new_n19246_, new_n19056_ );
nor  ( new_n19248_, new_n19247_, new_n19245_ );
and  ( new_n19249_, new_n19247_, new_n19245_ );
xor  ( new_n19250_, new_n18880_, new_n18874_ );
xnor ( new_n19251_, new_n19250_, new_n18886_ );
nor  ( new_n19252_, new_n19251_, new_n19249_ );
nor  ( new_n19253_, new_n19252_, new_n19248_ );
nor  ( new_n19254_, new_n19253_, new_n19243_ );
nor  ( new_n19255_, new_n19242_, new_n19240_ );
or   ( new_n19256_, new_n19255_, new_n19254_ );
xnor ( new_n19257_, new_n19122_, new_n19020_ );
xor  ( new_n19258_, new_n19257_, new_n19126_ );
nor  ( new_n19259_, new_n19258_, new_n19256_ );
nand ( new_n19260_, new_n19258_, new_n19256_ );
xnor ( new_n19261_, new_n19009_, new_n19007_ );
and  ( new_n19262_, new_n19261_, new_n19260_ );
or   ( new_n19263_, new_n19262_, new_n19259_ );
xor  ( new_n19264_, new_n18957_, new_n18946_ );
xor  ( new_n19265_, new_n19264_, new_n18977_ );
or   ( new_n19266_, new_n19265_, new_n19263_ );
and  ( new_n19267_, new_n19265_, new_n19263_ );
xnor ( new_n19268_, new_n19128_, new_n19010_ );
xor  ( new_n19269_, new_n19268_, new_n19132_ );
or   ( new_n19270_, new_n19269_, new_n19267_ );
and  ( new_n19271_, new_n19270_, new_n19266_ );
nor  ( new_n19272_, new_n19271_, new_n19145_ );
xor  ( new_n19273_, new_n19265_, new_n19263_ );
xor  ( new_n19274_, new_n19273_, new_n19269_ );
xor  ( new_n19275_, new_n19242_, new_n19240_ );
xor  ( new_n19276_, new_n19275_, new_n19253_ );
xnor ( new_n19277_, new_n19108_, new_n19058_ );
xnor ( new_n19278_, new_n19277_, new_n19120_ );
nor  ( new_n19279_, new_n19278_, new_n19276_ );
xor  ( new_n19280_, new_n19226_, new_n19199_ );
xor  ( new_n19281_, new_n19280_, new_n19237_ );
xnor ( new_n19282_, new_n19247_, new_n19245_ );
xnor ( new_n19283_, new_n19282_, new_n19251_ );
nor  ( new_n19284_, new_n19283_, new_n19281_ );
xor  ( new_n19285_, new_n19014_, new_n19012_ );
xor  ( new_n19286_, new_n19285_, new_n19018_ );
or   ( new_n19287_, new_n19286_, new_n19284_ );
and  ( new_n19288_, new_n19286_, new_n19284_ );
or   ( new_n19289_, new_n4302_, new_n10220_ );
or   ( new_n19290_, new_n4304_, new_n9679_ );
and  ( new_n19291_, new_n19290_, new_n19289_ );
xor  ( new_n19292_, new_n19291_, new_n3895_ );
or   ( new_n19293_, new_n6173_, new_n8115_ );
or   ( new_n19294_, new_n6175_, new_n8117_ );
and  ( new_n19295_, new_n19294_, new_n19293_ );
xor  ( new_n19296_, new_n19295_, new_n5597_ );
or   ( new_n19297_, new_n5604_, new_n8481_ );
or   ( new_n19298_, new_n5606_, new_n8352_ );
and  ( new_n19299_, new_n19298_, new_n19297_ );
xor  ( new_n19300_, new_n19299_, new_n5206_ );
or   ( new_n19301_, new_n19300_, new_n19296_ );
and  ( new_n19302_, new_n19300_, new_n19296_ );
or   ( new_n19303_, new_n5207_, new_n9099_ );
or   ( new_n19304_, new_n5209_, new_n8995_ );
and  ( new_n19305_, new_n19304_, new_n19303_ );
xor  ( new_n19306_, new_n19305_, new_n4708_ );
or   ( new_n19307_, new_n19306_, new_n19302_ );
and  ( new_n19308_, new_n19307_, new_n19301_ );
or   ( new_n19309_, new_n19308_, new_n19292_ );
nand ( new_n19310_, new_n19308_, new_n19292_ );
or   ( new_n19311_, new_n4709_, new_n9679_ );
or   ( new_n19312_, new_n4711_, new_n9681_ );
and  ( new_n19313_, new_n19312_, new_n19311_ );
xor  ( new_n19314_, new_n19313_, new_n4295_ );
or   ( new_n19315_, new_n4302_, new_n10541_ );
or   ( new_n19316_, new_n4304_, new_n10220_ );
and  ( new_n19317_, new_n19316_, new_n19315_ );
xor  ( new_n19318_, new_n19317_, new_n3895_ );
and  ( new_n19319_, new_n19318_, new_n19314_ );
nor  ( new_n19320_, new_n19318_, new_n19314_ );
and  ( new_n19321_, new_n3731_, RIbb31578_128 );
nor  ( new_n19322_, new_n19321_, new_n3460_ );
and  ( new_n19323_, new_n19321_, new_n3457_ );
nor  ( new_n19324_, new_n19323_, new_n19322_ );
nor  ( new_n19325_, new_n19324_, new_n19320_ );
nor  ( new_n19326_, new_n19325_, new_n19319_ );
nand ( new_n19327_, new_n19326_, new_n19310_ );
and  ( new_n19328_, new_n19327_, new_n19309_ );
or   ( new_n19329_, new_n7732_, new_n6425_ );
or   ( new_n19330_, new_n7734_, new_n6219_ );
and  ( new_n19331_, new_n19330_, new_n19329_ );
xor  ( new_n19332_, new_n19331_, new_n7177_ );
or   ( new_n19333_, new_n7184_, new_n6943_ );
or   ( new_n19334_, new_n7186_, new_n6589_ );
and  ( new_n19335_, new_n19334_, new_n19333_ );
xor  ( new_n19336_, new_n19335_, new_n6638_ );
nor  ( new_n19337_, new_n19336_, new_n19332_ );
and  ( new_n19338_, new_n19336_, new_n19332_ );
or   ( new_n19339_, new_n6645_, new_n7373_ );
or   ( new_n19340_, new_n6647_, new_n7149_ );
and  ( new_n19341_, new_n19340_, new_n19339_ );
xor  ( new_n19342_, new_n19341_, new_n6166_ );
nor  ( new_n19343_, new_n19342_, new_n19338_ );
nor  ( new_n19344_, new_n19343_, new_n19337_ );
or   ( new_n19345_, new_n10059_, new_n4603_ );
or   ( new_n19346_, new_n10061_, new_n4267_ );
and  ( new_n19347_, new_n19346_, new_n19345_ );
xor  ( new_n19348_, new_n19347_, new_n9421_ );
and  ( new_n19349_, RIbb2d888_64, RIbb2c6b8_102 );
or   ( new_n19350_, RIbb2d888_64, new_n4069_ );
and  ( new_n19351_, new_n19350_, RIbb2d900_63 );
or   ( new_n19352_, new_n19351_, new_n19349_ );
or   ( new_n19353_, new_n10770_, new_n3820_ );
and  ( new_n19354_, new_n19353_, new_n19352_ );
nor  ( new_n19355_, new_n19354_, new_n19348_ );
and  ( new_n19356_, new_n19354_, new_n19348_ );
nor  ( new_n19357_, new_n19356_, new_n3459_ );
nor  ( new_n19358_, new_n19357_, new_n19355_ );
or   ( new_n19359_, new_n9422_, new_n4859_ );
or   ( new_n19360_, new_n9424_, new_n4995_ );
and  ( new_n19361_, new_n19360_, new_n19359_ );
xor  ( new_n19362_, new_n19361_, new_n8873_ );
or   ( new_n19363_, new_n8874_, new_n5428_ );
or   ( new_n19364_, new_n8876_, new_n5171_ );
and  ( new_n19365_, new_n19364_, new_n19363_ );
xor  ( new_n19366_, new_n19365_, new_n8257_ );
or   ( new_n19367_, new_n19366_, new_n19362_ );
and  ( new_n19368_, new_n19366_, new_n19362_ );
or   ( new_n19369_, new_n8264_, new_n5899_ );
or   ( new_n19370_, new_n8266_, new_n5570_ );
and  ( new_n19371_, new_n19370_, new_n19369_ );
xor  ( new_n19372_, new_n19371_, new_n7725_ );
or   ( new_n19373_, new_n19372_, new_n19368_ );
and  ( new_n19374_, new_n19373_, new_n19367_ );
and  ( new_n19375_, new_n19374_, new_n19358_ );
or   ( new_n19376_, new_n19375_, new_n19344_ );
or   ( new_n19377_, new_n19374_, new_n19358_ );
and  ( new_n19378_, new_n19377_, new_n19376_ );
nor  ( new_n19379_, new_n19378_, new_n19328_ );
nand ( new_n19380_, new_n19378_, new_n19328_ );
or   ( new_n19381_, new_n3896_, new_n10841_ );
or   ( new_n19382_, new_n3898_, new_n10541_ );
and  ( new_n19383_, new_n19382_, new_n19381_ );
xor  ( new_n19384_, new_n19383_, new_n3459_ );
xnor ( new_n19385_, new_n19215_, new_n19211_ );
xor  ( new_n19386_, new_n19385_, new_n19221_ );
and  ( new_n19387_, new_n19386_, new_n19384_ );
or   ( new_n19388_, new_n19386_, new_n19384_ );
xor  ( new_n19389_, new_n19153_, new_n19149_ );
xnor ( new_n19390_, new_n19389_, new_n19159_ );
and  ( new_n19391_, new_n19390_, new_n19388_ );
or   ( new_n19392_, new_n19391_, new_n19387_ );
and  ( new_n19393_, new_n19392_, new_n19380_ );
or   ( new_n19394_, new_n19393_, new_n19379_ );
xor  ( new_n19395_, new_n19084_, new_n19078_ );
xnor ( new_n19396_, new_n19395_, new_n3116_ );
xnor ( new_n19397_, new_n19231_, new_n19229_ );
xor  ( new_n19398_, new_n19397_, new_n19235_ );
nand ( new_n19399_, new_n19398_, new_n19396_ );
nor  ( new_n19400_, new_n19398_, new_n19396_ );
xor  ( new_n19401_, new_n19205_, new_n19203_ );
xor  ( new_n19402_, new_n19401_, new_n19224_ );
or   ( new_n19403_, new_n19402_, new_n19400_ );
and  ( new_n19404_, new_n19403_, new_n19399_ );
and  ( new_n19405_, new_n19404_, new_n19394_ );
nor  ( new_n19406_, new_n19404_, new_n19394_ );
xnor ( new_n19407_, new_n19104_, new_n19088_ );
xnor ( new_n19408_, new_n19407_, new_n19074_ );
nor  ( new_n19409_, new_n19408_, new_n19406_ );
nor  ( new_n19410_, new_n19409_, new_n19405_ );
or   ( new_n19411_, new_n19410_, new_n19288_ );
and  ( new_n19412_, new_n19411_, new_n19287_ );
nand ( new_n19413_, new_n19412_, new_n19279_ );
nor  ( new_n19414_, new_n19412_, new_n19279_ );
xor  ( new_n19415_, new_n19258_, new_n19256_ );
xor  ( new_n19416_, new_n19415_, new_n19261_ );
or   ( new_n19417_, new_n19416_, new_n19414_ );
and  ( new_n19418_, new_n19417_, new_n19413_ );
nor  ( new_n19419_, new_n19418_, new_n19274_ );
xor  ( new_n19420_, new_n19412_, new_n19279_ );
xor  ( new_n19421_, new_n19420_, new_n19416_ );
xor  ( new_n19422_, new_n19179_, new_n19161_ );
xor  ( new_n19423_, new_n19422_, new_n19197_ );
xnor ( new_n19424_, new_n19171_, new_n19165_ );
xor  ( new_n19425_, new_n19424_, new_n19177_ );
xor  ( new_n19426_, new_n19189_, new_n19185_ );
xor  ( new_n19427_, new_n19426_, new_n19195_ );
or   ( new_n19428_, new_n19427_, new_n19425_ );
and  ( new_n19429_, new_n19427_, new_n19425_ );
xor  ( new_n19430_, new_n19386_, new_n19384_ );
xor  ( new_n19431_, new_n19430_, new_n19390_ );
or   ( new_n19432_, new_n19431_, new_n19429_ );
and  ( new_n19433_, new_n19432_, new_n19428_ );
or   ( new_n19434_, new_n19433_, new_n19423_ );
and  ( new_n19435_, new_n19433_, new_n19423_ );
or   ( new_n19436_, new_n10059_, new_n4995_ );
or   ( new_n19437_, new_n10061_, new_n4603_ );
and  ( new_n19438_, new_n19437_, new_n19436_ );
xor  ( new_n19439_, new_n19438_, new_n9421_ );
and  ( new_n19440_, RIbb2d888_64, RIbb2c640_103 );
or   ( new_n19441_, RIbb2d888_64, new_n4267_ );
and  ( new_n19442_, new_n19441_, RIbb2d900_63 );
or   ( new_n19443_, new_n19442_, new_n19440_ );
or   ( new_n19444_, new_n10770_, new_n4069_ );
and  ( new_n19445_, new_n19444_, new_n19443_ );
or   ( new_n19446_, new_n19445_, new_n19439_ );
and  ( new_n19447_, new_n19445_, new_n19439_ );
or   ( new_n19448_, new_n9422_, new_n5171_ );
or   ( new_n19449_, new_n9424_, new_n4859_ );
and  ( new_n19450_, new_n19449_, new_n19448_ );
xor  ( new_n19451_, new_n19450_, new_n8873_ );
or   ( new_n19452_, new_n19451_, new_n19447_ );
and  ( new_n19453_, new_n19452_, new_n19446_ );
or   ( new_n19454_, new_n8874_, new_n5570_ );
or   ( new_n19455_, new_n8876_, new_n5428_ );
and  ( new_n19456_, new_n19455_, new_n19454_ );
xor  ( new_n19457_, new_n19456_, new_n8257_ );
or   ( new_n19458_, new_n8264_, new_n6219_ );
or   ( new_n19459_, new_n8266_, new_n5899_ );
and  ( new_n19460_, new_n19459_, new_n19458_ );
xor  ( new_n19461_, new_n19460_, new_n7725_ );
or   ( new_n19462_, new_n19461_, new_n19457_ );
and  ( new_n19463_, new_n19461_, new_n19457_ );
or   ( new_n19464_, new_n7732_, new_n6589_ );
or   ( new_n19465_, new_n7734_, new_n6425_ );
and  ( new_n19466_, new_n19465_, new_n19464_ );
xor  ( new_n19467_, new_n19466_, new_n7177_ );
or   ( new_n19468_, new_n19467_, new_n19463_ );
and  ( new_n19469_, new_n19468_, new_n19462_ );
or   ( new_n19470_, new_n19469_, new_n19453_ );
and  ( new_n19471_, new_n19469_, new_n19453_ );
or   ( new_n19472_, new_n7184_, new_n7149_ );
or   ( new_n19473_, new_n7186_, new_n6943_ );
and  ( new_n19474_, new_n19473_, new_n19472_ );
xor  ( new_n19475_, new_n19474_, new_n6638_ );
or   ( new_n19476_, new_n6645_, new_n8117_ );
or   ( new_n19477_, new_n6647_, new_n7373_ );
and  ( new_n19478_, new_n19477_, new_n19476_ );
xor  ( new_n19479_, new_n19478_, new_n6166_ );
or   ( new_n19480_, new_n19479_, new_n19475_ );
and  ( new_n19481_, new_n19479_, new_n19475_ );
or   ( new_n19482_, new_n6173_, new_n8352_ );
or   ( new_n19483_, new_n6175_, new_n8115_ );
and  ( new_n19484_, new_n19483_, new_n19482_ );
xor  ( new_n19485_, new_n19484_, new_n5597_ );
or   ( new_n19486_, new_n19485_, new_n19481_ );
and  ( new_n19487_, new_n19486_, new_n19480_ );
or   ( new_n19488_, new_n19487_, new_n19471_ );
and  ( new_n19489_, new_n19488_, new_n19470_ );
xnor ( new_n19490_, new_n19318_, new_n19314_ );
xor  ( new_n19491_, new_n19490_, new_n19324_ );
or   ( new_n19492_, new_n5604_, new_n8995_ );
or   ( new_n19493_, new_n5606_, new_n8481_ );
and  ( new_n19494_, new_n19493_, new_n19492_ );
xor  ( new_n19495_, new_n19494_, new_n5206_ );
or   ( new_n19496_, new_n5207_, new_n9681_ );
or   ( new_n19497_, new_n5209_, new_n9099_ );
and  ( new_n19498_, new_n19497_, new_n19496_ );
xor  ( new_n19499_, new_n19498_, new_n4708_ );
or   ( new_n19500_, new_n19499_, new_n19495_ );
and  ( new_n19501_, new_n19499_, new_n19495_ );
or   ( new_n19502_, new_n4709_, new_n10220_ );
or   ( new_n19503_, new_n4711_, new_n9679_ );
and  ( new_n19504_, new_n19503_, new_n19502_ );
xor  ( new_n19505_, new_n19504_, new_n4295_ );
or   ( new_n19506_, new_n19505_, new_n19501_ );
and  ( new_n19507_, new_n19506_, new_n19500_ );
or   ( new_n19508_, new_n19507_, new_n19491_ );
nand ( new_n19509_, new_n19507_, new_n19491_ );
xor  ( new_n19510_, new_n19300_, new_n19296_ );
xnor ( new_n19511_, new_n19510_, new_n19306_ );
nand ( new_n19512_, new_n19511_, new_n19509_ );
and  ( new_n19513_, new_n19512_, new_n19508_ );
and  ( new_n19514_, new_n19513_, new_n19489_ );
nor  ( new_n19515_, new_n19513_, new_n19489_ );
xnor ( new_n19516_, new_n19336_, new_n19332_ );
xor  ( new_n19517_, new_n19516_, new_n19342_ );
xor  ( new_n19518_, new_n19354_, new_n19348_ );
xor  ( new_n19519_, new_n19518_, new_n3460_ );
nor  ( new_n19520_, new_n19519_, new_n19517_ );
and  ( new_n19521_, new_n19519_, new_n19517_ );
xor  ( new_n19522_, new_n19366_, new_n19362_ );
xnor ( new_n19523_, new_n19522_, new_n19372_ );
nor  ( new_n19524_, new_n19523_, new_n19521_ );
nor  ( new_n19525_, new_n19524_, new_n19520_ );
nor  ( new_n19526_, new_n19525_, new_n19515_ );
nor  ( new_n19527_, new_n19526_, new_n19514_ );
or   ( new_n19528_, new_n19527_, new_n19435_ );
and  ( new_n19529_, new_n19528_, new_n19434_ );
xnor ( new_n19530_, new_n19404_, new_n19394_ );
xor  ( new_n19531_, new_n19530_, new_n19408_ );
or   ( new_n19532_, new_n19531_, new_n19529_ );
and  ( new_n19533_, new_n19531_, new_n19529_ );
xnor ( new_n19534_, new_n19283_, new_n19281_ );
or   ( new_n19535_, new_n19534_, new_n19533_ );
and  ( new_n19536_, new_n19535_, new_n19532_ );
xnor ( new_n19537_, new_n19286_, new_n19284_ );
xor  ( new_n19538_, new_n19537_, new_n19410_ );
or   ( new_n19539_, new_n19538_, new_n19536_ );
and  ( new_n19540_, new_n19538_, new_n19536_ );
xnor ( new_n19541_, new_n19278_, new_n19276_ );
or   ( new_n19542_, new_n19541_, new_n19540_ );
and  ( new_n19543_, new_n19542_, new_n19539_ );
nor  ( new_n19544_, new_n19543_, new_n19421_ );
xor  ( new_n19545_, new_n19538_, new_n19536_ );
xor  ( new_n19546_, new_n19545_, new_n19541_ );
xor  ( new_n19547_, new_n19433_, new_n19423_ );
xnor ( new_n19548_, new_n19547_, new_n19527_ );
not  ( new_n19549_, new_n19548_ );
xor  ( new_n19550_, new_n19378_, new_n19328_ );
xor  ( new_n19551_, new_n19550_, new_n19392_ );
or   ( new_n19552_, new_n19551_, new_n19549_ );
xor  ( new_n19553_, new_n19374_, new_n19358_ );
xor  ( new_n19554_, new_n19553_, new_n19344_ );
xnor ( new_n19555_, new_n19513_, new_n19489_ );
xor  ( new_n19556_, new_n19555_, new_n19525_ );
or   ( new_n19557_, new_n19556_, new_n19554_ );
and  ( new_n19558_, new_n19556_, new_n19554_ );
xor  ( new_n19559_, new_n19427_, new_n19425_ );
xnor ( new_n19560_, new_n19559_, new_n19431_ );
or   ( new_n19561_, new_n19560_, new_n19558_ );
and  ( new_n19562_, new_n19561_, new_n19557_ );
xnor ( new_n19563_, new_n19398_, new_n19396_ );
xor  ( new_n19564_, new_n19563_, new_n19402_ );
nand ( new_n19565_, new_n19564_, new_n19562_ );
nor  ( new_n19566_, new_n19564_, new_n19562_ );
xor  ( new_n19567_, new_n19308_, new_n19292_ );
xor  ( new_n19568_, new_n19567_, new_n19326_ );
or   ( new_n19569_, new_n4709_, new_n10541_ );
or   ( new_n19570_, new_n4711_, new_n10220_ );
and  ( new_n19571_, new_n19570_, new_n19569_ );
xor  ( new_n19572_, new_n19571_, new_n4295_ );
not  ( new_n19573_, new_n19572_ );
and  ( new_n19574_, new_n4032_, RIbb31578_128 );
or   ( new_n19575_, new_n19574_, new_n3895_ );
nand ( new_n19576_, new_n19574_, new_n3892_ );
and  ( new_n19577_, new_n19576_, new_n19575_ );
nor  ( new_n19578_, new_n19577_, new_n19573_ );
or   ( new_n19579_, new_n4302_, new_n10841_ );
or   ( new_n19580_, new_n4304_, new_n10541_ );
and  ( new_n19581_, new_n19580_, new_n19579_ );
xor  ( new_n19582_, new_n19581_, new_n3895_ );
or   ( new_n19583_, new_n19582_, new_n19578_ );
and  ( new_n19584_, new_n19582_, new_n19578_ );
or   ( new_n19585_, new_n6173_, new_n8481_ );
or   ( new_n19586_, new_n6175_, new_n8352_ );
and  ( new_n19587_, new_n19586_, new_n19585_ );
xor  ( new_n19588_, new_n19587_, new_n5597_ );
or   ( new_n19589_, new_n5604_, new_n9099_ );
or   ( new_n19590_, new_n5606_, new_n8995_ );
and  ( new_n19591_, new_n19590_, new_n19589_ );
xor  ( new_n19592_, new_n19591_, new_n5206_ );
nor  ( new_n19593_, new_n19592_, new_n19588_ );
and  ( new_n19594_, new_n19592_, new_n19588_ );
or   ( new_n19595_, new_n5207_, new_n9679_ );
or   ( new_n19596_, new_n5209_, new_n9681_ );
and  ( new_n19597_, new_n19596_, new_n19595_ );
xor  ( new_n19598_, new_n19597_, new_n4708_ );
nor  ( new_n19599_, new_n19598_, new_n19594_ );
nor  ( new_n19600_, new_n19599_, new_n19593_ );
or   ( new_n19601_, new_n19600_, new_n19584_ );
and  ( new_n19602_, new_n19601_, new_n19583_ );
or   ( new_n19603_, new_n9422_, new_n5428_ );
or   ( new_n19604_, new_n9424_, new_n5171_ );
and  ( new_n19605_, new_n19604_, new_n19603_ );
xor  ( new_n19606_, new_n19605_, new_n8873_ );
or   ( new_n19607_, new_n8874_, new_n5899_ );
or   ( new_n19608_, new_n8876_, new_n5570_ );
and  ( new_n19609_, new_n19608_, new_n19607_ );
xor  ( new_n19610_, new_n19609_, new_n8257_ );
or   ( new_n19611_, new_n19610_, new_n19606_ );
and  ( new_n19612_, new_n19610_, new_n19606_ );
or   ( new_n19613_, new_n8264_, new_n6425_ );
or   ( new_n19614_, new_n8266_, new_n6219_ );
and  ( new_n19615_, new_n19614_, new_n19613_ );
xor  ( new_n19616_, new_n19615_, new_n7725_ );
or   ( new_n19617_, new_n19616_, new_n19612_ );
and  ( new_n19618_, new_n19617_, new_n19611_ );
or   ( new_n19619_, new_n10059_, new_n4859_ );
or   ( new_n19620_, new_n10061_, new_n4995_ );
and  ( new_n19621_, new_n19620_, new_n19619_ );
xor  ( new_n19622_, new_n19621_, new_n9421_ );
and  ( new_n19623_, RIbb2d888_64, RIbb2c5c8_104 );
or   ( new_n19624_, RIbb2d888_64, new_n4603_ );
and  ( new_n19625_, new_n19624_, RIbb2d900_63 );
or   ( new_n19626_, new_n19625_, new_n19623_ );
or   ( new_n19627_, new_n10770_, new_n4267_ );
and  ( new_n19628_, new_n19627_, new_n19626_ );
nor  ( new_n19629_, new_n19628_, new_n19622_ );
and  ( new_n19630_, new_n19628_, new_n19622_ );
nor  ( new_n19631_, new_n19630_, new_n3894_ );
nor  ( new_n19632_, new_n19631_, new_n19629_ );
or   ( new_n19633_, new_n7732_, new_n6943_ );
or   ( new_n19634_, new_n7734_, new_n6589_ );
and  ( new_n19635_, new_n19634_, new_n19633_ );
xor  ( new_n19636_, new_n19635_, new_n7177_ );
or   ( new_n19637_, new_n7184_, new_n7373_ );
or   ( new_n19638_, new_n7186_, new_n7149_ );
and  ( new_n19639_, new_n19638_, new_n19637_ );
xor  ( new_n19640_, new_n19639_, new_n6638_ );
or   ( new_n19641_, new_n19640_, new_n19636_ );
and  ( new_n19642_, new_n19640_, new_n19636_ );
or   ( new_n19643_, new_n6645_, new_n8115_ );
or   ( new_n19644_, new_n6647_, new_n8117_ );
and  ( new_n19645_, new_n19644_, new_n19643_ );
xor  ( new_n19646_, new_n19645_, new_n6166_ );
or   ( new_n19647_, new_n19646_, new_n19642_ );
and  ( new_n19648_, new_n19647_, new_n19641_ );
and  ( new_n19649_, new_n19648_, new_n19632_ );
or   ( new_n19650_, new_n19649_, new_n19618_ );
or   ( new_n19651_, new_n19648_, new_n19632_ );
and  ( new_n19652_, new_n19651_, new_n19650_ );
nand ( new_n19653_, new_n19652_, new_n19602_ );
nor  ( new_n19654_, new_n19652_, new_n19602_ );
xnor ( new_n19655_, new_n19461_, new_n19457_ );
xor  ( new_n19656_, new_n19655_, new_n19467_ );
xnor ( new_n19657_, new_n19499_, new_n19495_ );
xor  ( new_n19658_, new_n19657_, new_n19505_ );
nor  ( new_n19659_, new_n19658_, new_n19656_ );
and  ( new_n19660_, new_n19658_, new_n19656_ );
xor  ( new_n19661_, new_n19479_, new_n19475_ );
xnor ( new_n19662_, new_n19661_, new_n19485_ );
nor  ( new_n19663_, new_n19662_, new_n19660_ );
nor  ( new_n19664_, new_n19663_, new_n19659_ );
or   ( new_n19665_, new_n19664_, new_n19654_ );
and  ( new_n19666_, new_n19665_, new_n19653_ );
or   ( new_n19667_, new_n19666_, new_n19568_ );
and  ( new_n19668_, new_n19666_, new_n19568_ );
xor  ( new_n19669_, new_n19469_, new_n19453_ );
xor  ( new_n19670_, new_n19669_, new_n19487_ );
xnor ( new_n19671_, new_n19519_, new_n19517_ );
xor  ( new_n19672_, new_n19671_, new_n19523_ );
and  ( new_n19673_, new_n19672_, new_n19670_ );
nor  ( new_n19674_, new_n19672_, new_n19670_ );
xor  ( new_n19675_, new_n19507_, new_n19491_ );
xor  ( new_n19676_, new_n19675_, new_n19511_ );
nor  ( new_n19677_, new_n19676_, new_n19674_ );
nor  ( new_n19678_, new_n19677_, new_n19673_ );
or   ( new_n19679_, new_n19678_, new_n19668_ );
and  ( new_n19680_, new_n19679_, new_n19667_ );
or   ( new_n19681_, new_n19680_, new_n19566_ );
and  ( new_n19682_, new_n19681_, new_n19565_ );
or   ( new_n19683_, new_n19682_, new_n19552_ );
and  ( new_n19684_, new_n19682_, new_n19552_ );
xor  ( new_n19685_, new_n19531_, new_n19529_ );
xor  ( new_n19686_, new_n19685_, new_n19534_ );
or   ( new_n19687_, new_n19686_, new_n19684_ );
and  ( new_n19688_, new_n19687_, new_n19683_ );
nor  ( new_n19689_, new_n19688_, new_n19546_ );
xor  ( new_n19690_, new_n19682_, new_n19552_ );
xor  ( new_n19691_, new_n19690_, new_n19686_ );
xor  ( new_n19692_, new_n19564_, new_n19562_ );
xor  ( new_n19693_, new_n19692_, new_n19680_ );
xor  ( new_n19694_, new_n19672_, new_n19670_ );
xor  ( new_n19695_, new_n19694_, new_n19676_ );
xor  ( new_n19696_, new_n19658_, new_n19656_ );
xor  ( new_n19697_, new_n19696_, new_n19662_ );
xnor ( new_n19698_, new_n19582_, new_n19578_ );
xor  ( new_n19699_, new_n19698_, new_n19600_ );
or   ( new_n19700_, new_n19699_, new_n19697_ );
and  ( new_n19701_, new_n19699_, new_n19697_ );
xor  ( new_n19702_, new_n19445_, new_n19439_ );
xnor ( new_n19703_, new_n19702_, new_n19451_ );
or   ( new_n19704_, new_n19703_, new_n19701_ );
and  ( new_n19705_, new_n19704_, new_n19700_ );
nor  ( new_n19706_, new_n19705_, new_n19695_ );
nand ( new_n19707_, new_n19705_, new_n19695_ );
or   ( new_n19708_, new_n7184_, new_n8117_ );
or   ( new_n19709_, new_n7186_, new_n7373_ );
and  ( new_n19710_, new_n19709_, new_n19708_ );
xor  ( new_n19711_, new_n19710_, new_n6638_ );
or   ( new_n19712_, new_n6645_, new_n8352_ );
or   ( new_n19713_, new_n6647_, new_n8115_ );
and  ( new_n19714_, new_n19713_, new_n19712_ );
xor  ( new_n19715_, new_n19714_, new_n6166_ );
or   ( new_n19716_, new_n19715_, new_n19711_ );
and  ( new_n19717_, new_n19715_, new_n19711_ );
or   ( new_n19718_, new_n6173_, new_n8995_ );
or   ( new_n19719_, new_n6175_, new_n8481_ );
and  ( new_n19720_, new_n19719_, new_n19718_ );
xor  ( new_n19721_, new_n19720_, new_n5597_ );
or   ( new_n19722_, new_n19721_, new_n19717_ );
and  ( new_n19723_, new_n19722_, new_n19716_ );
or   ( new_n19724_, new_n8874_, new_n6219_ );
or   ( new_n19725_, new_n8876_, new_n5899_ );
and  ( new_n19726_, new_n19725_, new_n19724_ );
xor  ( new_n19727_, new_n19726_, new_n8257_ );
or   ( new_n19728_, new_n8264_, new_n6589_ );
or   ( new_n19729_, new_n8266_, new_n6425_ );
and  ( new_n19730_, new_n19729_, new_n19728_ );
xor  ( new_n19731_, new_n19730_, new_n7725_ );
or   ( new_n19732_, new_n19731_, new_n19727_ );
and  ( new_n19733_, new_n19731_, new_n19727_ );
or   ( new_n19734_, new_n7732_, new_n7149_ );
or   ( new_n19735_, new_n7734_, new_n6943_ );
and  ( new_n19736_, new_n19735_, new_n19734_ );
xor  ( new_n19737_, new_n19736_, new_n7177_ );
or   ( new_n19738_, new_n19737_, new_n19733_ );
and  ( new_n19739_, new_n19738_, new_n19732_ );
or   ( new_n19740_, new_n19739_, new_n19723_ );
and  ( new_n19741_, new_n19739_, new_n19723_ );
or   ( new_n19742_, new_n10059_, new_n5171_ );
or   ( new_n19743_, new_n10061_, new_n4859_ );
and  ( new_n19744_, new_n19743_, new_n19742_ );
xor  ( new_n19745_, new_n19744_, new_n9421_ );
and  ( new_n19746_, RIbb2d888_64, RIbb2c550_105 );
or   ( new_n19747_, RIbb2d888_64, new_n4995_ );
and  ( new_n19748_, new_n19747_, RIbb2d900_63 );
or   ( new_n19749_, new_n19748_, new_n19746_ );
or   ( new_n19750_, new_n10770_, new_n4603_ );
and  ( new_n19751_, new_n19750_, new_n19749_ );
or   ( new_n19752_, new_n19751_, new_n19745_ );
and  ( new_n19753_, new_n19751_, new_n19745_ );
or   ( new_n19754_, new_n9422_, new_n5570_ );
or   ( new_n19755_, new_n9424_, new_n5428_ );
and  ( new_n19756_, new_n19755_, new_n19754_ );
xor  ( new_n19757_, new_n19756_, new_n8873_ );
or   ( new_n19758_, new_n19757_, new_n19753_ );
and  ( new_n19759_, new_n19758_, new_n19752_ );
or   ( new_n19760_, new_n19759_, new_n19741_ );
and  ( new_n19761_, new_n19760_, new_n19740_ );
xor  ( new_n19762_, new_n19592_, new_n19588_ );
xor  ( new_n19763_, new_n19762_, new_n19598_ );
or   ( new_n19764_, new_n5604_, new_n9681_ );
or   ( new_n19765_, new_n5606_, new_n9099_ );
and  ( new_n19766_, new_n19765_, new_n19764_ );
xor  ( new_n19767_, new_n19766_, new_n5206_ );
or   ( new_n19768_, new_n5207_, new_n10220_ );
or   ( new_n19769_, new_n5209_, new_n9679_ );
and  ( new_n19770_, new_n19769_, new_n19768_ );
xor  ( new_n19771_, new_n19770_, new_n4708_ );
or   ( new_n19772_, new_n19771_, new_n19767_ );
and  ( new_n19773_, new_n19771_, new_n19767_ );
or   ( new_n19774_, new_n4709_, new_n10841_ );
or   ( new_n19775_, new_n4711_, new_n10541_ );
and  ( new_n19776_, new_n19775_, new_n19774_ );
xor  ( new_n19777_, new_n19776_, new_n4295_ );
or   ( new_n19778_, new_n19777_, new_n19773_ );
and  ( new_n19779_, new_n19778_, new_n19772_ );
or   ( new_n19780_, new_n19779_, new_n19763_ );
and  ( new_n19781_, new_n19779_, new_n19763_ );
xor  ( new_n19782_, new_n19577_, new_n19573_ );
or   ( new_n19783_, new_n19782_, new_n19781_ );
and  ( new_n19784_, new_n19783_, new_n19780_ );
and  ( new_n19785_, new_n19784_, new_n19761_ );
or   ( new_n19786_, new_n19784_, new_n19761_ );
xnor ( new_n19787_, new_n19610_, new_n19606_ );
xor  ( new_n19788_, new_n19787_, new_n19616_ );
xor  ( new_n19789_, new_n19628_, new_n19622_ );
xor  ( new_n19790_, new_n19789_, new_n3895_ );
nor  ( new_n19791_, new_n19790_, new_n19788_ );
and  ( new_n19792_, new_n19790_, new_n19788_ );
xor  ( new_n19793_, new_n19640_, new_n19636_ );
xnor ( new_n19794_, new_n19793_, new_n19646_ );
nor  ( new_n19795_, new_n19794_, new_n19792_ );
nor  ( new_n19796_, new_n19795_, new_n19791_ );
not  ( new_n19797_, new_n19796_ );
and  ( new_n19798_, new_n19797_, new_n19786_ );
or   ( new_n19799_, new_n19798_, new_n19785_ );
and  ( new_n19800_, new_n19799_, new_n19707_ );
or   ( new_n19801_, new_n19800_, new_n19706_ );
xnor ( new_n19802_, new_n19666_, new_n19568_ );
xor  ( new_n19803_, new_n19802_, new_n19678_ );
nand ( new_n19804_, new_n19803_, new_n19801_ );
nor  ( new_n19805_, new_n19803_, new_n19801_ );
xor  ( new_n19806_, new_n19556_, new_n19554_ );
xnor ( new_n19807_, new_n19806_, new_n19560_ );
or   ( new_n19808_, new_n19807_, new_n19805_ );
and  ( new_n19809_, new_n19808_, new_n19804_ );
or   ( new_n19810_, new_n19809_, new_n19693_ );
nand ( new_n19811_, new_n19809_, new_n19693_ );
xor  ( new_n19812_, new_n19551_, new_n19549_ );
nand ( new_n19813_, new_n19812_, new_n19811_ );
and  ( new_n19814_, new_n19813_, new_n19810_ );
nor  ( new_n19815_, new_n19814_, new_n19691_ );
xor  ( new_n19816_, new_n19784_, new_n19761_ );
xor  ( new_n19817_, new_n19816_, new_n19797_ );
xnor ( new_n19818_, new_n19699_, new_n19697_ );
xor  ( new_n19819_, new_n19818_, new_n19703_ );
nand ( new_n19820_, new_n19819_, new_n19817_ );
xnor ( new_n19821_, new_n19648_, new_n19632_ );
xor  ( new_n19822_, new_n19821_, new_n19618_ );
xor  ( new_n19823_, new_n19739_, new_n19723_ );
xor  ( new_n19824_, new_n19823_, new_n19759_ );
xnor ( new_n19825_, new_n19790_, new_n19788_ );
xor  ( new_n19826_, new_n19825_, new_n19794_ );
nand ( new_n19827_, new_n19826_, new_n19824_ );
nor  ( new_n19828_, new_n19826_, new_n19824_ );
xnor ( new_n19829_, new_n19779_, new_n19763_ );
xor  ( new_n19830_, new_n19829_, new_n19782_ );
or   ( new_n19831_, new_n19830_, new_n19828_ );
and  ( new_n19832_, new_n19831_, new_n19827_ );
or   ( new_n19833_, new_n19832_, new_n19822_ );
nand ( new_n19834_, new_n19832_, new_n19822_ );
xor  ( new_n19835_, new_n19731_, new_n19727_ );
xnor ( new_n19836_, new_n19835_, new_n19737_ );
xnor ( new_n19837_, new_n19751_, new_n19745_ );
xor  ( new_n19838_, new_n19837_, new_n19757_ );
nor  ( new_n19839_, new_n19838_, new_n19836_ );
or   ( new_n19840_, new_n9422_, new_n5899_ );
or   ( new_n19841_, new_n9424_, new_n5570_ );
and  ( new_n19842_, new_n19841_, new_n19840_ );
xor  ( new_n19843_, new_n19842_, new_n8873_ );
or   ( new_n19844_, new_n8874_, new_n6425_ );
or   ( new_n19845_, new_n8876_, new_n6219_ );
and  ( new_n19846_, new_n19845_, new_n19844_ );
xor  ( new_n19847_, new_n19846_, new_n8257_ );
or   ( new_n19848_, new_n19847_, new_n19843_ );
and  ( new_n19849_, new_n19847_, new_n19843_ );
or   ( new_n19850_, new_n8264_, new_n6943_ );
or   ( new_n19851_, new_n8266_, new_n6589_ );
and  ( new_n19852_, new_n19851_, new_n19850_ );
xor  ( new_n19853_, new_n19852_, new_n7725_ );
or   ( new_n19854_, new_n19853_, new_n19849_ );
and  ( new_n19855_, new_n19854_, new_n19848_ );
or   ( new_n19856_, new_n10059_, new_n5428_ );
or   ( new_n19857_, new_n10061_, new_n5171_ );
and  ( new_n19858_, new_n19857_, new_n19856_ );
xor  ( new_n19859_, new_n19858_, new_n9421_ );
and  ( new_n19860_, RIbb2d888_64, RIbb2c4d8_106 );
or   ( new_n19861_, RIbb2d888_64, new_n4859_ );
and  ( new_n19862_, new_n19861_, RIbb2d900_63 );
or   ( new_n19863_, new_n19862_, new_n19860_ );
or   ( new_n19864_, new_n10770_, new_n4995_ );
and  ( new_n19865_, new_n19864_, new_n19863_ );
nor  ( new_n19866_, new_n19865_, new_n19859_ );
and  ( new_n19867_, new_n19865_, new_n19859_ );
nor  ( new_n19868_, new_n19867_, new_n4294_ );
nor  ( new_n19869_, new_n19868_, new_n19866_ );
or   ( new_n19870_, new_n7732_, new_n7373_ );
or   ( new_n19871_, new_n7734_, new_n7149_ );
and  ( new_n19872_, new_n19871_, new_n19870_ );
xor  ( new_n19873_, new_n19872_, new_n7177_ );
or   ( new_n19874_, new_n7184_, new_n8115_ );
or   ( new_n19875_, new_n7186_, new_n8117_ );
and  ( new_n19876_, new_n19875_, new_n19874_ );
xor  ( new_n19877_, new_n19876_, new_n6638_ );
or   ( new_n19878_, new_n19877_, new_n19873_ );
and  ( new_n19879_, new_n19877_, new_n19873_ );
or   ( new_n19880_, new_n6645_, new_n8481_ );
or   ( new_n19881_, new_n6647_, new_n8352_ );
and  ( new_n19882_, new_n19881_, new_n19880_ );
xor  ( new_n19883_, new_n19882_, new_n6166_ );
or   ( new_n19884_, new_n19883_, new_n19879_ );
and  ( new_n19885_, new_n19884_, new_n19878_ );
and  ( new_n19886_, new_n19885_, new_n19869_ );
or   ( new_n19887_, new_n19886_, new_n19855_ );
or   ( new_n19888_, new_n19885_, new_n19869_ );
and  ( new_n19889_, new_n19888_, new_n19887_ );
nor  ( new_n19890_, new_n19889_, new_n19839_ );
and  ( new_n19891_, new_n19889_, new_n19839_ );
xor  ( new_n19892_, new_n19771_, new_n19767_ );
xor  ( new_n19893_, new_n19892_, new_n19777_ );
or   ( new_n19894_, new_n6173_, new_n9099_ );
or   ( new_n19895_, new_n6175_, new_n8995_ );
and  ( new_n19896_, new_n19895_, new_n19894_ );
xor  ( new_n19897_, new_n19896_, new_n5597_ );
or   ( new_n19898_, new_n5604_, new_n9679_ );
or   ( new_n19899_, new_n5606_, new_n9681_ );
and  ( new_n19900_, new_n19899_, new_n19898_ );
xor  ( new_n19901_, new_n19900_, new_n5206_ );
or   ( new_n19902_, new_n19901_, new_n19897_ );
and  ( new_n19903_, new_n19901_, new_n19897_ );
or   ( new_n19904_, new_n5207_, new_n10541_ );
or   ( new_n19905_, new_n5209_, new_n10220_ );
and  ( new_n19906_, new_n19905_, new_n19904_ );
xor  ( new_n19907_, new_n19906_, new_n4708_ );
or   ( new_n19908_, new_n19907_, new_n19903_ );
and  ( new_n19909_, new_n19908_, new_n19902_ );
nor  ( new_n19910_, new_n19909_, new_n19893_ );
and  ( new_n19911_, new_n19909_, new_n19893_ );
not  ( new_n19912_, new_n19911_ );
xor  ( new_n19913_, new_n19715_, new_n19711_ );
xnor ( new_n19914_, new_n19913_, new_n19721_ );
and  ( new_n19915_, new_n19914_, new_n19912_ );
nor  ( new_n19916_, new_n19915_, new_n19910_ );
nor  ( new_n19917_, new_n19916_, new_n19891_ );
nor  ( new_n19918_, new_n19917_, new_n19890_ );
nand ( new_n19919_, new_n19918_, new_n19834_ );
and  ( new_n19920_, new_n19919_, new_n19833_ );
nor  ( new_n19921_, new_n19920_, new_n19820_ );
nand ( new_n19922_, new_n19920_, new_n19820_ );
xor  ( new_n19923_, new_n19652_, new_n19602_ );
xnor ( new_n19924_, new_n19923_, new_n19664_ );
and  ( new_n19925_, new_n19924_, new_n19922_ );
or   ( new_n19926_, new_n19925_, new_n19921_ );
xnor ( new_n19927_, new_n19803_, new_n19801_ );
xor  ( new_n19928_, new_n19927_, new_n19807_ );
and  ( new_n19929_, new_n19928_, new_n19926_ );
xor  ( new_n19930_, new_n19809_, new_n19693_ );
xor  ( new_n19931_, new_n19930_, new_n19812_ );
and  ( new_n19932_, new_n19931_, new_n19929_ );
xor  ( new_n19933_, new_n19920_, new_n19820_ );
xnor ( new_n19934_, new_n19933_, new_n19924_ );
xor  ( new_n19935_, new_n19705_, new_n19695_ );
xnor ( new_n19936_, new_n19935_, new_n19799_ );
nor  ( new_n19937_, new_n19936_, new_n19934_ );
xor  ( new_n19938_, new_n19928_, new_n19926_ );
and  ( new_n19939_, new_n19938_, new_n19937_ );
xnor ( new_n19940_, new_n19936_, new_n19934_ );
xor  ( new_n19941_, new_n19826_, new_n19824_ );
xor  ( new_n19942_, new_n19941_, new_n19830_ );
xnor ( new_n19943_, new_n19885_, new_n19869_ );
xor  ( new_n19944_, new_n19943_, new_n19855_ );
xor  ( new_n19945_, new_n19909_, new_n19893_ );
xor  ( new_n19946_, new_n19945_, new_n19914_ );
or   ( new_n19947_, new_n19946_, new_n19944_ );
and  ( new_n19948_, new_n19946_, new_n19944_ );
xnor ( new_n19949_, new_n19838_, new_n19836_ );
or   ( new_n19950_, new_n19949_, new_n19948_ );
and  ( new_n19951_, new_n19950_, new_n19947_ );
nor  ( new_n19952_, new_n19951_, new_n19942_ );
and  ( new_n19953_, new_n19951_, new_n19942_ );
xor  ( new_n19954_, new_n19847_, new_n19843_ );
xnor ( new_n19955_, new_n19954_, new_n19853_ );
xor  ( new_n19956_, new_n19865_, new_n19859_ );
xor  ( new_n19957_, new_n19956_, new_n4295_ );
nor  ( new_n19958_, new_n19957_, new_n19955_ );
or   ( new_n19959_, new_n7184_, new_n8352_ );
or   ( new_n19960_, new_n7186_, new_n8115_ );
and  ( new_n19961_, new_n19960_, new_n19959_ );
xor  ( new_n19962_, new_n19961_, new_n6638_ );
or   ( new_n19963_, new_n6645_, new_n8995_ );
or   ( new_n19964_, new_n6647_, new_n8481_ );
and  ( new_n19965_, new_n19964_, new_n19963_ );
xor  ( new_n19966_, new_n19965_, new_n6166_ );
or   ( new_n19967_, new_n19966_, new_n19962_ );
and  ( new_n19968_, new_n19966_, new_n19962_ );
or   ( new_n19969_, new_n6173_, new_n9681_ );
or   ( new_n19970_, new_n6175_, new_n9099_ );
and  ( new_n19971_, new_n19970_, new_n19969_ );
xor  ( new_n19972_, new_n19971_, new_n5597_ );
or   ( new_n19973_, new_n19972_, new_n19968_ );
and  ( new_n19974_, new_n19973_, new_n19967_ );
or   ( new_n19975_, new_n10059_, new_n5570_ );
or   ( new_n19976_, new_n10061_, new_n5428_ );
and  ( new_n19977_, new_n19976_, new_n19975_ );
xor  ( new_n19978_, new_n19977_, new_n9421_ );
and  ( new_n19979_, RIbb2d888_64, RIbb2c460_107 );
or   ( new_n19980_, RIbb2d888_64, new_n5171_ );
and  ( new_n19981_, new_n19980_, RIbb2d900_63 );
or   ( new_n19982_, new_n19981_, new_n19979_ );
or   ( new_n19983_, new_n10770_, new_n4859_ );
and  ( new_n19984_, new_n19983_, new_n19982_ );
or   ( new_n19985_, new_n19984_, new_n19978_ );
and  ( new_n19986_, new_n19984_, new_n19978_ );
or   ( new_n19987_, new_n9422_, new_n6219_ );
or   ( new_n19988_, new_n9424_, new_n5899_ );
and  ( new_n19989_, new_n19988_, new_n19987_ );
xor  ( new_n19990_, new_n19989_, new_n8873_ );
or   ( new_n19991_, new_n19990_, new_n19986_ );
and  ( new_n19992_, new_n19991_, new_n19985_ );
or   ( new_n19993_, new_n19992_, new_n19974_ );
and  ( new_n19994_, new_n19992_, new_n19974_ );
or   ( new_n19995_, new_n8874_, new_n6589_ );
or   ( new_n19996_, new_n8876_, new_n6425_ );
and  ( new_n19997_, new_n19996_, new_n19995_ );
xor  ( new_n19998_, new_n19997_, new_n8257_ );
or   ( new_n19999_, new_n8264_, new_n7149_ );
or   ( new_n20000_, new_n8266_, new_n6943_ );
and  ( new_n20001_, new_n20000_, new_n19999_ );
xor  ( new_n20002_, new_n20001_, new_n7725_ );
or   ( new_n20003_, new_n20002_, new_n19998_ );
and  ( new_n20004_, new_n20002_, new_n19998_ );
or   ( new_n20005_, new_n7732_, new_n8117_ );
or   ( new_n20006_, new_n7734_, new_n7373_ );
and  ( new_n20007_, new_n20006_, new_n20005_ );
xor  ( new_n20008_, new_n20007_, new_n7177_ );
or   ( new_n20009_, new_n20008_, new_n20004_ );
and  ( new_n20010_, new_n20009_, new_n20003_ );
or   ( new_n20011_, new_n20010_, new_n19994_ );
and  ( new_n20012_, new_n20011_, new_n19993_ );
and  ( new_n20013_, new_n20012_, new_n19958_ );
nor  ( new_n20014_, new_n20012_, new_n19958_ );
and  ( new_n20015_, new_n4541_, RIbb31578_128 );
or   ( new_n20016_, new_n20015_, new_n4295_ );
nand ( new_n20017_, new_n20015_, new_n4292_ );
and  ( new_n20018_, new_n20017_, new_n20016_ );
xnor ( new_n20019_, new_n19901_, new_n19897_ );
xor  ( new_n20020_, new_n20019_, new_n19907_ );
nor  ( new_n20021_, new_n20020_, new_n20018_ );
and  ( new_n20022_, new_n20020_, new_n20018_ );
xor  ( new_n20023_, new_n19877_, new_n19873_ );
xnor ( new_n20024_, new_n20023_, new_n19883_ );
nor  ( new_n20025_, new_n20024_, new_n20022_ );
nor  ( new_n20026_, new_n20025_, new_n20021_ );
nor  ( new_n20027_, new_n20026_, new_n20014_ );
nor  ( new_n20028_, new_n20027_, new_n20013_ );
nor  ( new_n20029_, new_n20028_, new_n19953_ );
or   ( new_n20030_, new_n20029_, new_n19952_ );
xor  ( new_n20031_, new_n19832_, new_n19822_ );
xor  ( new_n20032_, new_n20031_, new_n19918_ );
nand ( new_n20033_, new_n20032_, new_n20030_ );
nor  ( new_n20034_, new_n20032_, new_n20030_ );
xnor ( new_n20035_, new_n19819_, new_n19817_ );
or   ( new_n20036_, new_n20035_, new_n20034_ );
and  ( new_n20037_, new_n20036_, new_n20033_ );
nor  ( new_n20038_, new_n20037_, new_n19940_ );
xor  ( new_n20039_, new_n20032_, new_n20030_ );
xor  ( new_n20040_, new_n20039_, new_n20035_ );
xor  ( new_n20041_, new_n19951_, new_n19942_ );
xor  ( new_n20042_, new_n20041_, new_n20028_ );
xnor ( new_n20043_, new_n19889_, new_n19839_ );
xor  ( new_n20044_, new_n20043_, new_n19916_ );
or   ( new_n20045_, new_n20044_, new_n20042_ );
and  ( new_n20046_, new_n20044_, new_n20042_ );
xor  ( new_n20047_, new_n19946_, new_n19944_ );
xor  ( new_n20048_, new_n20047_, new_n19949_ );
xor  ( new_n20049_, new_n19992_, new_n19974_ );
xor  ( new_n20050_, new_n20049_, new_n20010_ );
xnor ( new_n20051_, new_n20020_, new_n20018_ );
xor  ( new_n20052_, new_n20051_, new_n20024_ );
nand ( new_n20053_, new_n20052_, new_n20050_ );
or   ( new_n20054_, new_n20052_, new_n20050_ );
xor  ( new_n20055_, new_n19957_, new_n19955_ );
nand ( new_n20056_, new_n20055_, new_n20054_ );
and  ( new_n20057_, new_n20056_, new_n20053_ );
nor  ( new_n20058_, new_n20057_, new_n20048_ );
and  ( new_n20059_, new_n20057_, new_n20048_ );
or   ( new_n20060_, new_n10059_, new_n5899_ );
or   ( new_n20061_, new_n10061_, new_n5570_ );
and  ( new_n20062_, new_n20061_, new_n20060_ );
xor  ( new_n20063_, new_n20062_, new_n9421_ );
and  ( new_n20064_, RIbb2d888_64, RIbb2c3e8_108 );
or   ( new_n20065_, RIbb2d888_64, new_n5428_ );
and  ( new_n20066_, new_n20065_, RIbb2d900_63 );
or   ( new_n20067_, new_n20066_, new_n20064_ );
or   ( new_n20068_, new_n10770_, new_n5171_ );
and  ( new_n20069_, new_n20068_, new_n20067_ );
or   ( new_n20070_, new_n20069_, new_n20063_ );
and  ( new_n20071_, new_n20069_, new_n20063_ );
or   ( new_n20072_, new_n20071_, new_n4707_ );
and  ( new_n20073_, new_n20072_, new_n20070_ );
or   ( new_n20074_, new_n9422_, new_n6425_ );
or   ( new_n20075_, new_n9424_, new_n6219_ );
and  ( new_n20076_, new_n20075_, new_n20074_ );
xor  ( new_n20077_, new_n20076_, new_n8873_ );
or   ( new_n20078_, new_n8874_, new_n6943_ );
or   ( new_n20079_, new_n8876_, new_n6589_ );
and  ( new_n20080_, new_n20079_, new_n20078_ );
xor  ( new_n20081_, new_n20080_, new_n8257_ );
or   ( new_n20082_, new_n20081_, new_n20077_ );
and  ( new_n20083_, new_n20081_, new_n20077_ );
or   ( new_n20084_, new_n8264_, new_n7373_ );
or   ( new_n20085_, new_n8266_, new_n7149_ );
and  ( new_n20086_, new_n20085_, new_n20084_ );
xor  ( new_n20087_, new_n20086_, new_n7725_ );
or   ( new_n20088_, new_n20087_, new_n20083_ );
and  ( new_n20089_, new_n20088_, new_n20082_ );
nor  ( new_n20090_, new_n20089_, new_n20073_ );
nand ( new_n20091_, new_n20089_, new_n20073_ );
or   ( new_n20092_, new_n7732_, new_n8115_ );
or   ( new_n20093_, new_n7734_, new_n8117_ );
and  ( new_n20094_, new_n20093_, new_n20092_ );
xor  ( new_n20095_, new_n20094_, new_n7177_ );
or   ( new_n20096_, new_n7184_, new_n8481_ );
or   ( new_n20097_, new_n7186_, new_n8352_ );
and  ( new_n20098_, new_n20097_, new_n20096_ );
xor  ( new_n20099_, new_n20098_, new_n6638_ );
nor  ( new_n20100_, new_n20099_, new_n20095_ );
and  ( new_n20101_, new_n20099_, new_n20095_ );
or   ( new_n20102_, new_n6645_, new_n9099_ );
or   ( new_n20103_, new_n6647_, new_n8995_ );
and  ( new_n20104_, new_n20103_, new_n20102_ );
xor  ( new_n20105_, new_n20104_, new_n6166_ );
nor  ( new_n20106_, new_n20105_, new_n20101_ );
nor  ( new_n20107_, new_n20106_, new_n20100_ );
not  ( new_n20108_, new_n20107_ );
and  ( new_n20109_, new_n20108_, new_n20091_ );
or   ( new_n20110_, new_n20109_, new_n20090_ );
xnor ( new_n20111_, new_n19984_, new_n19978_ );
xor  ( new_n20112_, new_n20111_, new_n19990_ );
xnor ( new_n20113_, new_n19966_, new_n19962_ );
xor  ( new_n20114_, new_n20113_, new_n19972_ );
or   ( new_n20115_, new_n20114_, new_n20112_ );
and  ( new_n20116_, new_n20114_, new_n20112_ );
xor  ( new_n20117_, new_n20002_, new_n19998_ );
xnor ( new_n20118_, new_n20117_, new_n20008_ );
or   ( new_n20119_, new_n20118_, new_n20116_ );
and  ( new_n20120_, new_n20119_, new_n20115_ );
nor  ( new_n20121_, new_n20120_, new_n20110_ );
and  ( new_n20122_, new_n20120_, new_n20110_ );
or   ( new_n20123_, new_n5604_, new_n10220_ );
or   ( new_n20124_, new_n5606_, new_n9679_ );
and  ( new_n20125_, new_n20124_, new_n20123_ );
xor  ( new_n20126_, new_n20125_, new_n5205_ );
or   ( new_n20127_, new_n6173_, new_n9679_ );
or   ( new_n20128_, new_n6175_, new_n9681_ );
and  ( new_n20129_, new_n20128_, new_n20127_ );
xor  ( new_n20130_, new_n20129_, new_n5597_ );
or   ( new_n20131_, new_n5604_, new_n10541_ );
or   ( new_n20132_, new_n5606_, new_n10220_ );
and  ( new_n20133_, new_n20132_, new_n20131_ );
xor  ( new_n20134_, new_n20133_, new_n5206_ );
nand ( new_n20135_, new_n20134_, new_n20130_ );
nor  ( new_n20136_, new_n20134_, new_n20130_ );
and  ( new_n20137_, new_n4958_, RIbb31578_128 );
nor  ( new_n20138_, new_n20137_, new_n4708_ );
and  ( new_n20139_, new_n20137_, new_n4705_ );
nor  ( new_n20140_, new_n20139_, new_n20138_ );
or   ( new_n20141_, new_n20140_, new_n20136_ );
and  ( new_n20142_, new_n20141_, new_n20135_ );
nor  ( new_n20143_, new_n20142_, new_n20126_ );
and  ( new_n20144_, new_n20142_, new_n20126_ );
or   ( new_n20145_, new_n5207_, new_n10841_ );
or   ( new_n20146_, new_n5209_, new_n10541_ );
and  ( new_n20147_, new_n20146_, new_n20145_ );
xor  ( new_n20148_, new_n20147_, new_n4708_ );
not  ( new_n20149_, new_n20148_ );
nor  ( new_n20150_, new_n20149_, new_n20144_ );
nor  ( new_n20151_, new_n20150_, new_n20143_ );
nor  ( new_n20152_, new_n20151_, new_n20122_ );
nor  ( new_n20153_, new_n20152_, new_n20121_ );
nor  ( new_n20154_, new_n20153_, new_n20059_ );
nor  ( new_n20155_, new_n20154_, new_n20058_ );
or   ( new_n20156_, new_n20155_, new_n20046_ );
and  ( new_n20157_, new_n20156_, new_n20045_ );
nor  ( new_n20158_, new_n20157_, new_n20040_ );
xnor ( new_n20159_, new_n20057_, new_n20048_ );
xor  ( new_n20160_, new_n20159_, new_n20153_ );
xnor ( new_n20161_, new_n20012_, new_n19958_ );
xor  ( new_n20162_, new_n20161_, new_n20026_ );
and  ( new_n20163_, new_n20162_, new_n20160_ );
nor  ( new_n20164_, new_n20162_, new_n20160_ );
or   ( new_n20165_, new_n10059_, new_n6219_ );
or   ( new_n20166_, new_n10061_, new_n5899_ );
and  ( new_n20167_, new_n20166_, new_n20165_ );
xor  ( new_n20168_, new_n20167_, new_n9421_ );
and  ( new_n20169_, RIbb2d888_64, RIbb2c370_109 );
or   ( new_n20170_, RIbb2d888_64, new_n5570_ );
and  ( new_n20171_, new_n20170_, RIbb2d900_63 );
or   ( new_n20172_, new_n20171_, new_n20169_ );
or   ( new_n20173_, new_n10770_, new_n5428_ );
and  ( new_n20174_, new_n20173_, new_n20172_ );
or   ( new_n20175_, new_n20174_, new_n20168_ );
and  ( new_n20176_, new_n20174_, new_n20168_ );
or   ( new_n20177_, new_n9422_, new_n6589_ );
or   ( new_n20178_, new_n9424_, new_n6425_ );
and  ( new_n20179_, new_n20178_, new_n20177_ );
xor  ( new_n20180_, new_n20179_, new_n8873_ );
or   ( new_n20181_, new_n20180_, new_n20176_ );
and  ( new_n20182_, new_n20181_, new_n20175_ );
or   ( new_n20183_, new_n7184_, new_n8995_ );
or   ( new_n20184_, new_n7186_, new_n8481_ );
and  ( new_n20185_, new_n20184_, new_n20183_ );
xor  ( new_n20186_, new_n20185_, new_n6638_ );
or   ( new_n20187_, new_n6645_, new_n9681_ );
or   ( new_n20188_, new_n6647_, new_n9099_ );
and  ( new_n20189_, new_n20188_, new_n20187_ );
xor  ( new_n20190_, new_n20189_, new_n6166_ );
or   ( new_n20191_, new_n20190_, new_n20186_ );
and  ( new_n20192_, new_n20190_, new_n20186_ );
or   ( new_n20193_, new_n6173_, new_n10220_ );
or   ( new_n20194_, new_n6175_, new_n9679_ );
and  ( new_n20195_, new_n20194_, new_n20193_ );
xor  ( new_n20196_, new_n20195_, new_n5597_ );
or   ( new_n20197_, new_n20196_, new_n20192_ );
and  ( new_n20198_, new_n20197_, new_n20191_ );
or   ( new_n20199_, new_n20198_, new_n20182_ );
and  ( new_n20200_, new_n20198_, new_n20182_ );
or   ( new_n20201_, new_n8874_, new_n7149_ );
or   ( new_n20202_, new_n8876_, new_n6943_ );
and  ( new_n20203_, new_n20202_, new_n20201_ );
xor  ( new_n20204_, new_n20203_, new_n8257_ );
or   ( new_n20205_, new_n8264_, new_n8117_ );
or   ( new_n20206_, new_n8266_, new_n7373_ );
and  ( new_n20207_, new_n20206_, new_n20205_ );
xor  ( new_n20208_, new_n20207_, new_n7725_ );
nor  ( new_n20209_, new_n20208_, new_n20204_ );
and  ( new_n20210_, new_n20208_, new_n20204_ );
or   ( new_n20211_, new_n7732_, new_n8352_ );
or   ( new_n20212_, new_n7734_, new_n8115_ );
and  ( new_n20213_, new_n20212_, new_n20211_ );
xor  ( new_n20214_, new_n20213_, new_n7177_ );
nor  ( new_n20215_, new_n20214_, new_n20210_ );
nor  ( new_n20216_, new_n20215_, new_n20209_ );
or   ( new_n20217_, new_n20216_, new_n20200_ );
and  ( new_n20218_, new_n20217_, new_n20199_ );
xnor ( new_n20219_, new_n20114_, new_n20112_ );
xor  ( new_n20220_, new_n20219_, new_n20118_ );
or   ( new_n20221_, new_n20220_, new_n20218_ );
nand ( new_n20222_, new_n20220_, new_n20218_ );
xor  ( new_n20223_, new_n20081_, new_n20077_ );
xor  ( new_n20224_, new_n20223_, new_n20087_ );
xnor ( new_n20225_, new_n20134_, new_n20130_ );
xor  ( new_n20226_, new_n20225_, new_n20140_ );
and  ( new_n20227_, new_n20226_, new_n20224_ );
nor  ( new_n20228_, new_n20226_, new_n20224_ );
xor  ( new_n20229_, new_n20099_, new_n20095_ );
xnor ( new_n20230_, new_n20229_, new_n20105_ );
nor  ( new_n20231_, new_n20230_, new_n20228_ );
nor  ( new_n20232_, new_n20231_, new_n20227_ );
nand ( new_n20233_, new_n20232_, new_n20222_ );
and  ( new_n20234_, new_n20233_, new_n20221_ );
xnor ( new_n20235_, new_n20120_, new_n20110_ );
xor  ( new_n20236_, new_n20235_, new_n20151_ );
and  ( new_n20237_, new_n20236_, new_n20234_ );
nor  ( new_n20238_, new_n20236_, new_n20234_ );
xor  ( new_n20239_, new_n20052_, new_n20050_ );
xor  ( new_n20240_, new_n20239_, new_n20055_ );
not  ( new_n20241_, new_n20240_ );
nor  ( new_n20242_, new_n20241_, new_n20238_ );
nor  ( new_n20243_, new_n20242_, new_n20237_ );
nor  ( new_n20244_, new_n20243_, new_n20164_ );
or   ( new_n20245_, new_n20244_, new_n20163_ );
xnor ( new_n20246_, new_n20044_, new_n20042_ );
xor  ( new_n20247_, new_n20246_, new_n20155_ );
and  ( new_n20248_, new_n20247_, new_n20245_ );
xor  ( new_n20249_, new_n20162_, new_n20160_ );
xor  ( new_n20250_, new_n20249_, new_n20243_ );
xor  ( new_n20251_, new_n20089_, new_n20073_ );
xor  ( new_n20252_, new_n20251_, new_n20108_ );
xor  ( new_n20253_, new_n20220_, new_n20218_ );
xor  ( new_n20254_, new_n20253_, new_n20232_ );
or   ( new_n20255_, new_n20254_, new_n20252_ );
xor  ( new_n20256_, new_n20198_, new_n20182_ );
xnor ( new_n20257_, new_n20256_, new_n20216_ );
xnor ( new_n20258_, new_n20226_, new_n20224_ );
xnor ( new_n20259_, new_n20258_, new_n20230_ );
nor  ( new_n20260_, new_n20259_, new_n20257_ );
xor  ( new_n20261_, new_n20069_, new_n20063_ );
xor  ( new_n20262_, new_n20261_, new_n4707_ );
or   ( new_n20263_, new_n5604_, new_n10841_ );
or   ( new_n20264_, new_n5606_, new_n10541_ );
and  ( new_n20265_, new_n20264_, new_n20263_ );
xor  ( new_n20266_, new_n20265_, new_n5205_ );
xnor ( new_n20267_, new_n20190_, new_n20186_ );
xor  ( new_n20268_, new_n20267_, new_n20196_ );
nand ( new_n20269_, new_n20268_, new_n20266_ );
nor  ( new_n20270_, new_n20268_, new_n20266_ );
xor  ( new_n20271_, new_n20208_, new_n20204_ );
xor  ( new_n20272_, new_n20271_, new_n20214_ );
or   ( new_n20273_, new_n20272_, new_n20270_ );
and  ( new_n20274_, new_n20273_, new_n20269_ );
or   ( new_n20275_, new_n20274_, new_n20262_ );
and  ( new_n20276_, new_n20274_, new_n20262_ );
or   ( new_n20277_, new_n10059_, new_n6425_ );
or   ( new_n20278_, new_n10061_, new_n6219_ );
and  ( new_n20279_, new_n20278_, new_n20277_ );
xor  ( new_n20280_, new_n20279_, new_n9421_ );
and  ( new_n20281_, RIbb2d888_64, RIbb2c2f8_110 );
or   ( new_n20282_, RIbb2d888_64, new_n5899_ );
and  ( new_n20283_, new_n20282_, RIbb2d900_63 );
or   ( new_n20284_, new_n20283_, new_n20281_ );
or   ( new_n20285_, new_n10770_, new_n5570_ );
and  ( new_n20286_, new_n20285_, new_n20284_ );
or   ( new_n20287_, new_n20286_, new_n20280_ );
and  ( new_n20288_, new_n20286_, new_n20280_ );
or   ( new_n20289_, new_n20288_, new_n5205_ );
and  ( new_n20290_, new_n20289_, new_n20287_ );
or   ( new_n20291_, new_n7732_, new_n8481_ );
or   ( new_n20292_, new_n7734_, new_n8352_ );
and  ( new_n20293_, new_n20292_, new_n20291_ );
xor  ( new_n20294_, new_n20293_, new_n7177_ );
or   ( new_n20295_, new_n7184_, new_n9099_ );
or   ( new_n20296_, new_n7186_, new_n8995_ );
and  ( new_n20297_, new_n20296_, new_n20295_ );
xor  ( new_n20298_, new_n20297_, new_n6638_ );
or   ( new_n20299_, new_n20298_, new_n20294_ );
and  ( new_n20300_, new_n20298_, new_n20294_ );
or   ( new_n20301_, new_n6645_, new_n9679_ );
or   ( new_n20302_, new_n6647_, new_n9681_ );
and  ( new_n20303_, new_n20302_, new_n20301_ );
xor  ( new_n20304_, new_n20303_, new_n6166_ );
or   ( new_n20305_, new_n20304_, new_n20300_ );
and  ( new_n20306_, new_n20305_, new_n20299_ );
nor  ( new_n20307_, new_n20306_, new_n20290_ );
and  ( new_n20308_, new_n20306_, new_n20290_ );
or   ( new_n20309_, new_n9422_, new_n6943_ );
or   ( new_n20310_, new_n9424_, new_n6589_ );
and  ( new_n20311_, new_n20310_, new_n20309_ );
xor  ( new_n20312_, new_n20311_, new_n8873_ );
or   ( new_n20313_, new_n8874_, new_n7373_ );
or   ( new_n20314_, new_n8876_, new_n7149_ );
and  ( new_n20315_, new_n20314_, new_n20313_ );
xor  ( new_n20316_, new_n20315_, new_n8257_ );
nor  ( new_n20317_, new_n20316_, new_n20312_ );
and  ( new_n20318_, new_n20316_, new_n20312_ );
or   ( new_n20319_, new_n8264_, new_n8115_ );
or   ( new_n20320_, new_n8266_, new_n8117_ );
and  ( new_n20321_, new_n20320_, new_n20319_ );
xor  ( new_n20322_, new_n20321_, new_n7725_ );
nor  ( new_n20323_, new_n20322_, new_n20318_ );
nor  ( new_n20324_, new_n20323_, new_n20317_ );
nor  ( new_n20325_, new_n20324_, new_n20308_ );
nor  ( new_n20326_, new_n20325_, new_n20307_ );
or   ( new_n20327_, new_n20326_, new_n20276_ );
and  ( new_n20328_, new_n20327_, new_n20275_ );
nand ( new_n20329_, new_n20328_, new_n20260_ );
nor  ( new_n20330_, new_n20328_, new_n20260_ );
xor  ( new_n20331_, new_n20142_, new_n20126_ );
xor  ( new_n20332_, new_n20331_, new_n20149_ );
or   ( new_n20333_, new_n20332_, new_n20330_ );
and  ( new_n20334_, new_n20333_, new_n20329_ );
or   ( new_n20335_, new_n20334_, new_n20255_ );
and  ( new_n20336_, new_n20334_, new_n20255_ );
xor  ( new_n20337_, new_n20236_, new_n20234_ );
xor  ( new_n20338_, new_n20337_, new_n20241_ );
or   ( new_n20339_, new_n20338_, new_n20336_ );
and  ( new_n20340_, new_n20339_, new_n20335_ );
nor  ( new_n20341_, new_n20340_, new_n20250_ );
xor  ( new_n20342_, new_n20334_, new_n20255_ );
xor  ( new_n20343_, new_n20342_, new_n20338_ );
xor  ( new_n20344_, new_n20328_, new_n20260_ );
xor  ( new_n20345_, new_n20344_, new_n20332_ );
xor  ( new_n20346_, new_n20174_, new_n20168_ );
xor  ( new_n20347_, new_n20346_, new_n20180_ );
or   ( new_n20348_, new_n6173_, new_n10541_ );
or   ( new_n20349_, new_n6175_, new_n10220_ );
and  ( new_n20350_, new_n20349_, new_n20348_ );
xor  ( new_n20351_, new_n20350_, new_n5596_ );
and  ( new_n20352_, new_n5371_, RIbb31578_128 );
or   ( new_n20353_, new_n20352_, new_n5206_ );
nand ( new_n20354_, new_n20352_, new_n5203_ );
and  ( new_n20355_, new_n20354_, new_n20353_ );
nand ( new_n20356_, new_n20355_, new_n20351_ );
or   ( new_n20357_, new_n20355_, new_n20351_ );
xor  ( new_n20358_, new_n20298_, new_n20294_ );
xnor ( new_n20359_, new_n20358_, new_n20304_ );
nand ( new_n20360_, new_n20359_, new_n20357_ );
and  ( new_n20361_, new_n20360_, new_n20356_ );
nor  ( new_n20362_, new_n20361_, new_n20347_ );
nand ( new_n20363_, new_n20361_, new_n20347_ );
or   ( new_n20364_, new_n10059_, new_n6589_ );
or   ( new_n20365_, new_n10061_, new_n6425_ );
and  ( new_n20366_, new_n20365_, new_n20364_ );
xor  ( new_n20367_, new_n20366_, new_n9421_ );
and  ( new_n20368_, RIbb2d888_64, RIbb2c280_111 );
or   ( new_n20369_, RIbb2d888_64, new_n6219_ );
and  ( new_n20370_, new_n20369_, RIbb2d900_63 );
or   ( new_n20371_, new_n20370_, new_n20368_ );
or   ( new_n20372_, new_n10770_, new_n5899_ );
and  ( new_n20373_, new_n20372_, new_n20371_ );
or   ( new_n20374_, new_n20373_, new_n20367_ );
and  ( new_n20375_, new_n20373_, new_n20367_ );
or   ( new_n20376_, new_n9422_, new_n7149_ );
or   ( new_n20377_, new_n9424_, new_n6943_ );
and  ( new_n20378_, new_n20377_, new_n20376_ );
xor  ( new_n20379_, new_n20378_, new_n8873_ );
or   ( new_n20380_, new_n20379_, new_n20375_ );
and  ( new_n20381_, new_n20380_, new_n20374_ );
or   ( new_n20382_, new_n8874_, new_n8117_ );
or   ( new_n20383_, new_n8876_, new_n7373_ );
and  ( new_n20384_, new_n20383_, new_n20382_ );
xor  ( new_n20385_, new_n20384_, new_n8257_ );
or   ( new_n20386_, new_n8264_, new_n8352_ );
or   ( new_n20387_, new_n8266_, new_n8115_ );
and  ( new_n20388_, new_n20387_, new_n20386_ );
xor  ( new_n20389_, new_n20388_, new_n7725_ );
or   ( new_n20390_, new_n20389_, new_n20385_ );
and  ( new_n20391_, new_n20389_, new_n20385_ );
or   ( new_n20392_, new_n7732_, new_n8995_ );
or   ( new_n20393_, new_n7734_, new_n8481_ );
and  ( new_n20394_, new_n20393_, new_n20392_ );
xor  ( new_n20395_, new_n20394_, new_n7177_ );
or   ( new_n20396_, new_n20395_, new_n20391_ );
and  ( new_n20397_, new_n20396_, new_n20390_ );
nor  ( new_n20398_, new_n20397_, new_n20381_ );
nand ( new_n20399_, new_n20397_, new_n20381_ );
or   ( new_n20400_, new_n7184_, new_n9681_ );
or   ( new_n20401_, new_n7186_, new_n9099_ );
and  ( new_n20402_, new_n20401_, new_n20400_ );
xor  ( new_n20403_, new_n20402_, new_n6638_ );
or   ( new_n20404_, new_n6645_, new_n10220_ );
or   ( new_n20405_, new_n6647_, new_n9679_ );
and  ( new_n20406_, new_n20405_, new_n20404_ );
xor  ( new_n20407_, new_n20406_, new_n6166_ );
nor  ( new_n20408_, new_n20407_, new_n20403_ );
nand ( new_n20409_, new_n20407_, new_n20403_ );
or   ( new_n20410_, new_n6173_, new_n10841_ );
or   ( new_n20411_, new_n6175_, new_n10541_ );
and  ( new_n20412_, new_n20411_, new_n20410_ );
xor  ( new_n20413_, new_n20412_, new_n5597_ );
not  ( new_n20414_, new_n20413_ );
and  ( new_n20415_, new_n20414_, new_n20409_ );
or   ( new_n20416_, new_n20415_, new_n20408_ );
and  ( new_n20417_, new_n20416_, new_n20399_ );
or   ( new_n20418_, new_n20417_, new_n20398_ );
and  ( new_n20419_, new_n20418_, new_n20363_ );
or   ( new_n20420_, new_n20419_, new_n20362_ );
xnor ( new_n20421_, new_n20274_, new_n20262_ );
xor  ( new_n20422_, new_n20421_, new_n20326_ );
or   ( new_n20423_, new_n20422_, new_n20420_ );
and  ( new_n20424_, new_n20422_, new_n20420_ );
xnor ( new_n20425_, new_n20259_, new_n20257_ );
or   ( new_n20426_, new_n20425_, new_n20424_ );
and  ( new_n20427_, new_n20426_, new_n20423_ );
or   ( new_n20428_, new_n20427_, new_n20345_ );
and  ( new_n20429_, new_n20427_, new_n20345_ );
xnor ( new_n20430_, new_n20254_, new_n20252_ );
or   ( new_n20431_, new_n20430_, new_n20429_ );
and  ( new_n20432_, new_n20431_, new_n20428_ );
nor  ( new_n20433_, new_n20432_, new_n20343_ );
xor  ( new_n20434_, new_n20427_, new_n20345_ );
xor  ( new_n20435_, new_n20434_, new_n20430_ );
xor  ( new_n20436_, new_n20306_, new_n20290_ );
xnor ( new_n20437_, new_n20436_, new_n20324_ );
xor  ( new_n20438_, new_n20361_, new_n20347_ );
xor  ( new_n20439_, new_n20438_, new_n20418_ );
nor  ( new_n20440_, new_n20439_, new_n20437_ );
xor  ( new_n20441_, new_n20268_, new_n20266_ );
xor  ( new_n20442_, new_n20441_, new_n20272_ );
xor  ( new_n20443_, new_n20316_, new_n20312_ );
xor  ( new_n20444_, new_n20443_, new_n20322_ );
or   ( new_n20445_, new_n9422_, new_n7373_ );
or   ( new_n20446_, new_n9424_, new_n7149_ );
and  ( new_n20447_, new_n20446_, new_n20445_ );
xor  ( new_n20448_, new_n20447_, new_n8873_ );
or   ( new_n20449_, new_n8874_, new_n8115_ );
or   ( new_n20450_, new_n8876_, new_n8117_ );
and  ( new_n20451_, new_n20450_, new_n20449_ );
xor  ( new_n20452_, new_n20451_, new_n8257_ );
nor  ( new_n20453_, new_n20452_, new_n20448_ );
and  ( new_n20454_, new_n20452_, new_n20448_ );
or   ( new_n20455_, new_n8264_, new_n8481_ );
or   ( new_n20456_, new_n8266_, new_n8352_ );
and  ( new_n20457_, new_n20456_, new_n20455_ );
xor  ( new_n20458_, new_n20457_, new_n7725_ );
nor  ( new_n20459_, new_n20458_, new_n20454_ );
nor  ( new_n20460_, new_n20459_, new_n20453_ );
or   ( new_n20461_, new_n10059_, new_n6943_ );
or   ( new_n20462_, new_n10061_, new_n6589_ );
and  ( new_n20463_, new_n20462_, new_n20461_ );
xor  ( new_n20464_, new_n20463_, new_n9421_ );
and  ( new_n20465_, RIbb2d888_64, RIbb2c208_112 );
or   ( new_n20466_, RIbb2d888_64, new_n6425_ );
and  ( new_n20467_, new_n20466_, RIbb2d900_63 );
or   ( new_n20468_, new_n20467_, new_n20465_ );
or   ( new_n20469_, new_n10770_, new_n6219_ );
and  ( new_n20470_, new_n20469_, new_n20468_ );
nor  ( new_n20471_, new_n20470_, new_n20464_ );
and  ( new_n20472_, new_n20470_, new_n20464_ );
nor  ( new_n20473_, new_n20472_, new_n5596_ );
nor  ( new_n20474_, new_n20473_, new_n20471_ );
or   ( new_n20475_, new_n7732_, new_n9099_ );
or   ( new_n20476_, new_n7734_, new_n8995_ );
and  ( new_n20477_, new_n20476_, new_n20475_ );
xor  ( new_n20478_, new_n20477_, new_n7177_ );
or   ( new_n20479_, new_n7184_, new_n9679_ );
or   ( new_n20480_, new_n7186_, new_n9681_ );
and  ( new_n20481_, new_n20480_, new_n20479_ );
xor  ( new_n20482_, new_n20481_, new_n6638_ );
or   ( new_n20483_, new_n20482_, new_n20478_ );
and  ( new_n20484_, new_n20482_, new_n20478_ );
or   ( new_n20485_, new_n6645_, new_n10541_ );
or   ( new_n20486_, new_n6647_, new_n10220_ );
and  ( new_n20487_, new_n20486_, new_n20485_ );
xor  ( new_n20488_, new_n20487_, new_n6166_ );
or   ( new_n20489_, new_n20488_, new_n20484_ );
and  ( new_n20490_, new_n20489_, new_n20483_ );
and  ( new_n20491_, new_n20490_, new_n20474_ );
or   ( new_n20492_, new_n20491_, new_n20460_ );
or   ( new_n20493_, new_n20490_, new_n20474_ );
and  ( new_n20494_, new_n20493_, new_n20492_ );
or   ( new_n20495_, new_n20494_, new_n20444_ );
nand ( new_n20496_, new_n20494_, new_n20444_ );
xnor ( new_n20497_, new_n20389_, new_n20385_ );
xor  ( new_n20498_, new_n20497_, new_n20395_ );
xnor ( new_n20499_, new_n20373_, new_n20367_ );
xor  ( new_n20500_, new_n20499_, new_n20379_ );
nor  ( new_n20501_, new_n20500_, new_n20498_ );
and  ( new_n20502_, new_n20500_, new_n20498_ );
xor  ( new_n20503_, new_n20407_, new_n20403_ );
xor  ( new_n20504_, new_n20503_, new_n20414_ );
nor  ( new_n20505_, new_n20504_, new_n20502_ );
nor  ( new_n20506_, new_n20505_, new_n20501_ );
nand ( new_n20507_, new_n20506_, new_n20496_ );
and  ( new_n20508_, new_n20507_, new_n20495_ );
or   ( new_n20509_, new_n20508_, new_n20442_ );
nand ( new_n20510_, new_n20508_, new_n20442_ );
xor  ( new_n20511_, new_n20286_, new_n20280_ );
xor  ( new_n20512_, new_n20511_, new_n5206_ );
xor  ( new_n20513_, new_n20397_, new_n20381_ );
xor  ( new_n20514_, new_n20513_, new_n20416_ );
nor  ( new_n20515_, new_n20514_, new_n20512_ );
and  ( new_n20516_, new_n20514_, new_n20512_ );
xor  ( new_n20517_, new_n20355_, new_n20351_ );
xor  ( new_n20518_, new_n20517_, new_n20359_ );
nor  ( new_n20519_, new_n20518_, new_n20516_ );
nor  ( new_n20520_, new_n20519_, new_n20515_ );
nand ( new_n20521_, new_n20520_, new_n20510_ );
and  ( new_n20522_, new_n20521_, new_n20509_ );
nand ( new_n20523_, new_n20522_, new_n20440_ );
nor  ( new_n20524_, new_n20522_, new_n20440_ );
xor  ( new_n20525_, new_n20422_, new_n20420_ );
xor  ( new_n20526_, new_n20525_, new_n20425_ );
or   ( new_n20527_, new_n20526_, new_n20524_ );
and  ( new_n20528_, new_n20527_, new_n20523_ );
nor  ( new_n20529_, new_n20528_, new_n20435_ );
xor  ( new_n20530_, new_n20522_, new_n20440_ );
xor  ( new_n20531_, new_n20530_, new_n20526_ );
xor  ( new_n20532_, new_n20508_, new_n20442_ );
xor  ( new_n20533_, new_n20532_, new_n20520_ );
and  ( new_n20534_, new_n5915_, RIbb31578_128 );
or   ( new_n20535_, new_n20534_, new_n5597_ );
nand ( new_n20536_, new_n20534_, new_n5594_ );
and  ( new_n20537_, new_n20536_, new_n20535_ );
xnor ( new_n20538_, new_n20482_, new_n20478_ );
xor  ( new_n20539_, new_n20538_, new_n20488_ );
nor  ( new_n20540_, new_n20539_, new_n20537_ );
nand ( new_n20541_, new_n20539_, new_n20537_ );
xor  ( new_n20542_, new_n20452_, new_n20448_ );
xor  ( new_n20543_, new_n20542_, new_n20458_ );
and  ( new_n20544_, new_n20543_, new_n20541_ );
or   ( new_n20545_, new_n20544_, new_n20540_ );
xnor ( new_n20546_, new_n20500_, new_n20498_ );
xor  ( new_n20547_, new_n20546_, new_n20504_ );
nor  ( new_n20548_, new_n20547_, new_n20545_ );
nand ( new_n20549_, new_n20547_, new_n20545_ );
or   ( new_n20550_, new_n10059_, new_n7149_ );
or   ( new_n20551_, new_n10061_, new_n6943_ );
and  ( new_n20552_, new_n20551_, new_n20550_ );
xor  ( new_n20553_, new_n20552_, new_n9421_ );
and  ( new_n20554_, RIbb2d888_64, RIbb2c190_113 );
or   ( new_n20555_, RIbb2d888_64, new_n6589_ );
and  ( new_n20556_, new_n20555_, RIbb2d900_63 );
or   ( new_n20557_, new_n20556_, new_n20554_ );
or   ( new_n20558_, new_n10770_, new_n6425_ );
and  ( new_n20559_, new_n20558_, new_n20557_ );
nor  ( new_n20560_, new_n20559_, new_n20553_ );
nand ( new_n20561_, new_n20559_, new_n20553_ );
or   ( new_n20562_, new_n9422_, new_n8117_ );
or   ( new_n20563_, new_n9424_, new_n7373_ );
and  ( new_n20564_, new_n20563_, new_n20562_ );
xor  ( new_n20565_, new_n20564_, new_n8872_ );
and  ( new_n20566_, new_n20565_, new_n20561_ );
or   ( new_n20567_, new_n20566_, new_n20560_ );
or   ( new_n20568_, new_n7184_, new_n10220_ );
or   ( new_n20569_, new_n7186_, new_n9679_ );
and  ( new_n20570_, new_n20569_, new_n20568_ );
xor  ( new_n20571_, new_n20570_, new_n6638_ );
or   ( new_n20572_, new_n6645_, new_n10841_ );
or   ( new_n20573_, new_n6647_, new_n10541_ );
and  ( new_n20574_, new_n20573_, new_n20572_ );
xor  ( new_n20575_, new_n20574_, new_n6166_ );
and  ( new_n20576_, new_n20575_, new_n20571_ );
not  ( new_n20577_, new_n20576_ );
or   ( new_n20578_, new_n8874_, new_n8352_ );
or   ( new_n20579_, new_n8876_, new_n8115_ );
and  ( new_n20580_, new_n20579_, new_n20578_ );
xor  ( new_n20581_, new_n20580_, new_n8257_ );
or   ( new_n20582_, new_n8264_, new_n8995_ );
or   ( new_n20583_, new_n8266_, new_n8481_ );
and  ( new_n20584_, new_n20583_, new_n20582_ );
xor  ( new_n20585_, new_n20584_, new_n7725_ );
nor  ( new_n20586_, new_n20585_, new_n20581_ );
and  ( new_n20587_, new_n20585_, new_n20581_ );
or   ( new_n20588_, new_n7732_, new_n9681_ );
or   ( new_n20589_, new_n7734_, new_n9099_ );
and  ( new_n20590_, new_n20589_, new_n20588_ );
xor  ( new_n20591_, new_n20590_, new_n7177_ );
nor  ( new_n20592_, new_n20591_, new_n20587_ );
nor  ( new_n20593_, new_n20592_, new_n20586_ );
not  ( new_n20594_, new_n20593_ );
or   ( new_n20595_, new_n20594_, new_n20577_ );
and  ( new_n20596_, new_n20595_, new_n20567_ );
and  ( new_n20597_, new_n20594_, new_n20577_ );
or   ( new_n20598_, new_n20597_, new_n20596_ );
and  ( new_n20599_, new_n20598_, new_n20549_ );
or   ( new_n20600_, new_n20599_, new_n20548_ );
xor  ( new_n20601_, new_n20494_, new_n20444_ );
xor  ( new_n20602_, new_n20601_, new_n20506_ );
or   ( new_n20603_, new_n20602_, new_n20600_ );
and  ( new_n20604_, new_n20602_, new_n20600_ );
xor  ( new_n20605_, new_n20514_, new_n20512_ );
xor  ( new_n20606_, new_n20605_, new_n20518_ );
or   ( new_n20607_, new_n20606_, new_n20604_ );
and  ( new_n20608_, new_n20607_, new_n20603_ );
or   ( new_n20609_, new_n20608_, new_n20533_ );
nand ( new_n20610_, new_n20608_, new_n20533_ );
xor  ( new_n20611_, new_n20439_, new_n20437_ );
nand ( new_n20612_, new_n20611_, new_n20610_ );
and  ( new_n20613_, new_n20612_, new_n20609_ );
nor  ( new_n20614_, new_n20613_, new_n20531_ );
xor  ( new_n20615_, new_n20576_, new_n20567_ );
xor  ( new_n20616_, new_n20615_, new_n20593_ );
not  ( new_n20617_, new_n20616_ );
xor  ( new_n20618_, new_n20539_, new_n20537_ );
xor  ( new_n20619_, new_n20618_, new_n20543_ );
nand ( new_n20620_, new_n20619_, new_n20617_ );
xor  ( new_n20621_, new_n20470_, new_n20464_ );
xor  ( new_n20622_, new_n20621_, new_n5597_ );
xor  ( new_n20623_, new_n20559_, new_n20553_ );
xor  ( new_n20624_, new_n20623_, new_n20565_ );
xnor ( new_n20625_, new_n20585_, new_n20581_ );
xor  ( new_n20626_, new_n20625_, new_n20591_ );
or   ( new_n20627_, new_n20626_, new_n20624_ );
nand ( new_n20628_, new_n20626_, new_n20624_ );
xor  ( new_n20629_, new_n20575_, new_n20571_ );
nand ( new_n20630_, new_n20629_, new_n20628_ );
and  ( new_n20631_, new_n20630_, new_n20627_ );
or   ( new_n20632_, new_n20631_, new_n20622_ );
and  ( new_n20633_, new_n20631_, new_n20622_ );
or   ( new_n20634_, new_n10059_, new_n7373_ );
or   ( new_n20635_, new_n10061_, new_n7149_ );
and  ( new_n20636_, new_n20635_, new_n20634_ );
xor  ( new_n20637_, new_n20636_, new_n9421_ );
and  ( new_n20638_, RIbb2d888_64, RIbb2c118_114 );
or   ( new_n20639_, RIbb2d888_64, new_n6943_ );
and  ( new_n20640_, new_n20639_, RIbb2d900_63 );
or   ( new_n20641_, new_n20640_, new_n20638_ );
or   ( new_n20642_, new_n10770_, new_n6589_ );
and  ( new_n20643_, new_n20642_, new_n20641_ );
or   ( new_n20644_, new_n20643_, new_n20637_ );
and  ( new_n20645_, new_n20643_, new_n20637_ );
or   ( new_n20646_, new_n20645_, new_n6165_ );
and  ( new_n20647_, new_n20646_, new_n20644_ );
or   ( new_n20648_, new_n9422_, new_n8115_ );
or   ( new_n20649_, new_n9424_, new_n8117_ );
and  ( new_n20650_, new_n20649_, new_n20648_ );
xor  ( new_n20651_, new_n20650_, new_n8873_ );
or   ( new_n20652_, new_n8874_, new_n8481_ );
or   ( new_n20653_, new_n8876_, new_n8352_ );
and  ( new_n20654_, new_n20653_, new_n20652_ );
xor  ( new_n20655_, new_n20654_, new_n8257_ );
or   ( new_n20656_, new_n20655_, new_n20651_ );
and  ( new_n20657_, new_n20655_, new_n20651_ );
or   ( new_n20658_, new_n8264_, new_n9099_ );
or   ( new_n20659_, new_n8266_, new_n8995_ );
and  ( new_n20660_, new_n20659_, new_n20658_ );
xor  ( new_n20661_, new_n20660_, new_n7725_ );
or   ( new_n20662_, new_n20661_, new_n20657_ );
and  ( new_n20663_, new_n20662_, new_n20656_ );
and  ( new_n20664_, new_n20663_, new_n20647_ );
nor  ( new_n20665_, new_n20663_, new_n20647_ );
or   ( new_n20666_, new_n7732_, new_n9679_ );
or   ( new_n20667_, new_n7734_, new_n9681_ );
and  ( new_n20668_, new_n20667_, new_n20666_ );
xor  ( new_n20669_, new_n20668_, new_n7177_ );
or   ( new_n20670_, new_n7184_, new_n10541_ );
or   ( new_n20671_, new_n7186_, new_n10220_ );
and  ( new_n20672_, new_n20671_, new_n20670_ );
xor  ( new_n20673_, new_n20672_, new_n6638_ );
and  ( new_n20674_, new_n20673_, new_n20669_ );
nor  ( new_n20675_, new_n20673_, new_n20669_ );
and  ( new_n20676_, new_n6508_, RIbb31578_128 );
nor  ( new_n20677_, new_n20676_, new_n6166_ );
and  ( new_n20678_, new_n20676_, new_n6163_ );
nor  ( new_n20679_, new_n20678_, new_n20677_ );
nor  ( new_n20680_, new_n20679_, new_n20675_ );
nor  ( new_n20681_, new_n20680_, new_n20674_ );
nor  ( new_n20682_, new_n20681_, new_n20665_ );
nor  ( new_n20683_, new_n20682_, new_n20664_ );
or   ( new_n20684_, new_n20683_, new_n20633_ );
and  ( new_n20685_, new_n20684_, new_n20632_ );
or   ( new_n20686_, new_n20685_, new_n20620_ );
and  ( new_n20687_, new_n20685_, new_n20620_ );
xnor ( new_n20688_, new_n20490_, new_n20474_ );
xnor ( new_n20689_, new_n20688_, new_n20460_ );
not  ( new_n20690_, new_n20689_ );
or   ( new_n20691_, new_n20690_, new_n20687_ );
and  ( new_n20692_, new_n20691_, new_n20686_ );
xor  ( new_n20693_, new_n20602_, new_n20600_ );
xor  ( new_n20694_, new_n20693_, new_n20606_ );
nor  ( new_n20695_, new_n20694_, new_n20692_ );
xor  ( new_n20696_, new_n20608_, new_n20533_ );
xor  ( new_n20697_, new_n20696_, new_n20611_ );
and  ( new_n20698_, new_n20697_, new_n20695_ );
xor  ( new_n20699_, new_n20685_, new_n20620_ );
xor  ( new_n20700_, new_n20699_, new_n20690_ );
xor  ( new_n20701_, new_n20547_, new_n20545_ );
xor  ( new_n20702_, new_n20701_, new_n20598_ );
nor  ( new_n20703_, new_n20702_, new_n20700_ );
xor  ( new_n20704_, new_n20694_, new_n20692_ );
and  ( new_n20705_, new_n20704_, new_n20703_ );
xnor ( new_n20706_, new_n20702_, new_n20700_ );
xor  ( new_n20707_, new_n20643_, new_n20637_ );
xor  ( new_n20708_, new_n20707_, new_n6166_ );
xnor ( new_n20709_, new_n20655_, new_n20651_ );
xor  ( new_n20710_, new_n20709_, new_n20661_ );
nor  ( new_n20711_, new_n20710_, new_n20708_ );
xor  ( new_n20712_, new_n20626_, new_n20624_ );
xor  ( new_n20713_, new_n20712_, new_n20629_ );
or   ( new_n20714_, new_n20713_, new_n20711_ );
and  ( new_n20715_, new_n20713_, new_n20711_ );
xnor ( new_n20716_, new_n20673_, new_n20669_ );
xor  ( new_n20717_, new_n20716_, new_n20679_ );
or   ( new_n20718_, new_n10059_, new_n8117_ );
or   ( new_n20719_, new_n10061_, new_n7373_ );
and  ( new_n20720_, new_n20719_, new_n20718_ );
xor  ( new_n20721_, new_n20720_, new_n9421_ );
and  ( new_n20722_, RIbb2d888_64, RIbb2c0a0_115 );
or   ( new_n20723_, RIbb2d888_64, new_n7149_ );
and  ( new_n20724_, new_n20723_, RIbb2d900_63 );
or   ( new_n20725_, new_n20724_, new_n20722_ );
or   ( new_n20726_, new_n10770_, new_n6943_ );
and  ( new_n20727_, new_n20726_, new_n20725_ );
or   ( new_n20728_, new_n20727_, new_n20721_ );
and  ( new_n20729_, new_n20727_, new_n20721_ );
or   ( new_n20730_, new_n9422_, new_n8352_ );
or   ( new_n20731_, new_n9424_, new_n8115_ );
and  ( new_n20732_, new_n20731_, new_n20730_ );
xor  ( new_n20733_, new_n20732_, new_n8873_ );
or   ( new_n20734_, new_n20733_, new_n20729_ );
and  ( new_n20735_, new_n20734_, new_n20728_ );
nor  ( new_n20736_, new_n20735_, new_n20717_ );
and  ( new_n20737_, new_n20735_, new_n20717_ );
or   ( new_n20738_, new_n8874_, new_n8995_ );
or   ( new_n20739_, new_n8876_, new_n8481_ );
and  ( new_n20740_, new_n20739_, new_n20738_ );
xor  ( new_n20741_, new_n20740_, new_n8257_ );
or   ( new_n20742_, new_n8264_, new_n9681_ );
or   ( new_n20743_, new_n8266_, new_n9099_ );
and  ( new_n20744_, new_n20743_, new_n20742_ );
xor  ( new_n20745_, new_n20744_, new_n7725_ );
nor  ( new_n20746_, new_n20745_, new_n20741_ );
and  ( new_n20747_, new_n20745_, new_n20741_ );
or   ( new_n20748_, new_n7732_, new_n10220_ );
or   ( new_n20749_, new_n7734_, new_n9679_ );
and  ( new_n20750_, new_n20749_, new_n20748_ );
xor  ( new_n20751_, new_n20750_, new_n7177_ );
nor  ( new_n20752_, new_n20751_, new_n20747_ );
nor  ( new_n20753_, new_n20752_, new_n20746_ );
nor  ( new_n20754_, new_n20753_, new_n20737_ );
nor  ( new_n20755_, new_n20754_, new_n20736_ );
or   ( new_n20756_, new_n20755_, new_n20715_ );
and  ( new_n20757_, new_n20756_, new_n20714_ );
xnor ( new_n20758_, new_n20631_, new_n20622_ );
xor  ( new_n20759_, new_n20758_, new_n20683_ );
nand ( new_n20760_, new_n20759_, new_n20757_ );
or   ( new_n20761_, new_n20759_, new_n20757_ );
xor  ( new_n20762_, new_n20619_, new_n20617_ );
nand ( new_n20763_, new_n20762_, new_n20761_ );
and  ( new_n20764_, new_n20763_, new_n20760_ );
nor  ( new_n20765_, new_n20764_, new_n20706_ );
xor  ( new_n20766_, new_n20759_, new_n20757_ );
xor  ( new_n20767_, new_n20766_, new_n20762_ );
xnor ( new_n20768_, new_n20663_, new_n20647_ );
xor  ( new_n20769_, new_n20768_, new_n20681_ );
or   ( new_n20770_, new_n7184_, new_n10841_ );
or   ( new_n20771_, new_n7186_, new_n10541_ );
and  ( new_n20772_, new_n20771_, new_n20770_ );
xor  ( new_n20773_, new_n20772_, new_n6638_ );
or   ( new_n20774_, new_n10059_, new_n8115_ );
or   ( new_n20775_, new_n10061_, new_n8117_ );
and  ( new_n20776_, new_n20775_, new_n20774_ );
xor  ( new_n20777_, new_n20776_, new_n9421_ );
and  ( new_n20778_, RIbb2d888_64, RIbb2c028_116 );
or   ( new_n20779_, RIbb2d888_64, new_n7373_ );
and  ( new_n20780_, new_n20779_, RIbb2d900_63 );
or   ( new_n20781_, new_n20780_, new_n20778_ );
or   ( new_n20782_, new_n10770_, new_n7149_ );
and  ( new_n20783_, new_n20782_, new_n20781_ );
or   ( new_n20784_, new_n20783_, new_n20777_ );
and  ( new_n20785_, new_n20783_, new_n20777_ );
or   ( new_n20786_, new_n20785_, new_n6637_ );
and  ( new_n20787_, new_n20786_, new_n20784_ );
nor  ( new_n20788_, new_n20787_, new_n20773_ );
nand ( new_n20789_, new_n20787_, new_n20773_ );
or   ( new_n20790_, new_n9422_, new_n8481_ );
or   ( new_n20791_, new_n9424_, new_n8352_ );
and  ( new_n20792_, new_n20791_, new_n20790_ );
xor  ( new_n20793_, new_n20792_, new_n8873_ );
or   ( new_n20794_, new_n8874_, new_n9099_ );
or   ( new_n20795_, new_n8876_, new_n8995_ );
and  ( new_n20796_, new_n20795_, new_n20794_ );
xor  ( new_n20797_, new_n20796_, new_n8257_ );
nor  ( new_n20798_, new_n20797_, new_n20793_ );
nand ( new_n20799_, new_n20797_, new_n20793_ );
or   ( new_n20800_, new_n8264_, new_n9679_ );
or   ( new_n20801_, new_n8266_, new_n9681_ );
and  ( new_n20802_, new_n20801_, new_n20800_ );
xor  ( new_n20803_, new_n20802_, new_n7724_ );
and  ( new_n20804_, new_n20803_, new_n20799_ );
or   ( new_n20805_, new_n20804_, new_n20798_ );
and  ( new_n20806_, new_n20805_, new_n20789_ );
or   ( new_n20807_, new_n20806_, new_n20788_ );
xnor ( new_n20808_, new_n20735_, new_n20717_ );
xor  ( new_n20809_, new_n20808_, new_n20753_ );
nand ( new_n20810_, new_n20809_, new_n20807_ );
nor  ( new_n20811_, new_n20809_, new_n20807_ );
xor  ( new_n20812_, new_n20710_, new_n20708_ );
or   ( new_n20813_, new_n20812_, new_n20811_ );
and  ( new_n20814_, new_n20813_, new_n20810_ );
or   ( new_n20815_, new_n20814_, new_n20769_ );
nand ( new_n20816_, new_n20814_, new_n20769_ );
xor  ( new_n20817_, new_n20713_, new_n20711_ );
xnor ( new_n20818_, new_n20817_, new_n20755_ );
nand ( new_n20819_, new_n20818_, new_n20816_ );
and  ( new_n20820_, new_n20819_, new_n20815_ );
and  ( new_n20821_, new_n20820_, new_n20767_ );
xor  ( new_n20822_, new_n20727_, new_n20721_ );
xnor ( new_n20823_, new_n20822_, new_n20733_ );
xor  ( new_n20824_, new_n20787_, new_n20773_ );
xor  ( new_n20825_, new_n20824_, new_n20805_ );
or   ( new_n20826_, new_n20825_, new_n20823_ );
xnor ( new_n20827_, new_n20809_, new_n20807_ );
xor  ( new_n20828_, new_n20827_, new_n20812_ );
or   ( new_n20829_, new_n20828_, new_n20826_ );
nand ( new_n20830_, new_n20828_, new_n20826_ );
xor  ( new_n20831_, new_n20745_, new_n20741_ );
xor  ( new_n20832_, new_n20831_, new_n20751_ );
or   ( new_n20833_, new_n7732_, new_n10541_ );
or   ( new_n20834_, new_n7734_, new_n10220_ );
and  ( new_n20835_, new_n20834_, new_n20833_ );
xor  ( new_n20836_, new_n20835_, new_n7177_ );
or   ( new_n20837_, new_n8874_, new_n9681_ );
or   ( new_n20838_, new_n8876_, new_n9099_ );
and  ( new_n20839_, new_n20838_, new_n20837_ );
xor  ( new_n20840_, new_n20839_, new_n8257_ );
or   ( new_n20841_, new_n8264_, new_n10220_ );
or   ( new_n20842_, new_n8266_, new_n9679_ );
and  ( new_n20843_, new_n20842_, new_n20841_ );
xor  ( new_n20844_, new_n20843_, new_n7725_ );
or   ( new_n20845_, new_n20844_, new_n20840_ );
and  ( new_n20846_, new_n20844_, new_n20840_ );
or   ( new_n20847_, new_n7732_, new_n10841_ );
or   ( new_n20848_, new_n7734_, new_n10541_ );
and  ( new_n20849_, new_n20848_, new_n20847_ );
xor  ( new_n20850_, new_n20849_, new_n7177_ );
or   ( new_n20851_, new_n20850_, new_n20846_ );
and  ( new_n20852_, new_n20851_, new_n20845_ );
or   ( new_n20853_, new_n20852_, new_n20836_ );
and  ( new_n20854_, new_n20852_, new_n20836_ );
or   ( new_n20855_, new_n10059_, new_n8352_ );
or   ( new_n20856_, new_n10061_, new_n8115_ );
and  ( new_n20857_, new_n20856_, new_n20855_ );
xor  ( new_n20858_, new_n20857_, new_n9421_ );
and  ( new_n20859_, RIbb2d888_64, RIbb2bfb0_117 );
or   ( new_n20860_, RIbb2d888_64, new_n8117_ );
and  ( new_n20861_, new_n20860_, RIbb2d900_63 );
or   ( new_n20862_, new_n20861_, new_n20859_ );
or   ( new_n20863_, new_n10770_, new_n7373_ );
and  ( new_n20864_, new_n20863_, new_n20862_ );
nor  ( new_n20865_, new_n20864_, new_n20858_ );
and  ( new_n20866_, new_n20864_, new_n20858_ );
or   ( new_n20867_, new_n9422_, new_n8995_ );
or   ( new_n20868_, new_n9424_, new_n8481_ );
and  ( new_n20869_, new_n20868_, new_n20867_ );
xor  ( new_n20870_, new_n20869_, new_n8873_ );
nor  ( new_n20871_, new_n20870_, new_n20866_ );
nor  ( new_n20872_, new_n20871_, new_n20865_ );
or   ( new_n20873_, new_n20872_, new_n20854_ );
and  ( new_n20874_, new_n20873_, new_n20853_ );
nor  ( new_n20875_, new_n20874_, new_n20832_ );
and  ( new_n20876_, new_n20874_, new_n20832_ );
not  ( new_n20877_, new_n20876_ );
and  ( new_n20878_, new_n6908_, RIbb31578_128 );
or   ( new_n20879_, new_n20878_, new_n6638_ );
nand ( new_n20880_, new_n20878_, new_n6635_ );
and  ( new_n20881_, new_n20880_, new_n20879_ );
xor  ( new_n20882_, new_n20797_, new_n20793_ );
xor  ( new_n20883_, new_n20882_, new_n20803_ );
nor  ( new_n20884_, new_n20883_, new_n20881_ );
and  ( new_n20885_, new_n20883_, new_n20881_ );
xor  ( new_n20886_, new_n20783_, new_n20777_ );
xor  ( new_n20887_, new_n20886_, new_n6638_ );
nor  ( new_n20888_, new_n20887_, new_n20885_ );
nor  ( new_n20889_, new_n20888_, new_n20884_ );
and  ( new_n20890_, new_n20889_, new_n20877_ );
nor  ( new_n20891_, new_n20890_, new_n20875_ );
nand ( new_n20892_, new_n20891_, new_n20830_ );
and  ( new_n20893_, new_n20892_, new_n20829_ );
xor  ( new_n20894_, new_n20814_, new_n20769_ );
xor  ( new_n20895_, new_n20894_, new_n20818_ );
nor  ( new_n20896_, new_n20895_, new_n20893_ );
xor  ( new_n20897_, new_n20828_, new_n20826_ );
xor  ( new_n20898_, new_n20897_, new_n20891_ );
xnor ( new_n20899_, new_n20883_, new_n20881_ );
xor  ( new_n20900_, new_n20899_, new_n20887_ );
xor  ( new_n20901_, new_n20844_, new_n20840_ );
xor  ( new_n20902_, new_n20901_, new_n20850_ );
or   ( new_n20903_, new_n9422_, new_n9099_ );
or   ( new_n20904_, new_n9424_, new_n8995_ );
and  ( new_n20905_, new_n20904_, new_n20903_ );
xor  ( new_n20906_, new_n20905_, new_n8873_ );
or   ( new_n20907_, new_n8874_, new_n9679_ );
or   ( new_n20908_, new_n8876_, new_n9681_ );
and  ( new_n20909_, new_n20908_, new_n20907_ );
xor  ( new_n20910_, new_n20909_, new_n8257_ );
or   ( new_n20911_, new_n20910_, new_n20906_ );
and  ( new_n20912_, new_n20910_, new_n20906_ );
or   ( new_n20913_, new_n8264_, new_n10541_ );
or   ( new_n20914_, new_n8266_, new_n10220_ );
and  ( new_n20915_, new_n20914_, new_n20913_ );
xor  ( new_n20916_, new_n20915_, new_n7725_ );
or   ( new_n20917_, new_n20916_, new_n20912_ );
and  ( new_n20918_, new_n20917_, new_n20911_ );
or   ( new_n20919_, new_n20918_, new_n20902_ );
and  ( new_n20920_, new_n20918_, new_n20902_ );
or   ( new_n20921_, new_n10059_, new_n8481_ );
or   ( new_n20922_, new_n10061_, new_n8352_ );
and  ( new_n20923_, new_n20922_, new_n20921_ );
xor  ( new_n20924_, new_n20923_, new_n9421_ );
and  ( new_n20925_, RIbb2d888_64, RIbb2bf38_118 );
or   ( new_n20926_, RIbb2d888_64, new_n8115_ );
and  ( new_n20927_, new_n20926_, RIbb2d900_63 );
or   ( new_n20928_, new_n20927_, new_n20925_ );
or   ( new_n20929_, new_n10770_, new_n8117_ );
and  ( new_n20930_, new_n20929_, new_n20928_ );
nor  ( new_n20931_, new_n20930_, new_n20924_ );
and  ( new_n20932_, new_n20930_, new_n20924_ );
nor  ( new_n20933_, new_n20932_, new_n7176_ );
nor  ( new_n20934_, new_n20933_, new_n20931_ );
or   ( new_n20935_, new_n20934_, new_n20920_ );
and  ( new_n20936_, new_n20935_, new_n20919_ );
nor  ( new_n20937_, new_n20936_, new_n20900_ );
nand ( new_n20938_, new_n20936_, new_n20900_ );
xor  ( new_n20939_, new_n20852_, new_n20836_ );
xnor ( new_n20940_, new_n20939_, new_n20872_ );
and  ( new_n20941_, new_n20940_, new_n20938_ );
or   ( new_n20942_, new_n20941_, new_n20937_ );
xor  ( new_n20943_, new_n20874_, new_n20832_ );
xor  ( new_n20944_, new_n20943_, new_n20889_ );
nand ( new_n20945_, new_n20944_, new_n20942_ );
nor  ( new_n20946_, new_n20944_, new_n20942_ );
xor  ( new_n20947_, new_n20825_, new_n20823_ );
or   ( new_n20948_, new_n20947_, new_n20946_ );
and  ( new_n20949_, new_n20948_, new_n20945_ );
and  ( new_n20950_, new_n20949_, new_n20898_ );
and  ( new_n20951_, new_n7487_, RIbb31578_128 );
or   ( new_n20952_, new_n20951_, new_n7177_ );
nand ( new_n20953_, new_n20951_, new_n7174_ );
and  ( new_n20954_, new_n20953_, new_n20952_ );
xnor ( new_n20955_, new_n20910_, new_n20906_ );
xor  ( new_n20956_, new_n20955_, new_n20916_ );
or   ( new_n20957_, new_n20956_, new_n20954_ );
and  ( new_n20958_, new_n20956_, new_n20954_ );
or   ( new_n20959_, new_n10059_, new_n8995_ );
or   ( new_n20960_, new_n10061_, new_n8481_ );
and  ( new_n20961_, new_n20960_, new_n20959_ );
xor  ( new_n20962_, new_n20961_, new_n9421_ );
and  ( new_n20963_, RIbb2d888_64, RIbb2bec0_119 );
or   ( new_n20964_, RIbb2d888_64, new_n8352_ );
and  ( new_n20965_, new_n20964_, RIbb2d900_63 );
or   ( new_n20966_, new_n20965_, new_n20963_ );
or   ( new_n20967_, new_n10770_, new_n8115_ );
and  ( new_n20968_, new_n20967_, new_n20966_ );
nor  ( new_n20969_, new_n20968_, new_n20962_ );
and  ( new_n20970_, new_n20968_, new_n20962_ );
or   ( new_n20971_, new_n9422_, new_n9681_ );
or   ( new_n20972_, new_n9424_, new_n9099_ );
and  ( new_n20973_, new_n20972_, new_n20971_ );
xor  ( new_n20974_, new_n20973_, new_n8873_ );
nor  ( new_n20975_, new_n20974_, new_n20970_ );
nor  ( new_n20976_, new_n20975_, new_n20969_ );
not  ( new_n20977_, new_n20976_ );
or   ( new_n20978_, new_n20977_, new_n20958_ );
and  ( new_n20979_, new_n20978_, new_n20957_ );
xnor ( new_n20980_, new_n20864_, new_n20858_ );
xor  ( new_n20981_, new_n20980_, new_n20870_ );
nor  ( new_n20982_, new_n20981_, new_n20979_ );
and  ( new_n20983_, new_n20981_, new_n20979_ );
xor  ( new_n20984_, new_n20918_, new_n20902_ );
xnor ( new_n20985_, new_n20984_, new_n20934_ );
nor  ( new_n20986_, new_n20985_, new_n20983_ );
or   ( new_n20987_, new_n20986_, new_n20982_ );
xnor ( new_n20988_, new_n20936_, new_n20900_ );
xor  ( new_n20989_, new_n20988_, new_n20940_ );
nand ( new_n20990_, new_n20989_, new_n20987_ );
xnor ( new_n20991_, new_n20944_, new_n20942_ );
xor  ( new_n20992_, new_n20991_, new_n20947_ );
nor  ( new_n20993_, new_n20992_, new_n20990_ );
xor  ( new_n20994_, new_n20981_, new_n20979_ );
xor  ( new_n20995_, new_n20994_, new_n20985_ );
or   ( new_n20996_, new_n8264_, new_n10841_ );
or   ( new_n20997_, new_n8266_, new_n10541_ );
and  ( new_n20998_, new_n20997_, new_n20996_ );
xor  ( new_n20999_, new_n20998_, new_n7725_ );
not  ( new_n21000_, new_n20999_ );
xnor ( new_n21001_, new_n20968_, new_n20962_ );
xor  ( new_n21002_, new_n21001_, new_n20974_ );
or   ( new_n21003_, new_n21002_, new_n21000_ );
xor  ( new_n21004_, new_n20930_, new_n20924_ );
xor  ( new_n21005_, new_n21004_, new_n7177_ );
or   ( new_n21006_, new_n21005_, new_n21003_ );
and  ( new_n21007_, new_n21005_, new_n21003_ );
or   ( new_n21008_, new_n8874_, new_n10220_ );
or   ( new_n21009_, new_n8876_, new_n9679_ );
and  ( new_n21010_, new_n21009_, new_n21008_ );
xor  ( new_n21011_, new_n21010_, new_n8256_ );
or   ( new_n21012_, new_n9422_, new_n9679_ );
or   ( new_n21013_, new_n9424_, new_n9681_ );
and  ( new_n21014_, new_n21013_, new_n21012_ );
xor  ( new_n21015_, new_n21014_, new_n8873_ );
or   ( new_n21016_, new_n8874_, new_n10541_ );
or   ( new_n21017_, new_n8876_, new_n10220_ );
and  ( new_n21018_, new_n21017_, new_n21016_ );
xor  ( new_n21019_, new_n21018_, new_n8257_ );
nand ( new_n21020_, new_n21019_, new_n21015_ );
nor  ( new_n21021_, new_n21019_, new_n21015_ );
and  ( new_n21022_, new_n8040_, RIbb31578_128 );
nor  ( new_n21023_, new_n21022_, new_n7725_ );
and  ( new_n21024_, new_n21022_, new_n7722_ );
nor  ( new_n21025_, new_n21024_, new_n21023_ );
or   ( new_n21026_, new_n21025_, new_n21021_ );
and  ( new_n21027_, new_n21026_, new_n21020_ );
nor  ( new_n21028_, new_n21027_, new_n21011_ );
and  ( new_n21029_, new_n21027_, new_n21011_ );
not  ( new_n21030_, new_n21029_ );
or   ( new_n21031_, new_n10059_, new_n9099_ );
or   ( new_n21032_, new_n10061_, new_n8995_ );
and  ( new_n21033_, new_n21032_, new_n21031_ );
xor  ( new_n21034_, new_n21033_, new_n9421_ );
and  ( new_n21035_, RIbb2d888_64, RIbb2be48_120 );
or   ( new_n21036_, RIbb2d888_64, new_n8481_ );
and  ( new_n21037_, new_n21036_, RIbb2d900_63 );
or   ( new_n21038_, new_n21037_, new_n21035_ );
or   ( new_n21039_, new_n10770_, new_n8352_ );
and  ( new_n21040_, new_n21039_, new_n21038_ );
nor  ( new_n21041_, new_n21040_, new_n21034_ );
and  ( new_n21042_, new_n21040_, new_n21034_ );
nor  ( new_n21043_, new_n21042_, new_n7724_ );
nor  ( new_n21044_, new_n21043_, new_n21041_ );
and  ( new_n21045_, new_n21044_, new_n21030_ );
nor  ( new_n21046_, new_n21045_, new_n21028_ );
or   ( new_n21047_, new_n21046_, new_n21007_ );
and  ( new_n21048_, new_n21047_, new_n21006_ );
nor  ( new_n21049_, new_n21048_, new_n20995_ );
xor  ( new_n21050_, new_n20989_, new_n20987_ );
and  ( new_n21051_, new_n21050_, new_n21049_ );
xor  ( new_n21052_, new_n20956_, new_n20954_ );
xor  ( new_n21053_, new_n21052_, new_n20977_ );
xnor ( new_n21054_, new_n21005_, new_n21003_ );
xnor ( new_n21055_, new_n21054_, new_n21046_ );
nor  ( new_n21056_, new_n21055_, new_n21053_ );
xor  ( new_n21057_, new_n21048_, new_n20995_ );
and  ( new_n21058_, new_n21057_, new_n21056_ );
xnor ( new_n21059_, new_n21055_, new_n21053_ );
xor  ( new_n21060_, new_n21040_, new_n21034_ );
xor  ( new_n21061_, new_n21060_, new_n7724_ );
xnor ( new_n21062_, new_n21019_, new_n21015_ );
xor  ( new_n21063_, new_n21062_, new_n21025_ );
and  ( new_n21064_, new_n21063_, new_n21061_ );
or   ( new_n21065_, new_n21063_, new_n21061_ );
or   ( new_n21066_, new_n9422_, new_n10220_ );
or   ( new_n21067_, new_n9424_, new_n9679_ );
and  ( new_n21068_, new_n21067_, new_n21066_ );
xor  ( new_n21069_, new_n21068_, new_n8873_ );
or   ( new_n21070_, new_n10059_, new_n9681_ );
or   ( new_n21071_, new_n10061_, new_n9099_ );
and  ( new_n21072_, new_n21071_, new_n21070_ );
xor  ( new_n21073_, new_n21072_, new_n9421_ );
or   ( new_n21074_, new_n21073_, new_n21069_ );
and  ( new_n21075_, new_n21073_, new_n21069_ );
and  ( new_n21076_, RIbb2d888_64, RIbb2bdd0_121 );
not  ( new_n21077_, RIbb2d888_64 );
and  ( new_n21078_, new_n21077_, RIbb2bd58_122 );
nor  ( new_n21079_, new_n21078_, new_n10052_ );
nor  ( new_n21080_, new_n21079_, new_n21076_ );
and  ( new_n21081_, new_n10769_, RIbb2bdd0_121 );
nor  ( new_n21082_, new_n21081_, new_n21080_ );
or   ( new_n21083_, new_n21082_, new_n21075_ );
and  ( new_n21084_, new_n21083_, new_n21074_ );
and  ( new_n21085_, new_n21084_, new_n21065_ );
or   ( new_n21086_, new_n21085_, new_n21064_ );
xor  ( new_n21087_, new_n21027_, new_n21011_ );
xor  ( new_n21088_, new_n21087_, new_n21044_ );
nand ( new_n21089_, new_n21088_, new_n21086_ );
or   ( new_n21090_, new_n21088_, new_n21086_ );
xor  ( new_n21091_, new_n21002_, new_n21000_ );
nand ( new_n21092_, new_n21091_, new_n21090_ );
and  ( new_n21093_, new_n21092_, new_n21089_ );
nor  ( new_n21094_, new_n21093_, new_n21059_ );
or   ( new_n21095_, new_n9422_, new_n10541_ );
or   ( new_n21096_, new_n9424_, new_n10220_ );
and  ( new_n21097_, new_n21096_, new_n21095_ );
xor  ( new_n21098_, new_n21097_, new_n8873_ );
and  ( new_n21099_, new_n8649_, RIbb31578_128 );
or   ( new_n21100_, new_n21099_, new_n8257_ );
nand ( new_n21101_, new_n21099_, new_n8254_ );
nand ( new_n21102_, new_n21101_, new_n21100_ );
and  ( new_n21103_, new_n21102_, new_n21098_ );
or   ( new_n21104_, new_n10059_, new_n9679_ );
or   ( new_n21105_, new_n10061_, new_n9681_ );
and  ( new_n21106_, new_n21105_, new_n21104_ );
xor  ( new_n21107_, new_n21106_, new_n9421_ );
or   ( new_n21108_, new_n21107_, new_n8256_ );
and  ( new_n21109_, new_n21107_, new_n8256_ );
and  ( new_n21110_, RIbb2d888_64, RIbb2bd58_122 );
and  ( new_n21111_, new_n21077_, RIbb2bce0_123 );
nor  ( new_n21112_, new_n21111_, new_n10052_ );
nor  ( new_n21113_, new_n21112_, new_n21110_ );
and  ( new_n21114_, new_n10769_, RIbb2bd58_122 );
nor  ( new_n21115_, new_n21114_, new_n21113_ );
or   ( new_n21116_, new_n21115_, new_n21109_ );
and  ( new_n21117_, new_n21116_, new_n21108_ );
and  ( new_n21118_, new_n21117_, new_n21103_ );
or   ( new_n21119_, new_n21117_, new_n21103_ );
or   ( new_n21120_, new_n8874_, new_n10841_ );
or   ( new_n21121_, new_n8876_, new_n10541_ );
and  ( new_n21122_, new_n21121_, new_n21120_ );
xor  ( new_n21123_, new_n21122_, new_n8257_ );
and  ( new_n21124_, new_n21123_, new_n21119_ );
or   ( new_n21125_, new_n21124_, new_n21118_ );
xor  ( new_n21126_, new_n21063_, new_n21061_ );
xor  ( new_n21127_, new_n21126_, new_n21084_ );
and  ( new_n21128_, new_n21127_, new_n21125_ );
xor  ( new_n21129_, new_n21088_, new_n21086_ );
xor  ( new_n21130_, new_n21129_, new_n21091_ );
and  ( new_n21131_, new_n21130_, new_n21128_ );
xor  ( new_n21132_, new_n21117_, new_n21103_ );
xnor ( new_n21133_, new_n21132_, new_n21123_ );
xnor ( new_n21134_, new_n21073_, new_n21069_ );
xor  ( new_n21135_, new_n21134_, new_n21082_ );
nor  ( new_n21136_, new_n21135_, new_n21133_ );
xor  ( new_n21137_, new_n21127_, new_n21125_ );
and  ( new_n21138_, new_n21137_, new_n21136_ );
xnor ( new_n21139_, new_n21135_, new_n21133_ );
xnor ( new_n21140_, new_n21102_, new_n21098_ );
xor  ( new_n21141_, new_n21107_, new_n8257_ );
xor  ( new_n21142_, new_n21141_, new_n21115_ );
or   ( new_n21143_, new_n21142_, new_n21140_ );
nand ( new_n21144_, new_n21142_, new_n21140_ );
or   ( new_n21145_, new_n9422_, new_n10841_ );
or   ( new_n21146_, new_n9424_, new_n10541_ );
and  ( new_n21147_, new_n21146_, new_n21145_ );
xor  ( new_n21148_, new_n21147_, new_n8873_ );
or   ( new_n21149_, new_n10059_, new_n10220_ );
or   ( new_n21150_, new_n10061_, new_n9679_ );
and  ( new_n21151_, new_n21150_, new_n21149_ );
xor  ( new_n21152_, new_n21151_, new_n9421_ );
nor  ( new_n21153_, new_n21152_, new_n21148_ );
and  ( new_n21154_, new_n21152_, new_n21148_ );
and  ( new_n21155_, RIbb2d888_64, RIbb2bce0_123 );
and  ( new_n21156_, new_n21077_, RIbb2bc68_124 );
nor  ( new_n21157_, new_n21156_, new_n10052_ );
nor  ( new_n21158_, new_n21157_, new_n21155_ );
and  ( new_n21159_, new_n10769_, RIbb2bce0_123 );
nor  ( new_n21160_, new_n21159_, new_n21158_ );
nor  ( new_n21161_, new_n21160_, new_n21154_ );
nor  ( new_n21162_, new_n21161_, new_n21153_ );
nand ( new_n21163_, new_n21162_, new_n21144_ );
and  ( new_n21164_, new_n21163_, new_n21143_ );
nor  ( new_n21165_, new_n21164_, new_n21139_ );
or   ( new_n21166_, new_n10059_, new_n10541_ );
or   ( new_n21167_, new_n10061_, new_n10220_ );
and  ( new_n21168_, new_n21167_, new_n21166_ );
xor  ( new_n21169_, new_n21168_, new_n9421_ );
nor  ( new_n21170_, new_n21169_, new_n8872_ );
nand ( new_n21171_, new_n21169_, new_n8872_ );
or   ( new_n21172_, new_n21077_, new_n9681_ );
and  ( new_n21173_, new_n21077_, RIbb2bbf0_125 );
or   ( new_n21174_, new_n21173_, new_n10052_ );
and  ( new_n21175_, new_n21174_, new_n21172_ );
and  ( new_n21176_, new_n10769_, RIbb2bc68_124 );
or   ( new_n21177_, new_n21176_, new_n21175_ );
and  ( new_n21178_, new_n21177_, new_n21171_ );
or   ( new_n21179_, new_n21178_, new_n21170_ );
xnor ( new_n21180_, new_n21152_, new_n21148_ );
xor  ( new_n21181_, new_n21180_, new_n21160_ );
nor  ( new_n21182_, new_n21181_, new_n21179_ );
xor  ( new_n21183_, new_n21142_, new_n21140_ );
xor  ( new_n21184_, new_n21183_, new_n21162_ );
and  ( new_n21185_, new_n21184_, new_n21182_ );
and  ( new_n21186_, new_n9185_, RIbb31578_128 );
or   ( new_n21187_, new_n21186_, new_n8873_ );
nand ( new_n21188_, new_n21186_, new_n8870_ );
and  ( new_n21189_, new_n21188_, new_n21187_ );
xor  ( new_n21190_, new_n21169_, new_n8872_ );
xor  ( new_n21191_, new_n21190_, new_n21177_ );
nor  ( new_n21192_, new_n21191_, new_n21189_ );
xor  ( new_n21193_, new_n21181_, new_n21179_ );
and  ( new_n21194_, new_n21193_, new_n21192_ );
or   ( new_n21195_, new_n10059_, new_n10841_ );
or   ( new_n21196_, new_n10061_, new_n10541_ );
and  ( new_n21197_, new_n21196_, new_n21195_ );
xor  ( new_n21198_, new_n21197_, new_n9421_ );
and  ( new_n21199_, RIbb2d888_64, RIbb2bbf0_125 );
or   ( new_n21200_, RIbb2d888_64, new_n10220_ );
and  ( new_n21201_, new_n21200_, RIbb2d900_63 );
or   ( new_n21202_, new_n21201_, new_n21199_ );
or   ( new_n21203_, new_n10770_, new_n9679_ );
and  ( new_n21204_, new_n21203_, new_n21202_ );
and  ( new_n21205_, new_n21204_, new_n21198_ );
xor  ( new_n21206_, new_n21191_, new_n21189_ );
and  ( new_n21207_, new_n21206_, new_n21205_ );
and  ( new_n21208_, RIbb2d888_64, RIbb2bb78_126 );
or   ( new_n21209_, RIbb2d888_64, new_n10541_ );
and  ( new_n21210_, new_n21209_, RIbb2d900_63 );
or   ( new_n21211_, new_n21210_, new_n21208_ );
or   ( new_n21212_, new_n10770_, new_n10220_ );
and  ( new_n21213_, new_n21212_, new_n21211_ );
and  ( new_n21214_, new_n21213_, new_n9420_ );
xor  ( new_n21215_, new_n21204_, new_n21198_ );
and  ( new_n21216_, new_n21215_, new_n21214_ );
xor  ( new_n21217_, new_n21213_, new_n9421_ );
and  ( new_n21218_, new_n9738_, RIbb31578_128 );
or   ( new_n21219_, new_n21218_, new_n9421_ );
nand ( new_n21220_, new_n21218_, new_n9418_ );
and  ( new_n21221_, new_n21220_, new_n21219_ );
nor  ( new_n21222_, new_n21221_, new_n21217_ );
and  ( new_n21223_, RIbb31578_128, RIbb2d888_64 );
nor  ( new_n21224_, new_n21223_, new_n10052_ );
and  ( new_n21225_, RIbb2d888_64, RIbb31500_127 );
or   ( new_n21226_, new_n10841_, RIbb2d888_64 );
and  ( new_n21227_, new_n21226_, RIbb2d900_63 );
or   ( new_n21228_, new_n21227_, new_n21225_ );
or   ( new_n21229_, new_n10770_, new_n10541_ );
and  ( new_n21230_, new_n21229_, new_n21228_ );
and  ( new_n21231_, new_n21230_, new_n21224_ );
xor  ( new_n21232_, new_n21221_, new_n21217_ );
and  ( new_n21233_, new_n21232_, new_n21231_ );
nor  ( new_n21234_, new_n21233_, new_n21222_ );
not  ( new_n21235_, new_n21234_ );
xor  ( new_n21236_, new_n21215_, new_n21214_ );
and  ( new_n21237_, new_n21236_, new_n21235_ );
nor  ( new_n21238_, new_n21237_, new_n21216_ );
not  ( new_n21239_, new_n21238_ );
xor  ( new_n21240_, new_n21206_, new_n21205_ );
and  ( new_n21241_, new_n21240_, new_n21239_ );
nor  ( new_n21242_, new_n21241_, new_n21207_ );
not  ( new_n21243_, new_n21242_ );
xor  ( new_n21244_, new_n21193_, new_n21192_ );
and  ( new_n21245_, new_n21244_, new_n21243_ );
nor  ( new_n21246_, new_n21245_, new_n21194_ );
not  ( new_n21247_, new_n21246_ );
xor  ( new_n21248_, new_n21184_, new_n21182_ );
and  ( new_n21249_, new_n21248_, new_n21247_ );
nor  ( new_n21250_, new_n21249_, new_n21185_ );
not  ( new_n21251_, new_n21250_ );
xor  ( new_n21252_, new_n21164_, new_n21139_ );
and  ( new_n21253_, new_n21252_, new_n21251_ );
nor  ( new_n21254_, new_n21253_, new_n21165_ );
not  ( new_n21255_, new_n21254_ );
xor  ( new_n21256_, new_n21137_, new_n21136_ );
and  ( new_n21257_, new_n21256_, new_n21255_ );
nor  ( new_n21258_, new_n21257_, new_n21138_ );
not  ( new_n21259_, new_n21258_ );
xor  ( new_n21260_, new_n21130_, new_n21128_ );
and  ( new_n21261_, new_n21260_, new_n21259_ );
or   ( new_n21262_, new_n21261_, new_n21131_ );
xor  ( new_n21263_, new_n21093_, new_n21059_ );
and  ( new_n21264_, new_n21263_, new_n21262_ );
or   ( new_n21265_, new_n21264_, new_n21094_ );
xor  ( new_n21266_, new_n21057_, new_n21056_ );
and  ( new_n21267_, new_n21266_, new_n21265_ );
or   ( new_n21268_, new_n21267_, new_n21058_ );
xor  ( new_n21269_, new_n21050_, new_n21049_ );
and  ( new_n21270_, new_n21269_, new_n21268_ );
or   ( new_n21271_, new_n21270_, new_n21051_ );
xor  ( new_n21272_, new_n20992_, new_n20990_ );
and  ( new_n21273_, new_n21272_, new_n21271_ );
or   ( new_n21274_, new_n21273_, new_n20993_ );
xor  ( new_n21275_, new_n20949_, new_n20898_ );
and  ( new_n21276_, new_n21275_, new_n21274_ );
or   ( new_n21277_, new_n21276_, new_n20950_ );
xor  ( new_n21278_, new_n20895_, new_n20893_ );
and  ( new_n21279_, new_n21278_, new_n21277_ );
or   ( new_n21280_, new_n21279_, new_n20896_ );
xor  ( new_n21281_, new_n20820_, new_n20767_ );
and  ( new_n21282_, new_n21281_, new_n21280_ );
or   ( new_n21283_, new_n21282_, new_n20821_ );
xor  ( new_n21284_, new_n20764_, new_n20706_ );
and  ( new_n21285_, new_n21284_, new_n21283_ );
or   ( new_n21286_, new_n21285_, new_n20765_ );
xor  ( new_n21287_, new_n20704_, new_n20703_ );
and  ( new_n21288_, new_n21287_, new_n21286_ );
or   ( new_n21289_, new_n21288_, new_n20705_ );
xor  ( new_n21290_, new_n20697_, new_n20695_ );
and  ( new_n21291_, new_n21290_, new_n21289_ );
or   ( new_n21292_, new_n21291_, new_n20698_ );
xor  ( new_n21293_, new_n20613_, new_n20531_ );
and  ( new_n21294_, new_n21293_, new_n21292_ );
or   ( new_n21295_, new_n21294_, new_n20614_ );
xor  ( new_n21296_, new_n20528_, new_n20435_ );
and  ( new_n21297_, new_n21296_, new_n21295_ );
or   ( new_n21298_, new_n21297_, new_n20529_ );
xor  ( new_n21299_, new_n20432_, new_n20343_ );
and  ( new_n21300_, new_n21299_, new_n21298_ );
or   ( new_n21301_, new_n21300_, new_n20433_ );
xor  ( new_n21302_, new_n20340_, new_n20250_ );
and  ( new_n21303_, new_n21302_, new_n21301_ );
or   ( new_n21304_, new_n21303_, new_n20341_ );
xor  ( new_n21305_, new_n20247_, new_n20245_ );
and  ( new_n21306_, new_n21305_, new_n21304_ );
or   ( new_n21307_, new_n21306_, new_n20248_ );
xor  ( new_n21308_, new_n20157_, new_n20040_ );
and  ( new_n21309_, new_n21308_, new_n21307_ );
or   ( new_n21310_, new_n21309_, new_n20158_ );
xor  ( new_n21311_, new_n20037_, new_n19940_ );
and  ( new_n21312_, new_n21311_, new_n21310_ );
or   ( new_n21313_, new_n21312_, new_n20038_ );
xor  ( new_n21314_, new_n19938_, new_n19937_ );
and  ( new_n21315_, new_n21314_, new_n21313_ );
or   ( new_n21316_, new_n21315_, new_n19939_ );
xor  ( new_n21317_, new_n19931_, new_n19929_ );
and  ( new_n21318_, new_n21317_, new_n21316_ );
or   ( new_n21319_, new_n21318_, new_n19932_ );
xor  ( new_n21320_, new_n19814_, new_n19691_ );
and  ( new_n21321_, new_n21320_, new_n21319_ );
or   ( new_n21322_, new_n21321_, new_n19815_ );
xor  ( new_n21323_, new_n19688_, new_n19546_ );
and  ( new_n21324_, new_n21323_, new_n21322_ );
nor  ( new_n21325_, new_n21324_, new_n19689_ );
not  ( new_n21326_, new_n21325_ );
xor  ( new_n21327_, new_n19543_, new_n19421_ );
and  ( new_n21328_, new_n21327_, new_n21326_ );
or   ( new_n21329_, new_n21328_, new_n19544_ );
xor  ( new_n21330_, new_n19418_, new_n19274_ );
and  ( new_n21331_, new_n21330_, new_n21329_ );
or   ( new_n21332_, new_n21331_, new_n19419_ );
xor  ( new_n21333_, new_n19271_, new_n19145_ );
and  ( new_n21334_, new_n21333_, new_n21332_ );
or   ( new_n21335_, new_n21334_, new_n19272_ );
xor  ( new_n21336_, new_n19142_, new_n19005_ );
and  ( new_n21337_, new_n21336_, new_n21335_ );
or   ( new_n21338_, new_n21337_, new_n19143_ );
xor  ( new_n21339_, new_n19002_, new_n19000_ );
and  ( new_n21340_, new_n21339_, new_n21338_ );
or   ( new_n21341_, new_n21340_, new_n19003_ );
xor  ( new_n21342_, new_n18833_, new_n18682_ );
and  ( new_n21343_, new_n21342_, new_n21341_ );
or   ( new_n21344_, new_n21343_, new_n18834_ );
xor  ( new_n21345_, new_n18679_, new_n18538_ );
and  ( new_n21346_, new_n21345_, new_n21344_ );
or   ( new_n21347_, new_n21346_, new_n18680_ );
xor  ( new_n21348_, new_n18535_, new_n18359_ );
and  ( new_n21349_, new_n21348_, new_n21347_ );
or   ( new_n21350_, new_n21349_, new_n18536_ );
xor  ( new_n21351_, new_n18357_, new_n18356_ );
and  ( new_n21352_, new_n21351_, new_n21350_ );
or   ( new_n21353_, new_n21352_, new_n18358_ );
xor  ( new_n21354_, new_n18350_, new_n18349_ );
and  ( new_n21355_, new_n21354_, new_n21353_ );
or   ( new_n21356_, new_n21355_, new_n18351_ );
xor  ( new_n21357_, new_n18169_, new_n18167_ );
and  ( new_n21358_, new_n21357_, new_n21356_ );
or   ( new_n21359_, new_n21358_, new_n18170_ );
xor  ( new_n21360_, new_n17991_, new_n17799_ );
and  ( new_n21361_, new_n21360_, new_n21359_ );
or   ( new_n21362_, new_n21361_, new_n17992_ );
xor  ( new_n21363_, new_n17797_, new_n17795_ );
and  ( new_n21364_, new_n21363_, new_n21362_ );
or   ( new_n21365_, new_n21364_, new_n17798_ );
xor  ( new_n21366_, new_n17601_, new_n17414_ );
and  ( new_n21367_, new_n21366_, new_n21365_ );
or   ( new_n21368_, new_n21367_, new_n17602_ );
xor  ( new_n21369_, new_n17411_, new_n17199_ );
and  ( new_n21370_, new_n21369_, new_n21368_ );
or   ( new_n21371_, new_n21370_, new_n17412_ );
xor  ( new_n21372_, new_n17196_, new_n16997_ );
and  ( new_n21373_, new_n21372_, new_n21371_ );
or   ( new_n21374_, new_n21373_, new_n17197_ );
xor  ( new_n21375_, new_n16994_, new_n16798_ );
and  ( new_n21376_, new_n21375_, new_n21374_ );
or   ( new_n21377_, new_n21376_, new_n16995_ );
xor  ( new_n21378_, new_n16795_, new_n16584_ );
and  ( new_n21379_, new_n21378_, new_n21377_ );
or   ( new_n21380_, new_n21379_, new_n16796_ );
xor  ( new_n21381_, new_n16581_, new_n16368_ );
and  ( new_n21382_, new_n21381_, new_n21380_ );
or   ( new_n21383_, new_n21382_, new_n16582_ );
xor  ( new_n21384_, new_n16365_, new_n16363_ );
and  ( new_n21385_, new_n21384_, new_n21383_ );
or   ( new_n21386_, new_n21385_, new_n16366_ );
xor  ( new_n21387_, new_n16131_, new_n15895_ );
and  ( new_n21388_, new_n21387_, new_n21386_ );
or   ( new_n21389_, new_n21388_, new_n16132_ );
xor  ( new_n21390_, new_n15892_, new_n15669_ );
and  ( new_n21391_, new_n21390_, new_n21389_ );
or   ( new_n21392_, new_n21391_, new_n15893_ );
xor  ( new_n21393_, new_n15666_, new_n15442_ );
and  ( new_n21394_, new_n21393_, new_n21392_ );
or   ( new_n21395_, new_n21394_, new_n15667_ );
xor  ( new_n21396_, new_n15439_, new_n15188_ );
and  ( new_n21397_, new_n21396_, new_n21395_ );
or   ( new_n21398_, new_n21397_, new_n15440_ );
xor  ( new_n21399_, new_n15185_, new_n14954_ );
and  ( new_n21400_, new_n21399_, new_n21398_ );
or   ( new_n21401_, new_n21400_, new_n15186_ );
xor  ( new_n21402_, new_n14951_, new_n14704_ );
and  ( new_n21403_, new_n21402_, new_n21401_ );
or   ( new_n21404_, new_n21403_, new_n14952_ );
xor  ( new_n21405_, new_n14702_, new_n14701_ );
and  ( new_n21406_, new_n21405_, new_n21404_ );
or   ( new_n21407_, new_n21406_, new_n14703_ );
xor  ( new_n21408_, new_n14695_, new_n14694_ );
and  ( new_n21409_, new_n21408_, new_n21407_ );
or   ( new_n21410_, new_n21409_, new_n14696_ );
xor  ( new_n21411_, new_n14426_, new_n14425_ );
and  ( new_n21412_, new_n21411_, new_n21410_ );
or   ( new_n21413_, new_n21412_, new_n14427_ );
xor  ( new_n21414_, new_n14158_, new_n14156_ );
and  ( new_n21415_, new_n21414_, new_n21413_ );
or   ( new_n21416_, new_n21415_, new_n14159_ );
xor  ( new_n21417_, new_n13887_, new_n13607_ );
and  ( new_n21418_, new_n21417_, new_n21416_ );
nor  ( new_n21419_, new_n21418_, new_n13888_ );
not  ( new_n21420_, new_n21419_ );
xor  ( new_n21421_, new_n13605_, new_n13604_ );
and  ( new_n21422_, new_n21421_, new_n21420_ );
or   ( new_n21423_, new_n21422_, new_n13606_ );
xor  ( new_n21424_, new_n13327_, new_n13325_ );
and  ( new_n21425_, new_n21424_, new_n21423_ );
or   ( new_n21426_, new_n21425_, new_n13328_ );
xor  ( new_n21427_, new_n13053_, new_n12748_ );
and  ( new_n21428_, new_n21427_, new_n21426_ );
or   ( new_n21429_, new_n21428_, new_n13054_ );
xor  ( new_n21430_, new_n12746_, new_n12744_ );
and  ( new_n21431_, new_n21430_, new_n21429_ );
or   ( new_n21432_, new_n21431_, new_n12747_ );
xor  ( new_n21433_, new_n12463_, new_n12177_ );
and  ( new_n21434_, new_n21433_, new_n21432_ );
or   ( new_n21435_, new_n21434_, new_n12464_ );
xor  ( new_n21436_, new_n12174_, new_n11858_ );
and  ( new_n21437_, new_n21436_, new_n21435_ );
nor  ( new_n21438_, new_n21437_, new_n12175_ );
not  ( new_n21439_, new_n21438_ );
xor  ( new_n21440_, new_n11855_, new_n11553_ );
and  ( new_n21441_, new_n21440_, new_n21439_ );
or   ( new_n21442_, new_n21441_, new_n11856_ );
xor  ( new_n21443_, new_n11550_, new_n11233_ );
and  ( new_n21444_, new_n21443_, new_n21442_ );
nor  ( new_n21445_, new_n21444_, new_n11551_ );
not  ( new_n21446_, new_n21445_ );
xor  ( new_n21447_, new_n11230_, new_n10910_ );
and  ( new_n21448_, new_n21447_, new_n21446_ );
or   ( new_n21449_, new_n21448_, new_n11231_ );
xor  ( new_n21450_, new_n10907_, new_n10595_ );
and  ( new_n21451_, new_n21450_, new_n21449_ );
or   ( new_n21452_, new_n21451_, new_n10908_ );
xor  ( new_n21453_, new_n10592_, new_n10285_ );
and  ( new_n21454_, new_n21453_, new_n21452_ );
or   ( new_n21455_, new_n21454_, new_n10593_ );
xor  ( new_n21456_, new_n10283_, new_n10281_ );
and  ( new_n21457_, new_n21456_, new_n21455_ );
or   ( new_n21458_, new_n21457_, new_n10284_ );
xor  ( new_n21459_, new_n9963_, new_n9648_ );
and  ( new_n21460_, new_n21459_, new_n21458_ );
or   ( new_n21461_, new_n21460_, new_n9964_ );
xor  ( new_n21462_, new_n9646_, new_n9645_ );
and  ( new_n21463_, new_n21462_, new_n21461_ );
nor  ( new_n21464_, new_n21463_, new_n9647_ );
not  ( new_n21465_, new_n21464_ );
xor  ( new_n21466_, new_n9334_, new_n9332_ );
and  ( new_n21467_, new_n21466_, new_n21465_ );
nor  ( new_n21468_, new_n21467_, new_n9335_ );
not  ( new_n21469_, new_n21468_ );
xor  ( new_n21470_, new_n9042_, new_n8740_ );
and  ( new_n21471_, new_n21470_, new_n21469_ );
nor  ( new_n21472_, new_n21471_, new_n9043_ );
not  ( new_n21473_, new_n21472_ );
xor  ( new_n21474_, new_n8738_, new_n8737_ );
and  ( new_n21475_, new_n21474_, new_n21473_ );
or   ( new_n21476_, new_n21475_, new_n8739_ );
xor  ( new_n21477_, new_n8449_, new_n8448_ );
and  ( new_n21478_, new_n21477_, new_n21476_ );
or   ( new_n21479_, new_n21478_, new_n8450_ );
xor  ( new_n21480_, new_n8164_, new_n8163_ );
and  ( new_n21481_, new_n21480_, new_n21479_ );
or   ( new_n21482_, new_n21481_, new_n8165_ );
xor  ( new_n21483_, new_n7872_, new_n7871_ );
and  ( new_n21484_, new_n21483_, new_n21482_ );
or   ( new_n21485_, new_n21484_, new_n7873_ );
xor  ( new_n21486_, new_n7606_, new_n7605_ );
and  ( new_n21487_, new_n21486_, new_n21485_ );
nor  ( new_n21488_, new_n21487_, new_n7607_ );
not  ( new_n21489_, new_n21488_ );
xor  ( new_n21490_, new_n7341_, new_n7340_ );
and  ( new_n21491_, new_n21490_, new_n21489_ );
or   ( new_n21492_, new_n21491_, new_n7342_ );
xor  ( new_n21493_, new_n7079_, new_n7078_ );
and  ( new_n21494_, new_n21493_, new_n21492_ );
or   ( new_n21495_, new_n21494_, new_n7080_ );
xor  ( new_n21496_, new_n6815_, new_n6814_ );
and  ( new_n21497_, new_n21496_, new_n21495_ );
nor  ( new_n21498_, new_n21497_, new_n6816_ );
not  ( new_n21499_, new_n21498_ );
xor  ( new_n21500_, new_n6553_, new_n6552_ );
and  ( new_n21501_, new_n21500_, new_n21499_ );
or   ( new_n21502_, new_n21501_, new_n6554_ );
xor  ( new_n21503_, new_n6297_, new_n6296_ );
and  ( new_n21504_, new_n21503_, new_n21502_ );
or   ( new_n21505_, new_n21504_, new_n6298_ );
xor  ( new_n21506_, new_n6039_, new_n6038_ );
and  ( new_n21507_, new_n21506_, new_n21505_ );
or   ( new_n21508_, new_n21507_, new_n6040_ );
xor  ( new_n21509_, new_n5788_, new_n5787_ );
and  ( new_n21510_, new_n21509_, new_n21508_ );
nor  ( new_n21511_, new_n21510_, new_n5789_ );
not  ( new_n21512_, new_n21511_ );
xor  ( new_n21513_, new_n5538_, new_n5537_ );
and  ( new_n21514_, new_n21513_, new_n21512_ );
or   ( new_n21515_, new_n21514_, new_n5539_ );
xor  ( new_n21516_, new_n5308_, new_n5306_ );
and  ( new_n21517_, new_n21516_, new_n21515_ );
nor  ( new_n21518_, new_n21517_, new_n5309_ );
not  ( new_n21519_, new_n21518_ );
xor  ( new_n21520_, new_n5063_, new_n4636_ );
and  ( new_n21521_, new_n21520_, new_n21519_ );
nor  ( new_n21522_, new_n21521_, new_n5064_ );
not  ( new_n21523_, new_n21522_ );
xor  ( new_n21524_, new_n4633_, new_n4431_ );
and  ( new_n21525_, new_n21524_, new_n21523_ );
or   ( new_n21526_, new_n21525_, new_n4634_ );
xor  ( new_n21527_, new_n4428_, new_n4218_ );
and  ( new_n21528_, new_n21527_, new_n21526_ );
nor  ( new_n21529_, new_n21528_, new_n4429_ );
not  ( new_n21530_, new_n21529_ );
xor  ( new_n21531_, new_n4216_, new_n4215_ );
and  ( new_n21532_, new_n21531_, new_n21530_ );
nor  ( new_n21533_, new_n21532_, new_n4217_ );
not  ( new_n21534_, new_n21533_ );
xor  ( new_n21535_, new_n4007_, new_n4006_ );
and  ( new_n21536_, new_n21535_, new_n21534_ );
or   ( new_n21537_, new_n21536_, new_n4008_ );
xor  ( new_n21538_, new_n3805_, new_n3804_ );
and  ( new_n21539_, new_n21538_, new_n21537_ );
nor  ( new_n21540_, new_n21539_, new_n3806_ );
not  ( new_n21541_, new_n21540_ );
xor  ( new_n21542_, new_n3609_, new_n3608_ );
and  ( new_n21543_, new_n21542_, new_n21541_ );
or   ( new_n21544_, new_n21543_, new_n3610_ );
xor  ( new_n21545_, new_n3429_, new_n3428_ );
and  ( new_n21546_, new_n21545_, new_n21544_ );
or   ( new_n21547_, new_n21546_, new_n3430_ );
xor  ( new_n21548_, new_n3249_, new_n3248_ );
and  ( new_n21549_, new_n21548_, new_n21547_ );
nor  ( new_n21550_, new_n21549_, new_n3250_ );
not  ( new_n21551_, new_n21550_ );
xor  ( new_n21552_, new_n3077_, new_n3076_ );
and  ( new_n21553_, new_n21552_, new_n21551_ );
nor  ( new_n21554_, new_n21553_, new_n3078_ );
not  ( new_n21555_, new_n21554_ );
xor  ( new_n21556_, new_n2904_, new_n2903_ );
and  ( new_n21557_, new_n21556_, new_n21555_ );
or   ( new_n21558_, new_n21557_, new_n2905_ );
xor  ( new_n21559_, new_n2732_, new_n2731_ );
and  ( new_n21560_, new_n21559_, new_n21558_ );
nor  ( new_n21561_, new_n21560_, new_n2733_ );
not  ( new_n21562_, new_n21561_ );
xor  ( new_n21563_, new_n2565_, new_n2564_ );
and  ( new_n21564_, new_n21563_, new_n21562_ );
nor  ( new_n21565_, new_n21564_, new_n2566_ );
not  ( new_n21566_, new_n21565_ );
xor  ( new_n21567_, new_n2399_, new_n2397_ );
and  ( new_n21568_, new_n21567_, new_n21566_ );
nor  ( new_n21569_, new_n21568_, new_n2400_ );
not  ( new_n21570_, new_n21569_ );
xor  ( new_n21571_, new_n2228_, new_n1951_ );
and  ( new_n21572_, new_n21571_, new_n21570_ );
nor  ( new_n21573_, new_n21572_, new_n2229_ );
not  ( new_n21574_, new_n21573_ );
xor  ( new_n21575_, new_n1948_, new_n1813_ );
and  ( new_n21576_, new_n21575_, new_n21574_ );
nor  ( new_n21577_, new_n21576_, new_n1949_ );
not  ( new_n21578_, new_n21577_ );
xor  ( new_n21579_, new_n1811_, new_n1810_ );
and  ( new_n21580_, new_n21579_, new_n21578_ );
nor  ( new_n21581_, new_n21580_, new_n1812_ );
not  ( new_n21582_, new_n21581_ );
xor  ( new_n21583_, new_n1677_, new_n1676_ );
and  ( new_n21584_, new_n21583_, new_n21582_ );
nor  ( new_n21585_, new_n21584_, new_n1678_ );
not  ( new_n21586_, new_n21585_ );
xor  ( new_n21587_, new_n1557_, new_n1556_ );
and  ( new_n21588_, new_n21587_, new_n21586_ );
or   ( new_n21589_, new_n21588_, new_n1558_ );
xor  ( new_n21590_, new_n1432_, new_n1431_ );
and  ( new_n21591_, new_n21590_, new_n21589_ );
nor  ( new_n21592_, new_n21591_, new_n1433_ );
not  ( new_n21593_, new_n21592_ );
xor  ( new_n21594_, new_n1314_, new_n1313_ );
and  ( new_n21595_, new_n21594_, new_n21593_ );
or   ( new_n21596_, new_n21595_, new_n1315_ );
xor  ( new_n21597_, new_n1201_, new_n1200_ );
and  ( new_n21598_, new_n21597_, new_n21596_ );
nor  ( new_n21599_, new_n21598_, new_n1202_ );
not  ( new_n21600_, new_n21599_ );
xor  ( new_n21601_, new_n1087_, new_n1085_ );
and  ( new_n21602_, new_n21601_, new_n21600_ );
nor  ( new_n21603_, new_n21602_, new_n1088_ );
not  ( new_n21604_, new_n21603_ );
xor  ( new_n21605_, new_n976_, new_n798_ );
and  ( new_n21606_, new_n21605_, new_n21604_ );
or   ( new_n21607_, new_n21606_, new_n977_ );
xor  ( new_n21608_, new_n796_, new_n795_ );
and  ( new_n21609_, new_n21608_, new_n21607_ );
or   ( new_n21610_, new_n21609_, new_n797_ );
xor  ( new_n21611_, new_n716_, new_n715_ );
and  ( new_n21612_, new_n21611_, new_n21610_ );
nor  ( new_n21613_, new_n21612_, new_n717_ );
not  ( new_n21614_, new_n21613_ );
xor  ( new_n21615_, new_n637_, new_n578_ );
and  ( new_n21616_, new_n21615_, new_n21614_ );
nor  ( new_n21617_, new_n21616_, new_n638_ );
or   ( new_n21618_, new_n268_, new_n294_ );
or   ( new_n21619_, new_n271_, new_n301_ );
and  ( new_n21620_, new_n21619_, new_n21618_ );
and  ( new_n21621_, RIbb2f610_1, RIbb2d450_73 );
xor  ( new_n21622_, new_n21621_, new_n21620_ );
nor  ( new_n21623_, RIbb2f2c8_8, new_n309_ );
nor  ( new_n21624_, new_n332_, new_n21623_ );
and  ( new_n21625_, new_n332_, new_n311_ );
nor  ( new_n21626_, new_n21625_, new_n21624_ );
xor  ( new_n21627_, new_n21626_, new_n21622_ );
xnor ( new_n21628_, new_n21627_, new_n21617_ );
nand ( new_n21629_, new_n606_, new_n593_ );
or   ( new_n21630_, new_n616_, new_n611_ );
and  ( new_n21631_, new_n616_, new_n611_ );
or   ( new_n21632_, new_n628_, new_n21631_ );
and  ( new_n21633_, new_n21632_, new_n21630_ );
xor  ( new_n21634_, new_n21633_, new_n21629_ );
xor  ( new_n21635_, new_n292_, new_n263_ );
xor  ( new_n21636_, new_n21635_, new_n21634_ );
or   ( new_n21637_, new_n636_, new_n582_ );
and  ( new_n21638_, new_n298_, RIbb2d5b8_70 );
and  ( new_n21639_, new_n295_, RIbb2d630_69 );
or   ( new_n21640_, new_n21639_, new_n21638_ );
not  ( new_n21641_, new_n622_ );
not  ( new_n21642_, new_n626_ );
and  ( new_n21643_, new_n21642_, new_n21641_ );
or   ( new_n21644_, new_n21642_, new_n21641_ );
and  ( new_n21645_, new_n21644_, new_n618_ );
or   ( new_n21646_, new_n21645_, new_n21643_ );
or   ( new_n21647_, new_n604_, new_n601_ );
and  ( new_n21648_, new_n604_, new_n601_ );
or   ( new_n21649_, new_n21648_, new_n597_ );
and  ( new_n21650_, new_n21649_, new_n21647_ );
xor  ( new_n21651_, new_n21650_, new_n21646_ );
xor  ( new_n21652_, new_n21651_, new_n21640_ );
xor  ( new_n21653_, new_n21652_, new_n21637_ );
xor  ( new_n21654_, new_n21653_, new_n21636_ );
and  ( new_n21655_, new_n630_, new_n607_ );
nor  ( new_n21656_, new_n630_, new_n607_ );
nor  ( new_n21657_, new_n635_, new_n21656_ );
or   ( new_n21658_, new_n21657_, new_n21655_ );
nand ( new_n21659_, new_n591_, new_n587_ );
or   ( new_n21660_, new_n283_, new_n313_ );
or   ( new_n21661_, new_n286_, new_n319_ );
and  ( new_n21662_, new_n21661_, new_n21660_ );
or   ( new_n21663_, new_n317_, new_n333_ );
or   ( new_n21664_, new_n320_, new_n339_ );
and  ( new_n21665_, new_n21664_, new_n21663_ );
xor  ( new_n21666_, new_n21665_, new_n278_ );
xor  ( new_n21667_, new_n21666_, new_n21662_ );
xor  ( new_n21668_, new_n21667_, new_n21659_ );
xor  ( new_n21669_, new_n21668_, new_n21658_ );
xor  ( new_n21670_, new_n21669_, new_n21654_ );
xor  ( new_n21671_, new_n21670_, new_n21628_ );
not  ( new_n21672_, RIbb31848_134 );
or   ( new_n21673_, new_n283_, new_n21672_ );
not  ( new_n21674_, RIbb317d0_133 );
or   ( new_n21675_, new_n286_, new_n21674_ );
and  ( new_n21676_, new_n21675_, new_n21673_ );
xor  ( new_n21677_, new_n21676_, new_n278_ );
not  ( new_n21678_, RIbb31938_136 );
or   ( new_n21679_, new_n299_, new_n21678_ );
not  ( new_n21680_, RIbb318c0_135 );
or   ( new_n21681_, new_n302_, new_n21680_ );
and  ( new_n21682_, new_n21681_, new_n21679_ );
xor  ( new_n21683_, new_n21682_, new_n293_ );
nor  ( new_n21684_, new_n21683_, new_n21677_ );
not  ( new_n21685_, RIbb31a28_138 );
or   ( new_n21686_, new_n268_, new_n21685_ );
not  ( new_n21687_, RIbb319b0_137 );
or   ( new_n21688_, new_n271_, new_n21687_ );
and  ( new_n21689_, new_n21688_, new_n21686_ );
xor  ( new_n21690_, new_n21689_, new_n263_ );
and  ( new_n21691_, new_n21683_, new_n21677_ );
nor  ( new_n21692_, new_n21691_, new_n21690_ );
nor  ( new_n21693_, new_n21692_, new_n21684_ );
not  ( new_n21694_, RIbb31668_130 );
or   ( new_n21695_, new_n337_, new_n21694_ );
not  ( new_n21696_, RIbb315f0_129 );
or   ( new_n21697_, new_n340_, new_n21696_ );
and  ( new_n21698_, new_n21697_, new_n21695_ );
xor  ( new_n21699_, new_n21698_, new_n332_ );
and  ( new_n21700_, new_n21699_, new_n328_ );
not  ( new_n21701_, RIbb31758_132 );
or   ( new_n21702_, new_n317_, new_n21701_ );
not  ( new_n21703_, RIbb316e0_131 );
or   ( new_n21704_, new_n320_, new_n21703_ );
and  ( new_n21705_, new_n21704_, new_n21702_ );
xor  ( new_n21706_, new_n21705_, new_n312_ );
not  ( new_n21707_, new_n21706_ );
nor  ( new_n21708_, new_n21699_, new_n328_ );
nor  ( new_n21709_, new_n21708_, new_n21707_ );
nor  ( new_n21710_, new_n21709_, new_n21700_ );
xor  ( new_n21711_, new_n21710_, new_n21693_ );
or   ( new_n21712_, new_n283_, new_n21674_ );
or   ( new_n21713_, new_n286_, new_n21701_ );
and  ( new_n21714_, new_n21713_, new_n21712_ );
xor  ( new_n21715_, new_n21714_, new_n278_ );
or   ( new_n21716_, new_n317_, new_n21703_ );
or   ( new_n21717_, new_n320_, new_n21694_ );
and  ( new_n21718_, new_n21717_, new_n21716_ );
xor  ( new_n21719_, new_n21718_, new_n312_ );
and  ( new_n21720_, new_n336_, RIbb315f0_129 );
xor  ( new_n21721_, new_n21720_, new_n332_ );
not  ( new_n21722_, new_n21721_ );
xor  ( new_n21723_, new_n21722_, new_n21719_ );
xor  ( new_n21724_, new_n21723_, new_n21715_ );
nand ( new_n21725_, new_n21724_, new_n21711_ );
and  ( new_n21726_, RIbb31b18_140, RIbb2f610_1 );
or   ( new_n21727_, new_n337_, new_n21703_ );
or   ( new_n21728_, new_n340_, new_n21694_ );
and  ( new_n21729_, new_n21728_, new_n21727_ );
xor  ( new_n21730_, new_n21729_, new_n331_ );
and  ( new_n21731_, new_n373_, RIbb315f0_129 );
xor  ( new_n21732_, new_n21731_, new_n328_ );
nand ( new_n21733_, new_n21732_, new_n21730_ );
or   ( new_n21734_, new_n317_, new_n21674_ );
or   ( new_n21735_, new_n320_, new_n21701_ );
and  ( new_n21736_, new_n21735_, new_n21734_ );
xor  ( new_n21737_, new_n21736_, new_n312_ );
nor  ( new_n21738_, new_n21732_, new_n21730_ );
or   ( new_n21739_, new_n21738_, new_n21737_ );
and  ( new_n21740_, new_n21739_, new_n21733_ );
nor  ( new_n21741_, new_n21740_, new_n21726_ );
or   ( new_n21742_, new_n283_, new_n21680_ );
or   ( new_n21743_, new_n286_, new_n21672_ );
and  ( new_n21744_, new_n21743_, new_n21742_ );
xor  ( new_n21745_, new_n21744_, new_n278_ );
or   ( new_n21746_, new_n299_, new_n21687_ );
or   ( new_n21747_, new_n302_, new_n21678_ );
and  ( new_n21748_, new_n21747_, new_n21746_ );
xor  ( new_n21749_, new_n21748_, new_n293_ );
nor  ( new_n21750_, new_n21749_, new_n21745_ );
not  ( new_n21751_, RIbb31aa0_139 );
or   ( new_n21752_, new_n268_, new_n21751_ );
or   ( new_n21753_, new_n271_, new_n21685_ );
and  ( new_n21754_, new_n21753_, new_n21752_ );
xor  ( new_n21755_, new_n21754_, new_n263_ );
and  ( new_n21756_, new_n21749_, new_n21745_ );
nor  ( new_n21757_, new_n21756_, new_n21755_ );
nor  ( new_n21758_, new_n21757_, new_n21750_ );
and  ( new_n21759_, new_n21740_, new_n21726_ );
nor  ( new_n21760_, new_n21759_, new_n21758_ );
nor  ( new_n21761_, new_n21760_, new_n21741_ );
not  ( new_n21762_, new_n21761_ );
or   ( new_n21763_, new_n21751_, new_n260_ );
xnor ( new_n21764_, new_n21683_, new_n21677_ );
xor  ( new_n21765_, new_n21764_, new_n21690_ );
and  ( new_n21766_, new_n21765_, new_n21763_ );
nor  ( new_n21767_, new_n21765_, new_n21763_ );
not  ( new_n21768_, new_n21767_ );
xor  ( new_n21769_, new_n21699_, new_n328_ );
xor  ( new_n21770_, new_n21769_, new_n21707_ );
and  ( new_n21771_, new_n21770_, new_n21768_ );
nor  ( new_n21772_, new_n21771_, new_n21766_ );
not  ( new_n21773_, new_n21772_ );
or   ( new_n21774_, new_n21773_, new_n21762_ );
and  ( new_n21775_, new_n21773_, new_n21762_ );
or   ( new_n21776_, new_n21685_, new_n260_ );
or   ( new_n21777_, new_n299_, new_n21680_ );
or   ( new_n21778_, new_n302_, new_n21672_ );
and  ( new_n21779_, new_n21778_, new_n21777_ );
xor  ( new_n21780_, new_n21779_, new_n293_ );
or   ( new_n21781_, new_n268_, new_n21687_ );
or   ( new_n21782_, new_n271_, new_n21678_ );
and  ( new_n21783_, new_n21782_, new_n21781_ );
xor  ( new_n21784_, new_n21783_, new_n263_ );
xor  ( new_n21785_, new_n21784_, new_n21780_ );
xor  ( new_n21786_, new_n21785_, new_n21776_ );
or   ( new_n21787_, new_n21786_, new_n21775_ );
and  ( new_n21788_, new_n21787_, new_n21774_ );
xnor ( new_n21789_, new_n21788_, new_n21725_ );
xor  ( new_n21790_, new_n21789_, new_n21635_ );
xnor ( new_n21791_, new_n21790_, new_n21671_ );
not  ( new_n21792_, RIbb31b18_140 );
or   ( new_n21793_, new_n268_, new_n21792_ );
or   ( new_n21794_, new_n271_, new_n21751_ );
and  ( new_n21795_, new_n21794_, new_n21793_ );
xor  ( new_n21796_, new_n21795_, new_n263_ );
and  ( new_n21797_, RIbb31b90_141, RIbb2f610_1 );
nand ( new_n21798_, new_n21797_, new_n21796_ );
or   ( new_n21799_, new_n317_, new_n21672_ );
or   ( new_n21800_, new_n320_, new_n21674_ );
and  ( new_n21801_, new_n21800_, new_n21799_ );
xor  ( new_n21802_, new_n21801_, new_n312_ );
or   ( new_n21803_, new_n283_, new_n21678_ );
or   ( new_n21804_, new_n286_, new_n21680_ );
and  ( new_n21805_, new_n21804_, new_n21803_ );
xor  ( new_n21806_, new_n21805_, new_n278_ );
and  ( new_n21807_, new_n21806_, new_n21802_ );
or   ( new_n21808_, new_n21806_, new_n21802_ );
or   ( new_n21809_, new_n299_, new_n21685_ );
or   ( new_n21810_, new_n302_, new_n21687_ );
and  ( new_n21811_, new_n21810_, new_n21809_ );
xor  ( new_n21812_, new_n21811_, new_n293_ );
and  ( new_n21813_, new_n21812_, new_n21808_ );
nor  ( new_n21814_, new_n21813_, new_n21807_ );
or   ( new_n21815_, new_n337_, new_n21701_ );
or   ( new_n21816_, new_n340_, new_n21703_ );
and  ( new_n21817_, new_n21816_, new_n21815_ );
xor  ( new_n21818_, new_n21817_, new_n332_ );
and  ( new_n21819_, new_n21818_, new_n403_ );
or   ( new_n21820_, new_n21818_, new_n403_ );
or   ( new_n21821_, new_n409_, new_n21694_ );
or   ( new_n21822_, new_n411_, new_n21696_ );
and  ( new_n21823_, new_n21822_, new_n21821_ );
xor  ( new_n21824_, new_n21823_, new_n328_ );
and  ( new_n21825_, new_n21824_, new_n21820_ );
nor  ( new_n21826_, new_n21825_, new_n21819_ );
xor  ( new_n21827_, new_n21826_, new_n21814_ );
xor  ( new_n21828_, new_n21827_, new_n21798_ );
xor  ( new_n21829_, new_n21797_, new_n21796_ );
xor  ( new_n21830_, new_n21806_, new_n21802_ );
xor  ( new_n21831_, new_n21830_, new_n21812_ );
xor  ( new_n21832_, new_n21818_, new_n403_ );
xor  ( new_n21833_, new_n21832_, new_n21824_ );
xnor ( new_n21834_, new_n21833_, new_n21831_ );
xor  ( new_n21835_, new_n21834_, new_n21829_ );
or   ( new_n21836_, new_n299_, new_n21792_ );
or   ( new_n21837_, new_n302_, new_n21751_ );
and  ( new_n21838_, new_n21837_, new_n21836_ );
xor  ( new_n21839_, new_n21838_, new_n293_ );
not  ( new_n21840_, RIbb31c08_142 );
or   ( new_n21841_, new_n268_, new_n21840_ );
not  ( new_n21842_, RIbb31b90_141 );
or   ( new_n21843_, new_n271_, new_n21842_ );
and  ( new_n21844_, new_n21843_, new_n21841_ );
xor  ( new_n21845_, new_n21844_, new_n263_ );
nor  ( new_n21846_, new_n21845_, new_n21839_ );
not  ( new_n21847_, RIbb31c80_143 );
or   ( new_n21848_, new_n21847_, new_n260_ );
nand ( new_n21849_, new_n21845_, new_n21839_ );
and  ( new_n21850_, new_n21849_, new_n21848_ );
or   ( new_n21851_, new_n21850_, new_n21846_ );
or   ( new_n21852_, new_n524_, new_n21694_ );
or   ( new_n21853_, new_n526_, new_n21696_ );
and  ( new_n21854_, new_n21853_, new_n21852_ );
xor  ( new_n21855_, new_n21854_, new_n403_ );
nand ( new_n21856_, new_n21855_, new_n523_ );
nor  ( new_n21857_, new_n21855_, new_n523_ );
or   ( new_n21858_, new_n409_, new_n21701_ );
or   ( new_n21859_, new_n411_, new_n21703_ );
and  ( new_n21860_, new_n21859_, new_n21858_ );
xor  ( new_n21861_, new_n21860_, new_n327_ );
or   ( new_n21862_, new_n21861_, new_n21857_ );
and  ( new_n21863_, new_n21862_, new_n21856_ );
or   ( new_n21864_, new_n21863_, new_n21851_ );
and  ( new_n21865_, new_n21863_, new_n21851_ );
or   ( new_n21866_, new_n337_, new_n21672_ );
or   ( new_n21867_, new_n340_, new_n21674_ );
and  ( new_n21868_, new_n21867_, new_n21866_ );
xor  ( new_n21869_, new_n21868_, new_n332_ );
or   ( new_n21870_, new_n317_, new_n21678_ );
or   ( new_n21871_, new_n320_, new_n21680_ );
and  ( new_n21872_, new_n21871_, new_n21870_ );
xor  ( new_n21873_, new_n21872_, new_n312_ );
and  ( new_n21874_, new_n21873_, new_n21869_ );
nor  ( new_n21875_, new_n21873_, new_n21869_ );
or   ( new_n21876_, new_n283_, new_n21685_ );
or   ( new_n21877_, new_n286_, new_n21687_ );
and  ( new_n21878_, new_n21877_, new_n21876_ );
xor  ( new_n21879_, new_n21878_, new_n278_ );
not  ( new_n21880_, new_n21879_ );
nor  ( new_n21881_, new_n21880_, new_n21875_ );
nor  ( new_n21882_, new_n21881_, new_n21874_ );
or   ( new_n21883_, new_n21882_, new_n21865_ );
and  ( new_n21884_, new_n21883_, new_n21864_ );
or   ( new_n21885_, new_n21884_, new_n21835_ );
and  ( new_n21886_, new_n21884_, new_n21835_ );
or   ( new_n21887_, new_n337_, new_n21674_ );
or   ( new_n21888_, new_n340_, new_n21701_ );
and  ( new_n21889_, new_n21888_, new_n21887_ );
xor  ( new_n21890_, new_n21889_, new_n332_ );
or   ( new_n21891_, new_n409_, new_n21703_ );
or   ( new_n21892_, new_n411_, new_n21694_ );
and  ( new_n21893_, new_n21892_, new_n21891_ );
xor  ( new_n21894_, new_n21893_, new_n327_ );
and  ( new_n21895_, new_n456_, RIbb315f0_129 );
xor  ( new_n21896_, new_n21895_, new_n403_ );
xnor ( new_n21897_, new_n21896_, new_n21894_ );
xor  ( new_n21898_, new_n21897_, new_n21890_ );
or   ( new_n21899_, new_n299_, new_n21751_ );
or   ( new_n21900_, new_n302_, new_n21685_ );
and  ( new_n21901_, new_n21900_, new_n21899_ );
xor  ( new_n21902_, new_n21901_, new_n293_ );
or   ( new_n21903_, new_n317_, new_n21680_ );
or   ( new_n21904_, new_n320_, new_n21672_ );
and  ( new_n21905_, new_n21904_, new_n21903_ );
xor  ( new_n21906_, new_n21905_, new_n312_ );
or   ( new_n21907_, new_n283_, new_n21687_ );
or   ( new_n21908_, new_n286_, new_n21678_ );
and  ( new_n21909_, new_n21908_, new_n21907_ );
xor  ( new_n21910_, new_n21909_, new_n278_ );
xnor ( new_n21911_, new_n21910_, new_n21906_ );
xor  ( new_n21912_, new_n21911_, new_n21902_ );
or   ( new_n21913_, new_n21912_, new_n21898_ );
and  ( new_n21914_, new_n21912_, new_n21898_ );
or   ( new_n21915_, new_n268_, new_n21842_ );
or   ( new_n21916_, new_n271_, new_n21792_ );
and  ( new_n21917_, new_n21916_, new_n21915_ );
xor  ( new_n21918_, new_n21917_, new_n263_ );
and  ( new_n21919_, RIbb31c08_142, RIbb2f610_1 );
xor  ( new_n21920_, new_n21919_, new_n21918_ );
or   ( new_n21921_, new_n21920_, new_n21914_ );
and  ( new_n21922_, new_n21921_, new_n21913_ );
or   ( new_n21923_, new_n21922_, new_n21886_ );
and  ( new_n21924_, new_n21923_, new_n21885_ );
xnor ( new_n21925_, new_n21924_, new_n21828_ );
xnor ( new_n21926_, new_n21749_, new_n21745_ );
xor  ( new_n21927_, new_n21926_, new_n21755_ );
xnor ( new_n21928_, new_n21732_, new_n21730_ );
xor  ( new_n21929_, new_n21928_, new_n21737_ );
xor  ( new_n21930_, new_n21929_, new_n21927_ );
xnor ( new_n21931_, new_n21930_, new_n21726_ );
or   ( new_n21932_, new_n21919_, new_n21918_ );
nand ( new_n21933_, new_n21896_, new_n21894_ );
nor  ( new_n21934_, new_n21896_, new_n21894_ );
or   ( new_n21935_, new_n21934_, new_n21890_ );
and  ( new_n21936_, new_n21935_, new_n21933_ );
or   ( new_n21937_, new_n21936_, new_n21932_ );
and  ( new_n21938_, new_n21936_, new_n21932_ );
or   ( new_n21939_, new_n21910_, new_n21906_ );
and  ( new_n21940_, new_n21910_, new_n21906_ );
or   ( new_n21941_, new_n21940_, new_n21902_ );
and  ( new_n21942_, new_n21941_, new_n21939_ );
or   ( new_n21943_, new_n21942_, new_n21938_ );
and  ( new_n21944_, new_n21943_, new_n21937_ );
xor  ( new_n21945_, new_n21944_, new_n21931_ );
or   ( new_n21946_, new_n21833_, new_n21831_ );
and  ( new_n21947_, new_n21833_, new_n21831_ );
or   ( new_n21948_, new_n21947_, new_n21829_ );
and  ( new_n21949_, new_n21948_, new_n21946_ );
xor  ( new_n21950_, new_n21949_, new_n21945_ );
xor  ( new_n21951_, new_n21950_, new_n21925_ );
xor  ( new_n21952_, new_n21912_, new_n21898_ );
xor  ( new_n21953_, new_n21952_, new_n21920_ );
xor  ( new_n21954_, new_n21855_, new_n523_ );
xor  ( new_n21955_, new_n21954_, new_n21861_ );
xor  ( new_n21956_, new_n21845_, new_n21839_ );
xor  ( new_n21957_, new_n21956_, new_n21848_ );
or   ( new_n21958_, new_n21957_, new_n21955_ );
and  ( new_n21959_, new_n21957_, new_n21955_ );
xor  ( new_n21960_, new_n21873_, new_n21869_ );
xor  ( new_n21961_, new_n21960_, new_n21880_ );
or   ( new_n21962_, new_n21961_, new_n21959_ );
and  ( new_n21963_, new_n21962_, new_n21958_ );
nor  ( new_n21964_, new_n21963_, new_n21953_ );
nand ( new_n21965_, new_n21963_, new_n21953_ );
or   ( new_n21966_, new_n337_, new_n21680_ );
or   ( new_n21967_, new_n340_, new_n21672_ );
and  ( new_n21968_, new_n21967_, new_n21966_ );
xor  ( new_n21969_, new_n21968_, new_n332_ );
or   ( new_n21970_, new_n317_, new_n21687_ );
or   ( new_n21971_, new_n320_, new_n21678_ );
and  ( new_n21972_, new_n21971_, new_n21970_ );
xor  ( new_n21973_, new_n21972_, new_n312_ );
and  ( new_n21974_, new_n21973_, new_n21969_ );
or   ( new_n21975_, new_n21973_, new_n21969_ );
or   ( new_n21976_, new_n283_, new_n21751_ );
or   ( new_n21977_, new_n286_, new_n21685_ );
and  ( new_n21978_, new_n21977_, new_n21976_ );
xor  ( new_n21979_, new_n21978_, new_n278_ );
and  ( new_n21980_, new_n21979_, new_n21975_ );
or   ( new_n21981_, new_n21980_, new_n21974_ );
or   ( new_n21982_, new_n524_, new_n21703_ );
or   ( new_n21983_, new_n526_, new_n21694_ );
and  ( new_n21984_, new_n21983_, new_n21982_ );
xor  ( new_n21985_, new_n21984_, new_n402_ );
and  ( new_n21986_, new_n662_, RIbb315f0_129 );
xor  ( new_n21987_, new_n21986_, new_n523_ );
nand ( new_n21988_, new_n21987_, new_n21985_ );
nor  ( new_n21989_, new_n21987_, new_n21985_ );
or   ( new_n21990_, new_n409_, new_n21674_ );
or   ( new_n21991_, new_n411_, new_n21701_ );
and  ( new_n21992_, new_n21991_, new_n21990_ );
xor  ( new_n21993_, new_n21992_, new_n328_ );
or   ( new_n21994_, new_n21993_, new_n21989_ );
and  ( new_n21995_, new_n21994_, new_n21988_ );
and  ( new_n21996_, new_n21995_, new_n21981_ );
or   ( new_n21997_, new_n21995_, new_n21981_ );
or   ( new_n21998_, new_n299_, new_n21842_ );
or   ( new_n21999_, new_n302_, new_n21792_ );
and  ( new_n22000_, new_n21999_, new_n21998_ );
xor  ( new_n22001_, new_n22000_, new_n293_ );
or   ( new_n22002_, new_n268_, new_n21847_ );
or   ( new_n22003_, new_n271_, new_n21840_ );
and  ( new_n22004_, new_n22003_, new_n22002_ );
xor  ( new_n22005_, new_n22004_, new_n263_ );
or   ( new_n22006_, new_n22005_, new_n22001_ );
and  ( new_n22007_, RIbb31cf8_144, RIbb2f610_1 );
and  ( new_n22008_, new_n22005_, new_n22001_ );
or   ( new_n22009_, new_n22008_, new_n22007_ );
and  ( new_n22010_, new_n22009_, new_n22006_ );
and  ( new_n22011_, new_n22010_, new_n21997_ );
or   ( new_n22012_, new_n22011_, new_n21996_ );
and  ( new_n22013_, new_n22012_, new_n21965_ );
or   ( new_n22014_, new_n22013_, new_n21964_ );
xor  ( new_n22015_, new_n21936_, new_n21932_ );
xor  ( new_n22016_, new_n22015_, new_n21942_ );
nand ( new_n22017_, new_n22016_, new_n22014_ );
nor  ( new_n22018_, new_n22016_, new_n22014_ );
xor  ( new_n22019_, new_n21884_, new_n21835_ );
xor  ( new_n22020_, new_n22019_, new_n21922_ );
or   ( new_n22021_, new_n22020_, new_n22018_ );
and  ( new_n22022_, new_n22021_, new_n22017_ );
nor  ( new_n22023_, new_n22022_, new_n21951_ );
xor  ( new_n22024_, new_n21765_, new_n21763_ );
xor  ( new_n22025_, new_n22024_, new_n21770_ );
or   ( new_n22026_, new_n21929_, new_n21927_ );
and  ( new_n22027_, new_n21929_, new_n21927_ );
or   ( new_n22028_, new_n22027_, new_n21726_ );
and  ( new_n22029_, new_n22028_, new_n22026_ );
xor  ( new_n22030_, new_n22029_, new_n22025_ );
or   ( new_n22031_, new_n21826_, new_n21814_ );
and  ( new_n22032_, new_n21826_, new_n21814_ );
or   ( new_n22033_, new_n22032_, new_n21798_ );
and  ( new_n22034_, new_n22033_, new_n22031_ );
xor  ( new_n22035_, new_n22034_, new_n22030_ );
xnor ( new_n22036_, new_n21740_, new_n21726_ );
xor  ( new_n22037_, new_n22036_, new_n21758_ );
xor  ( new_n22038_, new_n22037_, new_n22035_ );
nor  ( new_n22039_, new_n21944_, new_n21931_ );
and  ( new_n22040_, new_n21944_, new_n21931_ );
nor  ( new_n22041_, new_n21949_, new_n22040_ );
nor  ( new_n22042_, new_n22041_, new_n22039_ );
not  ( new_n22043_, new_n22042_ );
xor  ( new_n22044_, new_n22043_, new_n22038_ );
nor  ( new_n22045_, new_n21924_, new_n21828_ );
nand ( new_n22046_, new_n21924_, new_n21828_ );
and  ( new_n22047_, new_n21950_, new_n22046_ );
nor  ( new_n22048_, new_n22047_, new_n22045_ );
xor  ( new_n22049_, new_n22048_, new_n22044_ );
and  ( new_n22050_, new_n22049_, new_n22023_ );
xor  ( new_n22051_, new_n21963_, new_n21953_ );
xor  ( new_n22052_, new_n22051_, new_n22012_ );
xor  ( new_n22053_, new_n22005_, new_n22001_ );
xnor ( new_n22054_, new_n22053_, new_n22007_ );
xnor ( new_n22055_, new_n21973_, new_n21969_ );
xor  ( new_n22056_, new_n22055_, new_n21979_ );
nand ( new_n22057_, new_n22056_, new_n22054_ );
or   ( new_n22058_, new_n409_, new_n21672_ );
or   ( new_n22059_, new_n411_, new_n21674_ );
and  ( new_n22060_, new_n22059_, new_n22058_ );
xor  ( new_n22061_, new_n22060_, new_n328_ );
or   ( new_n22062_, new_n337_, new_n21678_ );
or   ( new_n22063_, new_n340_, new_n21680_ );
and  ( new_n22064_, new_n22063_, new_n22062_ );
xor  ( new_n22065_, new_n22064_, new_n332_ );
nor  ( new_n22066_, new_n22065_, new_n22061_ );
nand ( new_n22067_, new_n22065_, new_n22061_ );
or   ( new_n22068_, new_n317_, new_n21685_ );
or   ( new_n22069_, new_n320_, new_n21687_ );
and  ( new_n22070_, new_n22069_, new_n22068_ );
xor  ( new_n22071_, new_n22070_, new_n311_ );
and  ( new_n22072_, new_n22071_, new_n22067_ );
or   ( new_n22073_, new_n22072_, new_n22066_ );
or   ( new_n22074_, new_n524_, new_n21701_ );
or   ( new_n22075_, new_n526_, new_n21703_ );
and  ( new_n22076_, new_n22075_, new_n22074_ );
xor  ( new_n22077_, new_n22076_, new_n403_ );
nand ( new_n22078_, new_n22077_, new_n748_ );
or   ( new_n22079_, new_n22077_, new_n748_ );
or   ( new_n22080_, new_n755_, new_n21694_ );
or   ( new_n22081_, new_n757_, new_n21696_ );
and  ( new_n22082_, new_n22081_, new_n22080_ );
xor  ( new_n22083_, new_n22082_, new_n523_ );
nand ( new_n22084_, new_n22083_, new_n22079_ );
and  ( new_n22085_, new_n22084_, new_n22078_ );
nand ( new_n22086_, new_n22085_, new_n22073_ );
nor  ( new_n22087_, new_n22085_, new_n22073_ );
or   ( new_n22088_, new_n283_, new_n21792_ );
or   ( new_n22089_, new_n286_, new_n21751_ );
and  ( new_n22090_, new_n22089_, new_n22088_ );
xor  ( new_n22091_, new_n22090_, new_n278_ );
or   ( new_n22092_, new_n299_, new_n21840_ );
or   ( new_n22093_, new_n302_, new_n21842_ );
and  ( new_n22094_, new_n22093_, new_n22092_ );
xor  ( new_n22095_, new_n22094_, new_n293_ );
nor  ( new_n22096_, new_n22095_, new_n22091_ );
and  ( new_n22097_, new_n22095_, new_n22091_ );
not  ( new_n22098_, RIbb31cf8_144 );
or   ( new_n22099_, new_n268_, new_n22098_ );
or   ( new_n22100_, new_n271_, new_n21847_ );
and  ( new_n22101_, new_n22100_, new_n22099_ );
xor  ( new_n22102_, new_n22101_, new_n263_ );
nor  ( new_n22103_, new_n22102_, new_n22097_ );
nor  ( new_n22104_, new_n22103_, new_n22096_ );
or   ( new_n22105_, new_n22104_, new_n22087_ );
and  ( new_n22106_, new_n22105_, new_n22086_ );
or   ( new_n22107_, new_n22106_, new_n22057_ );
and  ( new_n22108_, new_n22106_, new_n22057_ );
xor  ( new_n22109_, new_n21957_, new_n21955_ );
xnor ( new_n22110_, new_n22109_, new_n21961_ );
or   ( new_n22111_, new_n22110_, new_n22108_ );
and  ( new_n22112_, new_n22111_, new_n22107_ );
nor  ( new_n22113_, new_n22112_, new_n22052_ );
and  ( new_n22114_, new_n22112_, new_n22052_ );
xor  ( new_n22115_, new_n21863_, new_n21851_ );
xnor ( new_n22116_, new_n22115_, new_n21882_ );
nor  ( new_n22117_, new_n22116_, new_n22114_ );
nor  ( new_n22118_, new_n22117_, new_n22113_ );
xor  ( new_n22119_, new_n22016_, new_n22014_ );
xnor ( new_n22120_, new_n22119_, new_n22020_ );
and  ( new_n22121_, new_n22120_, new_n22118_ );
xor  ( new_n22122_, new_n22022_, new_n21951_ );
and  ( new_n22123_, new_n22122_, new_n22121_ );
xnor ( new_n22124_, new_n22120_, new_n22118_ );
xor  ( new_n22125_, new_n22085_, new_n22073_ );
xnor ( new_n22126_, new_n22125_, new_n22104_ );
xor  ( new_n22127_, new_n21987_, new_n21985_ );
xnor ( new_n22128_, new_n22127_, new_n21993_ );
not  ( new_n22129_, RIbb31d70_145 );
or   ( new_n22130_, new_n22129_, new_n260_ );
xor  ( new_n22131_, new_n22065_, new_n22061_ );
xor  ( new_n22132_, new_n22131_, new_n22071_ );
nand ( new_n22133_, new_n22132_, new_n22130_ );
nor  ( new_n22134_, new_n22132_, new_n22130_ );
xor  ( new_n22135_, new_n22095_, new_n22091_ );
xor  ( new_n22136_, new_n22135_, new_n22102_ );
or   ( new_n22137_, new_n22136_, new_n22134_ );
and  ( new_n22138_, new_n22137_, new_n22133_ );
xor  ( new_n22139_, new_n22138_, new_n22128_ );
or   ( new_n22140_, new_n755_, new_n21703_ );
or   ( new_n22141_, new_n757_, new_n21694_ );
and  ( new_n22142_, new_n22141_, new_n22140_ );
xor  ( new_n22143_, new_n22142_, new_n522_ );
and  ( new_n22144_, new_n822_, RIbb315f0_129 );
xor  ( new_n22145_, new_n22144_, new_n748_ );
nand ( new_n22146_, new_n22145_, new_n22143_ );
nor  ( new_n22147_, new_n22145_, new_n22143_ );
or   ( new_n22148_, new_n524_, new_n21674_ );
or   ( new_n22149_, new_n526_, new_n21701_ );
and  ( new_n22150_, new_n22149_, new_n22148_ );
xor  ( new_n22151_, new_n22150_, new_n403_ );
or   ( new_n22152_, new_n22151_, new_n22147_ );
and  ( new_n22153_, new_n22152_, new_n22146_ );
or   ( new_n22154_, new_n409_, new_n21680_ );
or   ( new_n22155_, new_n411_, new_n21672_ );
and  ( new_n22156_, new_n22155_, new_n22154_ );
xor  ( new_n22157_, new_n22156_, new_n328_ );
or   ( new_n22158_, new_n337_, new_n21687_ );
or   ( new_n22159_, new_n340_, new_n21678_ );
and  ( new_n22160_, new_n22159_, new_n22158_ );
xor  ( new_n22161_, new_n22160_, new_n332_ );
or   ( new_n22162_, new_n22161_, new_n22157_ );
and  ( new_n22163_, new_n22161_, new_n22157_ );
or   ( new_n22164_, new_n317_, new_n21751_ );
or   ( new_n22165_, new_n320_, new_n21685_ );
and  ( new_n22166_, new_n22165_, new_n22164_ );
xor  ( new_n22167_, new_n22166_, new_n312_ );
or   ( new_n22168_, new_n22167_, new_n22163_ );
and  ( new_n22169_, new_n22168_, new_n22162_ );
or   ( new_n22170_, new_n22169_, new_n22153_ );
and  ( new_n22171_, new_n22169_, new_n22153_ );
or   ( new_n22172_, new_n283_, new_n21842_ );
or   ( new_n22173_, new_n286_, new_n21792_ );
and  ( new_n22174_, new_n22173_, new_n22172_ );
xor  ( new_n22175_, new_n22174_, new_n278_ );
or   ( new_n22176_, new_n299_, new_n21847_ );
or   ( new_n22177_, new_n302_, new_n21840_ );
and  ( new_n22178_, new_n22177_, new_n22176_ );
xor  ( new_n22179_, new_n22178_, new_n293_ );
nor  ( new_n22180_, new_n22179_, new_n22175_ );
and  ( new_n22181_, new_n22179_, new_n22175_ );
or   ( new_n22182_, new_n268_, new_n22129_ );
or   ( new_n22183_, new_n271_, new_n22098_ );
and  ( new_n22184_, new_n22183_, new_n22182_ );
xor  ( new_n22185_, new_n22184_, new_n263_ );
nor  ( new_n22186_, new_n22185_, new_n22181_ );
nor  ( new_n22187_, new_n22186_, new_n22180_ );
or   ( new_n22188_, new_n22187_, new_n22171_ );
and  ( new_n22189_, new_n22188_, new_n22170_ );
xor  ( new_n22190_, new_n22189_, new_n22139_ );
nor  ( new_n22191_, new_n22190_, new_n22126_ );
xor  ( new_n22192_, new_n22132_, new_n22130_ );
xor  ( new_n22193_, new_n22192_, new_n22136_ );
xor  ( new_n22194_, new_n22077_, new_n748_ );
xor  ( new_n22195_, new_n22194_, new_n22083_ );
or   ( new_n22196_, new_n22195_, new_n22193_ );
nand ( new_n22197_, new_n22195_, new_n22193_ );
xor  ( new_n22198_, new_n22169_, new_n22153_ );
xnor ( new_n22199_, new_n22198_, new_n22187_ );
nand ( new_n22200_, new_n22199_, new_n22197_ );
and  ( new_n22201_, new_n22200_, new_n22196_ );
xor  ( new_n22202_, new_n22161_, new_n22157_ );
xnor ( new_n22203_, new_n22202_, new_n22167_ );
xnor ( new_n22204_, new_n22145_, new_n22143_ );
xor  ( new_n22205_, new_n22204_, new_n22151_ );
or   ( new_n22206_, new_n22205_, new_n22203_ );
not  ( new_n22207_, RIbb31de8_146 );
or   ( new_n22208_, new_n22207_, new_n260_ );
xnor ( new_n22209_, new_n22179_, new_n22175_ );
xor  ( new_n22210_, new_n22209_, new_n22185_ );
and  ( new_n22211_, new_n22210_, new_n22208_ );
nand ( new_n22212_, new_n22211_, new_n22206_ );
nor  ( new_n22213_, new_n22211_, new_n22206_ );
or   ( new_n22214_, new_n897_, new_n21694_ );
or   ( new_n22215_, new_n899_, new_n21696_ );
and  ( new_n22216_, new_n22215_, new_n22214_ );
xor  ( new_n22217_, new_n22216_, new_n748_ );
and  ( new_n22218_, new_n22217_, new_n896_ );
or   ( new_n22219_, new_n22217_, new_n896_ );
or   ( new_n22220_, new_n755_, new_n21701_ );
or   ( new_n22221_, new_n757_, new_n21703_ );
and  ( new_n22222_, new_n22221_, new_n22220_ );
xor  ( new_n22223_, new_n22222_, new_n523_ );
and  ( new_n22224_, new_n22223_, new_n22219_ );
or   ( new_n22225_, new_n22224_, new_n22218_ );
or   ( new_n22226_, new_n524_, new_n21672_ );
or   ( new_n22227_, new_n526_, new_n21674_ );
and  ( new_n22228_, new_n22227_, new_n22226_ );
xor  ( new_n22229_, new_n22228_, new_n403_ );
or   ( new_n22230_, new_n409_, new_n21678_ );
or   ( new_n22231_, new_n411_, new_n21680_ );
and  ( new_n22232_, new_n22231_, new_n22230_ );
xor  ( new_n22233_, new_n22232_, new_n328_ );
or   ( new_n22234_, new_n22233_, new_n22229_ );
and  ( new_n22235_, new_n22233_, new_n22229_ );
or   ( new_n22236_, new_n337_, new_n21685_ );
or   ( new_n22237_, new_n340_, new_n21687_ );
and  ( new_n22238_, new_n22237_, new_n22236_ );
xor  ( new_n22239_, new_n22238_, new_n332_ );
or   ( new_n22240_, new_n22239_, new_n22235_ );
and  ( new_n22241_, new_n22240_, new_n22234_ );
nor  ( new_n22242_, new_n22241_, new_n22225_ );
and  ( new_n22243_, new_n22241_, new_n22225_ );
or   ( new_n22244_, new_n317_, new_n21792_ );
or   ( new_n22245_, new_n320_, new_n21751_ );
and  ( new_n22246_, new_n22245_, new_n22244_ );
xor  ( new_n22247_, new_n22246_, new_n312_ );
or   ( new_n22248_, new_n283_, new_n21840_ );
or   ( new_n22249_, new_n286_, new_n21842_ );
and  ( new_n22250_, new_n22249_, new_n22248_ );
xor  ( new_n22251_, new_n22250_, new_n278_ );
nor  ( new_n22252_, new_n22251_, new_n22247_ );
and  ( new_n22253_, new_n22251_, new_n22247_ );
or   ( new_n22254_, new_n299_, new_n22098_ );
or   ( new_n22255_, new_n302_, new_n21847_ );
and  ( new_n22256_, new_n22255_, new_n22254_ );
xor  ( new_n22257_, new_n22256_, new_n293_ );
nor  ( new_n22258_, new_n22257_, new_n22253_ );
nor  ( new_n22259_, new_n22258_, new_n22252_ );
nor  ( new_n22260_, new_n22259_, new_n22243_ );
nor  ( new_n22261_, new_n22260_, new_n22242_ );
or   ( new_n22262_, new_n22261_, new_n22213_ );
and  ( new_n22263_, new_n22262_, new_n22212_ );
or   ( new_n22264_, new_n22263_, new_n22201_ );
and  ( new_n22265_, new_n22263_, new_n22201_ );
xnor ( new_n22266_, new_n22056_, new_n22054_ );
or   ( new_n22267_, new_n22266_, new_n22265_ );
and  ( new_n22268_, new_n22267_, new_n22264_ );
nand ( new_n22269_, new_n22268_, new_n22191_ );
nor  ( new_n22270_, new_n22268_, new_n22191_ );
not  ( new_n22271_, new_n22128_ );
and  ( new_n22272_, new_n22138_, new_n22271_ );
or   ( new_n22273_, new_n22138_, new_n22271_ );
and  ( new_n22274_, new_n22189_, new_n22273_ );
nor  ( new_n22275_, new_n22274_, new_n22272_ );
not  ( new_n22276_, new_n22275_ );
xor  ( new_n22277_, new_n21995_, new_n21981_ );
xor  ( new_n22278_, new_n22277_, new_n22010_ );
xor  ( new_n22279_, new_n22278_, new_n22276_ );
xnor ( new_n22280_, new_n22106_, new_n22057_ );
xor  ( new_n22281_, new_n22280_, new_n22110_ );
xor  ( new_n22282_, new_n22281_, new_n22279_ );
or   ( new_n22283_, new_n22282_, new_n22270_ );
and  ( new_n22284_, new_n22283_, new_n22269_ );
xnor ( new_n22285_, new_n22112_, new_n22052_ );
xor  ( new_n22286_, new_n22285_, new_n22116_ );
or   ( new_n22287_, new_n22286_, new_n22284_ );
and  ( new_n22288_, new_n22286_, new_n22284_ );
nand ( new_n22289_, new_n22278_, new_n22276_ );
nor  ( new_n22290_, new_n22278_, new_n22276_ );
or   ( new_n22291_, new_n22281_, new_n22290_ );
and  ( new_n22292_, new_n22291_, new_n22289_ );
or   ( new_n22293_, new_n22292_, new_n22288_ );
and  ( new_n22294_, new_n22293_, new_n22287_ );
nor  ( new_n22295_, new_n22294_, new_n22124_ );
xor  ( new_n22296_, new_n22210_, new_n22208_ );
xnor ( new_n22297_, new_n22241_, new_n22225_ );
xor  ( new_n22298_, new_n22297_, new_n22259_ );
nor  ( new_n22299_, new_n22298_, new_n22296_ );
nand ( new_n22300_, new_n22298_, new_n22296_ );
xor  ( new_n22301_, new_n22205_, new_n22203_ );
and  ( new_n22302_, new_n22301_, new_n22300_ );
or   ( new_n22303_, new_n22302_, new_n22299_ );
not  ( new_n22304_, RIbb31e60_147 );
or   ( new_n22305_, new_n268_, new_n22304_ );
or   ( new_n22306_, new_n271_, new_n22207_ );
and  ( new_n22307_, new_n22306_, new_n22305_ );
xor  ( new_n22308_, new_n22307_, new_n263_ );
and  ( new_n22309_, RIbb31ed8_148, RIbb2f610_1 );
or   ( new_n22310_, new_n22309_, new_n22308_ );
or   ( new_n22311_, new_n268_, new_n22207_ );
or   ( new_n22312_, new_n271_, new_n22129_ );
and  ( new_n22313_, new_n22312_, new_n22311_ );
xor  ( new_n22314_, new_n22313_, new_n263_ );
or   ( new_n22315_, new_n22314_, new_n22310_ );
and  ( new_n22316_, new_n22314_, new_n22310_ );
and  ( new_n22317_, RIbb31e60_147, RIbb2f610_1 );
or   ( new_n22318_, new_n22317_, new_n22316_ );
and  ( new_n22319_, new_n22318_, new_n22315_ );
or   ( new_n22320_, new_n524_, new_n21680_ );
or   ( new_n22321_, new_n526_, new_n21672_ );
and  ( new_n22322_, new_n22321_, new_n22320_ );
xor  ( new_n22323_, new_n22322_, new_n403_ );
or   ( new_n22324_, new_n409_, new_n21687_ );
or   ( new_n22325_, new_n411_, new_n21678_ );
and  ( new_n22326_, new_n22325_, new_n22324_ );
xor  ( new_n22327_, new_n22326_, new_n328_ );
or   ( new_n22328_, new_n22327_, new_n22323_ );
and  ( new_n22329_, new_n22327_, new_n22323_ );
or   ( new_n22330_, new_n337_, new_n21751_ );
or   ( new_n22331_, new_n340_, new_n21685_ );
and  ( new_n22332_, new_n22331_, new_n22330_ );
xor  ( new_n22333_, new_n22332_, new_n332_ );
or   ( new_n22334_, new_n22333_, new_n22329_ );
and  ( new_n22335_, new_n22334_, new_n22328_ );
or   ( new_n22336_, new_n317_, new_n21842_ );
or   ( new_n22337_, new_n320_, new_n21792_ );
and  ( new_n22338_, new_n22337_, new_n22336_ );
xor  ( new_n22339_, new_n22338_, new_n312_ );
or   ( new_n22340_, new_n283_, new_n21847_ );
or   ( new_n22341_, new_n286_, new_n21840_ );
and  ( new_n22342_, new_n22341_, new_n22340_ );
xor  ( new_n22343_, new_n22342_, new_n278_ );
or   ( new_n22344_, new_n22343_, new_n22339_ );
and  ( new_n22345_, new_n22343_, new_n22339_ );
or   ( new_n22346_, new_n299_, new_n22129_ );
or   ( new_n22347_, new_n302_, new_n22098_ );
and  ( new_n22348_, new_n22347_, new_n22346_ );
xor  ( new_n22349_, new_n22348_, new_n293_ );
or   ( new_n22350_, new_n22349_, new_n22345_ );
and  ( new_n22351_, new_n22350_, new_n22344_ );
or   ( new_n22352_, new_n22351_, new_n22335_ );
and  ( new_n22353_, new_n22351_, new_n22335_ );
or   ( new_n22354_, new_n897_, new_n21703_ );
or   ( new_n22355_, new_n899_, new_n21694_ );
and  ( new_n22356_, new_n22355_, new_n22354_ );
xor  ( new_n22357_, new_n22356_, new_n747_ );
and  ( new_n22358_, new_n1042_, RIbb315f0_129 );
xor  ( new_n22359_, new_n22358_, new_n896_ );
and  ( new_n22360_, new_n22359_, new_n22357_ );
nor  ( new_n22361_, new_n22359_, new_n22357_ );
or   ( new_n22362_, new_n755_, new_n21674_ );
or   ( new_n22363_, new_n757_, new_n21701_ );
and  ( new_n22364_, new_n22363_, new_n22362_ );
xor  ( new_n22365_, new_n22364_, new_n523_ );
nor  ( new_n22366_, new_n22365_, new_n22361_ );
nor  ( new_n22367_, new_n22366_, new_n22360_ );
or   ( new_n22368_, new_n22367_, new_n22353_ );
and  ( new_n22369_, new_n22368_, new_n22352_ );
or   ( new_n22370_, new_n22369_, new_n22319_ );
nand ( new_n22371_, new_n22369_, new_n22319_ );
xor  ( new_n22372_, new_n22217_, new_n895_ );
xor  ( new_n22373_, new_n22372_, new_n22223_ );
xnor ( new_n22374_, new_n22233_, new_n22229_ );
xor  ( new_n22375_, new_n22374_, new_n22239_ );
nor  ( new_n22376_, new_n22375_, new_n22373_ );
and  ( new_n22377_, new_n22375_, new_n22373_ );
xor  ( new_n22378_, new_n22251_, new_n22247_ );
xnor ( new_n22379_, new_n22378_, new_n22257_ );
nor  ( new_n22380_, new_n22379_, new_n22377_ );
nor  ( new_n22381_, new_n22380_, new_n22376_ );
nand ( new_n22382_, new_n22381_, new_n22371_ );
and  ( new_n22383_, new_n22382_, new_n22370_ );
or   ( new_n22384_, new_n22383_, new_n22303_ );
nand ( new_n22385_, new_n22383_, new_n22303_ );
xor  ( new_n22386_, new_n22195_, new_n22193_ );
xor  ( new_n22387_, new_n22386_, new_n22199_ );
nand ( new_n22388_, new_n22387_, new_n22385_ );
and  ( new_n22389_, new_n22388_, new_n22384_ );
xor  ( new_n22390_, new_n22263_, new_n22201_ );
xor  ( new_n22391_, new_n22390_, new_n22266_ );
or   ( new_n22392_, new_n22391_, new_n22389_ );
and  ( new_n22393_, new_n22391_, new_n22389_ );
xor  ( new_n22394_, new_n22190_, new_n22126_ );
or   ( new_n22395_, new_n22394_, new_n22393_ );
and  ( new_n22396_, new_n22395_, new_n22392_ );
xnor ( new_n22397_, new_n22268_, new_n22191_ );
xor  ( new_n22398_, new_n22397_, new_n22282_ );
nand ( new_n22399_, new_n22398_, new_n22396_ );
xor  ( new_n22400_, new_n22286_, new_n22284_ );
xor  ( new_n22401_, new_n22400_, new_n22292_ );
nor  ( new_n22402_, new_n22401_, new_n22399_ );
xnor ( new_n22403_, new_n22391_, new_n22389_ );
xor  ( new_n22404_, new_n22403_, new_n22394_ );
xnor ( new_n22405_, new_n22298_, new_n22296_ );
xor  ( new_n22406_, new_n22405_, new_n22301_ );
xnor ( new_n22407_, new_n22351_, new_n22335_ );
xor  ( new_n22408_, new_n22407_, new_n22367_ );
xnor ( new_n22409_, new_n22314_, new_n22310_ );
xor  ( new_n22410_, new_n22409_, new_n22317_ );
or   ( new_n22411_, new_n22410_, new_n22408_ );
and  ( new_n22412_, new_n22410_, new_n22408_ );
xor  ( new_n22413_, new_n22375_, new_n22373_ );
xor  ( new_n22414_, new_n22413_, new_n22379_ );
or   ( new_n22415_, new_n22414_, new_n22412_ );
and  ( new_n22416_, new_n22415_, new_n22411_ );
or   ( new_n22417_, new_n22416_, new_n22406_ );
and  ( new_n22418_, new_n22416_, new_n22406_ );
or   ( new_n22419_, new_n299_, new_n22207_ );
or   ( new_n22420_, new_n302_, new_n22129_ );
and  ( new_n22421_, new_n22420_, new_n22419_ );
xor  ( new_n22422_, new_n22421_, new_n293_ );
not  ( new_n22423_, RIbb31ed8_148 );
or   ( new_n22424_, new_n268_, new_n22423_ );
or   ( new_n22425_, new_n271_, new_n22304_ );
and  ( new_n22426_, new_n22425_, new_n22424_ );
xor  ( new_n22427_, new_n22426_, new_n263_ );
nor  ( new_n22428_, new_n22427_, new_n22422_ );
and  ( new_n22429_, RIbb31f50_149, RIbb2f610_1 );
not  ( new_n22430_, new_n22429_ );
nand ( new_n22431_, new_n22427_, new_n22422_ );
and  ( new_n22432_, new_n22431_, new_n22430_ );
or   ( new_n22433_, new_n22432_, new_n22428_ );
xnor ( new_n22434_, new_n22343_, new_n22339_ );
xor  ( new_n22435_, new_n22434_, new_n22349_ );
nor  ( new_n22436_, new_n22435_, new_n22433_ );
and  ( new_n22437_, new_n22435_, new_n22433_ );
xor  ( new_n22438_, new_n22309_, new_n22308_ );
nor  ( new_n22439_, new_n22438_, new_n22437_ );
or   ( new_n22440_, new_n22439_, new_n22436_ );
or   ( new_n22441_, new_n1135_, new_n21694_ );
or   ( new_n22442_, new_n1137_, new_n21696_ );
and  ( new_n22443_, new_n22442_, new_n22441_ );
xor  ( new_n22444_, new_n22443_, new_n896_ );
and  ( new_n22445_, new_n22444_, new_n1129_ );
or   ( new_n22446_, new_n22444_, new_n1129_ );
or   ( new_n22447_, new_n897_, new_n21701_ );
or   ( new_n22448_, new_n899_, new_n21703_ );
and  ( new_n22449_, new_n22448_, new_n22447_ );
xor  ( new_n22450_, new_n22449_, new_n748_ );
and  ( new_n22451_, new_n22450_, new_n22446_ );
or   ( new_n22452_, new_n22451_, new_n22445_ );
or   ( new_n22453_, new_n337_, new_n21792_ );
or   ( new_n22454_, new_n340_, new_n21751_ );
and  ( new_n22455_, new_n22454_, new_n22453_ );
xor  ( new_n22456_, new_n22455_, new_n332_ );
or   ( new_n22457_, new_n317_, new_n21840_ );
or   ( new_n22458_, new_n320_, new_n21842_ );
and  ( new_n22459_, new_n22458_, new_n22457_ );
xor  ( new_n22460_, new_n22459_, new_n312_ );
or   ( new_n22461_, new_n22460_, new_n22456_ );
and  ( new_n22462_, new_n22460_, new_n22456_ );
or   ( new_n22463_, new_n283_, new_n22098_ );
or   ( new_n22464_, new_n286_, new_n21847_ );
and  ( new_n22465_, new_n22464_, new_n22463_ );
xor  ( new_n22466_, new_n22465_, new_n278_ );
or   ( new_n22467_, new_n22466_, new_n22462_ );
and  ( new_n22468_, new_n22467_, new_n22461_ );
or   ( new_n22469_, new_n22468_, new_n22452_ );
and  ( new_n22470_, new_n22468_, new_n22452_ );
or   ( new_n22471_, new_n755_, new_n21672_ );
or   ( new_n22472_, new_n757_, new_n21674_ );
and  ( new_n22473_, new_n22472_, new_n22471_ );
xor  ( new_n22474_, new_n22473_, new_n523_ );
or   ( new_n22475_, new_n524_, new_n21678_ );
or   ( new_n22476_, new_n526_, new_n21680_ );
and  ( new_n22477_, new_n22476_, new_n22475_ );
xor  ( new_n22478_, new_n22477_, new_n403_ );
nor  ( new_n22479_, new_n22478_, new_n22474_ );
and  ( new_n22480_, new_n22478_, new_n22474_ );
or   ( new_n22481_, new_n409_, new_n21685_ );
or   ( new_n22482_, new_n411_, new_n21687_ );
and  ( new_n22483_, new_n22482_, new_n22481_ );
xor  ( new_n22484_, new_n22483_, new_n328_ );
nor  ( new_n22485_, new_n22484_, new_n22480_ );
nor  ( new_n22486_, new_n22485_, new_n22479_ );
or   ( new_n22487_, new_n22486_, new_n22470_ );
and  ( new_n22488_, new_n22487_, new_n22469_ );
nor  ( new_n22489_, new_n22488_, new_n22440_ );
and  ( new_n22490_, new_n22488_, new_n22440_ );
xor  ( new_n22491_, new_n22327_, new_n22323_ );
xnor ( new_n22492_, new_n22491_, new_n22333_ );
xnor ( new_n22493_, new_n22359_, new_n22357_ );
xor  ( new_n22494_, new_n22493_, new_n22365_ );
nor  ( new_n22495_, new_n22494_, new_n22492_ );
nor  ( new_n22496_, new_n22495_, new_n22490_ );
or   ( new_n22497_, new_n22496_, new_n22489_ );
or   ( new_n22498_, new_n22497_, new_n22418_ );
and  ( new_n22499_, new_n22498_, new_n22417_ );
xnor ( new_n22500_, new_n22211_, new_n22206_ );
xor  ( new_n22501_, new_n22500_, new_n22261_ );
or   ( new_n22502_, new_n22501_, new_n22499_ );
and  ( new_n22503_, new_n22501_, new_n22499_ );
xor  ( new_n22504_, new_n22383_, new_n22303_ );
xor  ( new_n22505_, new_n22504_, new_n22387_ );
or   ( new_n22506_, new_n22505_, new_n22503_ );
and  ( new_n22507_, new_n22506_, new_n22502_ );
nor  ( new_n22508_, new_n22507_, new_n22404_ );
xor  ( new_n22509_, new_n22398_, new_n22396_ );
and  ( new_n22510_, new_n22509_, new_n22508_ );
xor  ( new_n22511_, new_n22501_, new_n22499_ );
xor  ( new_n22512_, new_n22511_, new_n22505_ );
xor  ( new_n22513_, new_n22369_, new_n22319_ );
xor  ( new_n22514_, new_n22513_, new_n22381_ );
xor  ( new_n22515_, new_n22410_, new_n22408_ );
xor  ( new_n22516_, new_n22515_, new_n22414_ );
xnor ( new_n22517_, new_n22468_, new_n22452_ );
xor  ( new_n22518_, new_n22517_, new_n22486_ );
xor  ( new_n22519_, new_n22435_, new_n22433_ );
xor  ( new_n22520_, new_n22519_, new_n22438_ );
or   ( new_n22521_, new_n22520_, new_n22518_ );
and  ( new_n22522_, new_n22520_, new_n22518_ );
xnor ( new_n22523_, new_n22494_, new_n22492_ );
or   ( new_n22524_, new_n22523_, new_n22522_ );
and  ( new_n22525_, new_n22524_, new_n22521_ );
or   ( new_n22526_, new_n22525_, new_n22516_ );
and  ( new_n22527_, new_n22525_, new_n22516_ );
xor  ( new_n22528_, new_n22444_, new_n1129_ );
xor  ( new_n22529_, new_n22528_, new_n22450_ );
not  ( new_n22530_, new_n22529_ );
xnor ( new_n22531_, new_n22478_, new_n22474_ );
xor  ( new_n22532_, new_n22531_, new_n22484_ );
nor  ( new_n22533_, new_n22532_, new_n22530_ );
or   ( new_n22534_, new_n337_, new_n21842_ );
or   ( new_n22535_, new_n340_, new_n21792_ );
and  ( new_n22536_, new_n22535_, new_n22534_ );
xor  ( new_n22537_, new_n22536_, new_n332_ );
or   ( new_n22538_, new_n317_, new_n21847_ );
or   ( new_n22539_, new_n320_, new_n21840_ );
and  ( new_n22540_, new_n22539_, new_n22538_ );
xor  ( new_n22541_, new_n22540_, new_n312_ );
or   ( new_n22542_, new_n22541_, new_n22537_ );
and  ( new_n22543_, new_n22541_, new_n22537_ );
or   ( new_n22544_, new_n283_, new_n22129_ );
or   ( new_n22545_, new_n286_, new_n22098_ );
and  ( new_n22546_, new_n22545_, new_n22544_ );
xor  ( new_n22547_, new_n22546_, new_n278_ );
or   ( new_n22548_, new_n22547_, new_n22543_ );
and  ( new_n22549_, new_n22548_, new_n22542_ );
or   ( new_n22550_, new_n1135_, new_n21703_ );
or   ( new_n22551_, new_n1137_, new_n21694_ );
and  ( new_n22552_, new_n22551_, new_n22550_ );
xor  ( new_n22553_, new_n22552_, new_n895_ );
and  ( new_n22554_, new_n1253_, RIbb315f0_129 );
xor  ( new_n22555_, new_n22554_, new_n1129_ );
nand ( new_n22556_, new_n22555_, new_n22553_ );
nor  ( new_n22557_, new_n22555_, new_n22553_ );
or   ( new_n22558_, new_n897_, new_n21674_ );
or   ( new_n22559_, new_n899_, new_n21701_ );
and  ( new_n22560_, new_n22559_, new_n22558_ );
xor  ( new_n22561_, new_n22560_, new_n748_ );
or   ( new_n22562_, new_n22561_, new_n22557_ );
and  ( new_n22563_, new_n22562_, new_n22556_ );
or   ( new_n22564_, new_n22563_, new_n22549_ );
and  ( new_n22565_, new_n22563_, new_n22549_ );
or   ( new_n22566_, new_n755_, new_n21680_ );
or   ( new_n22567_, new_n757_, new_n21672_ );
and  ( new_n22568_, new_n22567_, new_n22566_ );
xor  ( new_n22569_, new_n22568_, new_n523_ );
or   ( new_n22570_, new_n524_, new_n21687_ );
or   ( new_n22571_, new_n526_, new_n21678_ );
and  ( new_n22572_, new_n22571_, new_n22570_ );
xor  ( new_n22573_, new_n22572_, new_n403_ );
nor  ( new_n22574_, new_n22573_, new_n22569_ );
and  ( new_n22575_, new_n22573_, new_n22569_ );
or   ( new_n22576_, new_n409_, new_n21751_ );
or   ( new_n22577_, new_n411_, new_n21685_ );
and  ( new_n22578_, new_n22577_, new_n22576_ );
xor  ( new_n22579_, new_n22578_, new_n328_ );
nor  ( new_n22580_, new_n22579_, new_n22575_ );
nor  ( new_n22581_, new_n22580_, new_n22574_ );
or   ( new_n22582_, new_n22581_, new_n22565_ );
and  ( new_n22583_, new_n22582_, new_n22564_ );
nor  ( new_n22584_, new_n22583_, new_n22533_ );
and  ( new_n22585_, new_n22583_, new_n22533_ );
or   ( new_n22586_, new_n299_, new_n22304_ );
or   ( new_n22587_, new_n302_, new_n22207_ );
and  ( new_n22588_, new_n22587_, new_n22586_ );
xor  ( new_n22589_, new_n22588_, new_n293_ );
not  ( new_n22590_, RIbb31f50_149 );
or   ( new_n22591_, new_n268_, new_n22590_ );
or   ( new_n22592_, new_n271_, new_n22423_ );
and  ( new_n22593_, new_n22592_, new_n22591_ );
xor  ( new_n22594_, new_n22593_, new_n263_ );
nor  ( new_n22595_, new_n22594_, new_n22589_ );
and  ( new_n22596_, RIbb31fc8_150, RIbb2f610_1 );
not  ( new_n22597_, new_n22596_ );
nand ( new_n22598_, new_n22594_, new_n22589_ );
and  ( new_n22599_, new_n22598_, new_n22597_ );
or   ( new_n22600_, new_n22599_, new_n22595_ );
xnor ( new_n22601_, new_n22460_, new_n22456_ );
xor  ( new_n22602_, new_n22601_, new_n22466_ );
and  ( new_n22603_, new_n22602_, new_n22600_ );
nor  ( new_n22604_, new_n22602_, new_n22600_ );
not  ( new_n22605_, new_n22604_ );
xor  ( new_n22606_, new_n22427_, new_n22422_ );
xor  ( new_n22607_, new_n22606_, new_n22430_ );
and  ( new_n22608_, new_n22607_, new_n22605_ );
nor  ( new_n22609_, new_n22608_, new_n22603_ );
nor  ( new_n22610_, new_n22609_, new_n22585_ );
nor  ( new_n22611_, new_n22610_, new_n22584_ );
not  ( new_n22612_, new_n22611_ );
or   ( new_n22613_, new_n22612_, new_n22527_ );
and  ( new_n22614_, new_n22613_, new_n22526_ );
or   ( new_n22615_, new_n22614_, new_n22514_ );
and  ( new_n22616_, new_n22614_, new_n22514_ );
xor  ( new_n22617_, new_n22416_, new_n22406_ );
xor  ( new_n22618_, new_n22617_, new_n22497_ );
or   ( new_n22619_, new_n22618_, new_n22616_ );
and  ( new_n22620_, new_n22619_, new_n22615_ );
nor  ( new_n22621_, new_n22620_, new_n22512_ );
xor  ( new_n22622_, new_n22507_, new_n22404_ );
and  ( new_n22623_, new_n22622_, new_n22621_ );
xor  ( new_n22624_, new_n22614_, new_n22514_ );
xor  ( new_n22625_, new_n22624_, new_n22618_ );
xor  ( new_n22626_, new_n22520_, new_n22518_ );
xor  ( new_n22627_, new_n22626_, new_n22523_ );
xor  ( new_n22628_, new_n22594_, new_n22589_ );
xor  ( new_n22629_, new_n22628_, new_n22597_ );
not  ( new_n22630_, new_n22629_ );
or   ( new_n22631_, new_n283_, new_n22207_ );
or   ( new_n22632_, new_n286_, new_n22129_ );
and  ( new_n22633_, new_n22632_, new_n22631_ );
xor  ( new_n22634_, new_n22633_, new_n278_ );
or   ( new_n22635_, new_n299_, new_n22423_ );
or   ( new_n22636_, new_n302_, new_n22304_ );
and  ( new_n22637_, new_n22636_, new_n22635_ );
xor  ( new_n22638_, new_n22637_, new_n293_ );
or   ( new_n22639_, new_n22638_, new_n22634_ );
and  ( new_n22640_, new_n22638_, new_n22634_ );
not  ( new_n22641_, RIbb31fc8_150 );
or   ( new_n22642_, new_n268_, new_n22641_ );
or   ( new_n22643_, new_n271_, new_n22590_ );
and  ( new_n22644_, new_n22643_, new_n22642_ );
xor  ( new_n22645_, new_n22644_, new_n263_ );
or   ( new_n22646_, new_n22645_, new_n22640_ );
and  ( new_n22647_, new_n22646_, new_n22639_ );
or   ( new_n22648_, new_n22647_, new_n22630_ );
or   ( new_n22649_, new_n1135_, new_n21701_ );
or   ( new_n22650_, new_n1137_, new_n21703_ );
and  ( new_n22651_, new_n22650_, new_n22649_ );
xor  ( new_n22652_, new_n22651_, new_n896_ );
and  ( new_n22653_, new_n22652_, new_n1358_ );
or   ( new_n22654_, new_n22652_, new_n1358_ );
or   ( new_n22655_, new_n1364_, new_n21694_ );
or   ( new_n22656_, new_n1366_, new_n21696_ );
and  ( new_n22657_, new_n22656_, new_n22655_ );
xor  ( new_n22658_, new_n22657_, new_n1129_ );
and  ( new_n22659_, new_n22658_, new_n22654_ );
or   ( new_n22660_, new_n22659_, new_n22653_ );
or   ( new_n22661_, new_n897_, new_n21672_ );
or   ( new_n22662_, new_n899_, new_n21674_ );
and  ( new_n22663_, new_n22662_, new_n22661_ );
xor  ( new_n22664_, new_n22663_, new_n748_ );
or   ( new_n22665_, new_n755_, new_n21678_ );
or   ( new_n22666_, new_n757_, new_n21680_ );
and  ( new_n22667_, new_n22666_, new_n22665_ );
xor  ( new_n22668_, new_n22667_, new_n523_ );
or   ( new_n22669_, new_n22668_, new_n22664_ );
and  ( new_n22670_, new_n22668_, new_n22664_ );
or   ( new_n22671_, new_n524_, new_n21685_ );
or   ( new_n22672_, new_n526_, new_n21687_ );
and  ( new_n22673_, new_n22672_, new_n22671_ );
xor  ( new_n22674_, new_n22673_, new_n403_ );
or   ( new_n22675_, new_n22674_, new_n22670_ );
and  ( new_n22676_, new_n22675_, new_n22669_ );
or   ( new_n22677_, new_n22676_, new_n22660_ );
and  ( new_n22678_, new_n22676_, new_n22660_ );
or   ( new_n22679_, new_n409_, new_n21792_ );
or   ( new_n22680_, new_n411_, new_n21751_ );
and  ( new_n22681_, new_n22680_, new_n22679_ );
xor  ( new_n22682_, new_n22681_, new_n328_ );
or   ( new_n22683_, new_n337_, new_n21840_ );
or   ( new_n22684_, new_n340_, new_n21842_ );
and  ( new_n22685_, new_n22684_, new_n22683_ );
xor  ( new_n22686_, new_n22685_, new_n332_ );
or   ( new_n22687_, new_n22686_, new_n22682_ );
and  ( new_n22688_, new_n22686_, new_n22682_ );
or   ( new_n22689_, new_n317_, new_n22098_ );
or   ( new_n22690_, new_n320_, new_n21847_ );
and  ( new_n22691_, new_n22690_, new_n22689_ );
xor  ( new_n22692_, new_n22691_, new_n312_ );
or   ( new_n22693_, new_n22692_, new_n22688_ );
and  ( new_n22694_, new_n22693_, new_n22687_ );
or   ( new_n22695_, new_n22694_, new_n22678_ );
and  ( new_n22696_, new_n22695_, new_n22677_ );
nand ( new_n22697_, new_n22696_, new_n22648_ );
nor  ( new_n22698_, new_n22696_, new_n22648_ );
xnor ( new_n22699_, new_n22555_, new_n22553_ );
xor  ( new_n22700_, new_n22699_, new_n22561_ );
xnor ( new_n22701_, new_n22541_, new_n22537_ );
xor  ( new_n22702_, new_n22701_, new_n22547_ );
nor  ( new_n22703_, new_n22702_, new_n22700_ );
and  ( new_n22704_, new_n22702_, new_n22700_ );
xor  ( new_n22705_, new_n22573_, new_n22569_ );
xnor ( new_n22706_, new_n22705_, new_n22579_ );
nor  ( new_n22707_, new_n22706_, new_n22704_ );
nor  ( new_n22708_, new_n22707_, new_n22703_ );
or   ( new_n22709_, new_n22708_, new_n22698_ );
and  ( new_n22710_, new_n22709_, new_n22697_ );
and  ( new_n22711_, new_n22710_, new_n22627_ );
xor  ( new_n22712_, new_n22602_, new_n22600_ );
xor  ( new_n22713_, new_n22712_, new_n22607_ );
xnor ( new_n22714_, new_n22563_, new_n22549_ );
xor  ( new_n22715_, new_n22714_, new_n22581_ );
nor  ( new_n22716_, new_n22715_, new_n22713_ );
and  ( new_n22717_, new_n22715_, new_n22713_ );
xor  ( new_n22718_, new_n22532_, new_n22530_ );
not  ( new_n22719_, new_n22718_ );
nor  ( new_n22720_, new_n22719_, new_n22717_ );
nor  ( new_n22721_, new_n22720_, new_n22716_ );
nor  ( new_n22722_, new_n22721_, new_n22711_ );
nor  ( new_n22723_, new_n22710_, new_n22627_ );
or   ( new_n22724_, new_n22723_, new_n22722_ );
xor  ( new_n22725_, new_n22488_, new_n22440_ );
xor  ( new_n22726_, new_n22725_, new_n22495_ );
nand ( new_n22727_, new_n22726_, new_n22724_ );
nor  ( new_n22728_, new_n22726_, new_n22724_ );
xor  ( new_n22729_, new_n22525_, new_n22516_ );
xor  ( new_n22730_, new_n22729_, new_n22612_ );
or   ( new_n22731_, new_n22730_, new_n22728_ );
and  ( new_n22732_, new_n22731_, new_n22727_ );
nor  ( new_n22733_, new_n22732_, new_n22625_ );
xor  ( new_n22734_, new_n22620_, new_n22512_ );
and  ( new_n22735_, new_n22734_, new_n22733_ );
xor  ( new_n22736_, new_n22710_, new_n22627_ );
xor  ( new_n22737_, new_n22736_, new_n22721_ );
xnor ( new_n22738_, new_n22583_, new_n22533_ );
xor  ( new_n22739_, new_n22738_, new_n22609_ );
nor  ( new_n22740_, new_n22739_, new_n22737_ );
nand ( new_n22741_, new_n22739_, new_n22737_ );
xor  ( new_n22742_, new_n22715_, new_n22713_ );
xor  ( new_n22743_, new_n22742_, new_n22719_ );
xor  ( new_n22744_, new_n22676_, new_n22660_ );
xor  ( new_n22745_, new_n22744_, new_n22694_ );
xnor ( new_n22746_, new_n22702_, new_n22700_ );
xor  ( new_n22747_, new_n22746_, new_n22706_ );
nand ( new_n22748_, new_n22747_, new_n22745_ );
nor  ( new_n22749_, new_n22747_, new_n22745_ );
xor  ( new_n22750_, new_n22647_, new_n22630_ );
or   ( new_n22751_, new_n22750_, new_n22749_ );
and  ( new_n22752_, new_n22751_, new_n22748_ );
nor  ( new_n22753_, new_n22752_, new_n22743_ );
nand ( new_n22754_, new_n22752_, new_n22743_ );
or   ( new_n22755_, new_n1364_, new_n21703_ );
or   ( new_n22756_, new_n1366_, new_n21694_ );
and  ( new_n22757_, new_n22756_, new_n22755_ );
xor  ( new_n22758_, new_n22757_, new_n1128_ );
and  ( new_n22759_, new_n1476_, RIbb315f0_129 );
xor  ( new_n22760_, new_n22759_, new_n1358_ );
nand ( new_n22761_, new_n22760_, new_n22758_ );
nor  ( new_n22762_, new_n22760_, new_n22758_ );
or   ( new_n22763_, new_n1135_, new_n21674_ );
or   ( new_n22764_, new_n1137_, new_n21701_ );
and  ( new_n22765_, new_n22764_, new_n22763_ );
xor  ( new_n22766_, new_n22765_, new_n896_ );
or   ( new_n22767_, new_n22766_, new_n22762_ );
and  ( new_n22768_, new_n22767_, new_n22761_ );
or   ( new_n22769_, new_n897_, new_n21680_ );
or   ( new_n22770_, new_n899_, new_n21672_ );
and  ( new_n22771_, new_n22770_, new_n22769_ );
xor  ( new_n22772_, new_n22771_, new_n748_ );
or   ( new_n22773_, new_n755_, new_n21687_ );
or   ( new_n22774_, new_n757_, new_n21678_ );
and  ( new_n22775_, new_n22774_, new_n22773_ );
xor  ( new_n22776_, new_n22775_, new_n523_ );
or   ( new_n22777_, new_n22776_, new_n22772_ );
and  ( new_n22778_, new_n22776_, new_n22772_ );
or   ( new_n22779_, new_n524_, new_n21751_ );
or   ( new_n22780_, new_n526_, new_n21685_ );
and  ( new_n22781_, new_n22780_, new_n22779_ );
xor  ( new_n22782_, new_n22781_, new_n403_ );
or   ( new_n22783_, new_n22782_, new_n22778_ );
and  ( new_n22784_, new_n22783_, new_n22777_ );
nor  ( new_n22785_, new_n22784_, new_n22768_ );
nand ( new_n22786_, new_n22784_, new_n22768_ );
or   ( new_n22787_, new_n409_, new_n21842_ );
or   ( new_n22788_, new_n411_, new_n21792_ );
and  ( new_n22789_, new_n22788_, new_n22787_ );
xor  ( new_n22790_, new_n22789_, new_n328_ );
or   ( new_n22791_, new_n337_, new_n21847_ );
or   ( new_n22792_, new_n340_, new_n21840_ );
and  ( new_n22793_, new_n22792_, new_n22791_ );
xor  ( new_n22794_, new_n22793_, new_n332_ );
nor  ( new_n22795_, new_n22794_, new_n22790_ );
and  ( new_n22796_, new_n22794_, new_n22790_ );
or   ( new_n22797_, new_n317_, new_n22129_ );
or   ( new_n22798_, new_n320_, new_n22098_ );
and  ( new_n22799_, new_n22798_, new_n22797_ );
xor  ( new_n22800_, new_n22799_, new_n312_ );
nor  ( new_n22801_, new_n22800_, new_n22796_ );
nor  ( new_n22802_, new_n22801_, new_n22795_ );
not  ( new_n22803_, new_n22802_ );
and  ( new_n22804_, new_n22803_, new_n22786_ );
or   ( new_n22805_, new_n22804_, new_n22785_ );
xnor ( new_n22806_, new_n22668_, new_n22664_ );
xor  ( new_n22807_, new_n22806_, new_n22674_ );
xnor ( new_n22808_, new_n22638_, new_n22634_ );
xor  ( new_n22809_, new_n22808_, new_n22645_ );
or   ( new_n22810_, new_n22809_, new_n22807_ );
and  ( new_n22811_, new_n22809_, new_n22807_ );
xor  ( new_n22812_, new_n22686_, new_n22682_ );
xnor ( new_n22813_, new_n22812_, new_n22692_ );
or   ( new_n22814_, new_n22813_, new_n22811_ );
and  ( new_n22815_, new_n22814_, new_n22810_ );
nor  ( new_n22816_, new_n22815_, new_n22805_ );
nand ( new_n22817_, new_n22815_, new_n22805_ );
and  ( new_n22818_, RIbb320b8_152, RIbb2f610_1 );
or   ( new_n22819_, new_n283_, new_n22304_ );
or   ( new_n22820_, new_n286_, new_n22207_ );
and  ( new_n22821_, new_n22820_, new_n22819_ );
xor  ( new_n22822_, new_n22821_, new_n278_ );
or   ( new_n22823_, new_n299_, new_n22590_ );
or   ( new_n22824_, new_n302_, new_n22423_ );
and  ( new_n22825_, new_n22824_, new_n22823_ );
xor  ( new_n22826_, new_n22825_, new_n293_ );
or   ( new_n22827_, new_n22826_, new_n22822_ );
and  ( new_n22828_, new_n22826_, new_n22822_ );
not  ( new_n22829_, RIbb32040_151 );
or   ( new_n22830_, new_n268_, new_n22829_ );
or   ( new_n22831_, new_n271_, new_n22641_ );
and  ( new_n22832_, new_n22831_, new_n22830_ );
xor  ( new_n22833_, new_n22832_, new_n263_ );
or   ( new_n22834_, new_n22833_, new_n22828_ );
and  ( new_n22835_, new_n22834_, new_n22827_ );
nor  ( new_n22836_, new_n22835_, new_n22818_ );
and  ( new_n22837_, new_n22835_, new_n22818_ );
and  ( new_n22838_, RIbb32040_151, RIbb2f610_1 );
nor  ( new_n22839_, new_n22838_, new_n22837_ );
nor  ( new_n22840_, new_n22839_, new_n22836_ );
and  ( new_n22841_, new_n22840_, new_n22817_ );
or   ( new_n22842_, new_n22841_, new_n22816_ );
and  ( new_n22843_, new_n22842_, new_n22754_ );
or   ( new_n22844_, new_n22843_, new_n22753_ );
and  ( new_n22845_, new_n22844_, new_n22741_ );
or   ( new_n22846_, new_n22845_, new_n22740_ );
xnor ( new_n22847_, new_n22726_, new_n22724_ );
xor  ( new_n22848_, new_n22847_, new_n22730_ );
and  ( new_n22849_, new_n22848_, new_n22846_ );
xor  ( new_n22850_, new_n22732_, new_n22625_ );
and  ( new_n22851_, new_n22850_, new_n22849_ );
xor  ( new_n22852_, new_n22752_, new_n22743_ );
xor  ( new_n22853_, new_n22852_, new_n22842_ );
xnor ( new_n22854_, new_n22747_, new_n22745_ );
xor  ( new_n22855_, new_n22854_, new_n22750_ );
or   ( new_n22856_, new_n1364_, new_n21701_ );
or   ( new_n22857_, new_n1366_, new_n21703_ );
and  ( new_n22858_, new_n22857_, new_n22856_ );
xor  ( new_n22859_, new_n22858_, new_n1129_ );
and  ( new_n22860_, new_n22859_, new_n1586_ );
or   ( new_n22861_, new_n22859_, new_n1586_ );
or   ( new_n22862_, new_n1593_, new_n21694_ );
or   ( new_n22863_, new_n1595_, new_n21696_ );
and  ( new_n22864_, new_n22863_, new_n22862_ );
xor  ( new_n22865_, new_n22864_, new_n1358_ );
and  ( new_n22866_, new_n22865_, new_n22861_ );
or   ( new_n22867_, new_n22866_, new_n22860_ );
or   ( new_n22868_, new_n524_, new_n21792_ );
or   ( new_n22869_, new_n526_, new_n21751_ );
and  ( new_n22870_, new_n22869_, new_n22868_ );
xor  ( new_n22871_, new_n22870_, new_n403_ );
or   ( new_n22872_, new_n409_, new_n21840_ );
or   ( new_n22873_, new_n411_, new_n21842_ );
and  ( new_n22874_, new_n22873_, new_n22872_ );
xor  ( new_n22875_, new_n22874_, new_n328_ );
or   ( new_n22876_, new_n22875_, new_n22871_ );
and  ( new_n22877_, new_n22875_, new_n22871_ );
or   ( new_n22878_, new_n337_, new_n22098_ );
or   ( new_n22879_, new_n340_, new_n21847_ );
and  ( new_n22880_, new_n22879_, new_n22878_ );
xor  ( new_n22881_, new_n22880_, new_n332_ );
or   ( new_n22882_, new_n22881_, new_n22877_ );
and  ( new_n22883_, new_n22882_, new_n22876_ );
nor  ( new_n22884_, new_n22883_, new_n22867_ );
nand ( new_n22885_, new_n22883_, new_n22867_ );
or   ( new_n22886_, new_n1135_, new_n21672_ );
or   ( new_n22887_, new_n1137_, new_n21674_ );
and  ( new_n22888_, new_n22887_, new_n22886_ );
xor  ( new_n22889_, new_n22888_, new_n896_ );
or   ( new_n22890_, new_n897_, new_n21678_ );
or   ( new_n22891_, new_n899_, new_n21680_ );
and  ( new_n22892_, new_n22891_, new_n22890_ );
xor  ( new_n22893_, new_n22892_, new_n748_ );
nor  ( new_n22894_, new_n22893_, new_n22889_ );
and  ( new_n22895_, new_n22893_, new_n22889_ );
or   ( new_n22896_, new_n755_, new_n21685_ );
or   ( new_n22897_, new_n757_, new_n21687_ );
and  ( new_n22898_, new_n22897_, new_n22896_ );
xor  ( new_n22899_, new_n22898_, new_n523_ );
nor  ( new_n22900_, new_n22899_, new_n22895_ );
or   ( new_n22901_, new_n22900_, new_n22894_ );
and  ( new_n22902_, new_n22901_, new_n22885_ );
or   ( new_n22903_, new_n22902_, new_n22884_ );
xnor ( new_n22904_, new_n22776_, new_n22772_ );
xor  ( new_n22905_, new_n22904_, new_n22782_ );
xnor ( new_n22906_, new_n22760_, new_n22758_ );
xor  ( new_n22907_, new_n22906_, new_n22766_ );
or   ( new_n22908_, new_n22907_, new_n22905_ );
and  ( new_n22909_, new_n22907_, new_n22905_ );
xnor ( new_n22910_, new_n22794_, new_n22790_ );
xor  ( new_n22911_, new_n22910_, new_n22800_ );
or   ( new_n22912_, new_n22911_, new_n22909_ );
and  ( new_n22913_, new_n22912_, new_n22908_ );
nand ( new_n22914_, new_n22913_, new_n22903_ );
nor  ( new_n22915_, new_n22913_, new_n22903_ );
not  ( new_n22916_, new_n22818_ );
or   ( new_n22917_, new_n317_, new_n22207_ );
or   ( new_n22918_, new_n320_, new_n22129_ );
and  ( new_n22919_, new_n22918_, new_n22917_ );
xor  ( new_n22920_, new_n22919_, new_n312_ );
or   ( new_n22921_, new_n283_, new_n22423_ );
or   ( new_n22922_, new_n286_, new_n22304_ );
and  ( new_n22923_, new_n22922_, new_n22921_ );
xor  ( new_n22924_, new_n22923_, new_n278_ );
or   ( new_n22925_, new_n22924_, new_n22920_ );
and  ( new_n22926_, new_n22924_, new_n22920_ );
or   ( new_n22927_, new_n299_, new_n22641_ );
or   ( new_n22928_, new_n302_, new_n22590_ );
and  ( new_n22929_, new_n22928_, new_n22927_ );
xor  ( new_n22930_, new_n22929_, new_n293_ );
or   ( new_n22931_, new_n22930_, new_n22926_ );
and  ( new_n22932_, new_n22931_, new_n22925_ );
nor  ( new_n22933_, new_n22932_, new_n22916_ );
and  ( new_n22934_, new_n22932_, new_n22916_ );
xor  ( new_n22935_, new_n22826_, new_n22822_ );
xnor ( new_n22936_, new_n22935_, new_n22833_ );
not  ( new_n22937_, new_n22936_ );
nor  ( new_n22938_, new_n22937_, new_n22934_ );
nor  ( new_n22939_, new_n22938_, new_n22933_ );
or   ( new_n22940_, new_n22939_, new_n22915_ );
and  ( new_n22941_, new_n22940_, new_n22914_ );
or   ( new_n22942_, new_n22941_, new_n22855_ );
and  ( new_n22943_, new_n22941_, new_n22855_ );
xnor ( new_n22944_, new_n22809_, new_n22807_ );
xor  ( new_n22945_, new_n22944_, new_n22813_ );
xor  ( new_n22946_, new_n22652_, new_n1358_ );
xor  ( new_n22947_, new_n22946_, new_n22658_ );
nor  ( new_n22948_, new_n22947_, new_n22945_ );
and  ( new_n22949_, new_n22947_, new_n22945_ );
not  ( new_n22950_, new_n22949_ );
xor  ( new_n22951_, new_n22835_, new_n22818_ );
xnor ( new_n22952_, new_n22951_, new_n22838_ );
and  ( new_n22953_, new_n22952_, new_n22950_ );
nor  ( new_n22954_, new_n22953_, new_n22948_ );
or   ( new_n22955_, new_n22954_, new_n22943_ );
and  ( new_n22956_, new_n22955_, new_n22942_ );
or   ( new_n22957_, new_n22956_, new_n22853_ );
and  ( new_n22958_, new_n22956_, new_n22853_ );
xor  ( new_n22959_, new_n22696_, new_n22648_ );
xnor ( new_n22960_, new_n22959_, new_n22708_ );
or   ( new_n22961_, new_n22960_, new_n22958_ );
and  ( new_n22962_, new_n22961_, new_n22957_ );
xor  ( new_n22963_, new_n22739_, new_n22737_ );
xor  ( new_n22964_, new_n22963_, new_n22844_ );
and  ( new_n22965_, new_n22964_, new_n22962_ );
xor  ( new_n22966_, new_n22848_, new_n22846_ );
and  ( new_n22967_, new_n22966_, new_n22965_ );
xor  ( new_n22968_, new_n22913_, new_n22903_ );
xnor ( new_n22969_, new_n22968_, new_n22939_ );
xor  ( new_n22970_, new_n22947_, new_n22945_ );
xor  ( new_n22971_, new_n22970_, new_n22952_ );
or   ( new_n22972_, new_n22971_, new_n22969_ );
not  ( new_n22973_, RIbb32130_153 );
or   ( new_n22974_, new_n268_, new_n22973_ );
not  ( new_n22975_, RIbb320b8_152 );
or   ( new_n22976_, new_n271_, new_n22975_ );
and  ( new_n22977_, new_n22976_, new_n22974_ );
xor  ( new_n22978_, new_n22977_, new_n263_ );
and  ( new_n22979_, RIbb321a8_154, RIbb2f610_1 );
or   ( new_n22980_, new_n22979_, new_n22978_ );
or   ( new_n22981_, new_n317_, new_n22304_ );
or   ( new_n22982_, new_n320_, new_n22207_ );
and  ( new_n22983_, new_n22982_, new_n22981_ );
xor  ( new_n22984_, new_n22983_, new_n312_ );
or   ( new_n22985_, new_n283_, new_n22590_ );
or   ( new_n22986_, new_n286_, new_n22423_ );
and  ( new_n22987_, new_n22986_, new_n22985_ );
xor  ( new_n22988_, new_n22987_, new_n278_ );
or   ( new_n22989_, new_n22988_, new_n22984_ );
and  ( new_n22990_, new_n22988_, new_n22984_ );
or   ( new_n22991_, new_n299_, new_n22829_ );
or   ( new_n22992_, new_n302_, new_n22641_ );
and  ( new_n22993_, new_n22992_, new_n22991_ );
xor  ( new_n22994_, new_n22993_, new_n293_ );
or   ( new_n22995_, new_n22994_, new_n22990_ );
and  ( new_n22996_, new_n22995_, new_n22989_ );
and  ( new_n22997_, new_n22996_, new_n22980_ );
or   ( new_n22998_, new_n22996_, new_n22980_ );
or   ( new_n22999_, new_n268_, new_n22975_ );
or   ( new_n23000_, new_n271_, new_n22829_ );
and  ( new_n23001_, new_n23000_, new_n22999_ );
xor  ( new_n23002_, new_n23001_, new_n263_ );
and  ( new_n23003_, new_n23002_, new_n22998_ );
or   ( new_n23004_, new_n23003_, new_n22997_ );
or   ( new_n23005_, new_n22973_, new_n260_ );
xnor ( new_n23006_, new_n22875_, new_n22871_ );
xor  ( new_n23007_, new_n23006_, new_n22881_ );
nand ( new_n23008_, new_n23007_, new_n23005_ );
nor  ( new_n23009_, new_n23007_, new_n23005_ );
xor  ( new_n23010_, new_n22924_, new_n22920_ );
xor  ( new_n23011_, new_n23010_, new_n22930_ );
or   ( new_n23012_, new_n23011_, new_n23009_ );
and  ( new_n23013_, new_n23012_, new_n23008_ );
nor  ( new_n23014_, new_n23013_, new_n23004_ );
nand ( new_n23015_, new_n23013_, new_n23004_ );
or   ( new_n23016_, new_n1135_, new_n21680_ );
or   ( new_n23017_, new_n1137_, new_n21672_ );
and  ( new_n23018_, new_n23017_, new_n23016_ );
xor  ( new_n23019_, new_n23018_, new_n896_ );
or   ( new_n23020_, new_n897_, new_n21687_ );
or   ( new_n23021_, new_n899_, new_n21678_ );
and  ( new_n23022_, new_n23021_, new_n23020_ );
xor  ( new_n23023_, new_n23022_, new_n748_ );
or   ( new_n23024_, new_n23023_, new_n23019_ );
and  ( new_n23025_, new_n23023_, new_n23019_ );
or   ( new_n23026_, new_n755_, new_n21751_ );
or   ( new_n23027_, new_n757_, new_n21685_ );
and  ( new_n23028_, new_n23027_, new_n23026_ );
xor  ( new_n23029_, new_n23028_, new_n523_ );
or   ( new_n23030_, new_n23029_, new_n23025_ );
and  ( new_n23031_, new_n23030_, new_n23024_ );
or   ( new_n23032_, new_n524_, new_n21842_ );
or   ( new_n23033_, new_n526_, new_n21792_ );
and  ( new_n23034_, new_n23033_, new_n23032_ );
xor  ( new_n23035_, new_n23034_, new_n403_ );
or   ( new_n23036_, new_n409_, new_n21847_ );
or   ( new_n23037_, new_n411_, new_n21840_ );
and  ( new_n23038_, new_n23037_, new_n23036_ );
xor  ( new_n23039_, new_n23038_, new_n328_ );
or   ( new_n23040_, new_n23039_, new_n23035_ );
and  ( new_n23041_, new_n23039_, new_n23035_ );
or   ( new_n23042_, new_n337_, new_n22129_ );
or   ( new_n23043_, new_n340_, new_n22098_ );
and  ( new_n23044_, new_n23043_, new_n23042_ );
xor  ( new_n23045_, new_n23044_, new_n332_ );
or   ( new_n23046_, new_n23045_, new_n23041_ );
and  ( new_n23047_, new_n23046_, new_n23040_ );
nor  ( new_n23048_, new_n23047_, new_n23031_ );
and  ( new_n23049_, new_n23047_, new_n23031_ );
or   ( new_n23050_, new_n1593_, new_n21703_ );
or   ( new_n23051_, new_n1595_, new_n21694_ );
and  ( new_n23052_, new_n23051_, new_n23050_ );
xor  ( new_n23053_, new_n23052_, new_n1357_ );
and  ( new_n23054_, new_n1741_, RIbb315f0_129 );
xor  ( new_n23055_, new_n23054_, new_n1586_ );
and  ( new_n23056_, new_n23055_, new_n23053_ );
nor  ( new_n23057_, new_n23055_, new_n23053_ );
or   ( new_n23058_, new_n1364_, new_n21674_ );
or   ( new_n23059_, new_n1366_, new_n21701_ );
and  ( new_n23060_, new_n23059_, new_n23058_ );
xor  ( new_n23061_, new_n23060_, new_n1129_ );
nor  ( new_n23062_, new_n23061_, new_n23057_ );
nor  ( new_n23063_, new_n23062_, new_n23056_ );
nor  ( new_n23064_, new_n23063_, new_n23049_ );
or   ( new_n23065_, new_n23064_, new_n23048_ );
and  ( new_n23066_, new_n23065_, new_n23015_ );
or   ( new_n23067_, new_n23066_, new_n23014_ );
xor  ( new_n23068_, new_n22907_, new_n22905_ );
xor  ( new_n23069_, new_n23068_, new_n22911_ );
xor  ( new_n23070_, new_n22883_, new_n22867_ );
xor  ( new_n23071_, new_n23070_, new_n22901_ );
or   ( new_n23072_, new_n23071_, new_n23069_ );
and  ( new_n23073_, new_n23071_, new_n23069_ );
xor  ( new_n23074_, new_n22932_, new_n22916_ );
xor  ( new_n23075_, new_n23074_, new_n22936_ );
or   ( new_n23076_, new_n23075_, new_n23073_ );
and  ( new_n23077_, new_n23076_, new_n23072_ );
or   ( new_n23078_, new_n23077_, new_n23067_ );
and  ( new_n23079_, new_n23077_, new_n23067_ );
xor  ( new_n23080_, new_n22784_, new_n22768_ );
xor  ( new_n23081_, new_n23080_, new_n22803_ );
or   ( new_n23082_, new_n23081_, new_n23079_ );
and  ( new_n23083_, new_n23082_, new_n23078_ );
nor  ( new_n23084_, new_n23083_, new_n22972_ );
and  ( new_n23085_, new_n23083_, new_n22972_ );
xor  ( new_n23086_, new_n22815_, new_n22805_ );
xor  ( new_n23087_, new_n23086_, new_n22840_ );
not  ( new_n23088_, new_n23087_ );
nor  ( new_n23089_, new_n23088_, new_n23085_ );
nor  ( new_n23090_, new_n23089_, new_n23084_ );
xnor ( new_n23091_, new_n22956_, new_n22853_ );
xor  ( new_n23092_, new_n23091_, new_n22960_ );
nor  ( new_n23093_, new_n23092_, new_n23090_ );
xor  ( new_n23094_, new_n22964_, new_n22962_ );
and  ( new_n23095_, new_n23094_, new_n23093_ );
xnor ( new_n23096_, new_n23092_, new_n23090_ );
xor  ( new_n23097_, new_n23083_, new_n22972_ );
xor  ( new_n23098_, new_n23097_, new_n23088_ );
xor  ( new_n23099_, new_n23007_, new_n23005_ );
xor  ( new_n23100_, new_n23099_, new_n23011_ );
xor  ( new_n23101_, new_n22859_, new_n1586_ );
xor  ( new_n23102_, new_n23101_, new_n22865_ );
and  ( new_n23103_, new_n23102_, new_n23100_ );
or   ( new_n23104_, new_n23102_, new_n23100_ );
xor  ( new_n23105_, new_n22893_, new_n22889_ );
xor  ( new_n23106_, new_n23105_, new_n22899_ );
and  ( new_n23107_, new_n23106_, new_n23104_ );
or   ( new_n23108_, new_n23107_, new_n23103_ );
xnor ( new_n23109_, new_n23071_, new_n23069_ );
xor  ( new_n23110_, new_n23109_, new_n23075_ );
and  ( new_n23111_, new_n23110_, new_n23108_ );
or   ( new_n23112_, new_n23110_, new_n23108_ );
or   ( new_n23113_, new_n1844_, new_n21694_ );
or   ( new_n23114_, new_n1846_, new_n21696_ );
and  ( new_n23115_, new_n23114_, new_n23113_ );
xor  ( new_n23116_, new_n23115_, new_n1586_ );
and  ( new_n23117_, new_n23116_, new_n1843_ );
or   ( new_n23118_, new_n23116_, new_n1843_ );
or   ( new_n23119_, new_n1593_, new_n21701_ );
or   ( new_n23120_, new_n1595_, new_n21703_ );
and  ( new_n23121_, new_n23120_, new_n23119_ );
xor  ( new_n23122_, new_n23121_, new_n1358_ );
and  ( new_n23123_, new_n23122_, new_n23118_ );
or   ( new_n23124_, new_n23123_, new_n23117_ );
or   ( new_n23125_, new_n1364_, new_n21672_ );
or   ( new_n23126_, new_n1366_, new_n21674_ );
and  ( new_n23127_, new_n23126_, new_n23125_ );
xor  ( new_n23128_, new_n23127_, new_n1129_ );
or   ( new_n23129_, new_n1135_, new_n21678_ );
or   ( new_n23130_, new_n1137_, new_n21680_ );
and  ( new_n23131_, new_n23130_, new_n23129_ );
xor  ( new_n23132_, new_n23131_, new_n896_ );
or   ( new_n23133_, new_n23132_, new_n23128_ );
and  ( new_n23134_, new_n23132_, new_n23128_ );
or   ( new_n23135_, new_n897_, new_n21685_ );
or   ( new_n23136_, new_n899_, new_n21687_ );
and  ( new_n23137_, new_n23136_, new_n23135_ );
xor  ( new_n23138_, new_n23137_, new_n748_ );
or   ( new_n23139_, new_n23138_, new_n23134_ );
and  ( new_n23140_, new_n23139_, new_n23133_ );
or   ( new_n23141_, new_n23140_, new_n23124_ );
and  ( new_n23142_, new_n23140_, new_n23124_ );
or   ( new_n23143_, new_n755_, new_n21792_ );
or   ( new_n23144_, new_n757_, new_n21751_ );
and  ( new_n23145_, new_n23144_, new_n23143_ );
xor  ( new_n23146_, new_n23145_, new_n523_ );
or   ( new_n23147_, new_n524_, new_n21840_ );
or   ( new_n23148_, new_n526_, new_n21842_ );
and  ( new_n23149_, new_n23148_, new_n23147_ );
xor  ( new_n23150_, new_n23149_, new_n403_ );
nor  ( new_n23151_, new_n23150_, new_n23146_ );
and  ( new_n23152_, new_n23150_, new_n23146_ );
or   ( new_n23153_, new_n409_, new_n22098_ );
or   ( new_n23154_, new_n411_, new_n21847_ );
and  ( new_n23155_, new_n23154_, new_n23153_ );
xor  ( new_n23156_, new_n23155_, new_n328_ );
nor  ( new_n23157_, new_n23156_, new_n23152_ );
nor  ( new_n23158_, new_n23157_, new_n23151_ );
or   ( new_n23159_, new_n23158_, new_n23142_ );
and  ( new_n23160_, new_n23159_, new_n23141_ );
xnor ( new_n23161_, new_n22979_, new_n22978_ );
or   ( new_n23162_, new_n299_, new_n22975_ );
or   ( new_n23163_, new_n302_, new_n22829_ );
and  ( new_n23164_, new_n23163_, new_n23162_ );
xor  ( new_n23165_, new_n23164_, new_n293_ );
not  ( new_n23166_, RIbb321a8_154 );
or   ( new_n23167_, new_n268_, new_n23166_ );
or   ( new_n23168_, new_n271_, new_n22973_ );
and  ( new_n23169_, new_n23168_, new_n23167_ );
xor  ( new_n23170_, new_n23169_, new_n263_ );
or   ( new_n23171_, new_n23170_, new_n23165_ );
and  ( new_n23172_, RIbb32220_155, RIbb2f610_1 );
and  ( new_n23173_, new_n23170_, new_n23165_ );
or   ( new_n23174_, new_n23173_, new_n23172_ );
and  ( new_n23175_, new_n23174_, new_n23171_ );
or   ( new_n23176_, new_n23175_, new_n23161_ );
and  ( new_n23177_, new_n23175_, new_n23161_ );
or   ( new_n23178_, new_n337_, new_n22207_ );
or   ( new_n23179_, new_n340_, new_n22129_ );
and  ( new_n23180_, new_n23179_, new_n23178_ );
xor  ( new_n23181_, new_n23180_, new_n332_ );
or   ( new_n23182_, new_n317_, new_n22423_ );
or   ( new_n23183_, new_n320_, new_n22304_ );
and  ( new_n23184_, new_n23183_, new_n23182_ );
xor  ( new_n23185_, new_n23184_, new_n312_ );
or   ( new_n23186_, new_n23185_, new_n23181_ );
and  ( new_n23187_, new_n23185_, new_n23181_ );
or   ( new_n23188_, new_n283_, new_n22641_ );
or   ( new_n23189_, new_n286_, new_n22590_ );
and  ( new_n23190_, new_n23189_, new_n23188_ );
xor  ( new_n23191_, new_n23190_, new_n278_ );
or   ( new_n23192_, new_n23191_, new_n23187_ );
and  ( new_n23193_, new_n23192_, new_n23186_ );
or   ( new_n23194_, new_n23193_, new_n23177_ );
and  ( new_n23195_, new_n23194_, new_n23176_ );
and  ( new_n23196_, new_n23195_, new_n23160_ );
or   ( new_n23197_, new_n23195_, new_n23160_ );
xnor ( new_n23198_, new_n23039_, new_n23035_ );
xor  ( new_n23199_, new_n23198_, new_n23045_ );
xnor ( new_n23200_, new_n23023_, new_n23019_ );
xor  ( new_n23201_, new_n23200_, new_n23029_ );
nor  ( new_n23202_, new_n23201_, new_n23199_ );
nand ( new_n23203_, new_n23201_, new_n23199_ );
xor  ( new_n23204_, new_n22988_, new_n22984_ );
xor  ( new_n23205_, new_n23204_, new_n22994_ );
and  ( new_n23206_, new_n23205_, new_n23203_ );
or   ( new_n23207_, new_n23206_, new_n23202_ );
and  ( new_n23208_, new_n23207_, new_n23197_ );
or   ( new_n23209_, new_n23208_, new_n23196_ );
and  ( new_n23210_, new_n23209_, new_n23112_ );
or   ( new_n23211_, new_n23210_, new_n23111_ );
xnor ( new_n23212_, new_n23077_, new_n23067_ );
xor  ( new_n23213_, new_n23212_, new_n23081_ );
nand ( new_n23214_, new_n23213_, new_n23211_ );
or   ( new_n23215_, new_n23213_, new_n23211_ );
xor  ( new_n23216_, new_n22971_, new_n22969_ );
nand ( new_n23217_, new_n23216_, new_n23215_ );
and  ( new_n23218_, new_n23217_, new_n23214_ );
or   ( new_n23219_, new_n23218_, new_n23098_ );
and  ( new_n23220_, new_n23218_, new_n23098_ );
xnor ( new_n23221_, new_n22941_, new_n22855_ );
xor  ( new_n23222_, new_n23221_, new_n22954_ );
or   ( new_n23223_, new_n23222_, new_n23220_ );
and  ( new_n23224_, new_n23223_, new_n23219_ );
nor  ( new_n23225_, new_n23224_, new_n23096_ );
xor  ( new_n23226_, new_n23218_, new_n23098_ );
xor  ( new_n23227_, new_n23226_, new_n23222_ );
xor  ( new_n23228_, new_n23213_, new_n23211_ );
xor  ( new_n23229_, new_n23228_, new_n23216_ );
xor  ( new_n23230_, new_n23110_, new_n23108_ );
xor  ( new_n23231_, new_n23230_, new_n23209_ );
xor  ( new_n23232_, new_n23047_, new_n23031_ );
xor  ( new_n23233_, new_n23232_, new_n23063_ );
xor  ( new_n23234_, new_n23195_, new_n23160_ );
xor  ( new_n23235_, new_n23234_, new_n23207_ );
xor  ( new_n23236_, new_n23235_, new_n23233_ );
xor  ( new_n23237_, new_n23102_, new_n23100_ );
xor  ( new_n23238_, new_n23237_, new_n23106_ );
xor  ( new_n23239_, new_n23238_, new_n23236_ );
xor  ( new_n23240_, new_n23132_, new_n23128_ );
xnor ( new_n23241_, new_n23240_, new_n23138_ );
xnor ( new_n23242_, new_n23185_, new_n23181_ );
xor  ( new_n23243_, new_n23242_, new_n23191_ );
xnor ( new_n23244_, new_n23243_, new_n23241_ );
xnor ( new_n23245_, new_n23150_, new_n23146_ );
xor  ( new_n23246_, new_n23245_, new_n23156_ );
xor  ( new_n23247_, new_n23246_, new_n23244_ );
or   ( new_n23248_, new_n299_, new_n22973_ );
or   ( new_n23249_, new_n302_, new_n22975_ );
and  ( new_n23250_, new_n23249_, new_n23248_ );
xor  ( new_n23251_, new_n23250_, new_n293_ );
not  ( new_n23252_, RIbb32220_155 );
or   ( new_n23253_, new_n268_, new_n23252_ );
or   ( new_n23254_, new_n271_, new_n23166_ );
and  ( new_n23255_, new_n23254_, new_n23253_ );
xor  ( new_n23256_, new_n23255_, new_n263_ );
or   ( new_n23257_, new_n23256_, new_n23251_ );
and  ( new_n23258_, RIbb32298_156, RIbb2f610_1 );
and  ( new_n23259_, new_n23256_, new_n23251_ );
or   ( new_n23260_, new_n23259_, new_n23258_ );
and  ( new_n23261_, new_n23260_, new_n23257_ );
xor  ( new_n23262_, new_n23170_, new_n23165_ );
xor  ( new_n23263_, new_n23262_, new_n23172_ );
or   ( new_n23264_, new_n337_, new_n22304_ );
or   ( new_n23265_, new_n340_, new_n22207_ );
and  ( new_n23266_, new_n23265_, new_n23264_ );
xor  ( new_n23267_, new_n23266_, new_n332_ );
or   ( new_n23268_, new_n317_, new_n22590_ );
or   ( new_n23269_, new_n320_, new_n22423_ );
and  ( new_n23270_, new_n23269_, new_n23268_ );
xor  ( new_n23271_, new_n23270_, new_n312_ );
or   ( new_n23272_, new_n23271_, new_n23267_ );
and  ( new_n23273_, new_n23271_, new_n23267_ );
or   ( new_n23274_, new_n283_, new_n22829_ );
or   ( new_n23275_, new_n286_, new_n22641_ );
and  ( new_n23276_, new_n23275_, new_n23274_ );
xor  ( new_n23277_, new_n23276_, new_n278_ );
or   ( new_n23278_, new_n23277_, new_n23273_ );
and  ( new_n23279_, new_n23278_, new_n23272_ );
xor  ( new_n23280_, new_n23279_, new_n23263_ );
xor  ( new_n23281_, new_n23280_, new_n23261_ );
or   ( new_n23282_, new_n23281_, new_n23247_ );
and  ( new_n23283_, new_n23281_, new_n23247_ );
xor  ( new_n23284_, new_n23116_, new_n1843_ );
xor  ( new_n23285_, new_n23284_, new_n23122_ );
or   ( new_n23286_, new_n23285_, new_n23283_ );
and  ( new_n23287_, new_n23286_, new_n23282_ );
or   ( new_n23288_, new_n1593_, new_n21672_ );
or   ( new_n23289_, new_n1595_, new_n21674_ );
and  ( new_n23290_, new_n23289_, new_n23288_ );
xor  ( new_n23291_, new_n23290_, new_n1358_ );
or   ( new_n23292_, new_n1364_, new_n21678_ );
or   ( new_n23293_, new_n1366_, new_n21680_ );
and  ( new_n23294_, new_n23293_, new_n23292_ );
xor  ( new_n23295_, new_n23294_, new_n1129_ );
nor  ( new_n23296_, new_n23295_, new_n23291_ );
and  ( new_n23297_, new_n23295_, new_n23291_ );
or   ( new_n23298_, new_n1135_, new_n21685_ );
or   ( new_n23299_, new_n1137_, new_n21687_ );
and  ( new_n23300_, new_n23299_, new_n23298_ );
xor  ( new_n23301_, new_n23300_, new_n896_ );
nor  ( new_n23302_, new_n23301_, new_n23297_ );
or   ( new_n23303_, new_n23302_, new_n23296_ );
or   ( new_n23304_, new_n2122_, new_n21694_ );
or   ( new_n23305_, new_n2124_, new_n21696_ );
and  ( new_n23306_, new_n23305_, new_n23304_ );
xor  ( new_n23307_, new_n23306_, new_n1843_ );
nand ( new_n23308_, new_n23307_, new_n2121_ );
or   ( new_n23309_, new_n23307_, new_n2121_ );
or   ( new_n23310_, new_n1844_, new_n21701_ );
or   ( new_n23311_, new_n1846_, new_n21703_ );
and  ( new_n23312_, new_n23311_, new_n23310_ );
xor  ( new_n23313_, new_n23312_, new_n1586_ );
nand ( new_n23314_, new_n23313_, new_n23309_ );
and  ( new_n23315_, new_n23314_, new_n23308_ );
and  ( new_n23316_, new_n23315_, new_n23303_ );
nor  ( new_n23317_, new_n23315_, new_n23303_ );
or   ( new_n23318_, new_n897_, new_n21792_ );
or   ( new_n23319_, new_n899_, new_n21751_ );
and  ( new_n23320_, new_n23319_, new_n23318_ );
xor  ( new_n23321_, new_n23320_, new_n748_ );
or   ( new_n23322_, new_n755_, new_n21840_ );
or   ( new_n23323_, new_n757_, new_n21842_ );
and  ( new_n23324_, new_n23323_, new_n23322_ );
xor  ( new_n23325_, new_n23324_, new_n523_ );
nor  ( new_n23326_, new_n23325_, new_n23321_ );
and  ( new_n23327_, new_n23325_, new_n23321_ );
or   ( new_n23328_, new_n524_, new_n22098_ );
or   ( new_n23329_, new_n526_, new_n21847_ );
and  ( new_n23330_, new_n23329_, new_n23328_ );
xor  ( new_n23331_, new_n23330_, new_n403_ );
nor  ( new_n23332_, new_n23331_, new_n23327_ );
nor  ( new_n23333_, new_n23332_, new_n23326_ );
nor  ( new_n23334_, new_n23333_, new_n23317_ );
or   ( new_n23335_, new_n23334_, new_n23316_ );
xnor ( new_n23336_, new_n23271_, new_n23267_ );
xor  ( new_n23337_, new_n23336_, new_n23277_ );
xnor ( new_n23338_, new_n23256_, new_n23251_ );
xor  ( new_n23339_, new_n23338_, new_n23258_ );
or   ( new_n23340_, new_n23339_, new_n23337_ );
and  ( new_n23341_, new_n23339_, new_n23337_ );
or   ( new_n23342_, new_n409_, new_n22129_ );
or   ( new_n23343_, new_n411_, new_n22098_ );
and  ( new_n23344_, new_n23343_, new_n23342_ );
xor  ( new_n23345_, new_n23344_, new_n328_ );
or   ( new_n23346_, new_n755_, new_n21842_ );
or   ( new_n23347_, new_n757_, new_n21792_ );
and  ( new_n23348_, new_n23347_, new_n23346_ );
xor  ( new_n23349_, new_n23348_, new_n523_ );
or   ( new_n23350_, new_n524_, new_n21847_ );
or   ( new_n23351_, new_n526_, new_n21840_ );
and  ( new_n23352_, new_n23351_, new_n23350_ );
xor  ( new_n23353_, new_n23352_, new_n403_ );
xnor ( new_n23354_, new_n23353_, new_n23349_ );
xor  ( new_n23355_, new_n23354_, new_n23345_ );
or   ( new_n23356_, new_n23355_, new_n23341_ );
and  ( new_n23357_, new_n23356_, new_n23340_ );
nand ( new_n23358_, new_n23357_, new_n23335_ );
or   ( new_n23359_, new_n23357_, new_n23335_ );
or   ( new_n23360_, new_n283_, new_n22975_ );
or   ( new_n23361_, new_n286_, new_n22829_ );
and  ( new_n23362_, new_n23361_, new_n23360_ );
xor  ( new_n23363_, new_n23362_, new_n278_ );
or   ( new_n23364_, new_n299_, new_n23166_ );
or   ( new_n23365_, new_n302_, new_n22973_ );
and  ( new_n23366_, new_n23365_, new_n23364_ );
xor  ( new_n23367_, new_n23366_, new_n293_ );
nor  ( new_n23368_, new_n23367_, new_n23363_ );
and  ( new_n23369_, new_n23367_, new_n23363_ );
not  ( new_n23370_, RIbb32298_156 );
or   ( new_n23371_, new_n268_, new_n23370_ );
or   ( new_n23372_, new_n271_, new_n23252_ );
and  ( new_n23373_, new_n23372_, new_n23371_ );
xor  ( new_n23374_, new_n23373_, new_n263_ );
nor  ( new_n23375_, new_n23374_, new_n23369_ );
nor  ( new_n23376_, new_n23375_, new_n23368_ );
or   ( new_n23377_, new_n409_, new_n22207_ );
or   ( new_n23378_, new_n411_, new_n22129_ );
and  ( new_n23379_, new_n23378_, new_n23377_ );
xor  ( new_n23380_, new_n23379_, new_n328_ );
or   ( new_n23381_, new_n337_, new_n22423_ );
or   ( new_n23382_, new_n340_, new_n22304_ );
and  ( new_n23383_, new_n23382_, new_n23381_ );
xor  ( new_n23384_, new_n23383_, new_n332_ );
or   ( new_n23385_, new_n23384_, new_n23380_ );
and  ( new_n23386_, new_n23384_, new_n23380_ );
or   ( new_n23387_, new_n317_, new_n22641_ );
or   ( new_n23388_, new_n320_, new_n22590_ );
and  ( new_n23389_, new_n23388_, new_n23387_ );
xor  ( new_n23390_, new_n23389_, new_n312_ );
or   ( new_n23391_, new_n23390_, new_n23386_ );
and  ( new_n23392_, new_n23391_, new_n23385_ );
nor  ( new_n23393_, new_n23392_, new_n23376_ );
nand ( new_n23394_, new_n23393_, new_n23359_ );
and  ( new_n23395_, new_n23394_, new_n23358_ );
or   ( new_n23396_, new_n23395_, new_n23287_ );
nand ( new_n23397_, new_n23395_, new_n23287_ );
xor  ( new_n23398_, new_n23140_, new_n23124_ );
xnor ( new_n23399_, new_n23398_, new_n23158_ );
nand ( new_n23400_, new_n23399_, new_n23397_ );
and  ( new_n23401_, new_n23400_, new_n23396_ );
or   ( new_n23402_, new_n23401_, new_n23239_ );
and  ( new_n23403_, new_n23401_, new_n23239_ );
or   ( new_n23404_, new_n23279_, new_n23263_ );
and  ( new_n23405_, new_n23279_, new_n23263_ );
or   ( new_n23406_, new_n23405_, new_n23261_ );
and  ( new_n23407_, new_n23406_, new_n23404_ );
or   ( new_n23408_, new_n1844_, new_n21703_ );
or   ( new_n23409_, new_n1846_, new_n21694_ );
and  ( new_n23410_, new_n23409_, new_n23408_ );
xor  ( new_n23411_, new_n23410_, new_n1585_ );
and  ( new_n23412_, new_n2002_, RIbb315f0_129 );
xor  ( new_n23413_, new_n23412_, new_n1843_ );
nand ( new_n23414_, new_n23413_, new_n23411_ );
nor  ( new_n23415_, new_n23413_, new_n23411_ );
or   ( new_n23416_, new_n1593_, new_n21674_ );
or   ( new_n23417_, new_n1595_, new_n21701_ );
and  ( new_n23418_, new_n23417_, new_n23416_ );
xor  ( new_n23419_, new_n23418_, new_n1358_ );
or   ( new_n23420_, new_n23419_, new_n23415_ );
and  ( new_n23421_, new_n23420_, new_n23414_ );
nor  ( new_n23422_, new_n23353_, new_n23349_ );
and  ( new_n23423_, new_n23353_, new_n23349_ );
nor  ( new_n23424_, new_n23423_, new_n23345_ );
nor  ( new_n23425_, new_n23424_, new_n23422_ );
or   ( new_n23426_, new_n1364_, new_n21680_ );
or   ( new_n23427_, new_n1366_, new_n21672_ );
and  ( new_n23428_, new_n23427_, new_n23426_ );
xor  ( new_n23429_, new_n23428_, new_n1129_ );
or   ( new_n23430_, new_n1135_, new_n21687_ );
or   ( new_n23431_, new_n1137_, new_n21678_ );
and  ( new_n23432_, new_n23431_, new_n23430_ );
xor  ( new_n23433_, new_n23432_, new_n896_ );
or   ( new_n23434_, new_n23433_, new_n23429_ );
and  ( new_n23435_, new_n23433_, new_n23429_ );
or   ( new_n23436_, new_n897_, new_n21751_ );
or   ( new_n23437_, new_n899_, new_n21685_ );
and  ( new_n23438_, new_n23437_, new_n23436_ );
xor  ( new_n23439_, new_n23438_, new_n748_ );
or   ( new_n23440_, new_n23439_, new_n23435_ );
and  ( new_n23441_, new_n23440_, new_n23434_ );
and  ( new_n23442_, new_n23441_, new_n23425_ );
or   ( new_n23443_, new_n23442_, new_n23421_ );
or   ( new_n23444_, new_n23441_, new_n23425_ );
and  ( new_n23445_, new_n23444_, new_n23443_ );
nor  ( new_n23446_, new_n23445_, new_n23407_ );
and  ( new_n23447_, new_n23445_, new_n23407_ );
nor  ( new_n23448_, new_n23243_, new_n23241_ );
and  ( new_n23449_, new_n23243_, new_n23241_ );
nor  ( new_n23450_, new_n23246_, new_n23449_ );
nor  ( new_n23451_, new_n23450_, new_n23448_ );
not  ( new_n23452_, new_n23451_ );
nor  ( new_n23453_, new_n23452_, new_n23447_ );
nor  ( new_n23454_, new_n23453_, new_n23446_ );
xor  ( new_n23455_, new_n23055_, new_n23053_ );
xor  ( new_n23456_, new_n23455_, new_n23061_ );
xor  ( new_n23457_, new_n23201_, new_n23199_ );
xor  ( new_n23458_, new_n23457_, new_n23205_ );
and  ( new_n23459_, new_n23458_, new_n23456_ );
or   ( new_n23460_, new_n23458_, new_n23456_ );
xor  ( new_n23461_, new_n23175_, new_n23161_ );
xor  ( new_n23462_, new_n23461_, new_n23193_ );
and  ( new_n23463_, new_n23462_, new_n23460_ );
or   ( new_n23464_, new_n23463_, new_n23459_ );
xor  ( new_n23465_, new_n22996_, new_n22980_ );
xor  ( new_n23466_, new_n23465_, new_n23002_ );
xor  ( new_n23467_, new_n23466_, new_n23464_ );
xor  ( new_n23468_, new_n23467_, new_n23454_ );
or   ( new_n23469_, new_n23468_, new_n23403_ );
and  ( new_n23470_, new_n23469_, new_n23402_ );
or   ( new_n23471_, new_n23470_, new_n23231_ );
nand ( new_n23472_, new_n23470_, new_n23231_ );
and  ( new_n23473_, new_n23235_, new_n23233_ );
or   ( new_n23474_, new_n23235_, new_n23233_ );
and  ( new_n23475_, new_n23238_, new_n23474_ );
nor  ( new_n23476_, new_n23475_, new_n23473_ );
xor  ( new_n23477_, new_n23013_, new_n23004_ );
xor  ( new_n23478_, new_n23477_, new_n23065_ );
xor  ( new_n23479_, new_n23478_, new_n23476_ );
or   ( new_n23480_, new_n23466_, new_n23464_ );
and  ( new_n23481_, new_n23466_, new_n23464_ );
or   ( new_n23482_, new_n23481_, new_n23454_ );
and  ( new_n23483_, new_n23482_, new_n23480_ );
xnor ( new_n23484_, new_n23483_, new_n23479_ );
nand ( new_n23485_, new_n23484_, new_n23472_ );
and  ( new_n23486_, new_n23485_, new_n23471_ );
nand ( new_n23487_, new_n23486_, new_n23229_ );
nor  ( new_n23488_, new_n23486_, new_n23229_ );
nor  ( new_n23489_, new_n23478_, new_n23476_ );
nand ( new_n23490_, new_n23478_, new_n23476_ );
and  ( new_n23491_, new_n23483_, new_n23490_ );
nor  ( new_n23492_, new_n23491_, new_n23489_ );
or   ( new_n23493_, new_n23492_, new_n23488_ );
and  ( new_n23494_, new_n23493_, new_n23487_ );
nor  ( new_n23495_, new_n23494_, new_n23227_ );
xor  ( new_n23496_, new_n23445_, new_n23407_ );
xor  ( new_n23497_, new_n23496_, new_n23452_ );
not  ( new_n23498_, new_n23497_ );
xor  ( new_n23499_, new_n23395_, new_n23287_ );
xor  ( new_n23500_, new_n23499_, new_n23399_ );
nor  ( new_n23501_, new_n23500_, new_n23498_ );
xor  ( new_n23502_, new_n23458_, new_n23456_ );
xor  ( new_n23503_, new_n23502_, new_n23462_ );
or   ( new_n23504_, new_n2122_, new_n21703_ );
or   ( new_n23505_, new_n2124_, new_n21694_ );
and  ( new_n23506_, new_n23505_, new_n23504_ );
xor  ( new_n23507_, new_n23506_, new_n1842_ );
and  ( new_n23508_, new_n2244_, RIbb315f0_129 );
xor  ( new_n23509_, new_n23508_, new_n2121_ );
nand ( new_n23510_, new_n23509_, new_n23507_ );
nor  ( new_n23511_, new_n23509_, new_n23507_ );
or   ( new_n23512_, new_n1844_, new_n21674_ );
or   ( new_n23513_, new_n1846_, new_n21701_ );
and  ( new_n23514_, new_n23513_, new_n23512_ );
xor  ( new_n23515_, new_n23514_, new_n1586_ );
or   ( new_n23516_, new_n23515_, new_n23511_ );
and  ( new_n23517_, new_n23516_, new_n23510_ );
or   ( new_n23518_, new_n1593_, new_n21680_ );
or   ( new_n23519_, new_n1595_, new_n21672_ );
and  ( new_n23520_, new_n23519_, new_n23518_ );
xor  ( new_n23521_, new_n23520_, new_n1358_ );
or   ( new_n23522_, new_n1364_, new_n21687_ );
or   ( new_n23523_, new_n1366_, new_n21678_ );
and  ( new_n23524_, new_n23523_, new_n23522_ );
xor  ( new_n23525_, new_n23524_, new_n1129_ );
or   ( new_n23526_, new_n23525_, new_n23521_ );
and  ( new_n23527_, new_n23525_, new_n23521_ );
or   ( new_n23528_, new_n1135_, new_n21751_ );
or   ( new_n23529_, new_n1137_, new_n21685_ );
and  ( new_n23530_, new_n23529_, new_n23528_ );
xor  ( new_n23531_, new_n23530_, new_n896_ );
or   ( new_n23532_, new_n23531_, new_n23527_ );
and  ( new_n23533_, new_n23532_, new_n23526_ );
or   ( new_n23534_, new_n23533_, new_n23517_ );
and  ( new_n23535_, new_n23533_, new_n23517_ );
or   ( new_n23536_, new_n897_, new_n21842_ );
or   ( new_n23537_, new_n899_, new_n21792_ );
and  ( new_n23538_, new_n23537_, new_n23536_ );
xor  ( new_n23539_, new_n23538_, new_n748_ );
or   ( new_n23540_, new_n755_, new_n21847_ );
or   ( new_n23541_, new_n757_, new_n21840_ );
and  ( new_n23542_, new_n23541_, new_n23540_ );
xor  ( new_n23543_, new_n23542_, new_n523_ );
nor  ( new_n23544_, new_n23543_, new_n23539_ );
and  ( new_n23545_, new_n23543_, new_n23539_ );
or   ( new_n23546_, new_n524_, new_n22129_ );
or   ( new_n23547_, new_n526_, new_n22098_ );
and  ( new_n23548_, new_n23547_, new_n23546_ );
xor  ( new_n23549_, new_n23548_, new_n403_ );
nor  ( new_n23550_, new_n23549_, new_n23545_ );
nor  ( new_n23551_, new_n23550_, new_n23544_ );
or   ( new_n23552_, new_n23551_, new_n23535_ );
and  ( new_n23553_, new_n23552_, new_n23534_ );
not  ( new_n23554_, RIbb32310_157 );
or   ( new_n23555_, new_n23554_, new_n260_ );
xnor ( new_n23556_, new_n23367_, new_n23363_ );
xor  ( new_n23557_, new_n23556_, new_n23374_ );
nand ( new_n23558_, new_n23557_, new_n23555_ );
or   ( new_n23559_, new_n23557_, new_n23555_ );
xor  ( new_n23560_, new_n23384_, new_n23380_ );
xnor ( new_n23561_, new_n23560_, new_n23390_ );
nand ( new_n23562_, new_n23561_, new_n23559_ );
and  ( new_n23563_, new_n23562_, new_n23558_ );
nor  ( new_n23564_, new_n23563_, new_n23553_ );
nand ( new_n23565_, new_n23563_, new_n23553_ );
or   ( new_n23566_, new_n283_, new_n22973_ );
or   ( new_n23567_, new_n286_, new_n22975_ );
and  ( new_n23568_, new_n23567_, new_n23566_ );
xor  ( new_n23569_, new_n23568_, new_n278_ );
or   ( new_n23570_, new_n299_, new_n23252_ );
or   ( new_n23571_, new_n302_, new_n23166_ );
and  ( new_n23572_, new_n23571_, new_n23570_ );
xor  ( new_n23573_, new_n23572_, new_n293_ );
nor  ( new_n23574_, new_n23573_, new_n23569_ );
nand ( new_n23575_, new_n23573_, new_n23569_ );
or   ( new_n23576_, new_n268_, new_n23554_ );
or   ( new_n23577_, new_n271_, new_n23370_ );
and  ( new_n23578_, new_n23577_, new_n23576_ );
xor  ( new_n23579_, new_n23578_, new_n262_ );
and  ( new_n23580_, new_n23579_, new_n23575_ );
or   ( new_n23581_, new_n23580_, new_n23574_ );
and  ( new_n23582_, RIbb32388_158, RIbb2f610_1 );
not  ( new_n23583_, new_n23582_ );
or   ( new_n23584_, new_n409_, new_n22304_ );
or   ( new_n23585_, new_n411_, new_n22207_ );
and  ( new_n23586_, new_n23585_, new_n23584_ );
xor  ( new_n23587_, new_n23586_, new_n328_ );
or   ( new_n23588_, new_n337_, new_n22590_ );
or   ( new_n23589_, new_n340_, new_n22423_ );
and  ( new_n23590_, new_n23589_, new_n23588_ );
xor  ( new_n23591_, new_n23590_, new_n332_ );
nor  ( new_n23592_, new_n23591_, new_n23587_ );
and  ( new_n23593_, new_n23591_, new_n23587_ );
or   ( new_n23594_, new_n317_, new_n22829_ );
or   ( new_n23595_, new_n320_, new_n22641_ );
and  ( new_n23596_, new_n23595_, new_n23594_ );
xor  ( new_n23597_, new_n23596_, new_n312_ );
nor  ( new_n23598_, new_n23597_, new_n23593_ );
nor  ( new_n23599_, new_n23598_, new_n23592_ );
not  ( new_n23600_, new_n23599_ );
or   ( new_n23601_, new_n23600_, new_n23583_ );
and  ( new_n23602_, new_n23601_, new_n23581_ );
and  ( new_n23603_, new_n23600_, new_n23583_ );
or   ( new_n23604_, new_n23603_, new_n23602_ );
and  ( new_n23605_, new_n23604_, new_n23565_ );
or   ( new_n23606_, new_n23605_, new_n23564_ );
xnor ( new_n23607_, new_n23413_, new_n23411_ );
xor  ( new_n23608_, new_n23607_, new_n23419_ );
xor  ( new_n23609_, new_n23295_, new_n23291_ );
xor  ( new_n23610_, new_n23609_, new_n23301_ );
xor  ( new_n23611_, new_n23307_, new_n2121_ );
xor  ( new_n23612_, new_n23611_, new_n23313_ );
nand ( new_n23613_, new_n23612_, new_n23610_ );
nor  ( new_n23614_, new_n23612_, new_n23610_ );
xnor ( new_n23615_, new_n23325_, new_n23321_ );
xor  ( new_n23616_, new_n23615_, new_n23331_ );
or   ( new_n23617_, new_n23616_, new_n23614_ );
and  ( new_n23618_, new_n23617_, new_n23613_ );
or   ( new_n23619_, new_n23618_, new_n23608_ );
and  ( new_n23620_, new_n23618_, new_n23608_ );
xnor ( new_n23621_, new_n23433_, new_n23429_ );
xor  ( new_n23622_, new_n23621_, new_n23439_ );
or   ( new_n23623_, new_n23622_, new_n23620_ );
and  ( new_n23624_, new_n23623_, new_n23619_ );
nand ( new_n23625_, new_n23624_, new_n23606_ );
or   ( new_n23626_, new_n23624_, new_n23606_ );
xor  ( new_n23627_, new_n23315_, new_n23303_ );
xor  ( new_n23628_, new_n23627_, new_n23333_ );
xnor ( new_n23629_, new_n23339_, new_n23337_ );
xor  ( new_n23630_, new_n23629_, new_n23355_ );
and  ( new_n23631_, new_n23630_, new_n23628_ );
nor  ( new_n23632_, new_n23630_, new_n23628_ );
xor  ( new_n23633_, new_n23392_, new_n23376_ );
nor  ( new_n23634_, new_n23633_, new_n23632_ );
nor  ( new_n23635_, new_n23634_, new_n23631_ );
nand ( new_n23636_, new_n23635_, new_n23626_ );
and  ( new_n23637_, new_n23636_, new_n23625_ );
or   ( new_n23638_, new_n23637_, new_n23503_ );
and  ( new_n23639_, new_n23637_, new_n23503_ );
xnor ( new_n23640_, new_n23441_, new_n23425_ );
xor  ( new_n23641_, new_n23640_, new_n23421_ );
xor  ( new_n23642_, new_n23357_, new_n23335_ );
xor  ( new_n23643_, new_n23642_, new_n23393_ );
nor  ( new_n23644_, new_n23643_, new_n23641_ );
nand ( new_n23645_, new_n23643_, new_n23641_ );
xor  ( new_n23646_, new_n23281_, new_n23247_ );
xnor ( new_n23647_, new_n23646_, new_n23285_ );
not  ( new_n23648_, new_n23647_ );
and  ( new_n23649_, new_n23648_, new_n23645_ );
or   ( new_n23650_, new_n23649_, new_n23644_ );
or   ( new_n23651_, new_n23650_, new_n23639_ );
and  ( new_n23652_, new_n23651_, new_n23638_ );
nand ( new_n23653_, new_n23652_, new_n23501_ );
nor  ( new_n23654_, new_n23652_, new_n23501_ );
xor  ( new_n23655_, new_n23401_, new_n23239_ );
xnor ( new_n23656_, new_n23655_, new_n23468_ );
or   ( new_n23657_, new_n23656_, new_n23654_ );
and  ( new_n23658_, new_n23657_, new_n23653_ );
xor  ( new_n23659_, new_n23470_, new_n23231_ );
xor  ( new_n23660_, new_n23659_, new_n23484_ );
nor  ( new_n23661_, new_n23660_, new_n23658_ );
xnor ( new_n23662_, new_n23486_, new_n23229_ );
xor  ( new_n23663_, new_n23662_, new_n23492_ );
and  ( new_n23664_, new_n23663_, new_n23661_ );
xnor ( new_n23665_, new_n23652_, new_n23501_ );
xor  ( new_n23666_, new_n23665_, new_n23656_ );
xor  ( new_n23667_, new_n23637_, new_n23503_ );
xor  ( new_n23668_, new_n23667_, new_n23650_ );
or   ( new_n23669_, new_n1135_, new_n21792_ );
or   ( new_n23670_, new_n1137_, new_n21751_ );
and  ( new_n23671_, new_n23670_, new_n23669_ );
xor  ( new_n23672_, new_n23671_, new_n896_ );
or   ( new_n23673_, new_n897_, new_n21840_ );
or   ( new_n23674_, new_n899_, new_n21842_ );
and  ( new_n23675_, new_n23674_, new_n23673_ );
xor  ( new_n23676_, new_n23675_, new_n748_ );
nor  ( new_n23677_, new_n23676_, new_n23672_ );
and  ( new_n23678_, new_n23676_, new_n23672_ );
or   ( new_n23679_, new_n755_, new_n22098_ );
or   ( new_n23680_, new_n757_, new_n21847_ );
and  ( new_n23681_, new_n23680_, new_n23679_ );
xor  ( new_n23682_, new_n23681_, new_n523_ );
nor  ( new_n23683_, new_n23682_, new_n23678_ );
or   ( new_n23684_, new_n23683_, new_n23677_ );
or   ( new_n23685_, new_n2425_, new_n21694_ );
or   ( new_n23686_, new_n2427_, new_n21696_ );
and  ( new_n23687_, new_n23686_, new_n23685_ );
xor  ( new_n23688_, new_n23687_, new_n2121_ );
nand ( new_n23689_, new_n23688_, new_n2424_ );
or   ( new_n23690_, new_n23688_, new_n2424_ );
or   ( new_n23691_, new_n2122_, new_n21701_ );
or   ( new_n23692_, new_n2124_, new_n21703_ );
and  ( new_n23693_, new_n23692_, new_n23691_ );
xor  ( new_n23694_, new_n23693_, new_n1843_ );
nand ( new_n23695_, new_n23694_, new_n23690_ );
and  ( new_n23696_, new_n23695_, new_n23689_ );
nand ( new_n23697_, new_n23696_, new_n23684_ );
nor  ( new_n23698_, new_n23696_, new_n23684_ );
or   ( new_n23699_, new_n1844_, new_n21672_ );
or   ( new_n23700_, new_n1846_, new_n21674_ );
and  ( new_n23701_, new_n23700_, new_n23699_ );
xor  ( new_n23702_, new_n23701_, new_n1586_ );
or   ( new_n23703_, new_n1593_, new_n21678_ );
or   ( new_n23704_, new_n1595_, new_n21680_ );
and  ( new_n23705_, new_n23704_, new_n23703_ );
xor  ( new_n23706_, new_n23705_, new_n1358_ );
nor  ( new_n23707_, new_n23706_, new_n23702_ );
and  ( new_n23708_, new_n23706_, new_n23702_ );
or   ( new_n23709_, new_n1364_, new_n21685_ );
or   ( new_n23710_, new_n1366_, new_n21687_ );
and  ( new_n23711_, new_n23710_, new_n23709_ );
xor  ( new_n23712_, new_n23711_, new_n1129_ );
nor  ( new_n23713_, new_n23712_, new_n23708_ );
nor  ( new_n23714_, new_n23713_, new_n23707_ );
or   ( new_n23715_, new_n23714_, new_n23698_ );
and  ( new_n23716_, new_n23715_, new_n23697_ );
or   ( new_n23717_, new_n317_, new_n22975_ );
or   ( new_n23718_, new_n320_, new_n22829_ );
and  ( new_n23719_, new_n23718_, new_n23717_ );
xor  ( new_n23720_, new_n23719_, new_n312_ );
or   ( new_n23721_, new_n283_, new_n23166_ );
or   ( new_n23722_, new_n286_, new_n22973_ );
and  ( new_n23723_, new_n23722_, new_n23721_ );
xor  ( new_n23724_, new_n23723_, new_n278_ );
nor  ( new_n23725_, new_n23724_, new_n23720_ );
and  ( new_n23726_, new_n23724_, new_n23720_ );
or   ( new_n23727_, new_n299_, new_n23370_ );
or   ( new_n23728_, new_n302_, new_n23252_ );
and  ( new_n23729_, new_n23728_, new_n23727_ );
xor  ( new_n23730_, new_n23729_, new_n293_ );
nor  ( new_n23731_, new_n23730_, new_n23726_ );
nor  ( new_n23732_, new_n23731_, new_n23725_ );
not  ( new_n23733_, RIbb32388_158 );
or   ( new_n23734_, new_n268_, new_n23733_ );
or   ( new_n23735_, new_n271_, new_n23554_ );
and  ( new_n23736_, new_n23735_, new_n23734_ );
xor  ( new_n23737_, new_n23736_, new_n263_ );
and  ( new_n23738_, RIbb32400_159, RIbb2f610_1 );
and  ( new_n23739_, new_n23738_, new_n23737_ );
or   ( new_n23740_, new_n524_, new_n22207_ );
or   ( new_n23741_, new_n526_, new_n22129_ );
and  ( new_n23742_, new_n23741_, new_n23740_ );
xor  ( new_n23743_, new_n23742_, new_n403_ );
or   ( new_n23744_, new_n409_, new_n22423_ );
or   ( new_n23745_, new_n411_, new_n22304_ );
and  ( new_n23746_, new_n23745_, new_n23744_ );
xor  ( new_n23747_, new_n23746_, new_n328_ );
or   ( new_n23748_, new_n23747_, new_n23743_ );
and  ( new_n23749_, new_n23747_, new_n23743_ );
or   ( new_n23750_, new_n337_, new_n22641_ );
or   ( new_n23751_, new_n340_, new_n22590_ );
and  ( new_n23752_, new_n23751_, new_n23750_ );
xor  ( new_n23753_, new_n23752_, new_n332_ );
or   ( new_n23754_, new_n23753_, new_n23749_ );
and  ( new_n23755_, new_n23754_, new_n23748_ );
and  ( new_n23756_, new_n23755_, new_n23739_ );
or   ( new_n23757_, new_n23756_, new_n23732_ );
or   ( new_n23758_, new_n23755_, new_n23739_ );
and  ( new_n23759_, new_n23758_, new_n23757_ );
nor  ( new_n23760_, new_n23759_, new_n23716_ );
nand ( new_n23761_, new_n23759_, new_n23716_ );
xor  ( new_n23762_, new_n23573_, new_n23569_ );
xor  ( new_n23763_, new_n23762_, new_n23579_ );
xnor ( new_n23764_, new_n23591_, new_n23587_ );
xor  ( new_n23765_, new_n23764_, new_n23597_ );
nor  ( new_n23766_, new_n23765_, new_n23763_ );
and  ( new_n23767_, new_n23765_, new_n23763_ );
nor  ( new_n23768_, new_n23767_, new_n23582_ );
nor  ( new_n23769_, new_n23768_, new_n23766_ );
and  ( new_n23770_, new_n23769_, new_n23761_ );
or   ( new_n23771_, new_n23770_, new_n23760_ );
xor  ( new_n23772_, new_n23612_, new_n23610_ );
xor  ( new_n23773_, new_n23772_, new_n23616_ );
xnor ( new_n23774_, new_n23525_, new_n23521_ );
xor  ( new_n23775_, new_n23774_, new_n23531_ );
xnor ( new_n23776_, new_n23509_, new_n23507_ );
xor  ( new_n23777_, new_n23776_, new_n23515_ );
or   ( new_n23778_, new_n23777_, new_n23775_ );
and  ( new_n23779_, new_n23777_, new_n23775_ );
xnor ( new_n23780_, new_n23543_, new_n23539_ );
xor  ( new_n23781_, new_n23780_, new_n23549_ );
or   ( new_n23782_, new_n23781_, new_n23779_ );
and  ( new_n23783_, new_n23782_, new_n23778_ );
or   ( new_n23784_, new_n23783_, new_n23773_ );
and  ( new_n23785_, new_n23783_, new_n23773_ );
xor  ( new_n23786_, new_n23557_, new_n23555_ );
xor  ( new_n23787_, new_n23786_, new_n23561_ );
or   ( new_n23788_, new_n23787_, new_n23785_ );
and  ( new_n23789_, new_n23788_, new_n23784_ );
and  ( new_n23790_, new_n23789_, new_n23771_ );
or   ( new_n23791_, new_n23789_, new_n23771_ );
xor  ( new_n23792_, new_n23533_, new_n23517_ );
xnor ( new_n23793_, new_n23792_, new_n23551_ );
not  ( new_n23794_, new_n23793_ );
xor  ( new_n23795_, new_n23599_, new_n23583_ );
xor  ( new_n23796_, new_n23795_, new_n23581_ );
and  ( new_n23797_, new_n23796_, new_n23794_ );
not  ( new_n23798_, new_n23797_ );
and  ( new_n23799_, new_n23798_, new_n23791_ );
or   ( new_n23800_, new_n23799_, new_n23790_ );
xor  ( new_n23801_, new_n23618_, new_n23608_ );
xor  ( new_n23802_, new_n23801_, new_n23622_ );
xor  ( new_n23803_, new_n23563_, new_n23553_ );
xor  ( new_n23804_, new_n23803_, new_n23604_ );
or   ( new_n23805_, new_n23804_, new_n23802_ );
and  ( new_n23806_, new_n23804_, new_n23802_ );
xor  ( new_n23807_, new_n23630_, new_n23628_ );
xor  ( new_n23808_, new_n23807_, new_n23633_ );
or   ( new_n23809_, new_n23808_, new_n23806_ );
and  ( new_n23810_, new_n23809_, new_n23805_ );
nand ( new_n23811_, new_n23810_, new_n23800_ );
nor  ( new_n23812_, new_n23810_, new_n23800_ );
xor  ( new_n23813_, new_n23643_, new_n23641_ );
xor  ( new_n23814_, new_n23813_, new_n23648_ );
or   ( new_n23815_, new_n23814_, new_n23812_ );
and  ( new_n23816_, new_n23815_, new_n23811_ );
or   ( new_n23817_, new_n23816_, new_n23668_ );
and  ( new_n23818_, new_n23816_, new_n23668_ );
xor  ( new_n23819_, new_n23500_, new_n23498_ );
or   ( new_n23820_, new_n23819_, new_n23818_ );
and  ( new_n23821_, new_n23820_, new_n23817_ );
and  ( new_n23822_, new_n23821_, new_n23666_ );
xor  ( new_n23823_, new_n23660_, new_n23658_ );
and  ( new_n23824_, new_n23823_, new_n23822_ );
xnor ( new_n23825_, new_n23759_, new_n23716_ );
xor  ( new_n23826_, new_n23825_, new_n23769_ );
xnor ( new_n23827_, new_n23783_, new_n23773_ );
xor  ( new_n23828_, new_n23827_, new_n23787_ );
nor  ( new_n23829_, new_n23828_, new_n23826_ );
nand ( new_n23830_, new_n23828_, new_n23826_ );
xor  ( new_n23831_, new_n23796_, new_n23794_ );
not  ( new_n23832_, new_n23831_ );
and  ( new_n23833_, new_n23832_, new_n23830_ );
or   ( new_n23834_, new_n23833_, new_n23829_ );
xor  ( new_n23835_, new_n23804_, new_n23802_ );
xor  ( new_n23836_, new_n23835_, new_n23808_ );
or   ( new_n23837_, new_n23836_, new_n23834_ );
and  ( new_n23838_, new_n23836_, new_n23834_ );
xor  ( new_n23839_, new_n23696_, new_n23684_ );
xnor ( new_n23840_, new_n23839_, new_n23714_ );
not  ( new_n23841_, new_n23840_ );
xor  ( new_n23842_, new_n23755_, new_n23739_ );
xor  ( new_n23843_, new_n23842_, new_n23732_ );
nand ( new_n23844_, new_n23843_, new_n23841_ );
or   ( new_n23845_, new_n1135_, new_n21842_ );
or   ( new_n23846_, new_n1137_, new_n21792_ );
and  ( new_n23847_, new_n23846_, new_n23845_ );
xor  ( new_n23848_, new_n23847_, new_n896_ );
or   ( new_n23849_, new_n897_, new_n21847_ );
or   ( new_n23850_, new_n899_, new_n21840_ );
and  ( new_n23851_, new_n23850_, new_n23849_ );
xor  ( new_n23852_, new_n23851_, new_n748_ );
or   ( new_n23853_, new_n23852_, new_n23848_ );
and  ( new_n23854_, new_n23852_, new_n23848_ );
or   ( new_n23855_, new_n755_, new_n22129_ );
or   ( new_n23856_, new_n757_, new_n22098_ );
and  ( new_n23857_, new_n23856_, new_n23855_ );
xor  ( new_n23858_, new_n23857_, new_n523_ );
or   ( new_n23859_, new_n23858_, new_n23854_ );
and  ( new_n23860_, new_n23859_, new_n23853_ );
or   ( new_n23861_, new_n2425_, new_n21703_ );
or   ( new_n23862_, new_n2427_, new_n21694_ );
and  ( new_n23863_, new_n23862_, new_n23861_ );
xor  ( new_n23864_, new_n23863_, new_n2120_ );
and  ( new_n23865_, new_n2615_, RIbb315f0_129 );
xor  ( new_n23866_, new_n23865_, new_n2424_ );
nand ( new_n23867_, new_n23866_, new_n23864_ );
nor  ( new_n23868_, new_n23866_, new_n23864_ );
or   ( new_n23869_, new_n2122_, new_n21674_ );
or   ( new_n23870_, new_n2124_, new_n21701_ );
and  ( new_n23871_, new_n23870_, new_n23869_ );
xor  ( new_n23872_, new_n23871_, new_n1843_ );
or   ( new_n23873_, new_n23872_, new_n23868_ );
and  ( new_n23874_, new_n23873_, new_n23867_ );
or   ( new_n23875_, new_n23874_, new_n23860_ );
and  ( new_n23876_, new_n23874_, new_n23860_ );
or   ( new_n23877_, new_n1844_, new_n21680_ );
or   ( new_n23878_, new_n1846_, new_n21672_ );
and  ( new_n23879_, new_n23878_, new_n23877_ );
xor  ( new_n23880_, new_n23879_, new_n1586_ );
or   ( new_n23881_, new_n1593_, new_n21687_ );
or   ( new_n23882_, new_n1595_, new_n21678_ );
and  ( new_n23883_, new_n23882_, new_n23881_ );
xor  ( new_n23884_, new_n23883_, new_n1358_ );
nor  ( new_n23885_, new_n23884_, new_n23880_ );
and  ( new_n23886_, new_n23884_, new_n23880_ );
or   ( new_n23887_, new_n1364_, new_n21751_ );
or   ( new_n23888_, new_n1366_, new_n21685_ );
and  ( new_n23889_, new_n23888_, new_n23887_ );
xor  ( new_n23890_, new_n23889_, new_n1129_ );
nor  ( new_n23891_, new_n23890_, new_n23886_ );
nor  ( new_n23892_, new_n23891_, new_n23885_ );
or   ( new_n23893_, new_n23892_, new_n23876_ );
and  ( new_n23894_, new_n23893_, new_n23875_ );
not  ( new_n23895_, RIbb32400_159 );
or   ( new_n23896_, new_n268_, new_n23895_ );
or   ( new_n23897_, new_n271_, new_n23733_ );
and  ( new_n23898_, new_n23897_, new_n23896_ );
xor  ( new_n23899_, new_n23898_, new_n263_ );
and  ( new_n23900_, RIbb32478_160, RIbb2f610_1 );
or   ( new_n23901_, new_n23900_, new_n23899_ );
or   ( new_n23902_, new_n317_, new_n22973_ );
or   ( new_n23903_, new_n320_, new_n22975_ );
and  ( new_n23904_, new_n23903_, new_n23902_ );
xor  ( new_n23905_, new_n23904_, new_n312_ );
or   ( new_n23906_, new_n283_, new_n23252_ );
or   ( new_n23907_, new_n286_, new_n23166_ );
and  ( new_n23908_, new_n23907_, new_n23906_ );
xor  ( new_n23909_, new_n23908_, new_n278_ );
or   ( new_n23910_, new_n23909_, new_n23905_ );
and  ( new_n23911_, new_n23909_, new_n23905_ );
or   ( new_n23912_, new_n299_, new_n23554_ );
or   ( new_n23913_, new_n302_, new_n23370_ );
and  ( new_n23914_, new_n23913_, new_n23912_ );
xor  ( new_n23915_, new_n23914_, new_n293_ );
or   ( new_n23916_, new_n23915_, new_n23911_ );
and  ( new_n23917_, new_n23916_, new_n23910_ );
or   ( new_n23918_, new_n23917_, new_n23901_ );
and  ( new_n23919_, new_n23917_, new_n23901_ );
or   ( new_n23920_, new_n524_, new_n22304_ );
or   ( new_n23921_, new_n526_, new_n22207_ );
and  ( new_n23922_, new_n23921_, new_n23920_ );
xor  ( new_n23923_, new_n23922_, new_n403_ );
or   ( new_n23924_, new_n409_, new_n22590_ );
or   ( new_n23925_, new_n411_, new_n22423_ );
and  ( new_n23926_, new_n23925_, new_n23924_ );
xor  ( new_n23927_, new_n23926_, new_n328_ );
nor  ( new_n23928_, new_n23927_, new_n23923_ );
and  ( new_n23929_, new_n23927_, new_n23923_ );
or   ( new_n23930_, new_n337_, new_n22829_ );
or   ( new_n23931_, new_n340_, new_n22641_ );
and  ( new_n23932_, new_n23931_, new_n23930_ );
xor  ( new_n23933_, new_n23932_, new_n332_ );
nor  ( new_n23934_, new_n23933_, new_n23929_ );
nor  ( new_n23935_, new_n23934_, new_n23928_ );
or   ( new_n23936_, new_n23935_, new_n23919_ );
and  ( new_n23937_, new_n23936_, new_n23918_ );
nand ( new_n23938_, new_n23937_, new_n23894_ );
nor  ( new_n23939_, new_n23937_, new_n23894_ );
xnor ( new_n23940_, new_n23724_, new_n23720_ );
xor  ( new_n23941_, new_n23940_, new_n23730_ );
xnor ( new_n23942_, new_n23747_, new_n23743_ );
xor  ( new_n23943_, new_n23942_, new_n23753_ );
nor  ( new_n23944_, new_n23943_, new_n23941_ );
and  ( new_n23945_, new_n23943_, new_n23941_ );
xor  ( new_n23946_, new_n23738_, new_n23737_ );
not  ( new_n23947_, new_n23946_ );
nor  ( new_n23948_, new_n23947_, new_n23945_ );
nor  ( new_n23949_, new_n23948_, new_n23944_ );
or   ( new_n23950_, new_n23949_, new_n23939_ );
and  ( new_n23951_, new_n23950_, new_n23938_ );
nor  ( new_n23952_, new_n23951_, new_n23844_ );
and  ( new_n23953_, new_n23951_, new_n23844_ );
xor  ( new_n23954_, new_n23777_, new_n23775_ );
xor  ( new_n23955_, new_n23954_, new_n23781_ );
xor  ( new_n23956_, new_n23676_, new_n23672_ );
xor  ( new_n23957_, new_n23956_, new_n23682_ );
xor  ( new_n23958_, new_n23688_, new_n2424_ );
xor  ( new_n23959_, new_n23958_, new_n23694_ );
nand ( new_n23960_, new_n23959_, new_n23957_ );
nor  ( new_n23961_, new_n23959_, new_n23957_ );
xnor ( new_n23962_, new_n23706_, new_n23702_ );
xor  ( new_n23963_, new_n23962_, new_n23712_ );
or   ( new_n23964_, new_n23963_, new_n23961_ );
and  ( new_n23965_, new_n23964_, new_n23960_ );
nor  ( new_n23966_, new_n23965_, new_n23955_ );
and  ( new_n23967_, new_n23965_, new_n23955_ );
xor  ( new_n23968_, new_n23765_, new_n23763_ );
xnor ( new_n23969_, new_n23968_, new_n23583_ );
nor  ( new_n23970_, new_n23969_, new_n23967_ );
nor  ( new_n23971_, new_n23970_, new_n23966_ );
nor  ( new_n23972_, new_n23971_, new_n23953_ );
nor  ( new_n23973_, new_n23972_, new_n23952_ );
or   ( new_n23974_, new_n23973_, new_n23838_ );
and  ( new_n23975_, new_n23974_, new_n23837_ );
xor  ( new_n23976_, new_n23624_, new_n23606_ );
xor  ( new_n23977_, new_n23976_, new_n23635_ );
or   ( new_n23978_, new_n23977_, new_n23975_ );
and  ( new_n23979_, new_n23977_, new_n23975_ );
xor  ( new_n23980_, new_n23810_, new_n23800_ );
xnor ( new_n23981_, new_n23980_, new_n23814_ );
or   ( new_n23982_, new_n23981_, new_n23979_ );
and  ( new_n23983_, new_n23982_, new_n23978_ );
xnor ( new_n23984_, new_n23816_, new_n23668_ );
xor  ( new_n23985_, new_n23984_, new_n23819_ );
nor  ( new_n23986_, new_n23985_, new_n23983_ );
xor  ( new_n23987_, new_n23821_, new_n23666_ );
and  ( new_n23988_, new_n23987_, new_n23986_ );
xnor ( new_n23989_, new_n23977_, new_n23975_ );
xor  ( new_n23990_, new_n23989_, new_n23981_ );
xnor ( new_n23991_, new_n23836_, new_n23834_ );
xor  ( new_n23992_, new_n23991_, new_n23973_ );
xnor ( new_n23993_, new_n23965_, new_n23955_ );
xor  ( new_n23994_, new_n23993_, new_n23969_ );
xnor ( new_n23995_, new_n23937_, new_n23894_ );
xor  ( new_n23996_, new_n23995_, new_n23949_ );
or   ( new_n23997_, new_n23996_, new_n23994_ );
and  ( new_n23998_, new_n23996_, new_n23994_ );
xor  ( new_n23999_, new_n23843_, new_n23841_ );
or   ( new_n24000_, new_n23999_, new_n23998_ );
and  ( new_n24001_, new_n24000_, new_n23997_ );
or   ( new_n24002_, new_n299_, new_n23733_ );
or   ( new_n24003_, new_n302_, new_n23554_ );
and  ( new_n24004_, new_n24003_, new_n24002_ );
xor  ( new_n24005_, new_n24004_, new_n293_ );
not  ( new_n24006_, RIbb32478_160 );
or   ( new_n24007_, new_n268_, new_n24006_ );
or   ( new_n24008_, new_n271_, new_n23895_ );
and  ( new_n24009_, new_n24008_, new_n24007_ );
xor  ( new_n24010_, new_n24009_, new_n263_ );
or   ( new_n24011_, new_n24010_, new_n24005_ );
and  ( new_n24012_, RIbb324f0_161, RIbb2f610_1 );
and  ( new_n24013_, new_n24010_, new_n24005_ );
or   ( new_n24014_, new_n24013_, new_n24012_ );
and  ( new_n24015_, new_n24014_, new_n24011_ );
or   ( new_n24016_, new_n337_, new_n22975_ );
or   ( new_n24017_, new_n340_, new_n22829_ );
and  ( new_n24018_, new_n24017_, new_n24016_ );
xor  ( new_n24019_, new_n24018_, new_n332_ );
or   ( new_n24020_, new_n317_, new_n23166_ );
or   ( new_n24021_, new_n320_, new_n22973_ );
and  ( new_n24022_, new_n24021_, new_n24020_ );
xor  ( new_n24023_, new_n24022_, new_n312_ );
or   ( new_n24024_, new_n24023_, new_n24019_ );
and  ( new_n24025_, new_n24023_, new_n24019_ );
or   ( new_n24026_, new_n283_, new_n23370_ );
or   ( new_n24027_, new_n286_, new_n23252_ );
and  ( new_n24028_, new_n24027_, new_n24026_ );
xor  ( new_n24029_, new_n24028_, new_n278_ );
or   ( new_n24030_, new_n24029_, new_n24025_ );
and  ( new_n24031_, new_n24030_, new_n24024_ );
or   ( new_n24032_, new_n24031_, new_n24015_ );
and  ( new_n24033_, new_n24031_, new_n24015_ );
or   ( new_n24034_, new_n755_, new_n22207_ );
or   ( new_n24035_, new_n757_, new_n22129_ );
and  ( new_n24036_, new_n24035_, new_n24034_ );
xor  ( new_n24037_, new_n24036_, new_n523_ );
or   ( new_n24038_, new_n524_, new_n22423_ );
or   ( new_n24039_, new_n526_, new_n22304_ );
and  ( new_n24040_, new_n24039_, new_n24038_ );
xor  ( new_n24041_, new_n24040_, new_n403_ );
nor  ( new_n24042_, new_n24041_, new_n24037_ );
and  ( new_n24043_, new_n24041_, new_n24037_ );
or   ( new_n24044_, new_n409_, new_n22641_ );
or   ( new_n24045_, new_n411_, new_n22590_ );
and  ( new_n24046_, new_n24045_, new_n24044_ );
xor  ( new_n24047_, new_n24046_, new_n328_ );
nor  ( new_n24048_, new_n24047_, new_n24043_ );
nor  ( new_n24049_, new_n24048_, new_n24042_ );
or   ( new_n24050_, new_n24049_, new_n24033_ );
and  ( new_n24051_, new_n24050_, new_n24032_ );
or   ( new_n24052_, new_n2425_, new_n21701_ );
or   ( new_n24053_, new_n2427_, new_n21703_ );
and  ( new_n24054_, new_n24053_, new_n24052_ );
xor  ( new_n24055_, new_n24054_, new_n2121_ );
and  ( new_n24056_, new_n24055_, new_n2800_ );
or   ( new_n24057_, new_n24055_, new_n2800_ );
or   ( new_n24058_, new_n2807_, new_n21694_ );
or   ( new_n24059_, new_n2809_, new_n21696_ );
and  ( new_n24060_, new_n24059_, new_n24058_ );
xor  ( new_n24061_, new_n24060_, new_n2424_ );
and  ( new_n24062_, new_n24061_, new_n24057_ );
or   ( new_n24063_, new_n24062_, new_n24056_ );
or   ( new_n24064_, new_n2122_, new_n21672_ );
or   ( new_n24065_, new_n2124_, new_n21674_ );
and  ( new_n24066_, new_n24065_, new_n24064_ );
xor  ( new_n24067_, new_n24066_, new_n1843_ );
or   ( new_n24068_, new_n1844_, new_n21678_ );
or   ( new_n24069_, new_n1846_, new_n21680_ );
and  ( new_n24070_, new_n24069_, new_n24068_ );
xor  ( new_n24071_, new_n24070_, new_n1586_ );
or   ( new_n24072_, new_n24071_, new_n24067_ );
and  ( new_n24073_, new_n24071_, new_n24067_ );
or   ( new_n24074_, new_n1593_, new_n21685_ );
or   ( new_n24075_, new_n1595_, new_n21687_ );
and  ( new_n24076_, new_n24075_, new_n24074_ );
xor  ( new_n24077_, new_n24076_, new_n1358_ );
or   ( new_n24078_, new_n24077_, new_n24073_ );
and  ( new_n24079_, new_n24078_, new_n24072_ );
or   ( new_n24080_, new_n24079_, new_n24063_ );
and  ( new_n24081_, new_n24079_, new_n24063_ );
or   ( new_n24082_, new_n1364_, new_n21792_ );
or   ( new_n24083_, new_n1366_, new_n21751_ );
and  ( new_n24084_, new_n24083_, new_n24082_ );
xor  ( new_n24085_, new_n24084_, new_n1129_ );
or   ( new_n24086_, new_n1135_, new_n21840_ );
or   ( new_n24087_, new_n1137_, new_n21842_ );
and  ( new_n24088_, new_n24087_, new_n24086_ );
xor  ( new_n24089_, new_n24088_, new_n896_ );
nor  ( new_n24090_, new_n24089_, new_n24085_ );
and  ( new_n24091_, new_n24089_, new_n24085_ );
or   ( new_n24092_, new_n897_, new_n22098_ );
or   ( new_n24093_, new_n899_, new_n21847_ );
and  ( new_n24094_, new_n24093_, new_n24092_ );
xor  ( new_n24095_, new_n24094_, new_n748_ );
nor  ( new_n24096_, new_n24095_, new_n24091_ );
nor  ( new_n24097_, new_n24096_, new_n24090_ );
or   ( new_n24098_, new_n24097_, new_n24081_ );
and  ( new_n24099_, new_n24098_, new_n24080_ );
nor  ( new_n24100_, new_n24099_, new_n24051_ );
nand ( new_n24101_, new_n24099_, new_n24051_ );
xnor ( new_n24102_, new_n23909_, new_n23905_ );
xor  ( new_n24103_, new_n24102_, new_n23915_ );
xnor ( new_n24104_, new_n23927_, new_n23923_ );
xor  ( new_n24105_, new_n24104_, new_n23933_ );
or   ( new_n24106_, new_n24105_, new_n24103_ );
and  ( new_n24107_, new_n24105_, new_n24103_ );
xor  ( new_n24108_, new_n23900_, new_n23899_ );
or   ( new_n24109_, new_n24108_, new_n24107_ );
and  ( new_n24110_, new_n24109_, new_n24106_ );
and  ( new_n24111_, new_n24110_, new_n24101_ );
or   ( new_n24112_, new_n24111_, new_n24100_ );
xor  ( new_n24113_, new_n23959_, new_n23957_ );
xor  ( new_n24114_, new_n24113_, new_n23963_ );
xnor ( new_n24115_, new_n23866_, new_n23864_ );
xor  ( new_n24116_, new_n24115_, new_n23872_ );
xnor ( new_n24117_, new_n23852_, new_n23848_ );
xor  ( new_n24118_, new_n24117_, new_n23858_ );
or   ( new_n24119_, new_n24118_, new_n24116_ );
and  ( new_n24120_, new_n24118_, new_n24116_ );
xnor ( new_n24121_, new_n23884_, new_n23880_ );
xor  ( new_n24122_, new_n24121_, new_n23890_ );
or   ( new_n24123_, new_n24122_, new_n24120_ );
and  ( new_n24124_, new_n24123_, new_n24119_ );
or   ( new_n24125_, new_n24124_, new_n24114_ );
and  ( new_n24126_, new_n24124_, new_n24114_ );
xor  ( new_n24127_, new_n23943_, new_n23941_ );
xor  ( new_n24128_, new_n24127_, new_n23947_ );
or   ( new_n24129_, new_n24128_, new_n24126_ );
and  ( new_n24130_, new_n24129_, new_n24125_ );
nand ( new_n24131_, new_n24130_, new_n24112_ );
nor  ( new_n24132_, new_n24130_, new_n24112_ );
xor  ( new_n24133_, new_n23874_, new_n23860_ );
xnor ( new_n24134_, new_n24133_, new_n23892_ );
xnor ( new_n24135_, new_n23917_, new_n23901_ );
xor  ( new_n24136_, new_n24135_, new_n23935_ );
nor  ( new_n24137_, new_n24136_, new_n24134_ );
or   ( new_n24138_, new_n24137_, new_n24132_ );
and  ( new_n24139_, new_n24138_, new_n24131_ );
or   ( new_n24140_, new_n24139_, new_n24001_ );
nand ( new_n24141_, new_n24139_, new_n24001_ );
xor  ( new_n24142_, new_n23828_, new_n23826_ );
xor  ( new_n24143_, new_n24142_, new_n23832_ );
nand ( new_n24144_, new_n24143_, new_n24141_ );
and  ( new_n24145_, new_n24144_, new_n24140_ );
or   ( new_n24146_, new_n24145_, new_n23992_ );
nand ( new_n24147_, new_n24145_, new_n23992_ );
xor  ( new_n24148_, new_n23789_, new_n23771_ );
xor  ( new_n24149_, new_n24148_, new_n23798_ );
nand ( new_n24150_, new_n24149_, new_n24147_ );
and  ( new_n24151_, new_n24150_, new_n24146_ );
and  ( new_n24152_, new_n24151_, new_n23990_ );
xor  ( new_n24153_, new_n23985_, new_n23983_ );
and  ( new_n24154_, new_n24153_, new_n24152_ );
xnor ( new_n24155_, new_n23996_, new_n23994_ );
xor  ( new_n24156_, new_n24155_, new_n23999_ );
xor  ( new_n24157_, new_n24099_, new_n24051_ );
xor  ( new_n24158_, new_n24157_, new_n24110_ );
xor  ( new_n24159_, new_n24124_, new_n24114_ );
xor  ( new_n24160_, new_n24159_, new_n24128_ );
or   ( new_n24161_, new_n24160_, new_n24158_ );
nand ( new_n24162_, new_n24160_, new_n24158_ );
xor  ( new_n24163_, new_n24136_, new_n24134_ );
nand ( new_n24164_, new_n24163_, new_n24162_ );
and  ( new_n24165_, new_n24164_, new_n24161_ );
nor  ( new_n24166_, new_n24165_, new_n24156_ );
nand ( new_n24167_, new_n24165_, new_n24156_ );
xnor ( new_n24168_, new_n24031_, new_n24015_ );
xor  ( new_n24169_, new_n24168_, new_n24049_ );
xnor ( new_n24170_, new_n24079_, new_n24063_ );
xor  ( new_n24171_, new_n24170_, new_n24097_ );
or   ( new_n24172_, new_n24171_, new_n24169_ );
or   ( new_n24173_, new_n2807_, new_n21703_ );
or   ( new_n24174_, new_n2809_, new_n21694_ );
and  ( new_n24175_, new_n24174_, new_n24173_ );
xor  ( new_n24176_, new_n24175_, new_n2423_ );
and  ( new_n24177_, new_n2930_, RIbb315f0_129 );
xor  ( new_n24178_, new_n24177_, new_n2800_ );
nand ( new_n24179_, new_n24178_, new_n24176_ );
nor  ( new_n24180_, new_n24178_, new_n24176_ );
or   ( new_n24181_, new_n2425_, new_n21674_ );
or   ( new_n24182_, new_n2427_, new_n21701_ );
and  ( new_n24183_, new_n24182_, new_n24181_ );
xor  ( new_n24184_, new_n24183_, new_n2121_ );
or   ( new_n24185_, new_n24184_, new_n24180_ );
and  ( new_n24186_, new_n24185_, new_n24179_ );
or   ( new_n24187_, new_n2122_, new_n21680_ );
or   ( new_n24188_, new_n2124_, new_n21672_ );
and  ( new_n24189_, new_n24188_, new_n24187_ );
xor  ( new_n24190_, new_n24189_, new_n1843_ );
or   ( new_n24191_, new_n1844_, new_n21687_ );
or   ( new_n24192_, new_n1846_, new_n21678_ );
and  ( new_n24193_, new_n24192_, new_n24191_ );
xor  ( new_n24194_, new_n24193_, new_n1586_ );
or   ( new_n24195_, new_n24194_, new_n24190_ );
and  ( new_n24196_, new_n24194_, new_n24190_ );
or   ( new_n24197_, new_n1593_, new_n21751_ );
or   ( new_n24198_, new_n1595_, new_n21685_ );
and  ( new_n24199_, new_n24198_, new_n24197_ );
xor  ( new_n24200_, new_n24199_, new_n1358_ );
or   ( new_n24201_, new_n24200_, new_n24196_ );
and  ( new_n24202_, new_n24201_, new_n24195_ );
nor  ( new_n24203_, new_n24202_, new_n24186_ );
nand ( new_n24204_, new_n24202_, new_n24186_ );
or   ( new_n24205_, new_n1364_, new_n21842_ );
or   ( new_n24206_, new_n1366_, new_n21792_ );
and  ( new_n24207_, new_n24206_, new_n24205_ );
xor  ( new_n24208_, new_n24207_, new_n1129_ );
or   ( new_n24209_, new_n1135_, new_n21847_ );
or   ( new_n24210_, new_n1137_, new_n21840_ );
and  ( new_n24211_, new_n24210_, new_n24209_ );
xor  ( new_n24212_, new_n24211_, new_n896_ );
nor  ( new_n24213_, new_n24212_, new_n24208_ );
nand ( new_n24214_, new_n24212_, new_n24208_ );
or   ( new_n24215_, new_n897_, new_n22129_ );
or   ( new_n24216_, new_n899_, new_n22098_ );
and  ( new_n24217_, new_n24216_, new_n24215_ );
xor  ( new_n24218_, new_n24217_, new_n747_ );
and  ( new_n24219_, new_n24218_, new_n24214_ );
or   ( new_n24220_, new_n24219_, new_n24213_ );
and  ( new_n24221_, new_n24220_, new_n24204_ );
or   ( new_n24222_, new_n24221_, new_n24203_ );
or   ( new_n24223_, new_n299_, new_n23895_ );
or   ( new_n24224_, new_n302_, new_n23733_ );
and  ( new_n24225_, new_n24224_, new_n24223_ );
xor  ( new_n24226_, new_n24225_, new_n293_ );
not  ( new_n24227_, RIbb324f0_161 );
or   ( new_n24228_, new_n268_, new_n24227_ );
or   ( new_n24229_, new_n271_, new_n24006_ );
and  ( new_n24230_, new_n24229_, new_n24228_ );
xor  ( new_n24231_, new_n24230_, new_n263_ );
or   ( new_n24232_, new_n24231_, new_n24226_ );
and  ( new_n24233_, RIbb32568_162, RIbb2f610_1 );
and  ( new_n24234_, new_n24231_, new_n24226_ );
or   ( new_n24235_, new_n24234_, new_n24233_ );
and  ( new_n24236_, new_n24235_, new_n24232_ );
or   ( new_n24237_, new_n337_, new_n22973_ );
or   ( new_n24238_, new_n340_, new_n22975_ );
and  ( new_n24239_, new_n24238_, new_n24237_ );
xor  ( new_n24240_, new_n24239_, new_n332_ );
or   ( new_n24241_, new_n317_, new_n23252_ );
or   ( new_n24242_, new_n320_, new_n23166_ );
and  ( new_n24243_, new_n24242_, new_n24241_ );
xor  ( new_n24244_, new_n24243_, new_n312_ );
or   ( new_n24245_, new_n24244_, new_n24240_ );
and  ( new_n24246_, new_n24244_, new_n24240_ );
or   ( new_n24247_, new_n283_, new_n23554_ );
or   ( new_n24248_, new_n286_, new_n23370_ );
and  ( new_n24249_, new_n24248_, new_n24247_ );
xor  ( new_n24250_, new_n24249_, new_n278_ );
or   ( new_n24251_, new_n24250_, new_n24246_ );
and  ( new_n24252_, new_n24251_, new_n24245_ );
nor  ( new_n24253_, new_n24252_, new_n24236_ );
and  ( new_n24254_, new_n24252_, new_n24236_ );
or   ( new_n24255_, new_n755_, new_n22304_ );
or   ( new_n24256_, new_n757_, new_n22207_ );
and  ( new_n24257_, new_n24256_, new_n24255_ );
xor  ( new_n24258_, new_n24257_, new_n523_ );
or   ( new_n24259_, new_n524_, new_n22590_ );
or   ( new_n24260_, new_n526_, new_n22423_ );
and  ( new_n24261_, new_n24260_, new_n24259_ );
xor  ( new_n24262_, new_n24261_, new_n403_ );
nor  ( new_n24263_, new_n24262_, new_n24258_ );
and  ( new_n24264_, new_n24262_, new_n24258_ );
or   ( new_n24265_, new_n409_, new_n22829_ );
or   ( new_n24266_, new_n411_, new_n22641_ );
and  ( new_n24267_, new_n24266_, new_n24265_ );
xor  ( new_n24268_, new_n24267_, new_n328_ );
nor  ( new_n24269_, new_n24268_, new_n24264_ );
nor  ( new_n24270_, new_n24269_, new_n24263_ );
nor  ( new_n24271_, new_n24270_, new_n24254_ );
nor  ( new_n24272_, new_n24271_, new_n24253_ );
not  ( new_n24273_, new_n24272_ );
or   ( new_n24274_, new_n24273_, new_n24222_ );
and  ( new_n24275_, new_n24273_, new_n24222_ );
xnor ( new_n24276_, new_n24010_, new_n24005_ );
xor  ( new_n24277_, new_n24276_, new_n24012_ );
xnor ( new_n24278_, new_n24023_, new_n24019_ );
xor  ( new_n24279_, new_n24278_, new_n24029_ );
or   ( new_n24280_, new_n24279_, new_n24277_ );
and  ( new_n24281_, new_n24279_, new_n24277_ );
xnor ( new_n24282_, new_n24041_, new_n24037_ );
xor  ( new_n24283_, new_n24282_, new_n24047_ );
or   ( new_n24284_, new_n24283_, new_n24281_ );
and  ( new_n24285_, new_n24284_, new_n24280_ );
or   ( new_n24286_, new_n24285_, new_n24275_ );
and  ( new_n24287_, new_n24286_, new_n24274_ );
nor  ( new_n24288_, new_n24287_, new_n24172_ );
nand ( new_n24289_, new_n24287_, new_n24172_ );
xor  ( new_n24290_, new_n24118_, new_n24116_ );
xor  ( new_n24291_, new_n24290_, new_n24122_ );
xnor ( new_n24292_, new_n24071_, new_n24067_ );
xor  ( new_n24293_, new_n24292_, new_n24077_ );
xnor ( new_n24294_, new_n24089_, new_n24085_ );
xor  ( new_n24295_, new_n24294_, new_n24095_ );
or   ( new_n24296_, new_n24295_, new_n24293_ );
and  ( new_n24297_, new_n24295_, new_n24293_ );
xor  ( new_n24298_, new_n24055_, new_n2799_ );
xor  ( new_n24299_, new_n24298_, new_n24061_ );
or   ( new_n24300_, new_n24299_, new_n24297_ );
and  ( new_n24301_, new_n24300_, new_n24296_ );
nor  ( new_n24302_, new_n24301_, new_n24291_ );
nand ( new_n24303_, new_n24301_, new_n24291_ );
xnor ( new_n24304_, new_n24105_, new_n24103_ );
xor  ( new_n24305_, new_n24304_, new_n24108_ );
and  ( new_n24306_, new_n24305_, new_n24303_ );
or   ( new_n24307_, new_n24306_, new_n24302_ );
and  ( new_n24308_, new_n24307_, new_n24289_ );
or   ( new_n24309_, new_n24308_, new_n24288_ );
and  ( new_n24310_, new_n24309_, new_n24167_ );
or   ( new_n24311_, new_n24310_, new_n24166_ );
xnor ( new_n24312_, new_n23951_, new_n23844_ );
xor  ( new_n24313_, new_n24312_, new_n23971_ );
nand ( new_n24314_, new_n24313_, new_n24311_ );
nor  ( new_n24315_, new_n24313_, new_n24311_ );
xor  ( new_n24316_, new_n24139_, new_n24001_ );
xor  ( new_n24317_, new_n24316_, new_n24143_ );
or   ( new_n24318_, new_n24317_, new_n24315_ );
and  ( new_n24319_, new_n24318_, new_n24314_ );
xor  ( new_n24320_, new_n24145_, new_n23992_ );
xor  ( new_n24321_, new_n24320_, new_n24149_ );
nor  ( new_n24322_, new_n24321_, new_n24319_ );
xor  ( new_n24323_, new_n24151_, new_n23990_ );
and  ( new_n24324_, new_n24323_, new_n24322_ );
xnor ( new_n24325_, new_n24313_, new_n24311_ );
xor  ( new_n24326_, new_n24325_, new_n24317_ );
xor  ( new_n24327_, new_n24165_, new_n24156_ );
xor  ( new_n24328_, new_n24327_, new_n24309_ );
xor  ( new_n24329_, new_n24272_, new_n24222_ );
xor  ( new_n24330_, new_n24329_, new_n24285_ );
xor  ( new_n24331_, new_n24301_, new_n24291_ );
xor  ( new_n24332_, new_n24331_, new_n24305_ );
or   ( new_n24333_, new_n24332_, new_n24330_ );
and  ( new_n24334_, new_n24332_, new_n24330_ );
xor  ( new_n24335_, new_n24171_, new_n24169_ );
or   ( new_n24336_, new_n24335_, new_n24334_ );
and  ( new_n24337_, new_n24336_, new_n24333_ );
xor  ( new_n24338_, new_n24231_, new_n24226_ );
xnor ( new_n24339_, new_n24338_, new_n24233_ );
xnor ( new_n24340_, new_n24244_, new_n24240_ );
xor  ( new_n24341_, new_n24340_, new_n24250_ );
nand ( new_n24342_, new_n24341_, new_n24339_ );
or   ( new_n24343_, new_n1593_, new_n21792_ );
or   ( new_n24344_, new_n1595_, new_n21751_ );
and  ( new_n24345_, new_n24344_, new_n24343_ );
xor  ( new_n24346_, new_n24345_, new_n1358_ );
or   ( new_n24347_, new_n1364_, new_n21840_ );
or   ( new_n24348_, new_n1366_, new_n21842_ );
and  ( new_n24349_, new_n24348_, new_n24347_ );
xor  ( new_n24350_, new_n24349_, new_n1129_ );
nor  ( new_n24351_, new_n24350_, new_n24346_ );
or   ( new_n24352_, new_n1135_, new_n22098_ );
or   ( new_n24353_, new_n1137_, new_n21847_ );
and  ( new_n24354_, new_n24353_, new_n24352_ );
xor  ( new_n24355_, new_n24354_, new_n895_ );
nand ( new_n24356_, new_n24350_, new_n24346_ );
and  ( new_n24357_, new_n24356_, new_n24355_ );
or   ( new_n24358_, new_n24357_, new_n24351_ );
or   ( new_n24359_, new_n3117_, new_n21694_ );
or   ( new_n24360_, new_n3119_, new_n21696_ );
and  ( new_n24361_, new_n24360_, new_n24359_ );
xor  ( new_n24362_, new_n24361_, new_n2800_ );
nand ( new_n24363_, new_n24362_, new_n3116_ );
or   ( new_n24364_, new_n2807_, new_n21701_ );
or   ( new_n24365_, new_n2809_, new_n21703_ );
and  ( new_n24366_, new_n24365_, new_n24364_ );
xor  ( new_n24367_, new_n24366_, new_n2423_ );
nor  ( new_n24368_, new_n24362_, new_n3116_ );
or   ( new_n24369_, new_n24368_, new_n24367_ );
and  ( new_n24370_, new_n24369_, new_n24363_ );
nand ( new_n24371_, new_n24370_, new_n24358_ );
nor  ( new_n24372_, new_n24370_, new_n24358_ );
or   ( new_n24373_, new_n2425_, new_n21672_ );
or   ( new_n24374_, new_n2427_, new_n21674_ );
and  ( new_n24375_, new_n24374_, new_n24373_ );
xor  ( new_n24376_, new_n24375_, new_n2121_ );
or   ( new_n24377_, new_n2122_, new_n21678_ );
or   ( new_n24378_, new_n2124_, new_n21680_ );
and  ( new_n24379_, new_n24378_, new_n24377_ );
xor  ( new_n24380_, new_n24379_, new_n1843_ );
nor  ( new_n24381_, new_n24380_, new_n24376_ );
or   ( new_n24382_, new_n1844_, new_n21685_ );
or   ( new_n24383_, new_n1846_, new_n21687_ );
and  ( new_n24384_, new_n24383_, new_n24382_ );
xor  ( new_n24385_, new_n24384_, new_n1586_ );
and  ( new_n24386_, new_n24380_, new_n24376_ );
nor  ( new_n24387_, new_n24386_, new_n24385_ );
nor  ( new_n24388_, new_n24387_, new_n24381_ );
or   ( new_n24389_, new_n24388_, new_n24372_ );
and  ( new_n24390_, new_n24389_, new_n24371_ );
nor  ( new_n24391_, new_n24390_, new_n24342_ );
nand ( new_n24392_, new_n24390_, new_n24342_ );
or   ( new_n24393_, new_n897_, new_n22207_ );
or   ( new_n24394_, new_n899_, new_n22129_ );
and  ( new_n24395_, new_n24394_, new_n24393_ );
xor  ( new_n24396_, new_n24395_, new_n748_ );
or   ( new_n24397_, new_n755_, new_n22423_ );
or   ( new_n24398_, new_n757_, new_n22304_ );
and  ( new_n24399_, new_n24398_, new_n24397_ );
xor  ( new_n24400_, new_n24399_, new_n523_ );
or   ( new_n24401_, new_n24400_, new_n24396_ );
or   ( new_n24402_, new_n524_, new_n22641_ );
or   ( new_n24403_, new_n526_, new_n22590_ );
and  ( new_n24404_, new_n24403_, new_n24402_ );
xor  ( new_n24405_, new_n24404_, new_n403_ );
and  ( new_n24406_, new_n24400_, new_n24396_ );
or   ( new_n24407_, new_n24406_, new_n24405_ );
and  ( new_n24408_, new_n24407_, new_n24401_ );
or   ( new_n24409_, new_n283_, new_n23733_ );
or   ( new_n24410_, new_n286_, new_n23554_ );
and  ( new_n24411_, new_n24410_, new_n24409_ );
xor  ( new_n24412_, new_n24411_, new_n278_ );
or   ( new_n24413_, new_n299_, new_n24006_ );
or   ( new_n24414_, new_n302_, new_n23895_ );
and  ( new_n24415_, new_n24414_, new_n24413_ );
xor  ( new_n24416_, new_n24415_, new_n293_ );
or   ( new_n24417_, new_n24416_, new_n24412_ );
not  ( new_n24418_, RIbb32568_162 );
or   ( new_n24419_, new_n268_, new_n24418_ );
or   ( new_n24420_, new_n271_, new_n24227_ );
and  ( new_n24421_, new_n24420_, new_n24419_ );
xor  ( new_n24422_, new_n24421_, new_n263_ );
and  ( new_n24423_, new_n24416_, new_n24412_ );
or   ( new_n24424_, new_n24423_, new_n24422_ );
and  ( new_n24425_, new_n24424_, new_n24417_ );
nor  ( new_n24426_, new_n24425_, new_n24408_ );
nand ( new_n24427_, new_n24425_, new_n24408_ );
or   ( new_n24428_, new_n409_, new_n22975_ );
or   ( new_n24429_, new_n411_, new_n22829_ );
and  ( new_n24430_, new_n24429_, new_n24428_ );
xor  ( new_n24431_, new_n24430_, new_n328_ );
or   ( new_n24432_, new_n337_, new_n23166_ );
or   ( new_n24433_, new_n340_, new_n22973_ );
and  ( new_n24434_, new_n24433_, new_n24432_ );
xor  ( new_n24435_, new_n24434_, new_n332_ );
nor  ( new_n24436_, new_n24435_, new_n24431_ );
or   ( new_n24437_, new_n317_, new_n23370_ );
or   ( new_n24438_, new_n320_, new_n23252_ );
and  ( new_n24439_, new_n24438_, new_n24437_ );
xor  ( new_n24440_, new_n24439_, new_n312_ );
not  ( new_n24441_, new_n24440_ );
nand ( new_n24442_, new_n24435_, new_n24431_ );
and  ( new_n24443_, new_n24442_, new_n24441_ );
or   ( new_n24444_, new_n24443_, new_n24436_ );
and  ( new_n24445_, new_n24444_, new_n24427_ );
or   ( new_n24446_, new_n24445_, new_n24426_ );
and  ( new_n24447_, new_n24446_, new_n24392_ );
or   ( new_n24448_, new_n24447_, new_n24391_ );
xor  ( new_n24449_, new_n24279_, new_n24277_ );
xor  ( new_n24450_, new_n24449_, new_n24283_ );
xnor ( new_n24451_, new_n24194_, new_n24190_ );
xor  ( new_n24452_, new_n24451_, new_n24200_ );
xor  ( new_n24453_, new_n24212_, new_n24208_ );
xor  ( new_n24454_, new_n24453_, new_n24218_ );
or   ( new_n24455_, new_n24454_, new_n24452_ );
and  ( new_n24456_, new_n24454_, new_n24452_ );
xnor ( new_n24457_, new_n24262_, new_n24258_ );
xor  ( new_n24458_, new_n24457_, new_n24268_ );
or   ( new_n24459_, new_n24458_, new_n24456_ );
and  ( new_n24460_, new_n24459_, new_n24455_ );
or   ( new_n24461_, new_n24460_, new_n24450_ );
and  ( new_n24462_, new_n24460_, new_n24450_ );
xor  ( new_n24463_, new_n24295_, new_n24293_ );
xor  ( new_n24464_, new_n24463_, new_n24299_ );
or   ( new_n24465_, new_n24464_, new_n24462_ );
and  ( new_n24466_, new_n24465_, new_n24461_ );
nand ( new_n24467_, new_n24466_, new_n24448_ );
nor  ( new_n24468_, new_n24466_, new_n24448_ );
xor  ( new_n24469_, new_n24252_, new_n24236_ );
xnor ( new_n24470_, new_n24469_, new_n24270_ );
xor  ( new_n24471_, new_n24202_, new_n24186_ );
xor  ( new_n24472_, new_n24471_, new_n24220_ );
nor  ( new_n24473_, new_n24472_, new_n24470_ );
or   ( new_n24474_, new_n24473_, new_n24468_ );
and  ( new_n24475_, new_n24474_, new_n24467_ );
or   ( new_n24476_, new_n24475_, new_n24337_ );
and  ( new_n24477_, new_n24475_, new_n24337_ );
xor  ( new_n24478_, new_n24160_, new_n24158_ );
xor  ( new_n24479_, new_n24478_, new_n24163_ );
or   ( new_n24480_, new_n24479_, new_n24477_ );
and  ( new_n24481_, new_n24480_, new_n24476_ );
or   ( new_n24482_, new_n24481_, new_n24328_ );
nand ( new_n24483_, new_n24481_, new_n24328_ );
xor  ( new_n24484_, new_n24130_, new_n24112_ );
xnor ( new_n24485_, new_n24484_, new_n24137_ );
nand ( new_n24486_, new_n24485_, new_n24483_ );
and  ( new_n24487_, new_n24486_, new_n24482_ );
and  ( new_n24488_, new_n24487_, new_n24326_ );
xor  ( new_n24489_, new_n24321_, new_n24319_ );
and  ( new_n24490_, new_n24489_, new_n24488_ );
xor  ( new_n24491_, new_n24332_, new_n24330_ );
xor  ( new_n24492_, new_n24491_, new_n24335_ );
or   ( new_n24493_, new_n2425_, new_n21680_ );
or   ( new_n24494_, new_n2427_, new_n21672_ );
and  ( new_n24495_, new_n24494_, new_n24493_ );
xor  ( new_n24496_, new_n24495_, new_n2121_ );
or   ( new_n24497_, new_n2122_, new_n21687_ );
or   ( new_n24498_, new_n2124_, new_n21678_ );
and  ( new_n24499_, new_n24498_, new_n24497_ );
xor  ( new_n24500_, new_n24499_, new_n1843_ );
or   ( new_n24501_, new_n24500_, new_n24496_ );
or   ( new_n24502_, new_n1844_, new_n21751_ );
or   ( new_n24503_, new_n1846_, new_n21685_ );
and  ( new_n24504_, new_n24503_, new_n24502_ );
xor  ( new_n24505_, new_n24504_, new_n1586_ );
and  ( new_n24506_, new_n24500_, new_n24496_ );
or   ( new_n24507_, new_n24506_, new_n24505_ );
and  ( new_n24508_, new_n24507_, new_n24501_ );
or   ( new_n24509_, new_n1593_, new_n21842_ );
or   ( new_n24510_, new_n1595_, new_n21792_ );
and  ( new_n24511_, new_n24510_, new_n24509_ );
xor  ( new_n24512_, new_n24511_, new_n1358_ );
or   ( new_n24513_, new_n1364_, new_n21847_ );
or   ( new_n24514_, new_n1366_, new_n21840_ );
and  ( new_n24515_, new_n24514_, new_n24513_ );
xor  ( new_n24516_, new_n24515_, new_n1129_ );
or   ( new_n24517_, new_n24516_, new_n24512_ );
or   ( new_n24518_, new_n1135_, new_n22129_ );
or   ( new_n24519_, new_n1137_, new_n22098_ );
and  ( new_n24520_, new_n24519_, new_n24518_ );
xor  ( new_n24521_, new_n24520_, new_n896_ );
and  ( new_n24522_, new_n24516_, new_n24512_ );
or   ( new_n24523_, new_n24522_, new_n24521_ );
and  ( new_n24524_, new_n24523_, new_n24517_ );
or   ( new_n24525_, new_n24524_, new_n24508_ );
and  ( new_n24526_, new_n24524_, new_n24508_ );
or   ( new_n24527_, new_n3117_, new_n21703_ );
or   ( new_n24528_, new_n3119_, new_n21694_ );
and  ( new_n24529_, new_n24528_, new_n24527_ );
xor  ( new_n24530_, new_n24529_, new_n2799_ );
and  ( new_n24531_, new_n3293_, RIbb315f0_129 );
xor  ( new_n24532_, new_n24531_, new_n3116_ );
and  ( new_n24533_, new_n24532_, new_n24530_ );
or   ( new_n24534_, new_n2807_, new_n21674_ );
or   ( new_n24535_, new_n2809_, new_n21701_ );
and  ( new_n24536_, new_n24535_, new_n24534_ );
xor  ( new_n24537_, new_n24536_, new_n2424_ );
nor  ( new_n24538_, new_n24532_, new_n24530_ );
nor  ( new_n24539_, new_n24538_, new_n24537_ );
nor  ( new_n24540_, new_n24539_, new_n24533_ );
or   ( new_n24541_, new_n24540_, new_n24526_ );
and  ( new_n24542_, new_n24541_, new_n24525_ );
not  ( new_n24543_, RIbb325e0_163 );
or   ( new_n24544_, new_n24543_, new_n260_ );
xnor ( new_n24545_, new_n24416_, new_n24412_ );
xor  ( new_n24546_, new_n24545_, new_n24422_ );
nand ( new_n24547_, new_n24546_, new_n24544_ );
or   ( new_n24548_, new_n24546_, new_n24544_ );
xor  ( new_n24549_, new_n24435_, new_n24431_ );
xor  ( new_n24550_, new_n24549_, new_n24441_ );
nand ( new_n24551_, new_n24550_, new_n24548_ );
and  ( new_n24552_, new_n24551_, new_n24547_ );
nor  ( new_n24553_, new_n24552_, new_n24542_ );
nand ( new_n24554_, new_n24552_, new_n24542_ );
or   ( new_n24555_, new_n283_, new_n23895_ );
or   ( new_n24556_, new_n286_, new_n23733_ );
and  ( new_n24557_, new_n24556_, new_n24555_ );
xor  ( new_n24558_, new_n24557_, new_n278_ );
or   ( new_n24559_, new_n299_, new_n24227_ );
or   ( new_n24560_, new_n302_, new_n24006_ );
and  ( new_n24561_, new_n24560_, new_n24559_ );
xor  ( new_n24562_, new_n24561_, new_n293_ );
or   ( new_n24563_, new_n24562_, new_n24558_ );
or   ( new_n24564_, new_n268_, new_n24543_ );
or   ( new_n24565_, new_n271_, new_n24418_ );
and  ( new_n24566_, new_n24565_, new_n24564_ );
xor  ( new_n24567_, new_n24566_, new_n263_ );
and  ( new_n24568_, new_n24562_, new_n24558_ );
or   ( new_n24569_, new_n24568_, new_n24567_ );
and  ( new_n24570_, new_n24569_, new_n24563_ );
or   ( new_n24571_, new_n897_, new_n22304_ );
or   ( new_n24572_, new_n899_, new_n22207_ );
and  ( new_n24573_, new_n24572_, new_n24571_ );
xor  ( new_n24574_, new_n24573_, new_n748_ );
or   ( new_n24575_, new_n755_, new_n22590_ );
or   ( new_n24576_, new_n757_, new_n22423_ );
and  ( new_n24577_, new_n24576_, new_n24575_ );
xor  ( new_n24578_, new_n24577_, new_n523_ );
or   ( new_n24579_, new_n24578_, new_n24574_ );
or   ( new_n24580_, new_n524_, new_n22829_ );
or   ( new_n24581_, new_n526_, new_n22641_ );
and  ( new_n24582_, new_n24581_, new_n24580_ );
xor  ( new_n24583_, new_n24582_, new_n403_ );
and  ( new_n24584_, new_n24578_, new_n24574_ );
or   ( new_n24585_, new_n24584_, new_n24583_ );
and  ( new_n24586_, new_n24585_, new_n24579_ );
nor  ( new_n24587_, new_n24586_, new_n24570_ );
nand ( new_n24588_, new_n24586_, new_n24570_ );
or   ( new_n24589_, new_n409_, new_n22973_ );
or   ( new_n24590_, new_n411_, new_n22975_ );
and  ( new_n24591_, new_n24590_, new_n24589_ );
xor  ( new_n24592_, new_n24591_, new_n328_ );
or   ( new_n24593_, new_n337_, new_n23252_ );
or   ( new_n24594_, new_n340_, new_n23166_ );
and  ( new_n24595_, new_n24594_, new_n24593_ );
xor  ( new_n24596_, new_n24595_, new_n332_ );
nor  ( new_n24597_, new_n24596_, new_n24592_ );
or   ( new_n24598_, new_n317_, new_n23554_ );
or   ( new_n24599_, new_n320_, new_n23370_ );
and  ( new_n24600_, new_n24599_, new_n24598_ );
xor  ( new_n24601_, new_n24600_, new_n312_ );
not  ( new_n24602_, new_n24601_ );
nand ( new_n24603_, new_n24596_, new_n24592_ );
and  ( new_n24604_, new_n24603_, new_n24602_ );
or   ( new_n24605_, new_n24604_, new_n24597_ );
and  ( new_n24606_, new_n24605_, new_n24588_ );
or   ( new_n24607_, new_n24606_, new_n24587_ );
and  ( new_n24608_, new_n24607_, new_n24554_ );
or   ( new_n24609_, new_n24608_, new_n24553_ );
xnor ( new_n24610_, new_n24178_, new_n24176_ );
xor  ( new_n24611_, new_n24610_, new_n24184_ );
xor  ( new_n24612_, new_n24350_, new_n24346_ );
xor  ( new_n24613_, new_n24612_, new_n24355_ );
xnor ( new_n24614_, new_n24400_, new_n24396_ );
xor  ( new_n24615_, new_n24614_, new_n24405_ );
or   ( new_n24616_, new_n24615_, new_n24613_ );
and  ( new_n24617_, new_n24615_, new_n24613_ );
xor  ( new_n24618_, new_n24380_, new_n24376_ );
xnor ( new_n24619_, new_n24618_, new_n24385_ );
or   ( new_n24620_, new_n24619_, new_n24617_ );
and  ( new_n24621_, new_n24620_, new_n24616_ );
or   ( new_n24622_, new_n24621_, new_n24611_ );
and  ( new_n24623_, new_n24621_, new_n24611_ );
xor  ( new_n24624_, new_n24454_, new_n24452_ );
xor  ( new_n24625_, new_n24624_, new_n24458_ );
or   ( new_n24626_, new_n24625_, new_n24623_ );
and  ( new_n24627_, new_n24626_, new_n24622_ );
nand ( new_n24628_, new_n24627_, new_n24609_ );
or   ( new_n24629_, new_n24627_, new_n24609_ );
xnor ( new_n24630_, new_n24370_, new_n24358_ );
xor  ( new_n24631_, new_n24630_, new_n24388_ );
xor  ( new_n24632_, new_n24425_, new_n24408_ );
xor  ( new_n24633_, new_n24632_, new_n24444_ );
nor  ( new_n24634_, new_n24633_, new_n24631_ );
and  ( new_n24635_, new_n24633_, new_n24631_ );
xor  ( new_n24636_, new_n24341_, new_n24339_ );
nor  ( new_n24637_, new_n24636_, new_n24635_ );
nor  ( new_n24638_, new_n24637_, new_n24634_ );
nand ( new_n24639_, new_n24638_, new_n24629_ );
and  ( new_n24640_, new_n24639_, new_n24628_ );
or   ( new_n24641_, new_n24640_, new_n24492_ );
nand ( new_n24642_, new_n24640_, new_n24492_ );
xor  ( new_n24643_, new_n24460_, new_n24450_ );
xor  ( new_n24644_, new_n24643_, new_n24464_ );
xor  ( new_n24645_, new_n24390_, new_n24342_ );
xor  ( new_n24646_, new_n24645_, new_n24446_ );
nor  ( new_n24647_, new_n24646_, new_n24644_ );
and  ( new_n24648_, new_n24646_, new_n24644_ );
not  ( new_n24649_, new_n24648_ );
xor  ( new_n24650_, new_n24472_, new_n24470_ );
and  ( new_n24651_, new_n24650_, new_n24649_ );
nor  ( new_n24652_, new_n24651_, new_n24647_ );
nand ( new_n24653_, new_n24652_, new_n24642_ );
and  ( new_n24654_, new_n24653_, new_n24641_ );
xor  ( new_n24655_, new_n24287_, new_n24172_ );
xor  ( new_n24656_, new_n24655_, new_n24307_ );
nand ( new_n24657_, new_n24656_, new_n24654_ );
nor  ( new_n24658_, new_n24656_, new_n24654_ );
xnor ( new_n24659_, new_n24475_, new_n24337_ );
xor  ( new_n24660_, new_n24659_, new_n24479_ );
or   ( new_n24661_, new_n24660_, new_n24658_ );
and  ( new_n24662_, new_n24661_, new_n24657_ );
xor  ( new_n24663_, new_n24481_, new_n24328_ );
xor  ( new_n24664_, new_n24663_, new_n24485_ );
nor  ( new_n24665_, new_n24664_, new_n24662_ );
xor  ( new_n24666_, new_n24487_, new_n24326_ );
and  ( new_n24667_, new_n24666_, new_n24665_ );
xor  ( new_n24668_, new_n24656_, new_n24654_ );
xor  ( new_n24669_, new_n24668_, new_n24660_ );
xor  ( new_n24670_, new_n24362_, new_n3116_ );
xor  ( new_n24671_, new_n24670_, new_n24367_ );
xnor ( new_n24672_, new_n24516_, new_n24512_ );
xor  ( new_n24673_, new_n24672_, new_n24521_ );
xnor ( new_n24674_, new_n24578_, new_n24574_ );
xor  ( new_n24675_, new_n24674_, new_n24583_ );
or   ( new_n24676_, new_n24675_, new_n24673_ );
and  ( new_n24677_, new_n24675_, new_n24673_ );
xor  ( new_n24678_, new_n24596_, new_n24592_ );
xor  ( new_n24679_, new_n24678_, new_n24602_ );
or   ( new_n24680_, new_n24679_, new_n24677_ );
and  ( new_n24681_, new_n24680_, new_n24676_ );
nor  ( new_n24682_, new_n24681_, new_n24671_ );
and  ( new_n24683_, new_n24681_, new_n24671_ );
xor  ( new_n24684_, new_n24615_, new_n24613_ );
xnor ( new_n24685_, new_n24684_, new_n24619_ );
not  ( new_n24686_, new_n24685_ );
nor  ( new_n24687_, new_n24686_, new_n24683_ );
nor  ( new_n24688_, new_n24687_, new_n24682_ );
and  ( new_n24689_, RIbb32658_164, RIbb2f610_1 );
not  ( new_n24690_, new_n24689_ );
xnor ( new_n24691_, new_n24562_, new_n24558_ );
xor  ( new_n24692_, new_n24691_, new_n24567_ );
nand ( new_n24693_, new_n24692_, new_n24690_ );
or   ( new_n24694_, new_n3461_, new_n21694_ );
or   ( new_n24695_, new_n3463_, new_n21696_ );
and  ( new_n24696_, new_n24695_, new_n24694_ );
xor  ( new_n24697_, new_n24696_, new_n3116_ );
and  ( new_n24698_, new_n24697_, new_n3460_ );
or   ( new_n24699_, new_n3117_, new_n21701_ );
or   ( new_n24700_, new_n3119_, new_n21703_ );
and  ( new_n24701_, new_n24700_, new_n24699_ );
xor  ( new_n24702_, new_n24701_, new_n2800_ );
or   ( new_n24703_, new_n24697_, new_n3460_ );
and  ( new_n24704_, new_n24703_, new_n24702_ );
or   ( new_n24705_, new_n24704_, new_n24698_ );
or   ( new_n24706_, new_n2807_, new_n21672_ );
or   ( new_n24707_, new_n2809_, new_n21674_ );
and  ( new_n24708_, new_n24707_, new_n24706_ );
xor  ( new_n24709_, new_n24708_, new_n2424_ );
or   ( new_n24710_, new_n2425_, new_n21678_ );
or   ( new_n24711_, new_n2427_, new_n21680_ );
and  ( new_n24712_, new_n24711_, new_n24710_ );
xor  ( new_n24713_, new_n24712_, new_n2121_ );
or   ( new_n24714_, new_n24713_, new_n24709_ );
or   ( new_n24715_, new_n2122_, new_n21685_ );
or   ( new_n24716_, new_n2124_, new_n21687_ );
and  ( new_n24717_, new_n24716_, new_n24715_ );
xor  ( new_n24718_, new_n24717_, new_n1843_ );
and  ( new_n24719_, new_n24713_, new_n24709_ );
or   ( new_n24720_, new_n24719_, new_n24718_ );
and  ( new_n24721_, new_n24720_, new_n24714_ );
or   ( new_n24722_, new_n24721_, new_n24705_ );
and  ( new_n24723_, new_n24721_, new_n24705_ );
or   ( new_n24724_, new_n1844_, new_n21792_ );
or   ( new_n24725_, new_n1846_, new_n21751_ );
and  ( new_n24726_, new_n24725_, new_n24724_ );
xor  ( new_n24727_, new_n24726_, new_n1586_ );
or   ( new_n24728_, new_n1593_, new_n21840_ );
or   ( new_n24729_, new_n1595_, new_n21842_ );
and  ( new_n24730_, new_n24729_, new_n24728_ );
xor  ( new_n24731_, new_n24730_, new_n1358_ );
nor  ( new_n24732_, new_n24731_, new_n24727_ );
or   ( new_n24733_, new_n1364_, new_n22098_ );
or   ( new_n24734_, new_n1366_, new_n21847_ );
and  ( new_n24735_, new_n24734_, new_n24733_ );
xor  ( new_n24736_, new_n24735_, new_n1129_ );
and  ( new_n24737_, new_n24731_, new_n24727_ );
nor  ( new_n24738_, new_n24737_, new_n24736_ );
nor  ( new_n24739_, new_n24738_, new_n24732_ );
or   ( new_n24740_, new_n24739_, new_n24723_ );
and  ( new_n24741_, new_n24740_, new_n24722_ );
and  ( new_n24742_, new_n24741_, new_n24693_ );
or   ( new_n24743_, new_n1135_, new_n22207_ );
or   ( new_n24744_, new_n1137_, new_n22129_ );
and  ( new_n24745_, new_n24744_, new_n24743_ );
xor  ( new_n24746_, new_n24745_, new_n896_ );
or   ( new_n24747_, new_n897_, new_n22423_ );
or   ( new_n24748_, new_n899_, new_n22304_ );
and  ( new_n24749_, new_n24748_, new_n24747_ );
xor  ( new_n24750_, new_n24749_, new_n748_ );
or   ( new_n24751_, new_n24750_, new_n24746_ );
or   ( new_n24752_, new_n755_, new_n22641_ );
or   ( new_n24753_, new_n757_, new_n22590_ );
and  ( new_n24754_, new_n24753_, new_n24752_ );
xor  ( new_n24755_, new_n24754_, new_n523_ );
and  ( new_n24756_, new_n24750_, new_n24746_ );
or   ( new_n24757_, new_n24756_, new_n24755_ );
and  ( new_n24758_, new_n24757_, new_n24751_ );
or   ( new_n24759_, new_n524_, new_n22975_ );
or   ( new_n24760_, new_n526_, new_n22829_ );
and  ( new_n24761_, new_n24760_, new_n24759_ );
xor  ( new_n24762_, new_n24761_, new_n403_ );
or   ( new_n24763_, new_n409_, new_n23166_ );
or   ( new_n24764_, new_n411_, new_n22973_ );
and  ( new_n24765_, new_n24764_, new_n24763_ );
xor  ( new_n24766_, new_n24765_, new_n328_ );
or   ( new_n24767_, new_n24766_, new_n24762_ );
or   ( new_n24768_, new_n337_, new_n23370_ );
or   ( new_n24769_, new_n340_, new_n23252_ );
and  ( new_n24770_, new_n24769_, new_n24768_ );
xor  ( new_n24771_, new_n24770_, new_n332_ );
and  ( new_n24772_, new_n24766_, new_n24762_ );
or   ( new_n24773_, new_n24772_, new_n24771_ );
and  ( new_n24774_, new_n24773_, new_n24767_ );
nor  ( new_n24775_, new_n24774_, new_n24758_ );
and  ( new_n24776_, new_n24774_, new_n24758_ );
or   ( new_n24777_, new_n317_, new_n23733_ );
or   ( new_n24778_, new_n320_, new_n23554_ );
and  ( new_n24779_, new_n24778_, new_n24777_ );
xor  ( new_n24780_, new_n24779_, new_n312_ );
or   ( new_n24781_, new_n283_, new_n24006_ );
or   ( new_n24782_, new_n286_, new_n23895_ );
and  ( new_n24783_, new_n24782_, new_n24781_ );
xor  ( new_n24784_, new_n24783_, new_n278_ );
nor  ( new_n24785_, new_n24784_, new_n24780_ );
or   ( new_n24786_, new_n299_, new_n24418_ );
or   ( new_n24787_, new_n302_, new_n24227_ );
and  ( new_n24788_, new_n24787_, new_n24786_ );
xor  ( new_n24789_, new_n24788_, new_n293_ );
and  ( new_n24790_, new_n24784_, new_n24780_ );
nor  ( new_n24791_, new_n24790_, new_n24789_ );
nor  ( new_n24792_, new_n24791_, new_n24785_ );
nor  ( new_n24793_, new_n24792_, new_n24776_ );
nor  ( new_n24794_, new_n24793_, new_n24775_ );
not  ( new_n24795_, new_n24794_ );
nor  ( new_n24796_, new_n24741_, new_n24693_ );
nor  ( new_n24797_, new_n24796_, new_n24795_ );
nor  ( new_n24798_, new_n24797_, new_n24742_ );
and  ( new_n24799_, new_n24798_, new_n24688_ );
not  ( new_n24800_, new_n24799_ );
xnor ( new_n24801_, new_n24524_, new_n24508_ );
xor  ( new_n24802_, new_n24801_, new_n24540_ );
xor  ( new_n24803_, new_n24586_, new_n24570_ );
xor  ( new_n24804_, new_n24803_, new_n24605_ );
nor  ( new_n24805_, new_n24804_, new_n24802_ );
and  ( new_n24806_, new_n24804_, new_n24802_ );
xor  ( new_n24807_, new_n24546_, new_n24544_ );
xor  ( new_n24808_, new_n24807_, new_n24550_ );
nor  ( new_n24809_, new_n24808_, new_n24806_ );
nor  ( new_n24810_, new_n24809_, new_n24805_ );
not  ( new_n24811_, new_n24810_ );
and  ( new_n24812_, new_n24811_, new_n24800_ );
nor  ( new_n24813_, new_n24798_, new_n24688_ );
or   ( new_n24814_, new_n24813_, new_n24812_ );
xor  ( new_n24815_, new_n24646_, new_n24644_ );
xor  ( new_n24816_, new_n24815_, new_n24650_ );
nor  ( new_n24817_, new_n24816_, new_n24814_ );
nand ( new_n24818_, new_n24816_, new_n24814_ );
xor  ( new_n24819_, new_n24621_, new_n24611_ );
xor  ( new_n24820_, new_n24819_, new_n24625_ );
xor  ( new_n24821_, new_n24552_, new_n24542_ );
xor  ( new_n24822_, new_n24821_, new_n24607_ );
or   ( new_n24823_, new_n24822_, new_n24820_ );
and  ( new_n24824_, new_n24822_, new_n24820_ );
xor  ( new_n24825_, new_n24633_, new_n24631_ );
xor  ( new_n24826_, new_n24825_, new_n24636_ );
or   ( new_n24827_, new_n24826_, new_n24824_ );
and  ( new_n24828_, new_n24827_, new_n24823_ );
and  ( new_n24829_, new_n24828_, new_n24818_ );
or   ( new_n24830_, new_n24829_, new_n24817_ );
xnor ( new_n24831_, new_n24466_, new_n24448_ );
xor  ( new_n24832_, new_n24831_, new_n24473_ );
or   ( new_n24833_, new_n24832_, new_n24830_ );
and  ( new_n24834_, new_n24832_, new_n24830_ );
xor  ( new_n24835_, new_n24640_, new_n24492_ );
xor  ( new_n24836_, new_n24835_, new_n24652_ );
or   ( new_n24837_, new_n24836_, new_n24834_ );
and  ( new_n24838_, new_n24837_, new_n24833_ );
nor  ( new_n24839_, new_n24838_, new_n24669_ );
xor  ( new_n24840_, new_n24664_, new_n24662_ );
and  ( new_n24841_, new_n24840_, new_n24839_ );
xor  ( new_n24842_, new_n24832_, new_n24830_ );
xor  ( new_n24843_, new_n24842_, new_n24836_ );
xnor ( new_n24844_, new_n24822_, new_n24820_ );
xor  ( new_n24845_, new_n24844_, new_n24826_ );
xnor ( new_n24846_, new_n24500_, new_n24496_ );
xor  ( new_n24847_, new_n24846_, new_n24505_ );
xor  ( new_n24848_, new_n24697_, new_n3459_ );
xor  ( new_n24849_, new_n24848_, new_n24702_ );
xnor ( new_n24850_, new_n24713_, new_n24709_ );
xor  ( new_n24851_, new_n24850_, new_n24718_ );
or   ( new_n24852_, new_n24851_, new_n24849_ );
and  ( new_n24853_, new_n24851_, new_n24849_ );
xnor ( new_n24854_, new_n24731_, new_n24727_ );
xor  ( new_n24855_, new_n24854_, new_n24736_ );
or   ( new_n24856_, new_n24855_, new_n24853_ );
and  ( new_n24857_, new_n24856_, new_n24852_ );
nor  ( new_n24858_, new_n24857_, new_n24847_ );
nand ( new_n24859_, new_n24857_, new_n24847_ );
xnor ( new_n24860_, new_n24766_, new_n24762_ );
xor  ( new_n24861_, new_n24860_, new_n24771_ );
xnor ( new_n24862_, new_n24750_, new_n24746_ );
xor  ( new_n24863_, new_n24862_, new_n24755_ );
nor  ( new_n24864_, new_n24863_, new_n24861_ );
and  ( new_n24865_, new_n24863_, new_n24861_ );
xor  ( new_n24866_, new_n24784_, new_n24780_ );
xnor ( new_n24867_, new_n24866_, new_n24789_ );
nor  ( new_n24868_, new_n24867_, new_n24865_ );
nor  ( new_n24869_, new_n24868_, new_n24864_ );
not  ( new_n24870_, new_n24869_ );
and  ( new_n24871_, new_n24870_, new_n24859_ );
or   ( new_n24872_, new_n24871_, new_n24858_ );
or   ( new_n24873_, new_n524_, new_n22973_ );
or   ( new_n24874_, new_n526_, new_n22975_ );
and  ( new_n24875_, new_n24874_, new_n24873_ );
xor  ( new_n24876_, new_n24875_, new_n403_ );
or   ( new_n24877_, new_n409_, new_n23252_ );
or   ( new_n24878_, new_n411_, new_n23166_ );
and  ( new_n24879_, new_n24878_, new_n24877_ );
xor  ( new_n24880_, new_n24879_, new_n328_ );
or   ( new_n24881_, new_n24880_, new_n24876_ );
or   ( new_n24882_, new_n337_, new_n23554_ );
or   ( new_n24883_, new_n340_, new_n23370_ );
and  ( new_n24884_, new_n24883_, new_n24882_ );
xor  ( new_n24885_, new_n24884_, new_n332_ );
and  ( new_n24886_, new_n24880_, new_n24876_ );
or   ( new_n24887_, new_n24886_, new_n24885_ );
and  ( new_n24888_, new_n24887_, new_n24881_ );
or   ( new_n24889_, new_n1135_, new_n22304_ );
or   ( new_n24890_, new_n1137_, new_n22207_ );
and  ( new_n24891_, new_n24890_, new_n24889_ );
xor  ( new_n24892_, new_n24891_, new_n896_ );
or   ( new_n24893_, new_n897_, new_n22590_ );
or   ( new_n24894_, new_n899_, new_n22423_ );
and  ( new_n24895_, new_n24894_, new_n24893_ );
xor  ( new_n24896_, new_n24895_, new_n748_ );
or   ( new_n24897_, new_n24896_, new_n24892_ );
or   ( new_n24898_, new_n755_, new_n22829_ );
or   ( new_n24899_, new_n757_, new_n22641_ );
and  ( new_n24900_, new_n24899_, new_n24898_ );
xor  ( new_n24901_, new_n24900_, new_n523_ );
and  ( new_n24902_, new_n24896_, new_n24892_ );
or   ( new_n24903_, new_n24902_, new_n24901_ );
and  ( new_n24904_, new_n24903_, new_n24897_ );
nor  ( new_n24905_, new_n24904_, new_n24888_ );
and  ( new_n24906_, new_n24904_, new_n24888_ );
or   ( new_n24907_, new_n317_, new_n23895_ );
or   ( new_n24908_, new_n320_, new_n23733_ );
and  ( new_n24909_, new_n24908_, new_n24907_ );
xor  ( new_n24910_, new_n24909_, new_n312_ );
or   ( new_n24911_, new_n283_, new_n24227_ );
or   ( new_n24912_, new_n286_, new_n24006_ );
and  ( new_n24913_, new_n24912_, new_n24911_ );
xor  ( new_n24914_, new_n24913_, new_n278_ );
nor  ( new_n24915_, new_n24914_, new_n24910_ );
or   ( new_n24916_, new_n299_, new_n24543_ );
or   ( new_n24917_, new_n302_, new_n24418_ );
and  ( new_n24918_, new_n24917_, new_n24916_ );
xor  ( new_n24919_, new_n24918_, new_n293_ );
and  ( new_n24920_, new_n24914_, new_n24910_ );
nor  ( new_n24921_, new_n24920_, new_n24919_ );
nor  ( new_n24922_, new_n24921_, new_n24915_ );
nor  ( new_n24923_, new_n24922_, new_n24906_ );
nor  ( new_n24924_, new_n24923_, new_n24905_ );
not  ( new_n24925_, RIbb326d0_165 );
or   ( new_n24926_, new_n268_, new_n24925_ );
not  ( new_n24927_, RIbb32658_164 );
or   ( new_n24928_, new_n271_, new_n24927_ );
and  ( new_n24929_, new_n24928_, new_n24926_ );
xor  ( new_n24930_, new_n24929_, new_n263_ );
and  ( new_n24931_, RIbb32748_166, RIbb2f610_1 );
or   ( new_n24932_, new_n24931_, new_n24930_ );
or   ( new_n24933_, new_n268_, new_n24927_ );
or   ( new_n24934_, new_n271_, new_n24543_ );
and  ( new_n24935_, new_n24934_, new_n24933_ );
xor  ( new_n24936_, new_n24935_, new_n263_ );
or   ( new_n24937_, new_n24936_, new_n24932_ );
and  ( new_n24938_, RIbb326d0_165, RIbb2f610_1 );
and  ( new_n24939_, new_n24936_, new_n24932_ );
or   ( new_n24940_, new_n24939_, new_n24938_ );
and  ( new_n24941_, new_n24940_, new_n24937_ );
or   ( new_n24942_, new_n2807_, new_n21680_ );
or   ( new_n24943_, new_n2809_, new_n21672_ );
and  ( new_n24944_, new_n24943_, new_n24942_ );
xor  ( new_n24945_, new_n24944_, new_n2424_ );
or   ( new_n24946_, new_n2425_, new_n21687_ );
or   ( new_n24947_, new_n2427_, new_n21678_ );
and  ( new_n24948_, new_n24947_, new_n24946_ );
xor  ( new_n24949_, new_n24948_, new_n2121_ );
or   ( new_n24950_, new_n24949_, new_n24945_ );
or   ( new_n24951_, new_n2122_, new_n21751_ );
or   ( new_n24952_, new_n2124_, new_n21685_ );
and  ( new_n24953_, new_n24952_, new_n24951_ );
xor  ( new_n24954_, new_n24953_, new_n1843_ );
and  ( new_n24955_, new_n24949_, new_n24945_ );
or   ( new_n24956_, new_n24955_, new_n24954_ );
and  ( new_n24957_, new_n24956_, new_n24950_ );
or   ( new_n24958_, new_n3461_, new_n21703_ );
or   ( new_n24959_, new_n3463_, new_n21694_ );
and  ( new_n24960_, new_n24959_, new_n24958_ );
xor  ( new_n24961_, new_n24960_, new_n3115_ );
and  ( new_n24962_, new_n3733_, RIbb315f0_129 );
xor  ( new_n24963_, new_n24962_, new_n3460_ );
nand ( new_n24964_, new_n24963_, new_n24961_ );
or   ( new_n24965_, new_n3117_, new_n21674_ );
or   ( new_n24966_, new_n3119_, new_n21701_ );
and  ( new_n24967_, new_n24966_, new_n24965_ );
xor  ( new_n24968_, new_n24967_, new_n2800_ );
nor  ( new_n24969_, new_n24963_, new_n24961_ );
or   ( new_n24970_, new_n24969_, new_n24968_ );
and  ( new_n24971_, new_n24970_, new_n24964_ );
or   ( new_n24972_, new_n24971_, new_n24957_ );
and  ( new_n24973_, new_n24971_, new_n24957_ );
or   ( new_n24974_, new_n1844_, new_n21842_ );
or   ( new_n24975_, new_n1846_, new_n21792_ );
and  ( new_n24976_, new_n24975_, new_n24974_ );
xor  ( new_n24977_, new_n24976_, new_n1586_ );
or   ( new_n24978_, new_n1593_, new_n21847_ );
or   ( new_n24979_, new_n1595_, new_n21840_ );
and  ( new_n24980_, new_n24979_, new_n24978_ );
xor  ( new_n24981_, new_n24980_, new_n1358_ );
nor  ( new_n24982_, new_n24981_, new_n24977_ );
or   ( new_n24983_, new_n1364_, new_n22129_ );
or   ( new_n24984_, new_n1366_, new_n22098_ );
and  ( new_n24985_, new_n24984_, new_n24983_ );
xor  ( new_n24986_, new_n24985_, new_n1129_ );
and  ( new_n24987_, new_n24981_, new_n24977_ );
nor  ( new_n24988_, new_n24987_, new_n24986_ );
nor  ( new_n24989_, new_n24988_, new_n24982_ );
or   ( new_n24990_, new_n24989_, new_n24973_ );
and  ( new_n24991_, new_n24990_, new_n24972_ );
and  ( new_n24992_, new_n24991_, new_n24941_ );
or   ( new_n24993_, new_n24992_, new_n24924_ );
or   ( new_n24994_, new_n24991_, new_n24941_ );
and  ( new_n24995_, new_n24994_, new_n24993_ );
or   ( new_n24996_, new_n24995_, new_n24872_ );
nand ( new_n24997_, new_n24995_, new_n24872_ );
xor  ( new_n24998_, new_n24532_, new_n24530_ );
xor  ( new_n24999_, new_n24998_, new_n24537_ );
xnor ( new_n25000_, new_n24675_, new_n24673_ );
xor  ( new_n25001_, new_n25000_, new_n24679_ );
and  ( new_n25002_, new_n25001_, new_n24999_ );
xor  ( new_n25003_, new_n24692_, new_n24690_ );
nor  ( new_n25004_, new_n25001_, new_n24999_ );
nor  ( new_n25005_, new_n25004_, new_n25003_ );
nor  ( new_n25006_, new_n25005_, new_n25002_ );
nand ( new_n25007_, new_n25006_, new_n24997_ );
and  ( new_n25008_, new_n25007_, new_n24996_ );
nor  ( new_n25009_, new_n25008_, new_n24845_ );
nand ( new_n25010_, new_n25008_, new_n24845_ );
xor  ( new_n25011_, new_n24741_, new_n24693_ );
xor  ( new_n25012_, new_n25011_, new_n24795_ );
xor  ( new_n25013_, new_n24681_, new_n24671_ );
xor  ( new_n25014_, new_n25013_, new_n24686_ );
nor  ( new_n25015_, new_n25014_, new_n25012_ );
and  ( new_n25016_, new_n25014_, new_n25012_ );
not  ( new_n25017_, new_n25016_ );
xor  ( new_n25018_, new_n24804_, new_n24802_ );
xnor ( new_n25019_, new_n25018_, new_n24808_ );
and  ( new_n25020_, new_n25019_, new_n25017_ );
nor  ( new_n25021_, new_n25020_, new_n25015_ );
and  ( new_n25022_, new_n25021_, new_n25010_ );
or   ( new_n25023_, new_n25022_, new_n25009_ );
xor  ( new_n25024_, new_n24627_, new_n24609_ );
xor  ( new_n25025_, new_n25024_, new_n24638_ );
or   ( new_n25026_, new_n25025_, new_n25023_ );
and  ( new_n25027_, new_n25025_, new_n25023_ );
xor  ( new_n25028_, new_n24816_, new_n24814_ );
xor  ( new_n25029_, new_n25028_, new_n24828_ );
or   ( new_n25030_, new_n25029_, new_n25027_ );
and  ( new_n25031_, new_n25030_, new_n25026_ );
nor  ( new_n25032_, new_n25031_, new_n24843_ );
xor  ( new_n25033_, new_n24838_, new_n24669_ );
and  ( new_n25034_, new_n25033_, new_n25032_ );
xor  ( new_n25035_, new_n25025_, new_n25023_ );
xor  ( new_n25036_, new_n25035_, new_n25029_ );
xor  ( new_n25037_, new_n24798_, new_n24688_ );
or   ( new_n25038_, new_n25037_, new_n24811_ );
not  ( new_n25039_, new_n24812_ );
or   ( new_n25040_, new_n24813_, new_n25039_ );
and  ( new_n25041_, new_n25040_, new_n25038_ );
xor  ( new_n25042_, new_n25014_, new_n25012_ );
xor  ( new_n25043_, new_n25042_, new_n25019_ );
or   ( new_n25044_, new_n299_, new_n24927_ );
or   ( new_n25045_, new_n302_, new_n24543_ );
and  ( new_n25046_, new_n25045_, new_n25044_ );
xor  ( new_n25047_, new_n25046_, new_n293_ );
not  ( new_n25048_, RIbb32748_166 );
or   ( new_n25049_, new_n268_, new_n25048_ );
or   ( new_n25050_, new_n271_, new_n24925_ );
and  ( new_n25051_, new_n25050_, new_n25049_ );
xor  ( new_n25052_, new_n25051_, new_n263_ );
nor  ( new_n25053_, new_n25052_, new_n25047_ );
and  ( new_n25054_, RIbb327c0_167, RIbb2f610_1 );
not  ( new_n25055_, new_n25054_ );
nand ( new_n25056_, new_n25052_, new_n25047_ );
and  ( new_n25057_, new_n25056_, new_n25055_ );
or   ( new_n25058_, new_n25057_, new_n25053_ );
xnor ( new_n25059_, new_n24914_, new_n24910_ );
xor  ( new_n25060_, new_n25059_, new_n24919_ );
nor  ( new_n25061_, new_n25060_, new_n25058_ );
xor  ( new_n25062_, new_n24931_, new_n24930_ );
and  ( new_n25063_, new_n25060_, new_n25058_ );
nor  ( new_n25064_, new_n25063_, new_n25062_ );
or   ( new_n25065_, new_n25064_, new_n25061_ );
or   ( new_n25066_, new_n1364_, new_n22207_ );
or   ( new_n25067_, new_n1366_, new_n22129_ );
and  ( new_n25068_, new_n25067_, new_n25066_ );
xor  ( new_n25069_, new_n25068_, new_n1129_ );
or   ( new_n25070_, new_n1135_, new_n22423_ );
or   ( new_n25071_, new_n1137_, new_n22304_ );
and  ( new_n25072_, new_n25071_, new_n25070_ );
xor  ( new_n25073_, new_n25072_, new_n896_ );
or   ( new_n25074_, new_n25073_, new_n25069_ );
and  ( new_n25075_, new_n25073_, new_n25069_ );
or   ( new_n25076_, new_n897_, new_n22641_ );
or   ( new_n25077_, new_n899_, new_n22590_ );
and  ( new_n25078_, new_n25077_, new_n25076_ );
xor  ( new_n25079_, new_n25078_, new_n748_ );
or   ( new_n25080_, new_n25079_, new_n25075_ );
and  ( new_n25081_, new_n25080_, new_n25074_ );
or   ( new_n25082_, new_n755_, new_n22975_ );
or   ( new_n25083_, new_n757_, new_n22829_ );
and  ( new_n25084_, new_n25083_, new_n25082_ );
xor  ( new_n25085_, new_n25084_, new_n523_ );
or   ( new_n25086_, new_n524_, new_n23166_ );
or   ( new_n25087_, new_n526_, new_n22973_ );
and  ( new_n25088_, new_n25087_, new_n25086_ );
xor  ( new_n25089_, new_n25088_, new_n403_ );
or   ( new_n25090_, new_n25089_, new_n25085_ );
and  ( new_n25091_, new_n25089_, new_n25085_ );
or   ( new_n25092_, new_n409_, new_n23370_ );
or   ( new_n25093_, new_n411_, new_n23252_ );
and  ( new_n25094_, new_n25093_, new_n25092_ );
xor  ( new_n25095_, new_n25094_, new_n328_ );
or   ( new_n25096_, new_n25095_, new_n25091_ );
and  ( new_n25097_, new_n25096_, new_n25090_ );
or   ( new_n25098_, new_n25097_, new_n25081_ );
and  ( new_n25099_, new_n25097_, new_n25081_ );
or   ( new_n25100_, new_n337_, new_n23733_ );
or   ( new_n25101_, new_n340_, new_n23554_ );
and  ( new_n25102_, new_n25101_, new_n25100_ );
xor  ( new_n25103_, new_n25102_, new_n332_ );
or   ( new_n25104_, new_n317_, new_n24006_ );
or   ( new_n25105_, new_n320_, new_n23895_ );
and  ( new_n25106_, new_n25105_, new_n25104_ );
xor  ( new_n25107_, new_n25106_, new_n312_ );
nor  ( new_n25108_, new_n25107_, new_n25103_ );
or   ( new_n25109_, new_n283_, new_n24418_ );
or   ( new_n25110_, new_n286_, new_n24227_ );
and  ( new_n25111_, new_n25110_, new_n25109_ );
xor  ( new_n25112_, new_n25111_, new_n278_ );
and  ( new_n25113_, new_n25107_, new_n25103_ );
nor  ( new_n25114_, new_n25113_, new_n25112_ );
nor  ( new_n25115_, new_n25114_, new_n25108_ );
or   ( new_n25116_, new_n25115_, new_n25099_ );
and  ( new_n25117_, new_n25116_, new_n25098_ );
nor  ( new_n25118_, new_n25117_, new_n25065_ );
nand ( new_n25119_, new_n25117_, new_n25065_ );
or   ( new_n25120_, new_n3896_, new_n21694_ );
or   ( new_n25121_, new_n3898_, new_n21696_ );
and  ( new_n25122_, new_n25121_, new_n25120_ );
xor  ( new_n25123_, new_n25122_, new_n3460_ );
and  ( new_n25124_, new_n25123_, new_n3895_ );
or   ( new_n25125_, new_n25123_, new_n3895_ );
or   ( new_n25126_, new_n3461_, new_n21701_ );
or   ( new_n25127_, new_n3463_, new_n21703_ );
and  ( new_n25128_, new_n25127_, new_n25126_ );
xor  ( new_n25129_, new_n25128_, new_n3116_ );
and  ( new_n25130_, new_n25129_, new_n25125_ );
or   ( new_n25131_, new_n25130_, new_n25124_ );
or   ( new_n25132_, new_n3117_, new_n21672_ );
or   ( new_n25133_, new_n3119_, new_n21674_ );
and  ( new_n25134_, new_n25133_, new_n25132_ );
xor  ( new_n25135_, new_n25134_, new_n2800_ );
or   ( new_n25136_, new_n2807_, new_n21678_ );
or   ( new_n25137_, new_n2809_, new_n21680_ );
and  ( new_n25138_, new_n25137_, new_n25136_ );
xor  ( new_n25139_, new_n25138_, new_n2424_ );
or   ( new_n25140_, new_n25139_, new_n25135_ );
and  ( new_n25141_, new_n25139_, new_n25135_ );
or   ( new_n25142_, new_n2425_, new_n21685_ );
or   ( new_n25143_, new_n2427_, new_n21687_ );
and  ( new_n25144_, new_n25143_, new_n25142_ );
xor  ( new_n25145_, new_n25144_, new_n2121_ );
or   ( new_n25146_, new_n25145_, new_n25141_ );
and  ( new_n25147_, new_n25146_, new_n25140_ );
nor  ( new_n25148_, new_n25147_, new_n25131_ );
and  ( new_n25149_, new_n25147_, new_n25131_ );
or   ( new_n25150_, new_n2122_, new_n21792_ );
or   ( new_n25151_, new_n2124_, new_n21751_ );
and  ( new_n25152_, new_n25151_, new_n25150_ );
xor  ( new_n25153_, new_n25152_, new_n1843_ );
or   ( new_n25154_, new_n1844_, new_n21840_ );
or   ( new_n25155_, new_n1846_, new_n21842_ );
and  ( new_n25156_, new_n25155_, new_n25154_ );
xor  ( new_n25157_, new_n25156_, new_n1586_ );
nor  ( new_n25158_, new_n25157_, new_n25153_ );
and  ( new_n25159_, new_n25157_, new_n25153_ );
or   ( new_n25160_, new_n1593_, new_n22098_ );
or   ( new_n25161_, new_n1595_, new_n21847_ );
and  ( new_n25162_, new_n25161_, new_n25160_ );
xor  ( new_n25163_, new_n25162_, new_n1358_ );
nor  ( new_n25164_, new_n25163_, new_n25159_ );
nor  ( new_n25165_, new_n25164_, new_n25158_ );
nor  ( new_n25166_, new_n25165_, new_n25149_ );
nor  ( new_n25167_, new_n25166_, new_n25148_ );
not  ( new_n25168_, new_n25167_ );
and  ( new_n25169_, new_n25168_, new_n25119_ );
or   ( new_n25170_, new_n25169_, new_n25118_ );
xor  ( new_n25171_, new_n24963_, new_n24961_ );
xnor ( new_n25172_, new_n25171_, new_n24968_ );
xnor ( new_n25173_, new_n24949_, new_n24945_ );
xor  ( new_n25174_, new_n25173_, new_n24954_ );
or   ( new_n25175_, new_n25174_, new_n25172_ );
xnor ( new_n25176_, new_n24896_, new_n24892_ );
xor  ( new_n25177_, new_n25176_, new_n24901_ );
xnor ( new_n25178_, new_n24880_, new_n24876_ );
xor  ( new_n25179_, new_n25178_, new_n24885_ );
or   ( new_n25180_, new_n25179_, new_n25177_ );
and  ( new_n25181_, new_n25179_, new_n25177_ );
xnor ( new_n25182_, new_n24981_, new_n24977_ );
xor  ( new_n25183_, new_n25182_, new_n24986_ );
or   ( new_n25184_, new_n25183_, new_n25181_ );
and  ( new_n25185_, new_n25184_, new_n25180_ );
or   ( new_n25186_, new_n25185_, new_n25175_ );
and  ( new_n25187_, new_n25185_, new_n25175_ );
xor  ( new_n25188_, new_n24851_, new_n24849_ );
xor  ( new_n25189_, new_n25188_, new_n24855_ );
or   ( new_n25190_, new_n25189_, new_n25187_ );
and  ( new_n25191_, new_n25190_, new_n25186_ );
nand ( new_n25192_, new_n25191_, new_n25170_ );
or   ( new_n25193_, new_n25191_, new_n25170_ );
xnor ( new_n25194_, new_n24904_, new_n24888_ );
xor  ( new_n25195_, new_n25194_, new_n24922_ );
xnor ( new_n25196_, new_n24936_, new_n24932_ );
xor  ( new_n25197_, new_n25196_, new_n24938_ );
nor  ( new_n25198_, new_n25197_, new_n25195_ );
and  ( new_n25199_, new_n25197_, new_n25195_ );
xor  ( new_n25200_, new_n24863_, new_n24861_ );
xnor ( new_n25201_, new_n25200_, new_n24867_ );
not  ( new_n25202_, new_n25201_ );
nor  ( new_n25203_, new_n25202_, new_n25199_ );
nor  ( new_n25204_, new_n25203_, new_n25198_ );
nand ( new_n25205_, new_n25204_, new_n25193_ );
and  ( new_n25206_, new_n25205_, new_n25192_ );
or   ( new_n25207_, new_n25206_, new_n25043_ );
nand ( new_n25208_, new_n25206_, new_n25043_ );
xnor ( new_n25209_, new_n24721_, new_n24705_ );
xor  ( new_n25210_, new_n25209_, new_n24739_ );
xnor ( new_n25211_, new_n24774_, new_n24758_ );
xor  ( new_n25212_, new_n25211_, new_n24792_ );
nor  ( new_n25213_, new_n25212_, new_n25210_ );
and  ( new_n25214_, new_n25212_, new_n25210_ );
xor  ( new_n25215_, new_n25001_, new_n24999_ );
xnor ( new_n25216_, new_n25215_, new_n25003_ );
not  ( new_n25217_, new_n25216_ );
nor  ( new_n25218_, new_n25217_, new_n25214_ );
nor  ( new_n25219_, new_n25218_, new_n25213_ );
nand ( new_n25220_, new_n25219_, new_n25208_ );
and  ( new_n25221_, new_n25220_, new_n25207_ );
nand ( new_n25222_, new_n25221_, new_n25041_ );
nor  ( new_n25223_, new_n25221_, new_n25041_ );
xor  ( new_n25224_, new_n25008_, new_n24845_ );
xor  ( new_n25225_, new_n25224_, new_n25021_ );
or   ( new_n25226_, new_n25225_, new_n25223_ );
and  ( new_n25227_, new_n25226_, new_n25222_ );
nor  ( new_n25228_, new_n25227_, new_n25036_ );
xor  ( new_n25229_, new_n25031_, new_n24843_ );
and  ( new_n25230_, new_n25229_, new_n25228_ );
xor  ( new_n25231_, new_n24995_, new_n24872_ );
xor  ( new_n25232_, new_n25231_, new_n25006_ );
not  ( new_n25233_, new_n25232_ );
or   ( new_n25234_, new_n3117_, new_n21680_ );
or   ( new_n25235_, new_n3119_, new_n21672_ );
and  ( new_n25236_, new_n25235_, new_n25234_ );
xor  ( new_n25237_, new_n25236_, new_n2800_ );
or   ( new_n25238_, new_n2807_, new_n21687_ );
or   ( new_n25239_, new_n2809_, new_n21678_ );
and  ( new_n25240_, new_n25239_, new_n25238_ );
xor  ( new_n25241_, new_n25240_, new_n2424_ );
or   ( new_n25242_, new_n25241_, new_n25237_ );
and  ( new_n25243_, new_n25241_, new_n25237_ );
or   ( new_n25244_, new_n2425_, new_n21751_ );
or   ( new_n25245_, new_n2427_, new_n21685_ );
and  ( new_n25246_, new_n25245_, new_n25244_ );
xor  ( new_n25247_, new_n25246_, new_n2121_ );
or   ( new_n25248_, new_n25247_, new_n25243_ );
and  ( new_n25249_, new_n25248_, new_n25242_ );
or   ( new_n25250_, new_n3896_, new_n21703_ );
or   ( new_n25251_, new_n3898_, new_n21694_ );
and  ( new_n25252_, new_n25251_, new_n25250_ );
xor  ( new_n25253_, new_n25252_, new_n3459_ );
and  ( new_n25254_, new_n4034_, RIbb315f0_129 );
xor  ( new_n25255_, new_n25254_, new_n3895_ );
nand ( new_n25256_, new_n25255_, new_n25253_ );
nor  ( new_n25257_, new_n25255_, new_n25253_ );
or   ( new_n25258_, new_n3461_, new_n21674_ );
or   ( new_n25259_, new_n3463_, new_n21701_ );
and  ( new_n25260_, new_n25259_, new_n25258_ );
xor  ( new_n25261_, new_n25260_, new_n3116_ );
or   ( new_n25262_, new_n25261_, new_n25257_ );
and  ( new_n25263_, new_n25262_, new_n25256_ );
or   ( new_n25264_, new_n25263_, new_n25249_ );
and  ( new_n25265_, new_n25263_, new_n25249_ );
or   ( new_n25266_, new_n2122_, new_n21842_ );
or   ( new_n25267_, new_n2124_, new_n21792_ );
and  ( new_n25268_, new_n25267_, new_n25266_ );
xor  ( new_n25269_, new_n25268_, new_n1843_ );
or   ( new_n25270_, new_n1844_, new_n21847_ );
or   ( new_n25271_, new_n1846_, new_n21840_ );
and  ( new_n25272_, new_n25271_, new_n25270_ );
xor  ( new_n25273_, new_n25272_, new_n1586_ );
nor  ( new_n25274_, new_n25273_, new_n25269_ );
and  ( new_n25275_, new_n25273_, new_n25269_ );
or   ( new_n25276_, new_n1593_, new_n22129_ );
or   ( new_n25277_, new_n1595_, new_n22098_ );
and  ( new_n25278_, new_n25277_, new_n25276_ );
xor  ( new_n25279_, new_n25278_, new_n1358_ );
nor  ( new_n25280_, new_n25279_, new_n25275_ );
nor  ( new_n25281_, new_n25280_, new_n25274_ );
or   ( new_n25282_, new_n25281_, new_n25265_ );
and  ( new_n25283_, new_n25282_, new_n25264_ );
or   ( new_n25284_, new_n299_, new_n24925_ );
or   ( new_n25285_, new_n302_, new_n24927_ );
and  ( new_n25286_, new_n25285_, new_n25284_ );
xor  ( new_n25287_, new_n25286_, new_n293_ );
not  ( new_n25288_, RIbb327c0_167 );
or   ( new_n25289_, new_n268_, new_n25288_ );
or   ( new_n25290_, new_n271_, new_n25048_ );
and  ( new_n25291_, new_n25290_, new_n25289_ );
xor  ( new_n25292_, new_n25291_, new_n263_ );
nor  ( new_n25293_, new_n25292_, new_n25287_ );
and  ( new_n25294_, RIbb32838_168, RIbb2f610_1 );
not  ( new_n25295_, new_n25294_ );
nand ( new_n25296_, new_n25292_, new_n25287_ );
and  ( new_n25297_, new_n25296_, new_n25295_ );
or   ( new_n25298_, new_n25297_, new_n25293_ );
xnor ( new_n25299_, new_n25107_, new_n25103_ );
xor  ( new_n25300_, new_n25299_, new_n25112_ );
nand ( new_n25301_, new_n25300_, new_n25298_ );
or   ( new_n25302_, new_n25300_, new_n25298_ );
xor  ( new_n25303_, new_n25052_, new_n25047_ );
xor  ( new_n25304_, new_n25303_, new_n25055_ );
nand ( new_n25305_, new_n25304_, new_n25302_ );
and  ( new_n25306_, new_n25305_, new_n25301_ );
nor  ( new_n25307_, new_n25306_, new_n25283_ );
nand ( new_n25308_, new_n25306_, new_n25283_ );
or   ( new_n25309_, new_n1364_, new_n22304_ );
or   ( new_n25310_, new_n1366_, new_n22207_ );
and  ( new_n25311_, new_n25310_, new_n25309_ );
xor  ( new_n25312_, new_n25311_, new_n1129_ );
or   ( new_n25313_, new_n1135_, new_n22590_ );
or   ( new_n25314_, new_n1137_, new_n22423_ );
and  ( new_n25315_, new_n25314_, new_n25313_ );
xor  ( new_n25316_, new_n25315_, new_n896_ );
or   ( new_n25317_, new_n25316_, new_n25312_ );
and  ( new_n25318_, new_n25316_, new_n25312_ );
or   ( new_n25319_, new_n897_, new_n22829_ );
or   ( new_n25320_, new_n899_, new_n22641_ );
and  ( new_n25321_, new_n25320_, new_n25319_ );
xor  ( new_n25322_, new_n25321_, new_n748_ );
or   ( new_n25323_, new_n25322_, new_n25318_ );
and  ( new_n25324_, new_n25323_, new_n25317_ );
or   ( new_n25325_, new_n337_, new_n23895_ );
or   ( new_n25326_, new_n340_, new_n23733_ );
and  ( new_n25327_, new_n25326_, new_n25325_ );
xor  ( new_n25328_, new_n25327_, new_n332_ );
or   ( new_n25329_, new_n317_, new_n24227_ );
or   ( new_n25330_, new_n320_, new_n24006_ );
and  ( new_n25331_, new_n25330_, new_n25329_ );
xor  ( new_n25332_, new_n25331_, new_n312_ );
or   ( new_n25333_, new_n25332_, new_n25328_ );
and  ( new_n25334_, new_n25332_, new_n25328_ );
or   ( new_n25335_, new_n283_, new_n24543_ );
or   ( new_n25336_, new_n286_, new_n24418_ );
and  ( new_n25337_, new_n25336_, new_n25335_ );
xor  ( new_n25338_, new_n25337_, new_n278_ );
or   ( new_n25339_, new_n25338_, new_n25334_ );
and  ( new_n25340_, new_n25339_, new_n25333_ );
nor  ( new_n25341_, new_n25340_, new_n25324_ );
nand ( new_n25342_, new_n25340_, new_n25324_ );
or   ( new_n25343_, new_n755_, new_n22973_ );
or   ( new_n25344_, new_n757_, new_n22975_ );
and  ( new_n25345_, new_n25344_, new_n25343_ );
xor  ( new_n25346_, new_n25345_, new_n523_ );
or   ( new_n25347_, new_n524_, new_n23252_ );
or   ( new_n25348_, new_n526_, new_n23166_ );
and  ( new_n25349_, new_n25348_, new_n25347_ );
xor  ( new_n25350_, new_n25349_, new_n403_ );
nor  ( new_n25351_, new_n25350_, new_n25346_ );
nand ( new_n25352_, new_n25350_, new_n25346_ );
or   ( new_n25353_, new_n409_, new_n23554_ );
or   ( new_n25354_, new_n411_, new_n23370_ );
and  ( new_n25355_, new_n25354_, new_n25353_ );
xor  ( new_n25356_, new_n25355_, new_n328_ );
not  ( new_n25357_, new_n25356_ );
and  ( new_n25358_, new_n25357_, new_n25352_ );
or   ( new_n25359_, new_n25358_, new_n25351_ );
and  ( new_n25360_, new_n25359_, new_n25342_ );
or   ( new_n25361_, new_n25360_, new_n25341_ );
and  ( new_n25362_, new_n25361_, new_n25308_ );
or   ( new_n25363_, new_n25362_, new_n25307_ );
xnor ( new_n25364_, new_n25097_, new_n25081_ );
xor  ( new_n25365_, new_n25364_, new_n25115_ );
xnor ( new_n25366_, new_n25147_, new_n25131_ );
xor  ( new_n25367_, new_n25366_, new_n25165_ );
or   ( new_n25368_, new_n25367_, new_n25365_ );
and  ( new_n25369_, new_n25367_, new_n25365_ );
xor  ( new_n25370_, new_n25060_, new_n25058_ );
xor  ( new_n25371_, new_n25370_, new_n25062_ );
or   ( new_n25372_, new_n25371_, new_n25369_ );
and  ( new_n25373_, new_n25372_, new_n25368_ );
and  ( new_n25374_, new_n25373_, new_n25363_ );
nor  ( new_n25375_, new_n25373_, new_n25363_ );
xor  ( new_n25376_, new_n25179_, new_n25177_ );
xor  ( new_n25377_, new_n25376_, new_n25183_ );
xnor ( new_n25378_, new_n25089_, new_n25085_ );
xor  ( new_n25379_, new_n25378_, new_n25095_ );
xnor ( new_n25380_, new_n25073_, new_n25069_ );
xor  ( new_n25381_, new_n25380_, new_n25079_ );
or   ( new_n25382_, new_n25381_, new_n25379_ );
and  ( new_n25383_, new_n25381_, new_n25379_ );
xor  ( new_n25384_, new_n25157_, new_n25153_ );
xnor ( new_n25385_, new_n25384_, new_n25163_ );
or   ( new_n25386_, new_n25385_, new_n25383_ );
and  ( new_n25387_, new_n25386_, new_n25382_ );
nor  ( new_n25388_, new_n25387_, new_n25377_ );
and  ( new_n25389_, new_n25387_, new_n25377_ );
xor  ( new_n25390_, new_n25174_, new_n25172_ );
not  ( new_n25391_, new_n25390_ );
nor  ( new_n25392_, new_n25391_, new_n25389_ );
nor  ( new_n25393_, new_n25392_, new_n25388_ );
not  ( new_n25394_, new_n25393_ );
nor  ( new_n25395_, new_n25394_, new_n25375_ );
nor  ( new_n25396_, new_n25395_, new_n25374_ );
xor  ( new_n25397_, new_n24857_, new_n24847_ );
xor  ( new_n25398_, new_n25397_, new_n24870_ );
and  ( new_n25399_, new_n25398_, new_n25396_ );
xnor ( new_n25400_, new_n24971_, new_n24957_ );
xor  ( new_n25401_, new_n25400_, new_n24989_ );
xor  ( new_n25402_, new_n25185_, new_n25175_ );
xor  ( new_n25403_, new_n25402_, new_n25189_ );
nor  ( new_n25404_, new_n25403_, new_n25401_ );
and  ( new_n25405_, new_n25403_, new_n25401_ );
xor  ( new_n25406_, new_n25197_, new_n25195_ );
xor  ( new_n25407_, new_n25406_, new_n25202_ );
nor  ( new_n25408_, new_n25407_, new_n25405_ );
nor  ( new_n25409_, new_n25408_, new_n25404_ );
not  ( new_n25410_, new_n25396_ );
not  ( new_n25411_, new_n25398_ );
and  ( new_n25412_, new_n25411_, new_n25410_ );
nor  ( new_n25413_, new_n25412_, new_n25409_ );
nor  ( new_n25414_, new_n25413_, new_n25399_ );
not  ( new_n25415_, new_n25414_ );
and  ( new_n25416_, new_n25415_, new_n25233_ );
not  ( new_n25417_, new_n25416_ );
and  ( new_n25418_, new_n25414_, new_n25232_ );
xnor ( new_n25419_, new_n24991_, new_n24924_ );
xor  ( new_n25420_, new_n25419_, new_n24941_ );
xor  ( new_n25421_, new_n25191_, new_n25170_ );
xor  ( new_n25422_, new_n25421_, new_n25204_ );
nor  ( new_n25423_, new_n25422_, new_n25420_ );
and  ( new_n25424_, new_n25422_, new_n25420_ );
xor  ( new_n25425_, new_n25212_, new_n25210_ );
xor  ( new_n25426_, new_n25425_, new_n25217_ );
nor  ( new_n25427_, new_n25426_, new_n25424_ );
nor  ( new_n25428_, new_n25427_, new_n25423_ );
nor  ( new_n25429_, new_n25428_, new_n25418_ );
not  ( new_n25430_, new_n25429_ );
and  ( new_n25431_, new_n25430_, new_n25417_ );
xnor ( new_n25432_, new_n25221_, new_n25041_ );
xnor ( new_n25433_, new_n25432_, new_n25225_ );
nor  ( new_n25434_, new_n25433_, new_n25431_ );
xor  ( new_n25435_, new_n25227_, new_n25036_ );
and  ( new_n25436_, new_n25435_, new_n25434_ );
xnor ( new_n25437_, new_n25433_, new_n25431_ );
xor  ( new_n25438_, new_n25373_, new_n25363_ );
xor  ( new_n25439_, new_n25438_, new_n25393_ );
not  ( new_n25440_, new_n25439_ );
xnor ( new_n25441_, new_n25403_, new_n25401_ );
xor  ( new_n25442_, new_n25441_, new_n25407_ );
and  ( new_n25443_, new_n25442_, new_n25440_ );
xnor ( new_n25444_, new_n25422_, new_n25420_ );
xor  ( new_n25445_, new_n25444_, new_n25426_ );
or   ( new_n25446_, new_n25445_, new_n25443_ );
and  ( new_n25447_, new_n25445_, new_n25443_ );
xnor ( new_n25448_, new_n25139_, new_n25135_ );
xor  ( new_n25449_, new_n25448_, new_n25145_ );
xnor ( new_n25450_, new_n25255_, new_n25253_ );
xor  ( new_n25451_, new_n25450_, new_n25261_ );
xnor ( new_n25452_, new_n25241_, new_n25237_ );
xor  ( new_n25453_, new_n25452_, new_n25247_ );
or   ( new_n25454_, new_n25453_, new_n25451_ );
and  ( new_n25455_, new_n25453_, new_n25451_ );
xnor ( new_n25456_, new_n25273_, new_n25269_ );
xor  ( new_n25457_, new_n25456_, new_n25279_ );
or   ( new_n25458_, new_n25457_, new_n25455_ );
and  ( new_n25459_, new_n25458_, new_n25454_ );
nor  ( new_n25460_, new_n25459_, new_n25449_ );
and  ( new_n25461_, new_n25459_, new_n25449_ );
xnor ( new_n25462_, new_n25332_, new_n25328_ );
xor  ( new_n25463_, new_n25462_, new_n25338_ );
xnor ( new_n25464_, new_n25316_, new_n25312_ );
xor  ( new_n25465_, new_n25464_, new_n25322_ );
nor  ( new_n25466_, new_n25465_, new_n25463_ );
and  ( new_n25467_, new_n25465_, new_n25463_ );
xor  ( new_n25468_, new_n25350_, new_n25346_ );
xor  ( new_n25469_, new_n25468_, new_n25357_ );
nor  ( new_n25470_, new_n25469_, new_n25467_ );
nor  ( new_n25471_, new_n25470_, new_n25466_ );
nor  ( new_n25472_, new_n25471_, new_n25461_ );
or   ( new_n25473_, new_n25472_, new_n25460_ );
xor  ( new_n25474_, new_n25292_, new_n25287_ );
xor  ( new_n25475_, new_n25474_, new_n25295_ );
not  ( new_n25476_, new_n25475_ );
or   ( new_n25477_, new_n283_, new_n24927_ );
or   ( new_n25478_, new_n286_, new_n24543_ );
and  ( new_n25479_, new_n25478_, new_n25477_ );
xor  ( new_n25480_, new_n25479_, new_n278_ );
or   ( new_n25481_, new_n299_, new_n25048_ );
or   ( new_n25482_, new_n302_, new_n24925_ );
and  ( new_n25483_, new_n25482_, new_n25481_ );
xor  ( new_n25484_, new_n25483_, new_n293_ );
or   ( new_n25485_, new_n25484_, new_n25480_ );
not  ( new_n25486_, RIbb32838_168 );
or   ( new_n25487_, new_n268_, new_n25486_ );
or   ( new_n25488_, new_n271_, new_n25288_ );
and  ( new_n25489_, new_n25488_, new_n25487_ );
xor  ( new_n25490_, new_n25489_, new_n263_ );
and  ( new_n25491_, new_n25484_, new_n25480_ );
or   ( new_n25492_, new_n25491_, new_n25490_ );
and  ( new_n25493_, new_n25492_, new_n25485_ );
or   ( new_n25494_, new_n25493_, new_n25476_ );
or   ( new_n25495_, new_n2425_, new_n21792_ );
or   ( new_n25496_, new_n2427_, new_n21751_ );
and  ( new_n25497_, new_n25496_, new_n25495_ );
xor  ( new_n25498_, new_n25497_, new_n2121_ );
or   ( new_n25499_, new_n2122_, new_n21840_ );
or   ( new_n25500_, new_n2124_, new_n21842_ );
and  ( new_n25501_, new_n25500_, new_n25499_ );
xor  ( new_n25502_, new_n25501_, new_n1843_ );
nor  ( new_n25503_, new_n25502_, new_n25498_ );
or   ( new_n25504_, new_n1844_, new_n22098_ );
or   ( new_n25505_, new_n1846_, new_n21847_ );
and  ( new_n25506_, new_n25505_, new_n25504_ );
xor  ( new_n25507_, new_n25506_, new_n1585_ );
nand ( new_n25508_, new_n25502_, new_n25498_ );
and  ( new_n25509_, new_n25508_, new_n25507_ );
or   ( new_n25510_, new_n25509_, new_n25503_ );
or   ( new_n25511_, new_n3896_, new_n21701_ );
or   ( new_n25512_, new_n3898_, new_n21703_ );
and  ( new_n25513_, new_n25512_, new_n25511_ );
xor  ( new_n25514_, new_n25513_, new_n3460_ );
nand ( new_n25515_, new_n25514_, new_n4295_ );
nor  ( new_n25516_, new_n25514_, new_n4295_ );
or   ( new_n25517_, new_n4302_, new_n21694_ );
or   ( new_n25518_, new_n4304_, new_n21696_ );
and  ( new_n25519_, new_n25518_, new_n25517_ );
xor  ( new_n25520_, new_n25519_, new_n3894_ );
or   ( new_n25521_, new_n25520_, new_n25516_ );
and  ( new_n25522_, new_n25521_, new_n25515_ );
nand ( new_n25523_, new_n25522_, new_n25510_ );
nor  ( new_n25524_, new_n25522_, new_n25510_ );
or   ( new_n25525_, new_n3461_, new_n21672_ );
or   ( new_n25526_, new_n3463_, new_n21674_ );
and  ( new_n25527_, new_n25526_, new_n25525_ );
xor  ( new_n25528_, new_n25527_, new_n3116_ );
or   ( new_n25529_, new_n3117_, new_n21678_ );
or   ( new_n25530_, new_n3119_, new_n21680_ );
and  ( new_n25531_, new_n25530_, new_n25529_ );
xor  ( new_n25532_, new_n25531_, new_n2800_ );
or   ( new_n25533_, new_n25532_, new_n25528_ );
or   ( new_n25534_, new_n2807_, new_n21685_ );
or   ( new_n25535_, new_n2809_, new_n21687_ );
and  ( new_n25536_, new_n25535_, new_n25534_ );
xor  ( new_n25537_, new_n25536_, new_n2424_ );
and  ( new_n25538_, new_n25532_, new_n25528_ );
or   ( new_n25539_, new_n25538_, new_n25537_ );
and  ( new_n25540_, new_n25539_, new_n25533_ );
or   ( new_n25541_, new_n25540_, new_n25524_ );
and  ( new_n25542_, new_n25541_, new_n25523_ );
or   ( new_n25543_, new_n25542_, new_n25494_ );
and  ( new_n25544_, new_n25542_, new_n25494_ );
or   ( new_n25545_, new_n1593_, new_n22207_ );
or   ( new_n25546_, new_n1595_, new_n22129_ );
and  ( new_n25547_, new_n25546_, new_n25545_ );
xor  ( new_n25548_, new_n25547_, new_n1358_ );
or   ( new_n25549_, new_n1364_, new_n22423_ );
or   ( new_n25550_, new_n1366_, new_n22304_ );
and  ( new_n25551_, new_n25550_, new_n25549_ );
xor  ( new_n25552_, new_n25551_, new_n1129_ );
or   ( new_n25553_, new_n25552_, new_n25548_ );
or   ( new_n25554_, new_n1135_, new_n22641_ );
or   ( new_n25555_, new_n1137_, new_n22590_ );
and  ( new_n25556_, new_n25555_, new_n25554_ );
xor  ( new_n25557_, new_n25556_, new_n896_ );
and  ( new_n25558_, new_n25552_, new_n25548_ );
or   ( new_n25559_, new_n25558_, new_n25557_ );
and  ( new_n25560_, new_n25559_, new_n25553_ );
or   ( new_n25561_, new_n409_, new_n23733_ );
or   ( new_n25562_, new_n411_, new_n23554_ );
and  ( new_n25563_, new_n25562_, new_n25561_ );
xor  ( new_n25564_, new_n25563_, new_n328_ );
or   ( new_n25565_, new_n337_, new_n24006_ );
or   ( new_n25566_, new_n340_, new_n23895_ );
and  ( new_n25567_, new_n25566_, new_n25565_ );
xor  ( new_n25568_, new_n25567_, new_n332_ );
or   ( new_n25569_, new_n25568_, new_n25564_ );
or   ( new_n25570_, new_n317_, new_n24418_ );
or   ( new_n25571_, new_n320_, new_n24227_ );
and  ( new_n25572_, new_n25571_, new_n25570_ );
xor  ( new_n25573_, new_n25572_, new_n312_ );
and  ( new_n25574_, new_n25568_, new_n25564_ );
or   ( new_n25575_, new_n25574_, new_n25573_ );
and  ( new_n25576_, new_n25575_, new_n25569_ );
nor  ( new_n25577_, new_n25576_, new_n25560_ );
and  ( new_n25578_, new_n25576_, new_n25560_ );
or   ( new_n25579_, new_n897_, new_n22975_ );
or   ( new_n25580_, new_n899_, new_n22829_ );
and  ( new_n25581_, new_n25580_, new_n25579_ );
xor  ( new_n25582_, new_n25581_, new_n748_ );
or   ( new_n25583_, new_n755_, new_n23166_ );
or   ( new_n25584_, new_n757_, new_n22973_ );
and  ( new_n25585_, new_n25584_, new_n25583_ );
xor  ( new_n25586_, new_n25585_, new_n523_ );
nor  ( new_n25587_, new_n25586_, new_n25582_ );
or   ( new_n25588_, new_n524_, new_n23370_ );
or   ( new_n25589_, new_n526_, new_n23252_ );
and  ( new_n25590_, new_n25589_, new_n25588_ );
xor  ( new_n25591_, new_n25590_, new_n403_ );
and  ( new_n25592_, new_n25586_, new_n25582_ );
nor  ( new_n25593_, new_n25592_, new_n25591_ );
nor  ( new_n25594_, new_n25593_, new_n25587_ );
nor  ( new_n25595_, new_n25594_, new_n25578_ );
nor  ( new_n25596_, new_n25595_, new_n25577_ );
or   ( new_n25597_, new_n25596_, new_n25544_ );
and  ( new_n25598_, new_n25597_, new_n25543_ );
nor  ( new_n25599_, new_n25598_, new_n25473_ );
nand ( new_n25600_, new_n25598_, new_n25473_ );
xor  ( new_n25601_, new_n25123_, new_n3895_ );
xor  ( new_n25602_, new_n25601_, new_n25129_ );
xnor ( new_n25603_, new_n25381_, new_n25379_ );
xor  ( new_n25604_, new_n25603_, new_n25385_ );
nor  ( new_n25605_, new_n25604_, new_n25602_ );
nand ( new_n25606_, new_n25604_, new_n25602_ );
xor  ( new_n25607_, new_n25300_, new_n25298_ );
xor  ( new_n25608_, new_n25607_, new_n25304_ );
and  ( new_n25609_, new_n25608_, new_n25606_ );
or   ( new_n25610_, new_n25609_, new_n25605_ );
and  ( new_n25611_, new_n25610_, new_n25600_ );
or   ( new_n25612_, new_n25611_, new_n25599_ );
xor  ( new_n25613_, new_n25367_, new_n25365_ );
xor  ( new_n25614_, new_n25613_, new_n25371_ );
xor  ( new_n25615_, new_n25306_, new_n25283_ );
xor  ( new_n25616_, new_n25615_, new_n25361_ );
or   ( new_n25617_, new_n25616_, new_n25614_ );
and  ( new_n25618_, new_n25616_, new_n25614_ );
xor  ( new_n25619_, new_n25387_, new_n25377_ );
xor  ( new_n25620_, new_n25619_, new_n25391_ );
or   ( new_n25621_, new_n25620_, new_n25618_ );
and  ( new_n25622_, new_n25621_, new_n25617_ );
and  ( new_n25623_, new_n25622_, new_n25612_ );
nor  ( new_n25624_, new_n25622_, new_n25612_ );
not  ( new_n25625_, new_n25624_ );
xor  ( new_n25626_, new_n25117_, new_n25065_ );
xor  ( new_n25627_, new_n25626_, new_n25168_ );
and  ( new_n25628_, new_n25627_, new_n25625_ );
nor  ( new_n25629_, new_n25628_, new_n25623_ );
or   ( new_n25630_, new_n25629_, new_n25447_ );
and  ( new_n25631_, new_n25630_, new_n25446_ );
xor  ( new_n25632_, new_n25414_, new_n25233_ );
nand ( new_n25633_, new_n25632_, new_n25428_ );
or   ( new_n25634_, new_n25430_, new_n25416_ );
and  ( new_n25635_, new_n25634_, new_n25633_ );
nand ( new_n25636_, new_n25635_, new_n25631_ );
nor  ( new_n25637_, new_n25635_, new_n25631_ );
xor  ( new_n25638_, new_n25206_, new_n25043_ );
xor  ( new_n25639_, new_n25638_, new_n25219_ );
or   ( new_n25640_, new_n25639_, new_n25637_ );
and  ( new_n25641_, new_n25640_, new_n25636_ );
nor  ( new_n25642_, new_n25641_, new_n25437_ );
xor  ( new_n25643_, new_n25635_, new_n25631_ );
xor  ( new_n25644_, new_n25643_, new_n25639_ );
xor  ( new_n25645_, new_n25409_, new_n25411_ );
xor  ( new_n25646_, new_n25645_, new_n25410_ );
xor  ( new_n25647_, new_n25616_, new_n25614_ );
xor  ( new_n25648_, new_n25647_, new_n25620_ );
xnor ( new_n25649_, new_n25263_, new_n25249_ );
xor  ( new_n25650_, new_n25649_, new_n25281_ );
xor  ( new_n25651_, new_n25340_, new_n25324_ );
xor  ( new_n25652_, new_n25651_, new_n25359_ );
or   ( new_n25653_, new_n25652_, new_n25650_ );
and  ( new_n25654_, new_n25652_, new_n25650_ );
xor  ( new_n25655_, new_n25604_, new_n25602_ );
xor  ( new_n25656_, new_n25655_, new_n25608_ );
or   ( new_n25657_, new_n25656_, new_n25654_ );
and  ( new_n25658_, new_n25657_, new_n25653_ );
or   ( new_n25659_, new_n25658_, new_n25648_ );
and  ( new_n25660_, new_n25658_, new_n25648_ );
xor  ( new_n25661_, new_n25453_, new_n25451_ );
xor  ( new_n25662_, new_n25661_, new_n25457_ );
xor  ( new_n25663_, new_n25502_, new_n25498_ );
xor  ( new_n25664_, new_n25663_, new_n25507_ );
xnor ( new_n25665_, new_n25552_, new_n25548_ );
xor  ( new_n25666_, new_n25665_, new_n25557_ );
or   ( new_n25667_, new_n25666_, new_n25664_ );
and  ( new_n25668_, new_n25666_, new_n25664_ );
xor  ( new_n25669_, new_n25532_, new_n25528_ );
xnor ( new_n25670_, new_n25669_, new_n25537_ );
or   ( new_n25671_, new_n25670_, new_n25668_ );
and  ( new_n25672_, new_n25671_, new_n25667_ );
or   ( new_n25673_, new_n25672_, new_n25662_ );
and  ( new_n25674_, new_n25672_, new_n25662_ );
xnor ( new_n25675_, new_n25568_, new_n25564_ );
xor  ( new_n25676_, new_n25675_, new_n25573_ );
xnor ( new_n25677_, new_n25586_, new_n25582_ );
xor  ( new_n25678_, new_n25677_, new_n25591_ );
nor  ( new_n25679_, new_n25678_, new_n25676_ );
and  ( new_n25680_, new_n25678_, new_n25676_ );
xor  ( new_n25681_, new_n25484_, new_n25480_ );
xnor ( new_n25682_, new_n25681_, new_n25490_ );
nor  ( new_n25683_, new_n25682_, new_n25680_ );
nor  ( new_n25684_, new_n25683_, new_n25679_ );
or   ( new_n25685_, new_n25684_, new_n25674_ );
and  ( new_n25686_, new_n25685_, new_n25673_ );
xor  ( new_n25687_, new_n25576_, new_n25560_ );
xor  ( new_n25688_, new_n25687_, new_n25594_ );
xnor ( new_n25689_, new_n25465_, new_n25463_ );
xor  ( new_n25690_, new_n25689_, new_n25469_ );
nand ( new_n25691_, new_n25690_, new_n25688_ );
nor  ( new_n25692_, new_n25690_, new_n25688_ );
xor  ( new_n25693_, new_n25493_, new_n25476_ );
or   ( new_n25694_, new_n25693_, new_n25692_ );
and  ( new_n25695_, new_n25694_, new_n25691_ );
and  ( new_n25696_, new_n25695_, new_n25686_ );
or   ( new_n25697_, new_n25695_, new_n25686_ );
or   ( new_n25698_, new_n897_, new_n22973_ );
or   ( new_n25699_, new_n899_, new_n22975_ );
and  ( new_n25700_, new_n25699_, new_n25698_ );
xor  ( new_n25701_, new_n25700_, new_n748_ );
or   ( new_n25702_, new_n755_, new_n23252_ );
or   ( new_n25703_, new_n757_, new_n23166_ );
and  ( new_n25704_, new_n25703_, new_n25702_ );
xor  ( new_n25705_, new_n25704_, new_n523_ );
or   ( new_n25706_, new_n25705_, new_n25701_ );
and  ( new_n25707_, new_n25705_, new_n25701_ );
or   ( new_n25708_, new_n524_, new_n23554_ );
or   ( new_n25709_, new_n526_, new_n23370_ );
and  ( new_n25710_, new_n25709_, new_n25708_ );
xor  ( new_n25711_, new_n25710_, new_n403_ );
or   ( new_n25712_, new_n25711_, new_n25707_ );
and  ( new_n25713_, new_n25712_, new_n25706_ );
or   ( new_n25714_, new_n409_, new_n23895_ );
or   ( new_n25715_, new_n411_, new_n23733_ );
and  ( new_n25716_, new_n25715_, new_n25714_ );
xor  ( new_n25717_, new_n25716_, new_n328_ );
or   ( new_n25718_, new_n337_, new_n24227_ );
or   ( new_n25719_, new_n340_, new_n24006_ );
and  ( new_n25720_, new_n25719_, new_n25718_ );
xor  ( new_n25721_, new_n25720_, new_n332_ );
or   ( new_n25722_, new_n25721_, new_n25717_ );
and  ( new_n25723_, new_n25721_, new_n25717_ );
or   ( new_n25724_, new_n317_, new_n24543_ );
or   ( new_n25725_, new_n320_, new_n24418_ );
and  ( new_n25726_, new_n25725_, new_n25724_ );
xor  ( new_n25727_, new_n25726_, new_n312_ );
or   ( new_n25728_, new_n25727_, new_n25723_ );
and  ( new_n25729_, new_n25728_, new_n25722_ );
or   ( new_n25730_, new_n25729_, new_n25713_ );
and  ( new_n25731_, new_n25729_, new_n25713_ );
or   ( new_n25732_, new_n1593_, new_n22304_ );
or   ( new_n25733_, new_n1595_, new_n22207_ );
and  ( new_n25734_, new_n25733_, new_n25732_ );
xor  ( new_n25735_, new_n25734_, new_n1358_ );
or   ( new_n25736_, new_n1364_, new_n22590_ );
or   ( new_n25737_, new_n1366_, new_n22423_ );
and  ( new_n25738_, new_n25737_, new_n25736_ );
xor  ( new_n25739_, new_n25738_, new_n1129_ );
nor  ( new_n25740_, new_n25739_, new_n25735_ );
and  ( new_n25741_, new_n25739_, new_n25735_ );
or   ( new_n25742_, new_n1135_, new_n22829_ );
or   ( new_n25743_, new_n1137_, new_n22641_ );
and  ( new_n25744_, new_n25743_, new_n25742_ );
xor  ( new_n25745_, new_n25744_, new_n896_ );
nor  ( new_n25746_, new_n25745_, new_n25741_ );
nor  ( new_n25747_, new_n25746_, new_n25740_ );
or   ( new_n25748_, new_n25747_, new_n25731_ );
and  ( new_n25749_, new_n25748_, new_n25730_ );
or   ( new_n25750_, new_n4302_, new_n21703_ );
or   ( new_n25751_, new_n4304_, new_n21694_ );
and  ( new_n25752_, new_n25751_, new_n25750_ );
xor  ( new_n25753_, new_n25752_, new_n3894_ );
and  ( new_n25754_, new_n4543_, RIbb315f0_129 );
xor  ( new_n25755_, new_n25754_, new_n4295_ );
nand ( new_n25756_, new_n25755_, new_n25753_ );
nor  ( new_n25757_, new_n25755_, new_n25753_ );
or   ( new_n25758_, new_n3896_, new_n21674_ );
or   ( new_n25759_, new_n3898_, new_n21701_ );
and  ( new_n25760_, new_n25759_, new_n25758_ );
xor  ( new_n25761_, new_n25760_, new_n3460_ );
or   ( new_n25762_, new_n25761_, new_n25757_ );
and  ( new_n25763_, new_n25762_, new_n25756_ );
or   ( new_n25764_, new_n2425_, new_n21842_ );
or   ( new_n25765_, new_n2427_, new_n21792_ );
and  ( new_n25766_, new_n25765_, new_n25764_ );
xor  ( new_n25767_, new_n25766_, new_n2121_ );
or   ( new_n25768_, new_n2122_, new_n21847_ );
or   ( new_n25769_, new_n2124_, new_n21840_ );
and  ( new_n25770_, new_n25769_, new_n25768_ );
xor  ( new_n25771_, new_n25770_, new_n1843_ );
or   ( new_n25772_, new_n25771_, new_n25767_ );
and  ( new_n25773_, new_n25771_, new_n25767_ );
or   ( new_n25774_, new_n1844_, new_n22129_ );
or   ( new_n25775_, new_n1846_, new_n22098_ );
and  ( new_n25776_, new_n25775_, new_n25774_ );
xor  ( new_n25777_, new_n25776_, new_n1586_ );
or   ( new_n25778_, new_n25777_, new_n25773_ );
and  ( new_n25779_, new_n25778_, new_n25772_ );
or   ( new_n25780_, new_n25779_, new_n25763_ );
and  ( new_n25781_, new_n25779_, new_n25763_ );
or   ( new_n25782_, new_n3461_, new_n21680_ );
or   ( new_n25783_, new_n3463_, new_n21672_ );
and  ( new_n25784_, new_n25783_, new_n25782_ );
xor  ( new_n25785_, new_n25784_, new_n3116_ );
or   ( new_n25786_, new_n3117_, new_n21687_ );
or   ( new_n25787_, new_n3119_, new_n21678_ );
and  ( new_n25788_, new_n25787_, new_n25786_ );
xor  ( new_n25789_, new_n25788_, new_n2800_ );
nor  ( new_n25790_, new_n25789_, new_n25785_ );
and  ( new_n25791_, new_n25789_, new_n25785_ );
or   ( new_n25792_, new_n2807_, new_n21751_ );
or   ( new_n25793_, new_n2809_, new_n21685_ );
and  ( new_n25794_, new_n25793_, new_n25792_ );
xor  ( new_n25795_, new_n25794_, new_n2424_ );
nor  ( new_n25796_, new_n25795_, new_n25791_ );
nor  ( new_n25797_, new_n25796_, new_n25790_ );
or   ( new_n25798_, new_n25797_, new_n25781_ );
and  ( new_n25799_, new_n25798_, new_n25780_ );
nor  ( new_n25800_, new_n25799_, new_n25749_ );
nand ( new_n25801_, new_n25799_, new_n25749_ );
and  ( new_n25802_, RIbb32928_170, RIbb2f610_1 );
or   ( new_n25803_, new_n283_, new_n24925_ );
or   ( new_n25804_, new_n286_, new_n24927_ );
and  ( new_n25805_, new_n25804_, new_n25803_ );
xor  ( new_n25806_, new_n25805_, new_n278_ );
or   ( new_n25807_, new_n299_, new_n25288_ );
or   ( new_n25808_, new_n302_, new_n25048_ );
and  ( new_n25809_, new_n25808_, new_n25807_ );
xor  ( new_n25810_, new_n25809_, new_n293_ );
or   ( new_n25811_, new_n25810_, new_n25806_ );
and  ( new_n25812_, new_n25810_, new_n25806_ );
not  ( new_n25813_, RIbb328b0_169 );
or   ( new_n25814_, new_n268_, new_n25813_ );
or   ( new_n25815_, new_n271_, new_n25486_ );
and  ( new_n25816_, new_n25815_, new_n25814_ );
xor  ( new_n25817_, new_n25816_, new_n263_ );
or   ( new_n25818_, new_n25817_, new_n25812_ );
and  ( new_n25819_, new_n25818_, new_n25811_ );
nor  ( new_n25820_, new_n25819_, new_n25802_ );
and  ( new_n25821_, new_n25819_, new_n25802_ );
and  ( new_n25822_, RIbb328b0_169, RIbb2f610_1 );
nor  ( new_n25823_, new_n25822_, new_n25821_ );
or   ( new_n25824_, new_n25823_, new_n25820_ );
and  ( new_n25825_, new_n25824_, new_n25801_ );
or   ( new_n25826_, new_n25825_, new_n25800_ );
and  ( new_n25827_, new_n25826_, new_n25697_ );
or   ( new_n25828_, new_n25827_, new_n25696_ );
or   ( new_n25829_, new_n25828_, new_n25660_ );
and  ( new_n25830_, new_n25829_, new_n25659_ );
xor  ( new_n25831_, new_n25622_, new_n25612_ );
xor  ( new_n25832_, new_n25831_, new_n25627_ );
or   ( new_n25833_, new_n25832_, new_n25830_ );
nand ( new_n25834_, new_n25832_, new_n25830_ );
xor  ( new_n25835_, new_n25442_, new_n25440_ );
nand ( new_n25836_, new_n25835_, new_n25834_ );
and  ( new_n25837_, new_n25836_, new_n25833_ );
or   ( new_n25838_, new_n25837_, new_n25646_ );
and  ( new_n25839_, new_n25837_, new_n25646_ );
xor  ( new_n25840_, new_n25445_, new_n25443_ );
xnor ( new_n25841_, new_n25840_, new_n25629_ );
or   ( new_n25842_, new_n25841_, new_n25839_ );
and  ( new_n25843_, new_n25842_, new_n25838_ );
nor  ( new_n25844_, new_n25843_, new_n25644_ );
xnor ( new_n25845_, new_n25837_, new_n25646_ );
xor  ( new_n25846_, new_n25845_, new_n25841_ );
or   ( new_n25847_, new_n524_, new_n23733_ );
or   ( new_n25848_, new_n526_, new_n23554_ );
and  ( new_n25849_, new_n25848_, new_n25847_ );
xor  ( new_n25850_, new_n25849_, new_n403_ );
or   ( new_n25851_, new_n409_, new_n24006_ );
or   ( new_n25852_, new_n411_, new_n23895_ );
and  ( new_n25853_, new_n25852_, new_n25851_ );
xor  ( new_n25854_, new_n25853_, new_n328_ );
or   ( new_n25855_, new_n25854_, new_n25850_ );
and  ( new_n25856_, new_n25854_, new_n25850_ );
or   ( new_n25857_, new_n337_, new_n24418_ );
or   ( new_n25858_, new_n340_, new_n24227_ );
and  ( new_n25859_, new_n25858_, new_n25857_ );
xor  ( new_n25860_, new_n25859_, new_n332_ );
or   ( new_n25861_, new_n25860_, new_n25856_ );
and  ( new_n25862_, new_n25861_, new_n25855_ );
or   ( new_n25863_, new_n1844_, new_n22207_ );
or   ( new_n25864_, new_n1846_, new_n22129_ );
and  ( new_n25865_, new_n25864_, new_n25863_ );
xor  ( new_n25866_, new_n25865_, new_n1586_ );
or   ( new_n25867_, new_n1593_, new_n22423_ );
or   ( new_n25868_, new_n1595_, new_n22304_ );
and  ( new_n25869_, new_n25868_, new_n25867_ );
xor  ( new_n25870_, new_n25869_, new_n1358_ );
or   ( new_n25871_, new_n25870_, new_n25866_ );
and  ( new_n25872_, new_n25870_, new_n25866_ );
or   ( new_n25873_, new_n1364_, new_n22641_ );
or   ( new_n25874_, new_n1366_, new_n22590_ );
and  ( new_n25875_, new_n25874_, new_n25873_ );
xor  ( new_n25876_, new_n25875_, new_n1129_ );
or   ( new_n25877_, new_n25876_, new_n25872_ );
and  ( new_n25878_, new_n25877_, new_n25871_ );
or   ( new_n25879_, new_n25878_, new_n25862_ );
and  ( new_n25880_, new_n25878_, new_n25862_ );
or   ( new_n25881_, new_n1135_, new_n22975_ );
or   ( new_n25882_, new_n1137_, new_n22829_ );
and  ( new_n25883_, new_n25882_, new_n25881_ );
xor  ( new_n25884_, new_n25883_, new_n896_ );
or   ( new_n25885_, new_n897_, new_n23166_ );
or   ( new_n25886_, new_n899_, new_n22973_ );
and  ( new_n25887_, new_n25886_, new_n25885_ );
xor  ( new_n25888_, new_n25887_, new_n748_ );
or   ( new_n25889_, new_n25888_, new_n25884_ );
and  ( new_n25890_, new_n25888_, new_n25884_ );
or   ( new_n25891_, new_n755_, new_n23370_ );
or   ( new_n25892_, new_n757_, new_n23252_ );
and  ( new_n25893_, new_n25892_, new_n25891_ );
xor  ( new_n25894_, new_n25893_, new_n523_ );
or   ( new_n25895_, new_n25894_, new_n25890_ );
and  ( new_n25896_, new_n25895_, new_n25889_ );
or   ( new_n25897_, new_n25896_, new_n25880_ );
and  ( new_n25898_, new_n25897_, new_n25879_ );
or   ( new_n25899_, new_n2807_, new_n21792_ );
or   ( new_n25900_, new_n2809_, new_n21751_ );
and  ( new_n25901_, new_n25900_, new_n25899_ );
xor  ( new_n25902_, new_n25901_, new_n2424_ );
or   ( new_n25903_, new_n2425_, new_n21840_ );
or   ( new_n25904_, new_n2427_, new_n21842_ );
and  ( new_n25905_, new_n25904_, new_n25903_ );
xor  ( new_n25906_, new_n25905_, new_n2121_ );
nor  ( new_n25907_, new_n25906_, new_n25902_ );
nand ( new_n25908_, new_n25906_, new_n25902_ );
or   ( new_n25909_, new_n2122_, new_n22098_ );
or   ( new_n25910_, new_n2124_, new_n21847_ );
and  ( new_n25911_, new_n25910_, new_n25909_ );
xor  ( new_n25912_, new_n25911_, new_n1842_ );
and  ( new_n25913_, new_n25912_, new_n25908_ );
or   ( new_n25914_, new_n25913_, new_n25907_ );
or   ( new_n25915_, new_n4709_, new_n21694_ );
or   ( new_n25916_, new_n4711_, new_n21696_ );
and  ( new_n25917_, new_n25916_, new_n25915_ );
xor  ( new_n25918_, new_n25917_, new_n4295_ );
nand ( new_n25919_, new_n25918_, new_n4708_ );
nor  ( new_n25920_, new_n25918_, new_n4708_ );
or   ( new_n25921_, new_n4302_, new_n21701_ );
or   ( new_n25922_, new_n4304_, new_n21703_ );
and  ( new_n25923_, new_n25922_, new_n25921_ );
xor  ( new_n25924_, new_n25923_, new_n3894_ );
or   ( new_n25925_, new_n25924_, new_n25920_ );
and  ( new_n25926_, new_n25925_, new_n25919_ );
nand ( new_n25927_, new_n25926_, new_n25914_ );
nor  ( new_n25928_, new_n25926_, new_n25914_ );
or   ( new_n25929_, new_n3896_, new_n21672_ );
or   ( new_n25930_, new_n3898_, new_n21674_ );
and  ( new_n25931_, new_n25930_, new_n25929_ );
xor  ( new_n25932_, new_n25931_, new_n3460_ );
or   ( new_n25933_, new_n3461_, new_n21678_ );
or   ( new_n25934_, new_n3463_, new_n21680_ );
and  ( new_n25935_, new_n25934_, new_n25933_ );
xor  ( new_n25936_, new_n25935_, new_n3116_ );
nor  ( new_n25937_, new_n25936_, new_n25932_ );
and  ( new_n25938_, new_n25936_, new_n25932_ );
or   ( new_n25939_, new_n3117_, new_n21685_ );
or   ( new_n25940_, new_n3119_, new_n21687_ );
and  ( new_n25941_, new_n25940_, new_n25939_ );
xor  ( new_n25942_, new_n25941_, new_n2800_ );
nor  ( new_n25943_, new_n25942_, new_n25938_ );
nor  ( new_n25944_, new_n25943_, new_n25937_ );
or   ( new_n25945_, new_n25944_, new_n25928_ );
and  ( new_n25946_, new_n25945_, new_n25927_ );
nor  ( new_n25947_, new_n25946_, new_n25898_ );
nand ( new_n25948_, new_n25946_, new_n25898_ );
not  ( new_n25949_, new_n25802_ );
or   ( new_n25950_, new_n317_, new_n24927_ );
or   ( new_n25951_, new_n320_, new_n24543_ );
and  ( new_n25952_, new_n25951_, new_n25950_ );
xor  ( new_n25953_, new_n25952_, new_n312_ );
or   ( new_n25954_, new_n283_, new_n25048_ );
or   ( new_n25955_, new_n286_, new_n24925_ );
and  ( new_n25956_, new_n25955_, new_n25954_ );
xor  ( new_n25957_, new_n25956_, new_n278_ );
or   ( new_n25958_, new_n25957_, new_n25953_ );
and  ( new_n25959_, new_n25957_, new_n25953_ );
or   ( new_n25960_, new_n299_, new_n25486_ );
or   ( new_n25961_, new_n302_, new_n25288_ );
and  ( new_n25962_, new_n25961_, new_n25960_ );
xor  ( new_n25963_, new_n25962_, new_n293_ );
or   ( new_n25964_, new_n25963_, new_n25959_ );
and  ( new_n25965_, new_n25964_, new_n25958_ );
nor  ( new_n25966_, new_n25965_, new_n25949_ );
nand ( new_n25967_, new_n25965_, new_n25949_ );
xor  ( new_n25968_, new_n25810_, new_n25806_ );
xnor ( new_n25969_, new_n25968_, new_n25817_ );
and  ( new_n25970_, new_n25969_, new_n25967_ );
or   ( new_n25971_, new_n25970_, new_n25966_ );
and  ( new_n25972_, new_n25971_, new_n25948_ );
or   ( new_n25973_, new_n25972_, new_n25947_ );
xor  ( new_n25974_, new_n25514_, new_n4295_ );
xor  ( new_n25975_, new_n25974_, new_n25520_ );
xnor ( new_n25976_, new_n25721_, new_n25717_ );
xor  ( new_n25977_, new_n25976_, new_n25727_ );
xnor ( new_n25978_, new_n25705_, new_n25701_ );
xor  ( new_n25979_, new_n25978_, new_n25711_ );
or   ( new_n25980_, new_n25979_, new_n25977_ );
and  ( new_n25981_, new_n25979_, new_n25977_ );
xor  ( new_n25982_, new_n25739_, new_n25735_ );
xnor ( new_n25983_, new_n25982_, new_n25745_ );
or   ( new_n25984_, new_n25983_, new_n25981_ );
and  ( new_n25985_, new_n25984_, new_n25980_ );
or   ( new_n25986_, new_n25985_, new_n25975_ );
and  ( new_n25987_, new_n25985_, new_n25975_ );
xnor ( new_n25988_, new_n25771_, new_n25767_ );
xor  ( new_n25989_, new_n25988_, new_n25777_ );
xnor ( new_n25990_, new_n25755_, new_n25753_ );
xor  ( new_n25991_, new_n25990_, new_n25761_ );
nor  ( new_n25992_, new_n25991_, new_n25989_ );
and  ( new_n25993_, new_n25991_, new_n25989_ );
xor  ( new_n25994_, new_n25789_, new_n25785_ );
xnor ( new_n25995_, new_n25994_, new_n25795_ );
nor  ( new_n25996_, new_n25995_, new_n25993_ );
nor  ( new_n25997_, new_n25996_, new_n25992_ );
or   ( new_n25998_, new_n25997_, new_n25987_ );
and  ( new_n25999_, new_n25998_, new_n25986_ );
or   ( new_n26000_, new_n25999_, new_n25973_ );
and  ( new_n26001_, new_n25999_, new_n25973_ );
xor  ( new_n26002_, new_n25819_, new_n25802_ );
xor  ( new_n26003_, new_n26002_, new_n25822_ );
xnor ( new_n26004_, new_n25678_, new_n25676_ );
xor  ( new_n26005_, new_n26004_, new_n25682_ );
and  ( new_n26006_, new_n26005_, new_n26003_ );
nor  ( new_n26007_, new_n26005_, new_n26003_ );
xor  ( new_n26008_, new_n25666_, new_n25664_ );
xnor ( new_n26009_, new_n26008_, new_n25670_ );
not  ( new_n26010_, new_n26009_ );
nor  ( new_n26011_, new_n26010_, new_n26007_ );
nor  ( new_n26012_, new_n26011_, new_n26006_ );
or   ( new_n26013_, new_n26012_, new_n26001_ );
and  ( new_n26014_, new_n26013_, new_n26000_ );
xor  ( new_n26015_, new_n25522_, new_n25510_ );
xor  ( new_n26016_, new_n26015_, new_n25540_ );
xnor ( new_n26017_, new_n25672_, new_n25662_ );
xor  ( new_n26018_, new_n26017_, new_n25684_ );
nand ( new_n26019_, new_n26018_, new_n26016_ );
or   ( new_n26020_, new_n26018_, new_n26016_ );
xor  ( new_n26021_, new_n25690_, new_n25688_ );
xnor ( new_n26022_, new_n26021_, new_n25693_ );
nand ( new_n26023_, new_n26022_, new_n26020_ );
and  ( new_n26024_, new_n26023_, new_n26019_ );
and  ( new_n26025_, new_n26024_, new_n26014_ );
or   ( new_n26026_, new_n26024_, new_n26014_ );
xor  ( new_n26027_, new_n25459_, new_n25449_ );
xor  ( new_n26028_, new_n26027_, new_n25471_ );
and  ( new_n26029_, new_n26028_, new_n26026_ );
or   ( new_n26030_, new_n26029_, new_n26025_ );
xor  ( new_n26031_, new_n25695_, new_n25686_ );
xor  ( new_n26032_, new_n26031_, new_n25826_ );
xnor ( new_n26033_, new_n25542_, new_n25494_ );
xor  ( new_n26034_, new_n26033_, new_n25596_ );
or   ( new_n26035_, new_n26034_, new_n26032_ );
and  ( new_n26036_, new_n26034_, new_n26032_ );
xor  ( new_n26037_, new_n25652_, new_n25650_ );
xor  ( new_n26038_, new_n26037_, new_n25656_ );
or   ( new_n26039_, new_n26038_, new_n26036_ );
and  ( new_n26040_, new_n26039_, new_n26035_ );
or   ( new_n26041_, new_n26040_, new_n26030_ );
and  ( new_n26042_, new_n26040_, new_n26030_ );
xor  ( new_n26043_, new_n25598_, new_n25473_ );
xor  ( new_n26044_, new_n26043_, new_n25610_ );
or   ( new_n26045_, new_n26044_, new_n26042_ );
and  ( new_n26046_, new_n26045_, new_n26041_ );
xor  ( new_n26047_, new_n26040_, new_n26030_ );
xor  ( new_n26048_, new_n26047_, new_n26044_ );
xor  ( new_n26049_, new_n25799_, new_n25749_ );
xor  ( new_n26050_, new_n26049_, new_n25824_ );
xnor ( new_n26051_, new_n25779_, new_n25763_ );
xor  ( new_n26052_, new_n26051_, new_n25797_ );
xnor ( new_n26053_, new_n25729_, new_n25713_ );
xor  ( new_n26054_, new_n26053_, new_n25747_ );
or   ( new_n26055_, new_n26054_, new_n26052_ );
and  ( new_n26056_, new_n26054_, new_n26052_ );
xor  ( new_n26057_, new_n26005_, new_n26003_ );
xor  ( new_n26058_, new_n26057_, new_n26010_ );
or   ( new_n26059_, new_n26058_, new_n26056_ );
and  ( new_n26060_, new_n26059_, new_n26055_ );
or   ( new_n26061_, new_n26060_, new_n26050_ );
and  ( new_n26062_, new_n26060_, new_n26050_ );
not  ( new_n26063_, RIbb329a0_171 );
or   ( new_n26064_, new_n26063_, new_n260_ );
xnor ( new_n26065_, new_n25957_, new_n25953_ );
xor  ( new_n26066_, new_n26065_, new_n25963_ );
and  ( new_n26067_, new_n26066_, new_n26064_ );
or   ( new_n26068_, new_n26066_, new_n26064_ );
xnor ( new_n26069_, new_n25854_, new_n25850_ );
xor  ( new_n26070_, new_n26069_, new_n25860_ );
and  ( new_n26071_, new_n26070_, new_n26068_ );
or   ( new_n26072_, new_n26071_, new_n26067_ );
xnor ( new_n26073_, new_n25870_, new_n25866_ );
xor  ( new_n26074_, new_n26073_, new_n25876_ );
xor  ( new_n26075_, new_n25906_, new_n25902_ );
xor  ( new_n26076_, new_n26075_, new_n25912_ );
or   ( new_n26077_, new_n26076_, new_n26074_ );
and  ( new_n26078_, new_n26076_, new_n26074_ );
xor  ( new_n26079_, new_n25888_, new_n25884_ );
xnor ( new_n26080_, new_n26079_, new_n25894_ );
or   ( new_n26081_, new_n26080_, new_n26078_ );
and  ( new_n26082_, new_n26081_, new_n26077_ );
and  ( new_n26083_, new_n26082_, new_n26072_ );
nor  ( new_n26084_, new_n26082_, new_n26072_ );
xor  ( new_n26085_, new_n25991_, new_n25989_ );
xnor ( new_n26086_, new_n26085_, new_n25995_ );
nor  ( new_n26087_, new_n26086_, new_n26084_ );
or   ( new_n26088_, new_n26087_, new_n26083_ );
or   ( new_n26089_, new_n1135_, new_n22973_ );
or   ( new_n26090_, new_n1137_, new_n22975_ );
and  ( new_n26091_, new_n26090_, new_n26089_ );
xor  ( new_n26092_, new_n26091_, new_n896_ );
or   ( new_n26093_, new_n897_, new_n23252_ );
or   ( new_n26094_, new_n899_, new_n23166_ );
and  ( new_n26095_, new_n26094_, new_n26093_ );
xor  ( new_n26096_, new_n26095_, new_n748_ );
or   ( new_n26097_, new_n26096_, new_n26092_ );
and  ( new_n26098_, new_n26096_, new_n26092_ );
or   ( new_n26099_, new_n755_, new_n23554_ );
or   ( new_n26100_, new_n757_, new_n23370_ );
and  ( new_n26101_, new_n26100_, new_n26099_ );
xor  ( new_n26102_, new_n26101_, new_n523_ );
or   ( new_n26103_, new_n26102_, new_n26098_ );
and  ( new_n26104_, new_n26103_, new_n26097_ );
or   ( new_n26105_, new_n1844_, new_n22304_ );
or   ( new_n26106_, new_n1846_, new_n22207_ );
and  ( new_n26107_, new_n26106_, new_n26105_ );
xor  ( new_n26108_, new_n26107_, new_n1586_ );
or   ( new_n26109_, new_n1593_, new_n22590_ );
or   ( new_n26110_, new_n1595_, new_n22423_ );
and  ( new_n26111_, new_n26110_, new_n26109_ );
xor  ( new_n26112_, new_n26111_, new_n1358_ );
or   ( new_n26113_, new_n26112_, new_n26108_ );
and  ( new_n26114_, new_n26112_, new_n26108_ );
or   ( new_n26115_, new_n1364_, new_n22829_ );
or   ( new_n26116_, new_n1366_, new_n22641_ );
and  ( new_n26117_, new_n26116_, new_n26115_ );
xor  ( new_n26118_, new_n26117_, new_n1129_ );
or   ( new_n26119_, new_n26118_, new_n26114_ );
and  ( new_n26120_, new_n26119_, new_n26113_ );
nor  ( new_n26121_, new_n26120_, new_n26104_ );
nand ( new_n26122_, new_n26120_, new_n26104_ );
or   ( new_n26123_, new_n524_, new_n23895_ );
or   ( new_n26124_, new_n526_, new_n23733_ );
and  ( new_n26125_, new_n26124_, new_n26123_ );
xor  ( new_n26126_, new_n26125_, new_n403_ );
or   ( new_n26127_, new_n409_, new_n24227_ );
or   ( new_n26128_, new_n411_, new_n24006_ );
and  ( new_n26129_, new_n26128_, new_n26127_ );
xor  ( new_n26130_, new_n26129_, new_n328_ );
nor  ( new_n26131_, new_n26130_, new_n26126_ );
and  ( new_n26132_, new_n26130_, new_n26126_ );
or   ( new_n26133_, new_n337_, new_n24543_ );
or   ( new_n26134_, new_n340_, new_n24418_ );
and  ( new_n26135_, new_n26134_, new_n26133_ );
xor  ( new_n26136_, new_n26135_, new_n332_ );
nor  ( new_n26137_, new_n26136_, new_n26132_ );
nor  ( new_n26138_, new_n26137_, new_n26131_ );
not  ( new_n26139_, new_n26138_ );
and  ( new_n26140_, new_n26139_, new_n26122_ );
or   ( new_n26141_, new_n26140_, new_n26121_ );
or   ( new_n26142_, new_n2807_, new_n21842_ );
or   ( new_n26143_, new_n2809_, new_n21792_ );
and  ( new_n26144_, new_n26143_, new_n26142_ );
xor  ( new_n26145_, new_n26144_, new_n2424_ );
or   ( new_n26146_, new_n2425_, new_n21847_ );
or   ( new_n26147_, new_n2427_, new_n21840_ );
and  ( new_n26148_, new_n26147_, new_n26146_ );
xor  ( new_n26149_, new_n26148_, new_n2121_ );
or   ( new_n26150_, new_n26149_, new_n26145_ );
and  ( new_n26151_, new_n26149_, new_n26145_ );
or   ( new_n26152_, new_n2122_, new_n22129_ );
or   ( new_n26153_, new_n2124_, new_n22098_ );
and  ( new_n26154_, new_n26153_, new_n26152_ );
xor  ( new_n26155_, new_n26154_, new_n1843_ );
or   ( new_n26156_, new_n26155_, new_n26151_ );
and  ( new_n26157_, new_n26156_, new_n26150_ );
or   ( new_n26158_, new_n4709_, new_n21703_ );
or   ( new_n26159_, new_n4711_, new_n21694_ );
and  ( new_n26160_, new_n26159_, new_n26158_ );
xor  ( new_n26161_, new_n26160_, new_n4294_ );
and  ( new_n26162_, new_n4960_, RIbb315f0_129 );
xor  ( new_n26163_, new_n26162_, new_n4708_ );
nand ( new_n26164_, new_n26163_, new_n26161_ );
nor  ( new_n26165_, new_n26163_, new_n26161_ );
or   ( new_n26166_, new_n4302_, new_n21674_ );
or   ( new_n26167_, new_n4304_, new_n21701_ );
and  ( new_n26168_, new_n26167_, new_n26166_ );
xor  ( new_n26169_, new_n26168_, new_n3895_ );
or   ( new_n26170_, new_n26169_, new_n26165_ );
and  ( new_n26171_, new_n26170_, new_n26164_ );
nor  ( new_n26172_, new_n26171_, new_n26157_ );
and  ( new_n26173_, new_n26171_, new_n26157_ );
or   ( new_n26174_, new_n3896_, new_n21680_ );
or   ( new_n26175_, new_n3898_, new_n21672_ );
and  ( new_n26176_, new_n26175_, new_n26174_ );
xor  ( new_n26177_, new_n26176_, new_n3460_ );
or   ( new_n26178_, new_n3461_, new_n21687_ );
or   ( new_n26179_, new_n3463_, new_n21678_ );
and  ( new_n26180_, new_n26179_, new_n26178_ );
xor  ( new_n26181_, new_n26180_, new_n3116_ );
nor  ( new_n26182_, new_n26181_, new_n26177_ );
and  ( new_n26183_, new_n26181_, new_n26177_ );
or   ( new_n26184_, new_n3117_, new_n21751_ );
or   ( new_n26185_, new_n3119_, new_n21685_ );
and  ( new_n26186_, new_n26185_, new_n26184_ );
xor  ( new_n26187_, new_n26186_, new_n2800_ );
nor  ( new_n26188_, new_n26187_, new_n26183_ );
nor  ( new_n26189_, new_n26188_, new_n26182_ );
nor  ( new_n26190_, new_n26189_, new_n26173_ );
nor  ( new_n26191_, new_n26190_, new_n26172_ );
not  ( new_n26192_, new_n26191_ );
or   ( new_n26193_, new_n26192_, new_n26141_ );
and  ( new_n26194_, new_n26192_, new_n26141_ );
or   ( new_n26195_, new_n268_, new_n26063_ );
not  ( new_n26196_, RIbb32928_170 );
or   ( new_n26197_, new_n271_, new_n26196_ );
and  ( new_n26198_, new_n26197_, new_n26195_ );
xor  ( new_n26199_, new_n26198_, new_n263_ );
and  ( new_n26200_, RIbb32a18_172, RIbb2f610_1 );
or   ( new_n26201_, new_n26200_, new_n26199_ );
or   ( new_n26202_, new_n317_, new_n24925_ );
or   ( new_n26203_, new_n320_, new_n24927_ );
and  ( new_n26204_, new_n26203_, new_n26202_ );
xor  ( new_n26205_, new_n26204_, new_n312_ );
or   ( new_n26206_, new_n283_, new_n25288_ );
or   ( new_n26207_, new_n286_, new_n25048_ );
and  ( new_n26208_, new_n26207_, new_n26206_ );
xor  ( new_n26209_, new_n26208_, new_n278_ );
or   ( new_n26210_, new_n26209_, new_n26205_ );
and  ( new_n26211_, new_n26209_, new_n26205_ );
or   ( new_n26212_, new_n299_, new_n25813_ );
or   ( new_n26213_, new_n302_, new_n25486_ );
and  ( new_n26214_, new_n26213_, new_n26212_ );
xor  ( new_n26215_, new_n26214_, new_n293_ );
or   ( new_n26216_, new_n26215_, new_n26211_ );
and  ( new_n26217_, new_n26216_, new_n26210_ );
and  ( new_n26218_, new_n26217_, new_n26201_ );
nor  ( new_n26219_, new_n26217_, new_n26201_ );
not  ( new_n26220_, new_n26219_ );
or   ( new_n26221_, new_n268_, new_n26196_ );
or   ( new_n26222_, new_n271_, new_n25813_ );
and  ( new_n26223_, new_n26222_, new_n26221_ );
xor  ( new_n26224_, new_n26223_, new_n263_ );
and  ( new_n26225_, new_n26224_, new_n26220_ );
nor  ( new_n26226_, new_n26225_, new_n26218_ );
or   ( new_n26227_, new_n26226_, new_n26194_ );
and  ( new_n26228_, new_n26227_, new_n26193_ );
nor  ( new_n26229_, new_n26228_, new_n26088_ );
and  ( new_n26230_, new_n26228_, new_n26088_ );
xor  ( new_n26231_, new_n25878_, new_n25862_ );
xor  ( new_n26232_, new_n26231_, new_n25896_ );
xnor ( new_n26233_, new_n25979_, new_n25977_ );
xor  ( new_n26234_, new_n26233_, new_n25983_ );
and  ( new_n26235_, new_n26234_, new_n26232_ );
nor  ( new_n26236_, new_n26234_, new_n26232_ );
xor  ( new_n26237_, new_n25965_, new_n25949_ );
xor  ( new_n26238_, new_n26237_, new_n25969_ );
nor  ( new_n26239_, new_n26238_, new_n26236_ );
nor  ( new_n26240_, new_n26239_, new_n26235_ );
nor  ( new_n26241_, new_n26240_, new_n26230_ );
nor  ( new_n26242_, new_n26241_, new_n26229_ );
or   ( new_n26243_, new_n26242_, new_n26062_ );
and  ( new_n26244_, new_n26243_, new_n26061_ );
xor  ( new_n26245_, new_n26024_, new_n26014_ );
xor  ( new_n26246_, new_n26245_, new_n26028_ );
or   ( new_n26247_, new_n26246_, new_n26244_ );
and  ( new_n26248_, new_n26246_, new_n26244_ );
xor  ( new_n26249_, new_n26034_, new_n26032_ );
xor  ( new_n26250_, new_n26249_, new_n26038_ );
or   ( new_n26251_, new_n26250_, new_n26248_ );
and  ( new_n26252_, new_n26251_, new_n26247_ );
or   ( new_n26253_, new_n26252_, new_n26048_ );
and  ( new_n26254_, new_n26252_, new_n26048_ );
xor  ( new_n26255_, new_n25658_, new_n25648_ );
xor  ( new_n26256_, new_n26255_, new_n25828_ );
or   ( new_n26257_, new_n26256_, new_n26254_ );
and  ( new_n26258_, new_n26257_, new_n26253_ );
nand ( new_n26259_, new_n26258_, new_n26046_ );
nor  ( new_n26260_, new_n26258_, new_n26046_ );
xor  ( new_n26261_, new_n25832_, new_n25830_ );
xor  ( new_n26262_, new_n26261_, new_n25835_ );
or   ( new_n26263_, new_n26262_, new_n26260_ );
and  ( new_n26264_, new_n26263_, new_n26259_ );
and  ( new_n26265_, new_n26264_, new_n25846_ );
xor  ( new_n26266_, new_n26252_, new_n26048_ );
xor  ( new_n26267_, new_n26266_, new_n26256_ );
xor  ( new_n26268_, new_n25999_, new_n25973_ );
xnor ( new_n26269_, new_n26268_, new_n26012_ );
xnor ( new_n26270_, new_n26060_, new_n26050_ );
xor  ( new_n26271_, new_n26270_, new_n26242_ );
and  ( new_n26272_, new_n26271_, new_n26269_ );
xor  ( new_n26273_, new_n26018_, new_n26016_ );
xor  ( new_n26274_, new_n26273_, new_n26022_ );
xor  ( new_n26275_, new_n26054_, new_n26052_ );
xor  ( new_n26276_, new_n26275_, new_n26058_ );
xor  ( new_n26277_, new_n25946_, new_n25898_ );
xor  ( new_n26278_, new_n26277_, new_n25971_ );
nand ( new_n26279_, new_n26278_, new_n26276_ );
nor  ( new_n26280_, new_n26278_, new_n26276_ );
xor  ( new_n26281_, new_n26228_, new_n26088_ );
xnor ( new_n26282_, new_n26281_, new_n26240_ );
or   ( new_n26283_, new_n26282_, new_n26280_ );
and  ( new_n26284_, new_n26283_, new_n26279_ );
or   ( new_n26285_, new_n26284_, new_n26274_ );
and  ( new_n26286_, new_n26284_, new_n26274_ );
xnor ( new_n26287_, new_n25985_, new_n25975_ );
xor  ( new_n26288_, new_n26287_, new_n25997_ );
xnor ( new_n26289_, new_n25936_, new_n25932_ );
xor  ( new_n26290_, new_n26289_, new_n25942_ );
xnor ( new_n26291_, new_n26112_, new_n26108_ );
xor  ( new_n26292_, new_n26291_, new_n26118_ );
xnor ( new_n26293_, new_n26149_, new_n26145_ );
xor  ( new_n26294_, new_n26293_, new_n26155_ );
or   ( new_n26295_, new_n26294_, new_n26292_ );
and  ( new_n26296_, new_n26294_, new_n26292_ );
xor  ( new_n26297_, new_n26181_, new_n26177_ );
xnor ( new_n26298_, new_n26297_, new_n26187_ );
or   ( new_n26299_, new_n26298_, new_n26296_ );
and  ( new_n26300_, new_n26299_, new_n26295_ );
nor  ( new_n26301_, new_n26300_, new_n26290_ );
nand ( new_n26302_, new_n26300_, new_n26290_ );
xnor ( new_n26303_, new_n26209_, new_n26205_ );
xor  ( new_n26304_, new_n26303_, new_n26215_ );
xnor ( new_n26305_, new_n26096_, new_n26092_ );
xor  ( new_n26306_, new_n26305_, new_n26102_ );
nor  ( new_n26307_, new_n26306_, new_n26304_ );
nand ( new_n26308_, new_n26306_, new_n26304_ );
xor  ( new_n26309_, new_n26130_, new_n26126_ );
xor  ( new_n26310_, new_n26309_, new_n26136_ );
and  ( new_n26311_, new_n26310_, new_n26308_ );
or   ( new_n26312_, new_n26311_, new_n26307_ );
and  ( new_n26313_, new_n26312_, new_n26302_ );
or   ( new_n26314_, new_n26313_, new_n26301_ );
or   ( new_n26315_, new_n1364_, new_n22975_ );
or   ( new_n26316_, new_n1366_, new_n22829_ );
and  ( new_n26317_, new_n26316_, new_n26315_ );
xor  ( new_n26318_, new_n26317_, new_n1129_ );
or   ( new_n26319_, new_n1135_, new_n23166_ );
or   ( new_n26320_, new_n1137_, new_n22973_ );
and  ( new_n26321_, new_n26320_, new_n26319_ );
xor  ( new_n26322_, new_n26321_, new_n896_ );
or   ( new_n26323_, new_n26322_, new_n26318_ );
and  ( new_n26324_, new_n26322_, new_n26318_ );
or   ( new_n26325_, new_n897_, new_n23370_ );
or   ( new_n26326_, new_n899_, new_n23252_ );
and  ( new_n26327_, new_n26326_, new_n26325_ );
xor  ( new_n26328_, new_n26327_, new_n748_ );
or   ( new_n26329_, new_n26328_, new_n26324_ );
and  ( new_n26330_, new_n26329_, new_n26323_ );
or   ( new_n26331_, new_n2122_, new_n22207_ );
or   ( new_n26332_, new_n2124_, new_n22129_ );
and  ( new_n26333_, new_n26332_, new_n26331_ );
xor  ( new_n26334_, new_n26333_, new_n1843_ );
or   ( new_n26335_, new_n1844_, new_n22423_ );
or   ( new_n26336_, new_n1846_, new_n22304_ );
and  ( new_n26337_, new_n26336_, new_n26335_ );
xor  ( new_n26338_, new_n26337_, new_n1586_ );
or   ( new_n26339_, new_n26338_, new_n26334_ );
and  ( new_n26340_, new_n26338_, new_n26334_ );
or   ( new_n26341_, new_n1593_, new_n22641_ );
or   ( new_n26342_, new_n1595_, new_n22590_ );
and  ( new_n26343_, new_n26342_, new_n26341_ );
xor  ( new_n26344_, new_n26343_, new_n1358_ );
or   ( new_n26345_, new_n26344_, new_n26340_ );
and  ( new_n26346_, new_n26345_, new_n26339_ );
or   ( new_n26347_, new_n26346_, new_n26330_ );
and  ( new_n26348_, new_n26346_, new_n26330_ );
or   ( new_n26349_, new_n755_, new_n23733_ );
or   ( new_n26350_, new_n757_, new_n23554_ );
and  ( new_n26351_, new_n26350_, new_n26349_ );
xor  ( new_n26352_, new_n26351_, new_n523_ );
or   ( new_n26353_, new_n524_, new_n24006_ );
or   ( new_n26354_, new_n526_, new_n23895_ );
and  ( new_n26355_, new_n26354_, new_n26353_ );
xor  ( new_n26356_, new_n26355_, new_n403_ );
nor  ( new_n26357_, new_n26356_, new_n26352_ );
and  ( new_n26358_, new_n26356_, new_n26352_ );
or   ( new_n26359_, new_n409_, new_n24418_ );
or   ( new_n26360_, new_n411_, new_n24227_ );
and  ( new_n26361_, new_n26360_, new_n26359_ );
xor  ( new_n26362_, new_n26361_, new_n328_ );
nor  ( new_n26363_, new_n26362_, new_n26358_ );
nor  ( new_n26364_, new_n26363_, new_n26357_ );
or   ( new_n26365_, new_n26364_, new_n26348_ );
and  ( new_n26366_, new_n26365_, new_n26347_ );
xnor ( new_n26367_, new_n26200_, new_n26199_ );
or   ( new_n26368_, new_n299_, new_n26196_ );
or   ( new_n26369_, new_n302_, new_n25813_ );
and  ( new_n26370_, new_n26369_, new_n26368_ );
xor  ( new_n26371_, new_n26370_, new_n293_ );
not  ( new_n26372_, RIbb32a18_172 );
or   ( new_n26373_, new_n268_, new_n26372_ );
or   ( new_n26374_, new_n271_, new_n26063_ );
and  ( new_n26375_, new_n26374_, new_n26373_ );
xor  ( new_n26376_, new_n26375_, new_n263_ );
or   ( new_n26377_, new_n26376_, new_n26371_ );
and  ( new_n26378_, RIbb32a90_173, RIbb2f610_1 );
and  ( new_n26379_, new_n26376_, new_n26371_ );
or   ( new_n26380_, new_n26379_, new_n26378_ );
and  ( new_n26381_, new_n26380_, new_n26377_ );
or   ( new_n26382_, new_n26381_, new_n26367_ );
and  ( new_n26383_, new_n26381_, new_n26367_ );
or   ( new_n26384_, new_n337_, new_n24927_ );
or   ( new_n26385_, new_n340_, new_n24543_ );
and  ( new_n26386_, new_n26385_, new_n26384_ );
xor  ( new_n26387_, new_n26386_, new_n332_ );
or   ( new_n26388_, new_n317_, new_n25048_ );
or   ( new_n26389_, new_n320_, new_n24925_ );
and  ( new_n26390_, new_n26389_, new_n26388_ );
xor  ( new_n26391_, new_n26390_, new_n312_ );
nor  ( new_n26392_, new_n26391_, new_n26387_ );
and  ( new_n26393_, new_n26391_, new_n26387_ );
or   ( new_n26394_, new_n283_, new_n25486_ );
or   ( new_n26395_, new_n286_, new_n25288_ );
and  ( new_n26396_, new_n26395_, new_n26394_ );
xor  ( new_n26397_, new_n26396_, new_n278_ );
nor  ( new_n26398_, new_n26397_, new_n26393_ );
nor  ( new_n26399_, new_n26398_, new_n26392_ );
or   ( new_n26400_, new_n26399_, new_n26383_ );
and  ( new_n26401_, new_n26400_, new_n26382_ );
or   ( new_n26402_, new_n26401_, new_n26366_ );
and  ( new_n26403_, new_n26401_, new_n26366_ );
or   ( new_n26404_, new_n5207_, new_n21694_ );
or   ( new_n26405_, new_n5209_, new_n21696_ );
and  ( new_n26406_, new_n26405_, new_n26404_ );
xor  ( new_n26407_, new_n26406_, new_n4708_ );
and  ( new_n26408_, new_n26407_, new_n5206_ );
or   ( new_n26409_, new_n26407_, new_n5206_ );
or   ( new_n26410_, new_n4709_, new_n21701_ );
or   ( new_n26411_, new_n4711_, new_n21703_ );
and  ( new_n26412_, new_n26411_, new_n26410_ );
xor  ( new_n26413_, new_n26412_, new_n4295_ );
and  ( new_n26414_, new_n26413_, new_n26409_ );
or   ( new_n26415_, new_n26414_, new_n26408_ );
or   ( new_n26416_, new_n4302_, new_n21672_ );
or   ( new_n26417_, new_n4304_, new_n21674_ );
and  ( new_n26418_, new_n26417_, new_n26416_ );
xor  ( new_n26419_, new_n26418_, new_n3895_ );
or   ( new_n26420_, new_n3896_, new_n21678_ );
or   ( new_n26421_, new_n3898_, new_n21680_ );
and  ( new_n26422_, new_n26421_, new_n26420_ );
xor  ( new_n26423_, new_n26422_, new_n3460_ );
or   ( new_n26424_, new_n26423_, new_n26419_ );
and  ( new_n26425_, new_n26423_, new_n26419_ );
or   ( new_n26426_, new_n3461_, new_n21685_ );
or   ( new_n26427_, new_n3463_, new_n21687_ );
and  ( new_n26428_, new_n26427_, new_n26426_ );
xor  ( new_n26429_, new_n26428_, new_n3116_ );
or   ( new_n26430_, new_n26429_, new_n26425_ );
and  ( new_n26431_, new_n26430_, new_n26424_ );
nor  ( new_n26432_, new_n26431_, new_n26415_ );
and  ( new_n26433_, new_n26431_, new_n26415_ );
or   ( new_n26434_, new_n3117_, new_n21792_ );
or   ( new_n26435_, new_n3119_, new_n21751_ );
and  ( new_n26436_, new_n26435_, new_n26434_ );
xor  ( new_n26437_, new_n26436_, new_n2800_ );
or   ( new_n26438_, new_n2807_, new_n21840_ );
or   ( new_n26439_, new_n2809_, new_n21842_ );
and  ( new_n26440_, new_n26439_, new_n26438_ );
xor  ( new_n26441_, new_n26440_, new_n2424_ );
nor  ( new_n26442_, new_n26441_, new_n26437_ );
and  ( new_n26443_, new_n26441_, new_n26437_ );
or   ( new_n26444_, new_n2425_, new_n22098_ );
or   ( new_n26445_, new_n2427_, new_n21847_ );
and  ( new_n26446_, new_n26445_, new_n26444_ );
xor  ( new_n26447_, new_n26446_, new_n2121_ );
nor  ( new_n26448_, new_n26447_, new_n26443_ );
nor  ( new_n26449_, new_n26448_, new_n26442_ );
nor  ( new_n26450_, new_n26449_, new_n26433_ );
nor  ( new_n26451_, new_n26450_, new_n26432_ );
or   ( new_n26452_, new_n26451_, new_n26403_ );
and  ( new_n26453_, new_n26452_, new_n26402_ );
or   ( new_n26454_, new_n26453_, new_n26314_ );
nand ( new_n26455_, new_n26453_, new_n26314_ );
xor  ( new_n26456_, new_n25918_, new_n4708_ );
xor  ( new_n26457_, new_n26456_, new_n25924_ );
xor  ( new_n26458_, new_n26066_, new_n26064_ );
xor  ( new_n26459_, new_n26458_, new_n26070_ );
nor  ( new_n26460_, new_n26459_, new_n26457_ );
and  ( new_n26461_, new_n26459_, new_n26457_ );
xor  ( new_n26462_, new_n26076_, new_n26074_ );
xnor ( new_n26463_, new_n26462_, new_n26080_ );
not  ( new_n26464_, new_n26463_ );
nor  ( new_n26465_, new_n26464_, new_n26461_ );
nor  ( new_n26466_, new_n26465_, new_n26460_ );
nand ( new_n26467_, new_n26466_, new_n26455_ );
and  ( new_n26468_, new_n26467_, new_n26454_ );
nor  ( new_n26469_, new_n26468_, new_n26288_ );
and  ( new_n26470_, new_n26468_, new_n26288_ );
xnor ( new_n26471_, new_n25926_, new_n25914_ );
xor  ( new_n26472_, new_n26471_, new_n25944_ );
xor  ( new_n26473_, new_n26171_, new_n26157_ );
xor  ( new_n26474_, new_n26473_, new_n26189_ );
xor  ( new_n26475_, new_n26217_, new_n26201_ );
xor  ( new_n26476_, new_n26475_, new_n26224_ );
nand ( new_n26477_, new_n26476_, new_n26474_ );
nor  ( new_n26478_, new_n26476_, new_n26474_ );
xor  ( new_n26479_, new_n26120_, new_n26104_ );
xor  ( new_n26480_, new_n26479_, new_n26139_ );
or   ( new_n26481_, new_n26480_, new_n26478_ );
and  ( new_n26482_, new_n26481_, new_n26477_ );
nor  ( new_n26483_, new_n26482_, new_n26472_ );
and  ( new_n26484_, new_n26482_, new_n26472_ );
xor  ( new_n26485_, new_n26234_, new_n26232_ );
xnor ( new_n26486_, new_n26485_, new_n26238_ );
not  ( new_n26487_, new_n26486_ );
nor  ( new_n26488_, new_n26487_, new_n26484_ );
nor  ( new_n26489_, new_n26488_, new_n26483_ );
not  ( new_n26490_, new_n26489_ );
nor  ( new_n26491_, new_n26490_, new_n26470_ );
nor  ( new_n26492_, new_n26491_, new_n26469_ );
or   ( new_n26493_, new_n26492_, new_n26286_ );
and  ( new_n26494_, new_n26493_, new_n26285_ );
nand ( new_n26495_, new_n26494_, new_n26272_ );
nor  ( new_n26496_, new_n26494_, new_n26272_ );
xor  ( new_n26497_, new_n26246_, new_n26244_ );
xor  ( new_n26498_, new_n26497_, new_n26250_ );
or   ( new_n26499_, new_n26498_, new_n26496_ );
and  ( new_n26500_, new_n26499_, new_n26495_ );
or   ( new_n26501_, new_n26500_, new_n26267_ );
xnor ( new_n26502_, new_n26258_, new_n26046_ );
xor  ( new_n26503_, new_n26502_, new_n26262_ );
nor  ( new_n26504_, new_n26503_, new_n26501_ );
xor  ( new_n26505_, new_n26494_, new_n26272_ );
xor  ( new_n26506_, new_n26505_, new_n26498_ );
xor  ( new_n26507_, new_n26192_, new_n26141_ );
xor  ( new_n26508_, new_n26507_, new_n26226_ );
xor  ( new_n26509_, new_n26453_, new_n26314_ );
xor  ( new_n26510_, new_n26509_, new_n26466_ );
nor  ( new_n26511_, new_n26510_, new_n26508_ );
nand ( new_n26512_, new_n26510_, new_n26508_ );
xor  ( new_n26513_, new_n26482_, new_n26472_ );
xor  ( new_n26514_, new_n26513_, new_n26487_ );
not  ( new_n26515_, new_n26514_ );
and  ( new_n26516_, new_n26515_, new_n26512_ );
or   ( new_n26517_, new_n26516_, new_n26511_ );
xor  ( new_n26518_, new_n26082_, new_n26072_ );
xor  ( new_n26519_, new_n26518_, new_n26086_ );
xnor ( new_n26520_, new_n26163_, new_n26161_ );
xor  ( new_n26521_, new_n26520_, new_n26169_ );
xnor ( new_n26522_, new_n26322_, new_n26318_ );
xor  ( new_n26523_, new_n26522_, new_n26328_ );
xnor ( new_n26524_, new_n26356_, new_n26352_ );
xor  ( new_n26525_, new_n26524_, new_n26362_ );
or   ( new_n26526_, new_n26525_, new_n26523_ );
and  ( new_n26527_, new_n26525_, new_n26523_ );
xor  ( new_n26528_, new_n26391_, new_n26387_ );
xnor ( new_n26529_, new_n26528_, new_n26397_ );
or   ( new_n26530_, new_n26529_, new_n26527_ );
and  ( new_n26531_, new_n26530_, new_n26526_ );
nor  ( new_n26532_, new_n26531_, new_n26521_ );
and  ( new_n26533_, new_n26531_, new_n26521_ );
xnor ( new_n26534_, new_n26338_, new_n26334_ );
xor  ( new_n26535_, new_n26534_, new_n26344_ );
xnor ( new_n26536_, new_n26423_, new_n26419_ );
xor  ( new_n26537_, new_n26536_, new_n26429_ );
nor  ( new_n26538_, new_n26537_, new_n26535_ );
and  ( new_n26539_, new_n26537_, new_n26535_ );
xor  ( new_n26540_, new_n26441_, new_n26437_ );
xnor ( new_n26541_, new_n26540_, new_n26447_ );
nor  ( new_n26542_, new_n26541_, new_n26539_ );
nor  ( new_n26543_, new_n26542_, new_n26538_ );
nor  ( new_n26544_, new_n26543_, new_n26533_ );
or   ( new_n26545_, new_n26544_, new_n26532_ );
or   ( new_n26546_, new_n4302_, new_n21680_ );
or   ( new_n26547_, new_n4304_, new_n21672_ );
and  ( new_n26548_, new_n26547_, new_n26546_ );
xor  ( new_n26549_, new_n26548_, new_n3895_ );
or   ( new_n26550_, new_n3896_, new_n21687_ );
or   ( new_n26551_, new_n3898_, new_n21678_ );
and  ( new_n26552_, new_n26551_, new_n26550_ );
xor  ( new_n26553_, new_n26552_, new_n3460_ );
or   ( new_n26554_, new_n26553_, new_n26549_ );
and  ( new_n26555_, new_n26553_, new_n26549_ );
or   ( new_n26556_, new_n3461_, new_n21751_ );
or   ( new_n26557_, new_n3463_, new_n21685_ );
and  ( new_n26558_, new_n26557_, new_n26556_ );
xor  ( new_n26559_, new_n26558_, new_n3116_ );
or   ( new_n26560_, new_n26559_, new_n26555_ );
and  ( new_n26561_, new_n26560_, new_n26554_ );
or   ( new_n26562_, new_n5207_, new_n21703_ );
or   ( new_n26563_, new_n5209_, new_n21694_ );
and  ( new_n26564_, new_n26563_, new_n26562_ );
xor  ( new_n26565_, new_n26564_, new_n4707_ );
and  ( new_n26566_, new_n5373_, RIbb315f0_129 );
xor  ( new_n26567_, new_n26566_, new_n5206_ );
nand ( new_n26568_, new_n26567_, new_n26565_ );
nor  ( new_n26569_, new_n26567_, new_n26565_ );
or   ( new_n26570_, new_n4709_, new_n21674_ );
or   ( new_n26571_, new_n4711_, new_n21701_ );
and  ( new_n26572_, new_n26571_, new_n26570_ );
xor  ( new_n26573_, new_n26572_, new_n4295_ );
or   ( new_n26574_, new_n26573_, new_n26569_ );
and  ( new_n26575_, new_n26574_, new_n26568_ );
or   ( new_n26576_, new_n26575_, new_n26561_ );
and  ( new_n26577_, new_n26575_, new_n26561_ );
or   ( new_n26578_, new_n3117_, new_n21842_ );
or   ( new_n26579_, new_n3119_, new_n21792_ );
and  ( new_n26580_, new_n26579_, new_n26578_ );
xor  ( new_n26581_, new_n26580_, new_n2800_ );
or   ( new_n26582_, new_n2807_, new_n21847_ );
or   ( new_n26583_, new_n2809_, new_n21840_ );
and  ( new_n26584_, new_n26583_, new_n26582_ );
xor  ( new_n26585_, new_n26584_, new_n2424_ );
nor  ( new_n26586_, new_n26585_, new_n26581_ );
and  ( new_n26587_, new_n26585_, new_n26581_ );
or   ( new_n26588_, new_n2425_, new_n22129_ );
or   ( new_n26589_, new_n2427_, new_n22098_ );
and  ( new_n26590_, new_n26589_, new_n26588_ );
xor  ( new_n26591_, new_n26590_, new_n2121_ );
nor  ( new_n26592_, new_n26591_, new_n26587_ );
nor  ( new_n26593_, new_n26592_, new_n26586_ );
or   ( new_n26594_, new_n26593_, new_n26577_ );
and  ( new_n26595_, new_n26594_, new_n26576_ );
xor  ( new_n26596_, new_n26376_, new_n26371_ );
xor  ( new_n26597_, new_n26596_, new_n26378_ );
or   ( new_n26598_, new_n337_, new_n24925_ );
or   ( new_n26599_, new_n340_, new_n24927_ );
and  ( new_n26600_, new_n26599_, new_n26598_ );
xor  ( new_n26601_, new_n26600_, new_n332_ );
or   ( new_n26602_, new_n317_, new_n25288_ );
or   ( new_n26603_, new_n320_, new_n25048_ );
and  ( new_n26604_, new_n26603_, new_n26602_ );
xor  ( new_n26605_, new_n26604_, new_n312_ );
or   ( new_n26606_, new_n26605_, new_n26601_ );
and  ( new_n26607_, new_n26605_, new_n26601_ );
or   ( new_n26608_, new_n283_, new_n25813_ );
or   ( new_n26609_, new_n286_, new_n25486_ );
and  ( new_n26610_, new_n26609_, new_n26608_ );
xor  ( new_n26611_, new_n26610_, new_n278_ );
or   ( new_n26612_, new_n26611_, new_n26607_ );
and  ( new_n26613_, new_n26612_, new_n26606_ );
or   ( new_n26614_, new_n26613_, new_n26597_ );
and  ( new_n26615_, new_n26613_, new_n26597_ );
or   ( new_n26616_, new_n299_, new_n26063_ );
or   ( new_n26617_, new_n302_, new_n26196_ );
and  ( new_n26618_, new_n26617_, new_n26616_ );
xor  ( new_n26619_, new_n26618_, new_n293_ );
not  ( new_n26620_, RIbb32a90_173 );
or   ( new_n26621_, new_n268_, new_n26620_ );
or   ( new_n26622_, new_n271_, new_n26372_ );
and  ( new_n26623_, new_n26622_, new_n26621_ );
xor  ( new_n26624_, new_n26623_, new_n263_ );
nor  ( new_n26625_, new_n26624_, new_n26619_ );
and  ( new_n26626_, RIbb32b08_174, RIbb2f610_1 );
and  ( new_n26627_, new_n26624_, new_n26619_ );
nor  ( new_n26628_, new_n26627_, new_n26626_ );
nor  ( new_n26629_, new_n26628_, new_n26625_ );
or   ( new_n26630_, new_n26629_, new_n26615_ );
and  ( new_n26631_, new_n26630_, new_n26614_ );
or   ( new_n26632_, new_n26631_, new_n26595_ );
and  ( new_n26633_, new_n26631_, new_n26595_ );
or   ( new_n26634_, new_n1364_, new_n22973_ );
or   ( new_n26635_, new_n1366_, new_n22975_ );
and  ( new_n26636_, new_n26635_, new_n26634_ );
xor  ( new_n26637_, new_n26636_, new_n1129_ );
or   ( new_n26638_, new_n1135_, new_n23252_ );
or   ( new_n26639_, new_n1137_, new_n23166_ );
and  ( new_n26640_, new_n26639_, new_n26638_ );
xor  ( new_n26641_, new_n26640_, new_n896_ );
or   ( new_n26642_, new_n26641_, new_n26637_ );
and  ( new_n26643_, new_n26641_, new_n26637_ );
or   ( new_n26644_, new_n897_, new_n23554_ );
or   ( new_n26645_, new_n899_, new_n23370_ );
and  ( new_n26646_, new_n26645_, new_n26644_ );
xor  ( new_n26647_, new_n26646_, new_n748_ );
or   ( new_n26648_, new_n26647_, new_n26643_ );
and  ( new_n26649_, new_n26648_, new_n26642_ );
or   ( new_n26650_, new_n2122_, new_n22304_ );
or   ( new_n26651_, new_n2124_, new_n22207_ );
and  ( new_n26652_, new_n26651_, new_n26650_ );
xor  ( new_n26653_, new_n26652_, new_n1843_ );
or   ( new_n26654_, new_n1844_, new_n22590_ );
or   ( new_n26655_, new_n1846_, new_n22423_ );
and  ( new_n26656_, new_n26655_, new_n26654_ );
xor  ( new_n26657_, new_n26656_, new_n1586_ );
or   ( new_n26658_, new_n26657_, new_n26653_ );
and  ( new_n26659_, new_n26657_, new_n26653_ );
or   ( new_n26660_, new_n1593_, new_n22829_ );
or   ( new_n26661_, new_n1595_, new_n22641_ );
and  ( new_n26662_, new_n26661_, new_n26660_ );
xor  ( new_n26663_, new_n26662_, new_n1358_ );
or   ( new_n26664_, new_n26663_, new_n26659_ );
and  ( new_n26665_, new_n26664_, new_n26658_ );
nor  ( new_n26666_, new_n26665_, new_n26649_ );
and  ( new_n26667_, new_n26665_, new_n26649_ );
or   ( new_n26668_, new_n755_, new_n23895_ );
or   ( new_n26669_, new_n757_, new_n23733_ );
and  ( new_n26670_, new_n26669_, new_n26668_ );
xor  ( new_n26671_, new_n26670_, new_n523_ );
or   ( new_n26672_, new_n524_, new_n24227_ );
or   ( new_n26673_, new_n526_, new_n24006_ );
and  ( new_n26674_, new_n26673_, new_n26672_ );
xor  ( new_n26675_, new_n26674_, new_n403_ );
nor  ( new_n26676_, new_n26675_, new_n26671_ );
and  ( new_n26677_, new_n26675_, new_n26671_ );
or   ( new_n26678_, new_n409_, new_n24543_ );
or   ( new_n26679_, new_n411_, new_n24418_ );
and  ( new_n26680_, new_n26679_, new_n26678_ );
xor  ( new_n26681_, new_n26680_, new_n328_ );
nor  ( new_n26682_, new_n26681_, new_n26677_ );
nor  ( new_n26683_, new_n26682_, new_n26676_ );
nor  ( new_n26684_, new_n26683_, new_n26667_ );
nor  ( new_n26685_, new_n26684_, new_n26666_ );
or   ( new_n26686_, new_n26685_, new_n26633_ );
and  ( new_n26687_, new_n26686_, new_n26632_ );
or   ( new_n26688_, new_n26687_, new_n26545_ );
nand ( new_n26689_, new_n26687_, new_n26545_ );
xor  ( new_n26690_, new_n26306_, new_n26304_ );
xor  ( new_n26691_, new_n26690_, new_n26310_ );
xnor ( new_n26692_, new_n26294_, new_n26292_ );
xor  ( new_n26693_, new_n26692_, new_n26298_ );
and  ( new_n26694_, new_n26693_, new_n26691_ );
nor  ( new_n26695_, new_n26693_, new_n26691_ );
xor  ( new_n26696_, new_n26381_, new_n26367_ );
xnor ( new_n26697_, new_n26696_, new_n26399_ );
nor  ( new_n26698_, new_n26697_, new_n26695_ );
nor  ( new_n26699_, new_n26698_, new_n26694_ );
nand ( new_n26700_, new_n26699_, new_n26689_ );
and  ( new_n26701_, new_n26700_, new_n26688_ );
or   ( new_n26702_, new_n26701_, new_n26519_ );
nand ( new_n26703_, new_n26701_, new_n26519_ );
xor  ( new_n26704_, new_n26300_, new_n26290_ );
xor  ( new_n26705_, new_n26704_, new_n26312_ );
xnor ( new_n26706_, new_n26476_, new_n26474_ );
xor  ( new_n26707_, new_n26706_, new_n26480_ );
and  ( new_n26708_, new_n26707_, new_n26705_ );
nor  ( new_n26709_, new_n26707_, new_n26705_ );
xor  ( new_n26710_, new_n26459_, new_n26457_ );
xor  ( new_n26711_, new_n26710_, new_n26464_ );
nor  ( new_n26712_, new_n26711_, new_n26709_ );
nor  ( new_n26713_, new_n26712_, new_n26708_ );
nand ( new_n26714_, new_n26713_, new_n26703_ );
and  ( new_n26715_, new_n26714_, new_n26702_ );
nor  ( new_n26716_, new_n26715_, new_n26517_ );
nand ( new_n26717_, new_n26715_, new_n26517_ );
xor  ( new_n26718_, new_n26278_, new_n26276_ );
xnor ( new_n26719_, new_n26718_, new_n26282_ );
and  ( new_n26720_, new_n26719_, new_n26717_ );
or   ( new_n26721_, new_n26720_, new_n26716_ );
xnor ( new_n26722_, new_n26284_, new_n26274_ );
xor  ( new_n26723_, new_n26722_, new_n26492_ );
or   ( new_n26724_, new_n26723_, new_n26721_ );
nand ( new_n26725_, new_n26723_, new_n26721_ );
xor  ( new_n26726_, new_n26271_, new_n26269_ );
nand ( new_n26727_, new_n26726_, new_n26725_ );
and  ( new_n26728_, new_n26727_, new_n26724_ );
nor  ( new_n26729_, new_n26728_, new_n26506_ );
xor  ( new_n26730_, new_n26500_, new_n26267_ );
and  ( new_n26731_, new_n26730_, new_n26729_ );
xor  ( new_n26732_, new_n26723_, new_n26721_ );
xor  ( new_n26733_, new_n26732_, new_n26726_ );
xnor ( new_n26734_, new_n26715_, new_n26517_ );
xor  ( new_n26735_, new_n26734_, new_n26719_ );
or   ( new_n26736_, new_n409_, new_n24927_ );
or   ( new_n26737_, new_n411_, new_n24543_ );
and  ( new_n26738_, new_n26737_, new_n26736_ );
xor  ( new_n26739_, new_n26738_, new_n328_ );
or   ( new_n26740_, new_n337_, new_n25048_ );
or   ( new_n26741_, new_n340_, new_n24925_ );
and  ( new_n26742_, new_n26741_, new_n26740_ );
xor  ( new_n26743_, new_n26742_, new_n332_ );
nor  ( new_n26744_, new_n26743_, new_n26739_ );
and  ( new_n26745_, new_n26743_, new_n26739_ );
or   ( new_n26746_, new_n317_, new_n25486_ );
or   ( new_n26747_, new_n320_, new_n25288_ );
and  ( new_n26748_, new_n26747_, new_n26746_ );
xor  ( new_n26749_, new_n26748_, new_n312_ );
nor  ( new_n26750_, new_n26749_, new_n26745_ );
nor  ( new_n26751_, new_n26750_, new_n26744_ );
or   ( new_n26752_, new_n283_, new_n26196_ );
or   ( new_n26753_, new_n286_, new_n25813_ );
and  ( new_n26754_, new_n26753_, new_n26752_ );
xor  ( new_n26755_, new_n26754_, new_n278_ );
or   ( new_n26756_, new_n299_, new_n26372_ );
or   ( new_n26757_, new_n302_, new_n26063_ );
and  ( new_n26758_, new_n26757_, new_n26756_ );
xor  ( new_n26759_, new_n26758_, new_n293_ );
or   ( new_n26760_, new_n26759_, new_n26755_ );
and  ( new_n26761_, new_n26759_, new_n26755_ );
not  ( new_n26762_, RIbb32b08_174 );
or   ( new_n26763_, new_n268_, new_n26762_ );
or   ( new_n26764_, new_n271_, new_n26620_ );
and  ( new_n26765_, new_n26764_, new_n26763_ );
xor  ( new_n26766_, new_n26765_, new_n263_ );
or   ( new_n26767_, new_n26766_, new_n26761_ );
and  ( new_n26768_, new_n26767_, new_n26760_ );
or   ( new_n26769_, new_n26768_, new_n26751_ );
or   ( new_n26770_, new_n4709_, new_n21672_ );
or   ( new_n26771_, new_n4711_, new_n21674_ );
and  ( new_n26772_, new_n26771_, new_n26770_ );
xor  ( new_n26773_, new_n26772_, new_n4295_ );
or   ( new_n26774_, new_n4302_, new_n21678_ );
or   ( new_n26775_, new_n4304_, new_n21680_ );
and  ( new_n26776_, new_n26775_, new_n26774_ );
xor  ( new_n26777_, new_n26776_, new_n3895_ );
nor  ( new_n26778_, new_n26777_, new_n26773_ );
and  ( new_n26779_, new_n26777_, new_n26773_ );
or   ( new_n26780_, new_n3896_, new_n21685_ );
or   ( new_n26781_, new_n3898_, new_n21687_ );
and  ( new_n26782_, new_n26781_, new_n26780_ );
xor  ( new_n26783_, new_n26782_, new_n3460_ );
nor  ( new_n26784_, new_n26783_, new_n26779_ );
or   ( new_n26785_, new_n26784_, new_n26778_ );
or   ( new_n26786_, new_n5207_, new_n21701_ );
or   ( new_n26787_, new_n5209_, new_n21703_ );
and  ( new_n26788_, new_n26787_, new_n26786_ );
xor  ( new_n26789_, new_n26788_, new_n4708_ );
nand ( new_n26790_, new_n26789_, new_n5597_ );
or   ( new_n26791_, new_n26789_, new_n5597_ );
or   ( new_n26792_, new_n5604_, new_n21694_ );
or   ( new_n26793_, new_n5606_, new_n21696_ );
and  ( new_n26794_, new_n26793_, new_n26792_ );
xor  ( new_n26795_, new_n26794_, new_n5206_ );
nand ( new_n26796_, new_n26795_, new_n26791_ );
and  ( new_n26797_, new_n26796_, new_n26790_ );
nand ( new_n26798_, new_n26797_, new_n26785_ );
nor  ( new_n26799_, new_n26797_, new_n26785_ );
or   ( new_n26800_, new_n3461_, new_n21792_ );
or   ( new_n26801_, new_n3463_, new_n21751_ );
and  ( new_n26802_, new_n26801_, new_n26800_ );
xor  ( new_n26803_, new_n26802_, new_n3116_ );
or   ( new_n26804_, new_n3117_, new_n21840_ );
or   ( new_n26805_, new_n3119_, new_n21842_ );
and  ( new_n26806_, new_n26805_, new_n26804_ );
xor  ( new_n26807_, new_n26806_, new_n2800_ );
nor  ( new_n26808_, new_n26807_, new_n26803_ );
and  ( new_n26809_, new_n26807_, new_n26803_ );
or   ( new_n26810_, new_n2807_, new_n22098_ );
or   ( new_n26811_, new_n2809_, new_n21847_ );
and  ( new_n26812_, new_n26811_, new_n26810_ );
xor  ( new_n26813_, new_n26812_, new_n2424_ );
nor  ( new_n26814_, new_n26813_, new_n26809_ );
nor  ( new_n26815_, new_n26814_, new_n26808_ );
or   ( new_n26816_, new_n26815_, new_n26799_ );
and  ( new_n26817_, new_n26816_, new_n26798_ );
nor  ( new_n26818_, new_n26817_, new_n26769_ );
nand ( new_n26819_, new_n26817_, new_n26769_ );
or   ( new_n26820_, new_n1593_, new_n22975_ );
or   ( new_n26821_, new_n1595_, new_n22829_ );
and  ( new_n26822_, new_n26821_, new_n26820_ );
xor  ( new_n26823_, new_n26822_, new_n1358_ );
or   ( new_n26824_, new_n1364_, new_n23166_ );
or   ( new_n26825_, new_n1366_, new_n22973_ );
and  ( new_n26826_, new_n26825_, new_n26824_ );
xor  ( new_n26827_, new_n26826_, new_n1129_ );
or   ( new_n26828_, new_n26827_, new_n26823_ );
and  ( new_n26829_, new_n26827_, new_n26823_ );
or   ( new_n26830_, new_n1135_, new_n23370_ );
or   ( new_n26831_, new_n1137_, new_n23252_ );
and  ( new_n26832_, new_n26831_, new_n26830_ );
xor  ( new_n26833_, new_n26832_, new_n896_ );
or   ( new_n26834_, new_n26833_, new_n26829_ );
and  ( new_n26835_, new_n26834_, new_n26828_ );
or   ( new_n26836_, new_n897_, new_n23733_ );
or   ( new_n26837_, new_n899_, new_n23554_ );
and  ( new_n26838_, new_n26837_, new_n26836_ );
xor  ( new_n26839_, new_n26838_, new_n748_ );
or   ( new_n26840_, new_n755_, new_n24006_ );
or   ( new_n26841_, new_n757_, new_n23895_ );
and  ( new_n26842_, new_n26841_, new_n26840_ );
xor  ( new_n26843_, new_n26842_, new_n523_ );
or   ( new_n26844_, new_n26843_, new_n26839_ );
and  ( new_n26845_, new_n26843_, new_n26839_ );
or   ( new_n26846_, new_n524_, new_n24418_ );
or   ( new_n26847_, new_n526_, new_n24227_ );
and  ( new_n26848_, new_n26847_, new_n26846_ );
xor  ( new_n26849_, new_n26848_, new_n403_ );
or   ( new_n26850_, new_n26849_, new_n26845_ );
and  ( new_n26851_, new_n26850_, new_n26844_ );
nor  ( new_n26852_, new_n26851_, new_n26835_ );
and  ( new_n26853_, new_n26851_, new_n26835_ );
or   ( new_n26854_, new_n2425_, new_n22207_ );
or   ( new_n26855_, new_n2427_, new_n22129_ );
and  ( new_n26856_, new_n26855_, new_n26854_ );
xor  ( new_n26857_, new_n26856_, new_n2121_ );
or   ( new_n26858_, new_n2122_, new_n22423_ );
or   ( new_n26859_, new_n2124_, new_n22304_ );
and  ( new_n26860_, new_n26859_, new_n26858_ );
xor  ( new_n26861_, new_n26860_, new_n1843_ );
nor  ( new_n26862_, new_n26861_, new_n26857_ );
and  ( new_n26863_, new_n26861_, new_n26857_ );
or   ( new_n26864_, new_n1844_, new_n22641_ );
or   ( new_n26865_, new_n1846_, new_n22590_ );
and  ( new_n26866_, new_n26865_, new_n26864_ );
xor  ( new_n26867_, new_n26866_, new_n1586_ );
nor  ( new_n26868_, new_n26867_, new_n26863_ );
nor  ( new_n26869_, new_n26868_, new_n26862_ );
nor  ( new_n26870_, new_n26869_, new_n26853_ );
nor  ( new_n26871_, new_n26870_, new_n26852_ );
not  ( new_n26872_, new_n26871_ );
and  ( new_n26873_, new_n26872_, new_n26819_ );
or   ( new_n26874_, new_n26873_, new_n26818_ );
xor  ( new_n26875_, new_n26567_, new_n26565_ );
xnor ( new_n26876_, new_n26875_, new_n26573_ );
xnor ( new_n26877_, new_n26553_, new_n26549_ );
xor  ( new_n26878_, new_n26877_, new_n26559_ );
or   ( new_n26879_, new_n26878_, new_n26876_ );
xnor ( new_n26880_, new_n26657_, new_n26653_ );
xor  ( new_n26881_, new_n26880_, new_n26663_ );
xnor ( new_n26882_, new_n26641_, new_n26637_ );
xor  ( new_n26883_, new_n26882_, new_n26647_ );
or   ( new_n26884_, new_n26883_, new_n26881_ );
and  ( new_n26885_, new_n26883_, new_n26881_ );
xor  ( new_n26886_, new_n26585_, new_n26581_ );
xnor ( new_n26887_, new_n26886_, new_n26591_ );
or   ( new_n26888_, new_n26887_, new_n26885_ );
and  ( new_n26889_, new_n26888_, new_n26884_ );
or   ( new_n26890_, new_n26889_, new_n26879_ );
and  ( new_n26891_, new_n26889_, new_n26879_ );
xnor ( new_n26892_, new_n26675_, new_n26671_ );
xor  ( new_n26893_, new_n26892_, new_n26681_ );
xnor ( new_n26894_, new_n26605_, new_n26601_ );
xor  ( new_n26895_, new_n26894_, new_n26611_ );
nor  ( new_n26896_, new_n26895_, new_n26893_ );
and  ( new_n26897_, new_n26895_, new_n26893_ );
xor  ( new_n26898_, new_n26624_, new_n26619_ );
xnor ( new_n26899_, new_n26898_, new_n26626_ );
nor  ( new_n26900_, new_n26899_, new_n26897_ );
nor  ( new_n26901_, new_n26900_, new_n26896_ );
or   ( new_n26902_, new_n26901_, new_n26891_ );
and  ( new_n26903_, new_n26902_, new_n26890_ );
or   ( new_n26904_, new_n26903_, new_n26874_ );
nand ( new_n26905_, new_n26903_, new_n26874_ );
xor  ( new_n26906_, new_n26407_, new_n5206_ );
xor  ( new_n26907_, new_n26906_, new_n26413_ );
xnor ( new_n26908_, new_n26537_, new_n26535_ );
xor  ( new_n26909_, new_n26908_, new_n26541_ );
nor  ( new_n26910_, new_n26909_, new_n26907_ );
and  ( new_n26911_, new_n26909_, new_n26907_ );
xor  ( new_n26912_, new_n26525_, new_n26523_ );
xnor ( new_n26913_, new_n26912_, new_n26529_ );
nor  ( new_n26914_, new_n26913_, new_n26911_ );
nor  ( new_n26915_, new_n26914_, new_n26910_ );
nand ( new_n26916_, new_n26915_, new_n26905_ );
and  ( new_n26917_, new_n26916_, new_n26904_ );
xnor ( new_n26918_, new_n26431_, new_n26415_ );
xor  ( new_n26919_, new_n26918_, new_n26449_ );
xnor ( new_n26920_, new_n26575_, new_n26561_ );
xor  ( new_n26921_, new_n26920_, new_n26593_ );
xnor ( new_n26922_, new_n26665_, new_n26649_ );
xor  ( new_n26923_, new_n26922_, new_n26683_ );
or   ( new_n26924_, new_n26923_, new_n26921_ );
and  ( new_n26925_, new_n26923_, new_n26921_ );
xnor ( new_n26926_, new_n26613_, new_n26597_ );
xor  ( new_n26927_, new_n26926_, new_n26629_ );
or   ( new_n26928_, new_n26927_, new_n26925_ );
and  ( new_n26929_, new_n26928_, new_n26924_ );
or   ( new_n26930_, new_n26929_, new_n26919_ );
and  ( new_n26931_, new_n26929_, new_n26919_ );
xor  ( new_n26932_, new_n26346_, new_n26330_ );
xnor ( new_n26933_, new_n26932_, new_n26364_ );
or   ( new_n26934_, new_n26933_, new_n26931_ );
and  ( new_n26935_, new_n26934_, new_n26930_ );
or   ( new_n26936_, new_n26935_, new_n26917_ );
and  ( new_n26937_, new_n26935_, new_n26917_ );
xor  ( new_n26938_, new_n26531_, new_n26521_ );
xor  ( new_n26939_, new_n26938_, new_n26543_ );
xnor ( new_n26940_, new_n26631_, new_n26595_ );
xor  ( new_n26941_, new_n26940_, new_n26685_ );
nor  ( new_n26942_, new_n26941_, new_n26939_ );
and  ( new_n26943_, new_n26941_, new_n26939_ );
xor  ( new_n26944_, new_n26693_, new_n26691_ );
xnor ( new_n26945_, new_n26944_, new_n26697_ );
not  ( new_n26946_, new_n26945_ );
nor  ( new_n26947_, new_n26946_, new_n26943_ );
nor  ( new_n26948_, new_n26947_, new_n26942_ );
or   ( new_n26949_, new_n26948_, new_n26937_ );
and  ( new_n26950_, new_n26949_, new_n26936_ );
xor  ( new_n26951_, new_n26687_, new_n26545_ );
xor  ( new_n26952_, new_n26951_, new_n26699_ );
xnor ( new_n26953_, new_n26401_, new_n26366_ );
xor  ( new_n26954_, new_n26953_, new_n26451_ );
or   ( new_n26955_, new_n26954_, new_n26952_ );
and  ( new_n26956_, new_n26954_, new_n26952_ );
xor  ( new_n26957_, new_n26707_, new_n26705_ );
xor  ( new_n26958_, new_n26957_, new_n26711_ );
or   ( new_n26959_, new_n26958_, new_n26956_ );
and  ( new_n26960_, new_n26959_, new_n26955_ );
nand ( new_n26961_, new_n26960_, new_n26950_ );
nor  ( new_n26962_, new_n26960_, new_n26950_ );
xor  ( new_n26963_, new_n26510_, new_n26508_ );
xor  ( new_n26964_, new_n26963_, new_n26515_ );
or   ( new_n26965_, new_n26964_, new_n26962_ );
and  ( new_n26966_, new_n26965_, new_n26961_ );
or   ( new_n26967_, new_n26966_, new_n26735_ );
nand ( new_n26968_, new_n26966_, new_n26735_ );
xor  ( new_n26969_, new_n26468_, new_n26288_ );
xor  ( new_n26970_, new_n26969_, new_n26489_ );
nand ( new_n26971_, new_n26970_, new_n26968_ );
and  ( new_n26972_, new_n26971_, new_n26967_ );
and  ( new_n26973_, new_n26972_, new_n26733_ );
xor  ( new_n26974_, new_n26728_, new_n26506_ );
and  ( new_n26975_, new_n26974_, new_n26973_ );
xor  ( new_n26976_, new_n26954_, new_n26952_ );
xor  ( new_n26977_, new_n26976_, new_n26958_ );
xor  ( new_n26978_, new_n26903_, new_n26874_ );
xor  ( new_n26979_, new_n26978_, new_n26915_ );
xnor ( new_n26980_, new_n26929_, new_n26919_ );
xor  ( new_n26981_, new_n26980_, new_n26933_ );
nand ( new_n26982_, new_n26981_, new_n26979_ );
nor  ( new_n26983_, new_n26981_, new_n26979_ );
xor  ( new_n26984_, new_n26941_, new_n26939_ );
xor  ( new_n26985_, new_n26984_, new_n26946_ );
or   ( new_n26986_, new_n26985_, new_n26983_ );
and  ( new_n26987_, new_n26986_, new_n26982_ );
or   ( new_n26988_, new_n26987_, new_n26977_ );
and  ( new_n26989_, new_n26987_, new_n26977_ );
xor  ( new_n26990_, new_n26817_, new_n26769_ );
xor  ( new_n26991_, new_n26990_, new_n26872_ );
not  ( new_n26992_, new_n26991_ );
xnor ( new_n26993_, new_n26889_, new_n26879_ );
xor  ( new_n26994_, new_n26993_, new_n26901_ );
nand ( new_n26995_, new_n26994_, new_n26992_ );
xnor ( new_n26996_, new_n26883_, new_n26881_ );
xor  ( new_n26997_, new_n26996_, new_n26887_ );
xnor ( new_n26998_, new_n26895_, new_n26893_ );
xor  ( new_n26999_, new_n26998_, new_n26899_ );
nor  ( new_n27000_, new_n26999_, new_n26997_ );
nand ( new_n27001_, new_n26999_, new_n26997_ );
xor  ( new_n27002_, new_n26878_, new_n26876_ );
not  ( new_n27003_, new_n27002_ );
and  ( new_n27004_, new_n27003_, new_n27001_ );
or   ( new_n27005_, new_n27004_, new_n27000_ );
or   ( new_n27006_, new_n2425_, new_n22304_ );
or   ( new_n27007_, new_n2427_, new_n22207_ );
and  ( new_n27008_, new_n27007_, new_n27006_ );
xor  ( new_n27009_, new_n27008_, new_n2121_ );
or   ( new_n27010_, new_n2122_, new_n22590_ );
or   ( new_n27011_, new_n2124_, new_n22423_ );
and  ( new_n27012_, new_n27011_, new_n27010_ );
xor  ( new_n27013_, new_n27012_, new_n1843_ );
or   ( new_n27014_, new_n27013_, new_n27009_ );
and  ( new_n27015_, new_n27013_, new_n27009_ );
or   ( new_n27016_, new_n1844_, new_n22829_ );
or   ( new_n27017_, new_n1846_, new_n22641_ );
and  ( new_n27018_, new_n27017_, new_n27016_ );
xor  ( new_n27019_, new_n27018_, new_n1586_ );
or   ( new_n27020_, new_n27019_, new_n27015_ );
and  ( new_n27021_, new_n27020_, new_n27014_ );
or   ( new_n27022_, new_n1593_, new_n22973_ );
or   ( new_n27023_, new_n1595_, new_n22975_ );
and  ( new_n27024_, new_n27023_, new_n27022_ );
xor  ( new_n27025_, new_n27024_, new_n1358_ );
or   ( new_n27026_, new_n1364_, new_n23252_ );
or   ( new_n27027_, new_n1366_, new_n23166_ );
and  ( new_n27028_, new_n27027_, new_n27026_ );
xor  ( new_n27029_, new_n27028_, new_n1129_ );
or   ( new_n27030_, new_n27029_, new_n27025_ );
and  ( new_n27031_, new_n27029_, new_n27025_ );
or   ( new_n27032_, new_n1135_, new_n23554_ );
or   ( new_n27033_, new_n1137_, new_n23370_ );
and  ( new_n27034_, new_n27033_, new_n27032_ );
xor  ( new_n27035_, new_n27034_, new_n896_ );
or   ( new_n27036_, new_n27035_, new_n27031_ );
and  ( new_n27037_, new_n27036_, new_n27030_ );
or   ( new_n27038_, new_n27037_, new_n27021_ );
and  ( new_n27039_, new_n27037_, new_n27021_ );
or   ( new_n27040_, new_n897_, new_n23895_ );
or   ( new_n27041_, new_n899_, new_n23733_ );
and  ( new_n27042_, new_n27041_, new_n27040_ );
xor  ( new_n27043_, new_n27042_, new_n748_ );
or   ( new_n27044_, new_n755_, new_n24227_ );
or   ( new_n27045_, new_n757_, new_n24006_ );
and  ( new_n27046_, new_n27045_, new_n27044_ );
xor  ( new_n27047_, new_n27046_, new_n523_ );
nor  ( new_n27048_, new_n27047_, new_n27043_ );
and  ( new_n27049_, new_n27047_, new_n27043_ );
or   ( new_n27050_, new_n524_, new_n24543_ );
or   ( new_n27051_, new_n526_, new_n24418_ );
and  ( new_n27052_, new_n27051_, new_n27050_ );
xor  ( new_n27053_, new_n27052_, new_n403_ );
nor  ( new_n27054_, new_n27053_, new_n27049_ );
nor  ( new_n27055_, new_n27054_, new_n27048_ );
or   ( new_n27056_, new_n27055_, new_n27039_ );
and  ( new_n27057_, new_n27056_, new_n27038_ );
or   ( new_n27058_, new_n409_, new_n24925_ );
or   ( new_n27059_, new_n411_, new_n24927_ );
and  ( new_n27060_, new_n27059_, new_n27058_ );
xor  ( new_n27061_, new_n27060_, new_n328_ );
or   ( new_n27062_, new_n337_, new_n25288_ );
or   ( new_n27063_, new_n340_, new_n25048_ );
and  ( new_n27064_, new_n27063_, new_n27062_ );
xor  ( new_n27065_, new_n27064_, new_n332_ );
or   ( new_n27066_, new_n27065_, new_n27061_ );
and  ( new_n27067_, new_n27065_, new_n27061_ );
or   ( new_n27068_, new_n317_, new_n25813_ );
or   ( new_n27069_, new_n320_, new_n25486_ );
and  ( new_n27070_, new_n27069_, new_n27068_ );
xor  ( new_n27071_, new_n27070_, new_n312_ );
or   ( new_n27072_, new_n27071_, new_n27067_ );
and  ( new_n27073_, new_n27072_, new_n27066_ );
and  ( new_n27074_, RIbb32bf8_176, RIbb2f610_1 );
or   ( new_n27075_, new_n283_, new_n26063_ );
or   ( new_n27076_, new_n286_, new_n26196_ );
and  ( new_n27077_, new_n27076_, new_n27075_ );
xor  ( new_n27078_, new_n27077_, new_n278_ );
or   ( new_n27079_, new_n299_, new_n26620_ );
or   ( new_n27080_, new_n302_, new_n26372_ );
and  ( new_n27081_, new_n27080_, new_n27079_ );
xor  ( new_n27082_, new_n27081_, new_n293_ );
or   ( new_n27083_, new_n27082_, new_n27078_ );
and  ( new_n27084_, new_n27082_, new_n27078_ );
not  ( new_n27085_, RIbb32b80_175 );
or   ( new_n27086_, new_n268_, new_n27085_ );
or   ( new_n27087_, new_n271_, new_n26762_ );
and  ( new_n27088_, new_n27087_, new_n27086_ );
xor  ( new_n27089_, new_n27088_, new_n263_ );
or   ( new_n27090_, new_n27089_, new_n27084_ );
and  ( new_n27091_, new_n27090_, new_n27083_ );
and  ( new_n27092_, new_n27091_, new_n27074_ );
or   ( new_n27093_, new_n27092_, new_n27073_ );
or   ( new_n27094_, new_n27091_, new_n27074_ );
and  ( new_n27095_, new_n27094_, new_n27093_ );
nor  ( new_n27096_, new_n27095_, new_n27057_ );
or   ( new_n27097_, new_n5604_, new_n21703_ );
or   ( new_n27098_, new_n5606_, new_n21694_ );
and  ( new_n27099_, new_n27098_, new_n27097_ );
xor  ( new_n27100_, new_n27099_, new_n5205_ );
and  ( new_n27101_, new_n5917_, RIbb315f0_129 );
xor  ( new_n27102_, new_n27101_, new_n5597_ );
nand ( new_n27103_, new_n27102_, new_n27100_ );
nor  ( new_n27104_, new_n27102_, new_n27100_ );
or   ( new_n27105_, new_n5207_, new_n21674_ );
or   ( new_n27106_, new_n5209_, new_n21701_ );
and  ( new_n27107_, new_n27106_, new_n27105_ );
xor  ( new_n27108_, new_n27107_, new_n4708_ );
or   ( new_n27109_, new_n27108_, new_n27104_ );
and  ( new_n27110_, new_n27109_, new_n27103_ );
or   ( new_n27111_, new_n4709_, new_n21680_ );
or   ( new_n27112_, new_n4711_, new_n21672_ );
and  ( new_n27113_, new_n27112_, new_n27111_ );
xor  ( new_n27114_, new_n27113_, new_n4295_ );
or   ( new_n27115_, new_n4302_, new_n21687_ );
or   ( new_n27116_, new_n4304_, new_n21678_ );
and  ( new_n27117_, new_n27116_, new_n27115_ );
xor  ( new_n27118_, new_n27117_, new_n3895_ );
or   ( new_n27119_, new_n27118_, new_n27114_ );
and  ( new_n27120_, new_n27118_, new_n27114_ );
or   ( new_n27121_, new_n3896_, new_n21751_ );
or   ( new_n27122_, new_n3898_, new_n21685_ );
and  ( new_n27123_, new_n27122_, new_n27121_ );
xor  ( new_n27124_, new_n27123_, new_n3460_ );
or   ( new_n27125_, new_n27124_, new_n27120_ );
and  ( new_n27126_, new_n27125_, new_n27119_ );
nor  ( new_n27127_, new_n27126_, new_n27110_ );
and  ( new_n27128_, new_n27126_, new_n27110_ );
or   ( new_n27129_, new_n3461_, new_n21842_ );
or   ( new_n27130_, new_n3463_, new_n21792_ );
and  ( new_n27131_, new_n27130_, new_n27129_ );
xor  ( new_n27132_, new_n27131_, new_n3116_ );
or   ( new_n27133_, new_n3117_, new_n21847_ );
or   ( new_n27134_, new_n3119_, new_n21840_ );
and  ( new_n27135_, new_n27134_, new_n27133_ );
xor  ( new_n27136_, new_n27135_, new_n2800_ );
nor  ( new_n27137_, new_n27136_, new_n27132_ );
and  ( new_n27138_, new_n27136_, new_n27132_ );
or   ( new_n27139_, new_n2807_, new_n22129_ );
or   ( new_n27140_, new_n2809_, new_n22098_ );
and  ( new_n27141_, new_n27140_, new_n27139_ );
xor  ( new_n27142_, new_n27141_, new_n2424_ );
nor  ( new_n27143_, new_n27142_, new_n27138_ );
nor  ( new_n27144_, new_n27143_, new_n27137_ );
nor  ( new_n27145_, new_n27144_, new_n27128_ );
nor  ( new_n27146_, new_n27145_, new_n27127_ );
and  ( new_n27147_, new_n27095_, new_n27057_ );
nor  ( new_n27148_, new_n27147_, new_n27146_ );
nor  ( new_n27149_, new_n27148_, new_n27096_ );
not  ( new_n27150_, new_n27149_ );
or   ( new_n27151_, new_n27150_, new_n27005_ );
and  ( new_n27152_, new_n27150_, new_n27005_ );
xor  ( new_n27153_, new_n26807_, new_n26803_ );
xor  ( new_n27154_, new_n27153_, new_n26813_ );
xor  ( new_n27155_, new_n26789_, new_n5597_ );
xor  ( new_n27156_, new_n27155_, new_n26795_ );
and  ( new_n27157_, new_n27156_, new_n27154_ );
or   ( new_n27158_, new_n27156_, new_n27154_ );
xor  ( new_n27159_, new_n26777_, new_n26773_ );
xor  ( new_n27160_, new_n27159_, new_n26783_ );
and  ( new_n27161_, new_n27160_, new_n27158_ );
or   ( new_n27162_, new_n27161_, new_n27157_ );
or   ( new_n27163_, new_n27085_, new_n260_ );
xnor ( new_n27164_, new_n26743_, new_n26739_ );
xor  ( new_n27165_, new_n27164_, new_n26749_ );
nand ( new_n27166_, new_n27165_, new_n27163_ );
or   ( new_n27167_, new_n27165_, new_n27163_ );
xor  ( new_n27168_, new_n26759_, new_n26755_ );
xnor ( new_n27169_, new_n27168_, new_n26766_ );
nand ( new_n27170_, new_n27169_, new_n27167_ );
and  ( new_n27171_, new_n27170_, new_n27166_ );
nand ( new_n27172_, new_n27171_, new_n27162_ );
nor  ( new_n27173_, new_n27171_, new_n27162_ );
xnor ( new_n27174_, new_n26843_, new_n26839_ );
xor  ( new_n27175_, new_n27174_, new_n26849_ );
xnor ( new_n27176_, new_n26827_, new_n26823_ );
xor  ( new_n27177_, new_n27176_, new_n26833_ );
nor  ( new_n27178_, new_n27177_, new_n27175_ );
and  ( new_n27179_, new_n27177_, new_n27175_ );
xor  ( new_n27180_, new_n26861_, new_n26857_ );
xnor ( new_n27181_, new_n27180_, new_n26867_ );
nor  ( new_n27182_, new_n27181_, new_n27179_ );
nor  ( new_n27183_, new_n27182_, new_n27178_ );
or   ( new_n27184_, new_n27183_, new_n27173_ );
and  ( new_n27185_, new_n27184_, new_n27172_ );
or   ( new_n27186_, new_n27185_, new_n27152_ );
and  ( new_n27187_, new_n27186_, new_n27151_ );
or   ( new_n27188_, new_n27187_, new_n26995_ );
and  ( new_n27189_, new_n27187_, new_n26995_ );
xor  ( new_n27190_, new_n26923_, new_n26921_ );
xor  ( new_n27191_, new_n27190_, new_n26927_ );
xnor ( new_n27192_, new_n26909_, new_n26907_ );
xor  ( new_n27193_, new_n27192_, new_n26913_ );
nor  ( new_n27194_, new_n27193_, new_n27191_ );
and  ( new_n27195_, new_n27193_, new_n27191_ );
xnor ( new_n27196_, new_n26797_, new_n26785_ );
xor  ( new_n27197_, new_n27196_, new_n26815_ );
xnor ( new_n27198_, new_n26851_, new_n26835_ );
xor  ( new_n27199_, new_n27198_, new_n26869_ );
nor  ( new_n27200_, new_n27199_, new_n27197_ );
and  ( new_n27201_, new_n27199_, new_n27197_ );
xor  ( new_n27202_, new_n26768_, new_n26751_ );
nor  ( new_n27203_, new_n27202_, new_n27201_ );
nor  ( new_n27204_, new_n27203_, new_n27200_ );
nor  ( new_n27205_, new_n27204_, new_n27195_ );
nor  ( new_n27206_, new_n27205_, new_n27194_ );
or   ( new_n27207_, new_n27206_, new_n27189_ );
and  ( new_n27208_, new_n27207_, new_n27188_ );
or   ( new_n27209_, new_n27208_, new_n26989_ );
and  ( new_n27210_, new_n27209_, new_n26988_ );
xor  ( new_n27211_, new_n26701_, new_n26519_ );
xor  ( new_n27212_, new_n27211_, new_n26713_ );
or   ( new_n27213_, new_n27212_, new_n27210_ );
and  ( new_n27214_, new_n27212_, new_n27210_ );
xnor ( new_n27215_, new_n26960_, new_n26950_ );
xor  ( new_n27216_, new_n27215_, new_n26964_ );
or   ( new_n27217_, new_n27216_, new_n27214_ );
and  ( new_n27218_, new_n27217_, new_n27213_ );
xor  ( new_n27219_, new_n26966_, new_n26735_ );
xor  ( new_n27220_, new_n27219_, new_n26970_ );
nor  ( new_n27221_, new_n27220_, new_n27218_ );
xor  ( new_n27222_, new_n26972_, new_n26733_ );
and  ( new_n27223_, new_n27222_, new_n27221_ );
xor  ( new_n27224_, new_n27212_, new_n27210_ );
xor  ( new_n27225_, new_n27224_, new_n27216_ );
xor  ( new_n27226_, new_n27149_, new_n27005_ );
xor  ( new_n27227_, new_n27226_, new_n27185_ );
xnor ( new_n27228_, new_n27193_, new_n27191_ );
xor  ( new_n27229_, new_n27228_, new_n27204_ );
or   ( new_n27230_, new_n27229_, new_n27227_ );
and  ( new_n27231_, new_n27229_, new_n27227_ );
xor  ( new_n27232_, new_n26994_, new_n26992_ );
or   ( new_n27233_, new_n27232_, new_n27231_ );
and  ( new_n27234_, new_n27233_, new_n27230_ );
xnor ( new_n27235_, new_n26981_, new_n26979_ );
xor  ( new_n27236_, new_n27235_, new_n26985_ );
and  ( new_n27237_, new_n27236_, new_n27234_ );
or   ( new_n27238_, new_n27236_, new_n27234_ );
xor  ( new_n27239_, new_n27095_, new_n27057_ );
xnor ( new_n27240_, new_n27239_, new_n27146_ );
xnor ( new_n27241_, new_n27171_, new_n27162_ );
xnor ( new_n27242_, new_n27241_, new_n27183_ );
or   ( new_n27243_, new_n27242_, new_n27240_ );
xnor ( new_n27244_, new_n27118_, new_n27114_ );
xor  ( new_n27245_, new_n27244_, new_n27124_ );
xnor ( new_n27246_, new_n27102_, new_n27100_ );
xor  ( new_n27247_, new_n27246_, new_n27108_ );
or   ( new_n27248_, new_n27247_, new_n27245_ );
and  ( new_n27249_, new_n27247_, new_n27245_ );
xor  ( new_n27250_, new_n27136_, new_n27132_ );
xnor ( new_n27251_, new_n27250_, new_n27142_ );
or   ( new_n27252_, new_n27251_, new_n27249_ );
and  ( new_n27253_, new_n27252_, new_n27248_ );
xnor ( new_n27254_, new_n27065_, new_n27061_ );
xor  ( new_n27255_, new_n27254_, new_n27071_ );
xnor ( new_n27256_, new_n27082_, new_n27078_ );
xor  ( new_n27257_, new_n27256_, new_n27089_ );
or   ( new_n27258_, new_n27257_, new_n27255_ );
and  ( new_n27259_, new_n27257_, new_n27255_ );
or   ( new_n27260_, new_n27259_, new_n27074_ );
and  ( new_n27261_, new_n27260_, new_n27258_ );
nor  ( new_n27262_, new_n27261_, new_n27253_ );
nand ( new_n27263_, new_n27261_, new_n27253_ );
xnor ( new_n27264_, new_n27029_, new_n27025_ );
xor  ( new_n27265_, new_n27264_, new_n27035_ );
xnor ( new_n27266_, new_n27013_, new_n27009_ );
xor  ( new_n27267_, new_n27266_, new_n27019_ );
nor  ( new_n27268_, new_n27267_, new_n27265_ );
and  ( new_n27269_, new_n27267_, new_n27265_ );
xor  ( new_n27270_, new_n27047_, new_n27043_ );
xnor ( new_n27271_, new_n27270_, new_n27053_ );
nor  ( new_n27272_, new_n27271_, new_n27269_ );
nor  ( new_n27273_, new_n27272_, new_n27268_ );
not  ( new_n27274_, new_n27273_ );
and  ( new_n27275_, new_n27274_, new_n27263_ );
or   ( new_n27276_, new_n27275_, new_n27262_ );
or   ( new_n27277_, new_n1844_, new_n22975_ );
or   ( new_n27278_, new_n1846_, new_n22829_ );
and  ( new_n27279_, new_n27278_, new_n27277_ );
xor  ( new_n27280_, new_n27279_, new_n1586_ );
or   ( new_n27281_, new_n1593_, new_n23166_ );
or   ( new_n27282_, new_n1595_, new_n22973_ );
and  ( new_n27283_, new_n27282_, new_n27281_ );
xor  ( new_n27284_, new_n27283_, new_n1358_ );
or   ( new_n27285_, new_n27284_, new_n27280_ );
and  ( new_n27286_, new_n27284_, new_n27280_ );
or   ( new_n27287_, new_n1364_, new_n23370_ );
or   ( new_n27288_, new_n1366_, new_n23252_ );
and  ( new_n27289_, new_n27288_, new_n27287_ );
xor  ( new_n27290_, new_n27289_, new_n1129_ );
or   ( new_n27291_, new_n27290_, new_n27286_ );
and  ( new_n27292_, new_n27291_, new_n27285_ );
or   ( new_n27293_, new_n2807_, new_n22207_ );
or   ( new_n27294_, new_n2809_, new_n22129_ );
and  ( new_n27295_, new_n27294_, new_n27293_ );
xor  ( new_n27296_, new_n27295_, new_n2424_ );
or   ( new_n27297_, new_n2425_, new_n22423_ );
or   ( new_n27298_, new_n2427_, new_n22304_ );
and  ( new_n27299_, new_n27298_, new_n27297_ );
xor  ( new_n27300_, new_n27299_, new_n2121_ );
or   ( new_n27301_, new_n27300_, new_n27296_ );
and  ( new_n27302_, new_n27300_, new_n27296_ );
or   ( new_n27303_, new_n2122_, new_n22641_ );
or   ( new_n27304_, new_n2124_, new_n22590_ );
and  ( new_n27305_, new_n27304_, new_n27303_ );
xor  ( new_n27306_, new_n27305_, new_n1843_ );
or   ( new_n27307_, new_n27306_, new_n27302_ );
and  ( new_n27308_, new_n27307_, new_n27301_ );
or   ( new_n27309_, new_n27308_, new_n27292_ );
and  ( new_n27310_, new_n27308_, new_n27292_ );
or   ( new_n27311_, new_n1135_, new_n23733_ );
or   ( new_n27312_, new_n1137_, new_n23554_ );
and  ( new_n27313_, new_n27312_, new_n27311_ );
xor  ( new_n27314_, new_n27313_, new_n896_ );
or   ( new_n27315_, new_n897_, new_n24006_ );
or   ( new_n27316_, new_n899_, new_n23895_ );
and  ( new_n27317_, new_n27316_, new_n27315_ );
xor  ( new_n27318_, new_n27317_, new_n748_ );
nor  ( new_n27319_, new_n27318_, new_n27314_ );
and  ( new_n27320_, new_n27318_, new_n27314_ );
or   ( new_n27321_, new_n755_, new_n24418_ );
or   ( new_n27322_, new_n757_, new_n24227_ );
and  ( new_n27323_, new_n27322_, new_n27321_ );
xor  ( new_n27324_, new_n27323_, new_n523_ );
nor  ( new_n27325_, new_n27324_, new_n27320_ );
nor  ( new_n27326_, new_n27325_, new_n27319_ );
or   ( new_n27327_, new_n27326_, new_n27310_ );
and  ( new_n27328_, new_n27327_, new_n27309_ );
or   ( new_n27329_, new_n5207_, new_n21672_ );
or   ( new_n27330_, new_n5209_, new_n21674_ );
and  ( new_n27331_, new_n27330_, new_n27329_ );
xor  ( new_n27332_, new_n27331_, new_n4708_ );
or   ( new_n27333_, new_n4709_, new_n21678_ );
or   ( new_n27334_, new_n4711_, new_n21680_ );
and  ( new_n27335_, new_n27334_, new_n27333_ );
xor  ( new_n27336_, new_n27335_, new_n4295_ );
nor  ( new_n27337_, new_n27336_, new_n27332_ );
nand ( new_n27338_, new_n27336_, new_n27332_ );
or   ( new_n27339_, new_n4302_, new_n21685_ );
or   ( new_n27340_, new_n4304_, new_n21687_ );
and  ( new_n27341_, new_n27340_, new_n27339_ );
xor  ( new_n27342_, new_n27341_, new_n3895_ );
not  ( new_n27343_, new_n27342_ );
and  ( new_n27344_, new_n27343_, new_n27338_ );
or   ( new_n27345_, new_n27344_, new_n27337_ );
or   ( new_n27346_, new_n5604_, new_n21701_ );
or   ( new_n27347_, new_n5606_, new_n21703_ );
and  ( new_n27348_, new_n27347_, new_n27346_ );
xor  ( new_n27349_, new_n27348_, new_n5206_ );
nand ( new_n27350_, new_n27349_, new_n6166_ );
or   ( new_n27351_, new_n27349_, new_n6166_ );
or   ( new_n27352_, new_n6173_, new_n21694_ );
or   ( new_n27353_, new_n6175_, new_n21696_ );
and  ( new_n27354_, new_n27353_, new_n27352_ );
xor  ( new_n27355_, new_n27354_, new_n5597_ );
nand ( new_n27356_, new_n27355_, new_n27351_ );
and  ( new_n27357_, new_n27356_, new_n27350_ );
nand ( new_n27358_, new_n27357_, new_n27345_ );
nor  ( new_n27359_, new_n27357_, new_n27345_ );
or   ( new_n27360_, new_n3896_, new_n21792_ );
or   ( new_n27361_, new_n3898_, new_n21751_ );
and  ( new_n27362_, new_n27361_, new_n27360_ );
xor  ( new_n27363_, new_n27362_, new_n3460_ );
or   ( new_n27364_, new_n3461_, new_n21840_ );
or   ( new_n27365_, new_n3463_, new_n21842_ );
and  ( new_n27366_, new_n27365_, new_n27364_ );
xor  ( new_n27367_, new_n27366_, new_n3116_ );
or   ( new_n27368_, new_n27367_, new_n27363_ );
and  ( new_n27369_, new_n27367_, new_n27363_ );
or   ( new_n27370_, new_n3117_, new_n22098_ );
or   ( new_n27371_, new_n3119_, new_n21847_ );
and  ( new_n27372_, new_n27371_, new_n27370_ );
xor  ( new_n27373_, new_n27372_, new_n2800_ );
or   ( new_n27374_, new_n27373_, new_n27369_ );
and  ( new_n27375_, new_n27374_, new_n27368_ );
or   ( new_n27376_, new_n27375_, new_n27359_ );
and  ( new_n27377_, new_n27376_, new_n27358_ );
or   ( new_n27378_, new_n27377_, new_n27328_ );
and  ( new_n27379_, new_n27377_, new_n27328_ );
or   ( new_n27380_, new_n524_, new_n24927_ );
or   ( new_n27381_, new_n526_, new_n24543_ );
and  ( new_n27382_, new_n27381_, new_n27380_ );
xor  ( new_n27383_, new_n27382_, new_n403_ );
or   ( new_n27384_, new_n409_, new_n25048_ );
or   ( new_n27385_, new_n411_, new_n24925_ );
and  ( new_n27386_, new_n27385_, new_n27384_ );
xor  ( new_n27387_, new_n27386_, new_n328_ );
nor  ( new_n27388_, new_n27387_, new_n27383_ );
and  ( new_n27389_, new_n27387_, new_n27383_ );
or   ( new_n27390_, new_n337_, new_n25486_ );
or   ( new_n27391_, new_n340_, new_n25288_ );
and  ( new_n27392_, new_n27391_, new_n27390_ );
xor  ( new_n27393_, new_n27392_, new_n332_ );
nor  ( new_n27394_, new_n27393_, new_n27389_ );
nor  ( new_n27395_, new_n27394_, new_n27388_ );
not  ( new_n27396_, RIbb32bf8_176 );
or   ( new_n27397_, new_n268_, new_n27396_ );
or   ( new_n27398_, new_n271_, new_n27085_ );
and  ( new_n27399_, new_n27398_, new_n27397_ );
xor  ( new_n27400_, new_n27399_, new_n263_ );
and  ( new_n27401_, RIbb32c70_177, RIbb2f610_1 );
and  ( new_n27402_, new_n27401_, new_n27400_ );
or   ( new_n27403_, new_n317_, new_n26196_ );
or   ( new_n27404_, new_n320_, new_n25813_ );
and  ( new_n27405_, new_n27404_, new_n27403_ );
xor  ( new_n27406_, new_n27405_, new_n312_ );
or   ( new_n27407_, new_n283_, new_n26372_ );
or   ( new_n27408_, new_n286_, new_n26063_ );
and  ( new_n27409_, new_n27408_, new_n27407_ );
xor  ( new_n27410_, new_n27409_, new_n278_ );
nor  ( new_n27411_, new_n27410_, new_n27406_ );
and  ( new_n27412_, new_n27410_, new_n27406_ );
or   ( new_n27413_, new_n299_, new_n26762_ );
or   ( new_n27414_, new_n302_, new_n26620_ );
and  ( new_n27415_, new_n27414_, new_n27413_ );
xor  ( new_n27416_, new_n27415_, new_n293_ );
nor  ( new_n27417_, new_n27416_, new_n27412_ );
nor  ( new_n27418_, new_n27417_, new_n27411_ );
and  ( new_n27419_, new_n27418_, new_n27402_ );
nor  ( new_n27420_, new_n27419_, new_n27395_ );
nor  ( new_n27421_, new_n27418_, new_n27402_ );
nor  ( new_n27422_, new_n27421_, new_n27420_ );
or   ( new_n27423_, new_n27422_, new_n27379_ );
and  ( new_n27424_, new_n27423_, new_n27378_ );
nand ( new_n27425_, new_n27424_, new_n27276_ );
nor  ( new_n27426_, new_n27424_, new_n27276_ );
xnor ( new_n27427_, new_n27177_, new_n27175_ );
xor  ( new_n27428_, new_n27427_, new_n27181_ );
xor  ( new_n27429_, new_n27156_, new_n27154_ );
xor  ( new_n27430_, new_n27429_, new_n27160_ );
and  ( new_n27431_, new_n27430_, new_n27428_ );
nor  ( new_n27432_, new_n27430_, new_n27428_ );
xor  ( new_n27433_, new_n27165_, new_n27163_ );
xor  ( new_n27434_, new_n27433_, new_n27169_ );
nor  ( new_n27435_, new_n27434_, new_n27432_ );
nor  ( new_n27436_, new_n27435_, new_n27431_ );
or   ( new_n27437_, new_n27436_, new_n27426_ );
and  ( new_n27438_, new_n27437_, new_n27425_ );
nor  ( new_n27439_, new_n27438_, new_n27243_ );
and  ( new_n27440_, new_n27438_, new_n27243_ );
xor  ( new_n27441_, new_n27199_, new_n27197_ );
xor  ( new_n27442_, new_n27441_, new_n27202_ );
not  ( new_n27443_, new_n27074_ );
xor  ( new_n27444_, new_n27091_, new_n27443_ );
xor  ( new_n27445_, new_n27444_, new_n27073_ );
xnor ( new_n27446_, new_n27037_, new_n27021_ );
xor  ( new_n27447_, new_n27446_, new_n27055_ );
or   ( new_n27448_, new_n27447_, new_n27445_ );
and  ( new_n27449_, new_n27447_, new_n27445_ );
xor  ( new_n27450_, new_n27126_, new_n27110_ );
xnor ( new_n27451_, new_n27450_, new_n27144_ );
or   ( new_n27452_, new_n27451_, new_n27449_ );
and  ( new_n27453_, new_n27452_, new_n27448_ );
nor  ( new_n27454_, new_n27453_, new_n27442_ );
and  ( new_n27455_, new_n27453_, new_n27442_ );
xor  ( new_n27456_, new_n26999_, new_n26997_ );
xor  ( new_n27457_, new_n27456_, new_n27003_ );
nor  ( new_n27458_, new_n27457_, new_n27455_ );
nor  ( new_n27459_, new_n27458_, new_n27454_ );
nor  ( new_n27460_, new_n27459_, new_n27440_ );
nor  ( new_n27461_, new_n27460_, new_n27439_ );
not  ( new_n27462_, new_n27461_ );
and  ( new_n27463_, new_n27462_, new_n27238_ );
or   ( new_n27464_, new_n27463_, new_n27237_ );
xnor ( new_n27465_, new_n26935_, new_n26917_ );
xor  ( new_n27466_, new_n27465_, new_n26948_ );
nand ( new_n27467_, new_n27466_, new_n27464_ );
nor  ( new_n27468_, new_n27466_, new_n27464_ );
xor  ( new_n27469_, new_n26987_, new_n26977_ );
xor  ( new_n27470_, new_n27469_, new_n27208_ );
or   ( new_n27471_, new_n27470_, new_n27468_ );
and  ( new_n27472_, new_n27471_, new_n27467_ );
nor  ( new_n27473_, new_n27472_, new_n27225_ );
xor  ( new_n27474_, new_n27220_, new_n27218_ );
and  ( new_n27475_, new_n27474_, new_n27473_ );
xor  ( new_n27476_, new_n27466_, new_n27464_ );
xor  ( new_n27477_, new_n27476_, new_n27470_ );
xnor ( new_n27478_, new_n27453_, new_n27442_ );
xor  ( new_n27479_, new_n27478_, new_n27457_ );
xnor ( new_n27480_, new_n27424_, new_n27276_ );
xor  ( new_n27481_, new_n27480_, new_n27436_ );
nor  ( new_n27482_, new_n27481_, new_n27479_ );
nand ( new_n27483_, new_n27481_, new_n27479_ );
xnor ( new_n27484_, new_n27242_, new_n27240_ );
and  ( new_n27485_, new_n27484_, new_n27483_ );
or   ( new_n27486_, new_n27485_, new_n27482_ );
xnor ( new_n27487_, new_n27229_, new_n27227_ );
xor  ( new_n27488_, new_n27487_, new_n27232_ );
nor  ( new_n27489_, new_n27488_, new_n27486_ );
nand ( new_n27490_, new_n27488_, new_n27486_ );
xor  ( new_n27491_, new_n27261_, new_n27253_ );
xor  ( new_n27492_, new_n27491_, new_n27274_ );
xnor ( new_n27493_, new_n27377_, new_n27328_ );
xnor ( new_n27494_, new_n27493_, new_n27422_ );
nand ( new_n27495_, new_n27494_, new_n27492_ );
xnor ( new_n27496_, new_n27430_, new_n27428_ );
xor  ( new_n27497_, new_n27496_, new_n27434_ );
xnor ( new_n27498_, new_n27447_, new_n27445_ );
xor  ( new_n27499_, new_n27498_, new_n27451_ );
nand ( new_n27500_, new_n27499_, new_n27497_ );
nor  ( new_n27501_, new_n27499_, new_n27497_ );
xor  ( new_n27502_, new_n27357_, new_n27345_ );
xor  ( new_n27503_, new_n27502_, new_n27375_ );
xor  ( new_n27504_, new_n27418_, new_n27402_ );
xor  ( new_n27505_, new_n27504_, new_n27395_ );
and  ( new_n27506_, new_n27505_, new_n27503_ );
nor  ( new_n27507_, new_n27505_, new_n27503_ );
xor  ( new_n27508_, new_n27308_, new_n27292_ );
xnor ( new_n27509_, new_n27508_, new_n27326_ );
nor  ( new_n27510_, new_n27509_, new_n27507_ );
nor  ( new_n27511_, new_n27510_, new_n27506_ );
or   ( new_n27512_, new_n27511_, new_n27501_ );
and  ( new_n27513_, new_n27512_, new_n27500_ );
nor  ( new_n27514_, new_n27513_, new_n27495_ );
and  ( new_n27515_, new_n27513_, new_n27495_ );
xor  ( new_n27516_, new_n27367_, new_n27363_ );
xor  ( new_n27517_, new_n27516_, new_n27373_ );
xor  ( new_n27518_, new_n27349_, new_n6166_ );
xor  ( new_n27519_, new_n27518_, new_n27355_ );
nand ( new_n27520_, new_n27519_, new_n27517_ );
nor  ( new_n27521_, new_n27519_, new_n27517_ );
xor  ( new_n27522_, new_n27336_, new_n27332_ );
xor  ( new_n27523_, new_n27522_, new_n27343_ );
or   ( new_n27524_, new_n27523_, new_n27521_ );
and  ( new_n27525_, new_n27524_, new_n27520_ );
xnor ( new_n27526_, new_n27387_, new_n27383_ );
xor  ( new_n27527_, new_n27526_, new_n27393_ );
xnor ( new_n27528_, new_n27410_, new_n27406_ );
xor  ( new_n27529_, new_n27528_, new_n27416_ );
or   ( new_n27530_, new_n27529_, new_n27527_ );
nand ( new_n27531_, new_n27529_, new_n27527_ );
xor  ( new_n27532_, new_n27401_, new_n27400_ );
nand ( new_n27533_, new_n27532_, new_n27531_ );
and  ( new_n27534_, new_n27533_, new_n27530_ );
nor  ( new_n27535_, new_n27534_, new_n27525_ );
nand ( new_n27536_, new_n27534_, new_n27525_ );
xnor ( new_n27537_, new_n27300_, new_n27296_ );
xor  ( new_n27538_, new_n27537_, new_n27306_ );
xnor ( new_n27539_, new_n27284_, new_n27280_ );
xor  ( new_n27540_, new_n27539_, new_n27290_ );
nor  ( new_n27541_, new_n27540_, new_n27538_ );
and  ( new_n27542_, new_n27540_, new_n27538_ );
xor  ( new_n27543_, new_n27318_, new_n27314_ );
xnor ( new_n27544_, new_n27543_, new_n27324_ );
nor  ( new_n27545_, new_n27544_, new_n27542_ );
nor  ( new_n27546_, new_n27545_, new_n27541_ );
not  ( new_n27547_, new_n27546_ );
and  ( new_n27548_, new_n27547_, new_n27536_ );
or   ( new_n27549_, new_n27548_, new_n27535_ );
or   ( new_n27550_, new_n1135_, new_n23895_ );
or   ( new_n27551_, new_n1137_, new_n23733_ );
and  ( new_n27552_, new_n27551_, new_n27550_ );
xor  ( new_n27553_, new_n27552_, new_n896_ );
or   ( new_n27554_, new_n897_, new_n24227_ );
or   ( new_n27555_, new_n899_, new_n24006_ );
and  ( new_n27556_, new_n27555_, new_n27554_ );
xor  ( new_n27557_, new_n27556_, new_n748_ );
or   ( new_n27558_, new_n27557_, new_n27553_ );
and  ( new_n27559_, new_n27557_, new_n27553_ );
or   ( new_n27560_, new_n755_, new_n24543_ );
or   ( new_n27561_, new_n757_, new_n24418_ );
and  ( new_n27562_, new_n27561_, new_n27560_ );
xor  ( new_n27563_, new_n27562_, new_n523_ );
or   ( new_n27564_, new_n27563_, new_n27559_ );
and  ( new_n27565_, new_n27564_, new_n27558_ );
or   ( new_n27566_, new_n1844_, new_n22973_ );
or   ( new_n27567_, new_n1846_, new_n22975_ );
and  ( new_n27568_, new_n27567_, new_n27566_ );
xor  ( new_n27569_, new_n27568_, new_n1586_ );
or   ( new_n27570_, new_n1593_, new_n23252_ );
or   ( new_n27571_, new_n1595_, new_n23166_ );
and  ( new_n27572_, new_n27571_, new_n27570_ );
xor  ( new_n27573_, new_n27572_, new_n1358_ );
or   ( new_n27574_, new_n27573_, new_n27569_ );
and  ( new_n27575_, new_n27573_, new_n27569_ );
or   ( new_n27576_, new_n1364_, new_n23554_ );
or   ( new_n27577_, new_n1366_, new_n23370_ );
and  ( new_n27578_, new_n27577_, new_n27576_ );
xor  ( new_n27579_, new_n27578_, new_n1129_ );
or   ( new_n27580_, new_n27579_, new_n27575_ );
and  ( new_n27581_, new_n27580_, new_n27574_ );
or   ( new_n27582_, new_n27581_, new_n27565_ );
and  ( new_n27583_, new_n27581_, new_n27565_ );
or   ( new_n27584_, new_n2807_, new_n22304_ );
or   ( new_n27585_, new_n2809_, new_n22207_ );
and  ( new_n27586_, new_n27585_, new_n27584_ );
xor  ( new_n27587_, new_n27586_, new_n2424_ );
or   ( new_n27588_, new_n2425_, new_n22590_ );
or   ( new_n27589_, new_n2427_, new_n22423_ );
and  ( new_n27590_, new_n27589_, new_n27588_ );
xor  ( new_n27591_, new_n27590_, new_n2121_ );
nor  ( new_n27592_, new_n27591_, new_n27587_ );
and  ( new_n27593_, new_n27591_, new_n27587_ );
or   ( new_n27594_, new_n2122_, new_n22829_ );
or   ( new_n27595_, new_n2124_, new_n22641_ );
and  ( new_n27596_, new_n27595_, new_n27594_ );
xor  ( new_n27597_, new_n27596_, new_n1843_ );
nor  ( new_n27598_, new_n27597_, new_n27593_ );
nor  ( new_n27599_, new_n27598_, new_n27592_ );
or   ( new_n27600_, new_n27599_, new_n27583_ );
and  ( new_n27601_, new_n27600_, new_n27582_ );
not  ( new_n27602_, RIbb32c70_177 );
or   ( new_n27603_, new_n268_, new_n27602_ );
or   ( new_n27604_, new_n271_, new_n27396_ );
and  ( new_n27605_, new_n27604_, new_n27603_ );
xor  ( new_n27606_, new_n27605_, new_n263_ );
and  ( new_n27607_, RIbb32ce8_178, RIbb2f610_1 );
or   ( new_n27608_, new_n27607_, new_n27606_ );
or   ( new_n27609_, new_n524_, new_n24925_ );
or   ( new_n27610_, new_n526_, new_n24927_ );
and  ( new_n27611_, new_n27610_, new_n27609_ );
xor  ( new_n27612_, new_n27611_, new_n403_ );
or   ( new_n27613_, new_n409_, new_n25288_ );
or   ( new_n27614_, new_n411_, new_n25048_ );
and  ( new_n27615_, new_n27614_, new_n27613_ );
xor  ( new_n27616_, new_n27615_, new_n328_ );
or   ( new_n27617_, new_n27616_, new_n27612_ );
and  ( new_n27618_, new_n27616_, new_n27612_ );
or   ( new_n27619_, new_n337_, new_n25813_ );
or   ( new_n27620_, new_n340_, new_n25486_ );
and  ( new_n27621_, new_n27620_, new_n27619_ );
xor  ( new_n27622_, new_n27621_, new_n332_ );
or   ( new_n27623_, new_n27622_, new_n27618_ );
and  ( new_n27624_, new_n27623_, new_n27617_ );
or   ( new_n27625_, new_n27624_, new_n27608_ );
and  ( new_n27626_, new_n27624_, new_n27608_ );
or   ( new_n27627_, new_n317_, new_n26063_ );
or   ( new_n27628_, new_n320_, new_n26196_ );
and  ( new_n27629_, new_n27628_, new_n27627_ );
xor  ( new_n27630_, new_n27629_, new_n312_ );
or   ( new_n27631_, new_n283_, new_n26620_ );
or   ( new_n27632_, new_n286_, new_n26372_ );
and  ( new_n27633_, new_n27632_, new_n27631_ );
xor  ( new_n27634_, new_n27633_, new_n278_ );
nor  ( new_n27635_, new_n27634_, new_n27630_ );
and  ( new_n27636_, new_n27634_, new_n27630_ );
or   ( new_n27637_, new_n299_, new_n27085_ );
or   ( new_n27638_, new_n302_, new_n26762_ );
and  ( new_n27639_, new_n27638_, new_n27637_ );
xor  ( new_n27640_, new_n27639_, new_n293_ );
nor  ( new_n27641_, new_n27640_, new_n27636_ );
nor  ( new_n27642_, new_n27641_, new_n27635_ );
or   ( new_n27643_, new_n27642_, new_n27626_ );
and  ( new_n27644_, new_n27643_, new_n27625_ );
or   ( new_n27645_, new_n27644_, new_n27601_ );
and  ( new_n27646_, new_n27644_, new_n27601_ );
or   ( new_n27647_, new_n5207_, new_n21680_ );
or   ( new_n27648_, new_n5209_, new_n21672_ );
and  ( new_n27649_, new_n27648_, new_n27647_ );
xor  ( new_n27650_, new_n27649_, new_n4708_ );
or   ( new_n27651_, new_n4709_, new_n21687_ );
or   ( new_n27652_, new_n4711_, new_n21678_ );
and  ( new_n27653_, new_n27652_, new_n27651_ );
xor  ( new_n27654_, new_n27653_, new_n4295_ );
or   ( new_n27655_, new_n27654_, new_n27650_ );
and  ( new_n27656_, new_n27654_, new_n27650_ );
or   ( new_n27657_, new_n4302_, new_n21751_ );
or   ( new_n27658_, new_n4304_, new_n21685_ );
and  ( new_n27659_, new_n27658_, new_n27657_ );
xor  ( new_n27660_, new_n27659_, new_n3895_ );
or   ( new_n27661_, new_n27660_, new_n27656_ );
and  ( new_n27662_, new_n27661_, new_n27655_ );
or   ( new_n27663_, new_n3896_, new_n21842_ );
or   ( new_n27664_, new_n3898_, new_n21792_ );
and  ( new_n27665_, new_n27664_, new_n27663_ );
xor  ( new_n27666_, new_n27665_, new_n3460_ );
or   ( new_n27667_, new_n3461_, new_n21847_ );
or   ( new_n27668_, new_n3463_, new_n21840_ );
and  ( new_n27669_, new_n27668_, new_n27667_ );
xor  ( new_n27670_, new_n27669_, new_n3116_ );
or   ( new_n27671_, new_n27670_, new_n27666_ );
and  ( new_n27672_, new_n27670_, new_n27666_ );
or   ( new_n27673_, new_n3117_, new_n22129_ );
or   ( new_n27674_, new_n3119_, new_n22098_ );
and  ( new_n27675_, new_n27674_, new_n27673_ );
xor  ( new_n27676_, new_n27675_, new_n2800_ );
or   ( new_n27677_, new_n27676_, new_n27672_ );
and  ( new_n27678_, new_n27677_, new_n27671_ );
nor  ( new_n27679_, new_n27678_, new_n27662_ );
and  ( new_n27680_, new_n27678_, new_n27662_ );
or   ( new_n27681_, new_n6173_, new_n21703_ );
or   ( new_n27682_, new_n6175_, new_n21694_ );
and  ( new_n27683_, new_n27682_, new_n27681_ );
xor  ( new_n27684_, new_n27683_, new_n5596_ );
and  ( new_n27685_, new_n6510_, RIbb315f0_129 );
xor  ( new_n27686_, new_n27685_, new_n6166_ );
and  ( new_n27687_, new_n27686_, new_n27684_ );
nor  ( new_n27688_, new_n27686_, new_n27684_ );
or   ( new_n27689_, new_n5604_, new_n21674_ );
or   ( new_n27690_, new_n5606_, new_n21701_ );
and  ( new_n27691_, new_n27690_, new_n27689_ );
xor  ( new_n27692_, new_n27691_, new_n5206_ );
nor  ( new_n27693_, new_n27692_, new_n27688_ );
nor  ( new_n27694_, new_n27693_, new_n27687_ );
nor  ( new_n27695_, new_n27694_, new_n27680_ );
nor  ( new_n27696_, new_n27695_, new_n27679_ );
or   ( new_n27697_, new_n27696_, new_n27646_ );
and  ( new_n27698_, new_n27697_, new_n27645_ );
and  ( new_n27699_, new_n27698_, new_n27549_ );
nor  ( new_n27700_, new_n27698_, new_n27549_ );
xnor ( new_n27701_, new_n27267_, new_n27265_ );
xor  ( new_n27702_, new_n27701_, new_n27271_ );
xnor ( new_n27703_, new_n27247_, new_n27245_ );
xor  ( new_n27704_, new_n27703_, new_n27251_ );
and  ( new_n27705_, new_n27704_, new_n27702_ );
nor  ( new_n27706_, new_n27704_, new_n27702_ );
xor  ( new_n27707_, new_n27257_, new_n27255_ );
xnor ( new_n27708_, new_n27707_, new_n27443_ );
nor  ( new_n27709_, new_n27708_, new_n27706_ );
nor  ( new_n27710_, new_n27709_, new_n27705_ );
nor  ( new_n27711_, new_n27710_, new_n27700_ );
nor  ( new_n27712_, new_n27711_, new_n27699_ );
nor  ( new_n27713_, new_n27712_, new_n27515_ );
nor  ( new_n27714_, new_n27713_, new_n27514_ );
not  ( new_n27715_, new_n27714_ );
and  ( new_n27716_, new_n27715_, new_n27490_ );
or   ( new_n27717_, new_n27716_, new_n27489_ );
xnor ( new_n27718_, new_n27187_, new_n26995_ );
xor  ( new_n27719_, new_n27718_, new_n27206_ );
nand ( new_n27720_, new_n27719_, new_n27717_ );
or   ( new_n27721_, new_n27719_, new_n27717_ );
xor  ( new_n27722_, new_n27236_, new_n27234_ );
xor  ( new_n27723_, new_n27722_, new_n27462_ );
nand ( new_n27724_, new_n27723_, new_n27721_ );
and  ( new_n27725_, new_n27724_, new_n27720_ );
nor  ( new_n27726_, new_n27725_, new_n27477_ );
xor  ( new_n27727_, new_n27472_, new_n27225_ );
and  ( new_n27728_, new_n27727_, new_n27726_ );
xnor ( new_n27729_, new_n27438_, new_n27243_ );
xor  ( new_n27730_, new_n27729_, new_n27459_ );
xnor ( new_n27731_, new_n27698_, new_n27549_ );
xor  ( new_n27732_, new_n27731_, new_n27710_ );
xnor ( new_n27733_, new_n27499_, new_n27497_ );
xor  ( new_n27734_, new_n27733_, new_n27511_ );
nor  ( new_n27735_, new_n27734_, new_n27732_ );
nand ( new_n27736_, new_n27734_, new_n27732_ );
xnor ( new_n27737_, new_n27494_, new_n27492_ );
and  ( new_n27738_, new_n27737_, new_n27736_ );
or   ( new_n27739_, new_n27738_, new_n27735_ );
xor  ( new_n27740_, new_n27481_, new_n27479_ );
xor  ( new_n27741_, new_n27740_, new_n27484_ );
nand ( new_n27742_, new_n27741_, new_n27739_ );
nor  ( new_n27743_, new_n27741_, new_n27739_ );
xor  ( new_n27744_, new_n27534_, new_n27525_ );
xor  ( new_n27745_, new_n27744_, new_n27547_ );
xnor ( new_n27746_, new_n27644_, new_n27601_ );
xnor ( new_n27747_, new_n27746_, new_n27696_ );
and  ( new_n27748_, new_n27747_, new_n27745_ );
xnor ( new_n27749_, new_n27540_, new_n27538_ );
xor  ( new_n27750_, new_n27749_, new_n27544_ );
xnor ( new_n27751_, new_n27519_, new_n27517_ );
xor  ( new_n27752_, new_n27751_, new_n27523_ );
or   ( new_n27753_, new_n27752_, new_n27750_ );
and  ( new_n27754_, new_n27752_, new_n27750_ );
xor  ( new_n27755_, new_n27529_, new_n27527_ );
xor  ( new_n27756_, new_n27755_, new_n27532_ );
or   ( new_n27757_, new_n27756_, new_n27754_ );
and  ( new_n27758_, new_n27757_, new_n27753_ );
or   ( new_n27759_, new_n299_, new_n27396_ );
or   ( new_n27760_, new_n302_, new_n27085_ );
and  ( new_n27761_, new_n27760_, new_n27759_ );
xor  ( new_n27762_, new_n27761_, new_n293_ );
not  ( new_n27763_, RIbb32ce8_178 );
or   ( new_n27764_, new_n268_, new_n27763_ );
or   ( new_n27765_, new_n271_, new_n27602_ );
and  ( new_n27766_, new_n27765_, new_n27764_ );
xor  ( new_n27767_, new_n27766_, new_n263_ );
or   ( new_n27768_, new_n27767_, new_n27762_ );
and  ( new_n27769_, RIbb32d60_179, RIbb2f610_1 );
and  ( new_n27770_, new_n27767_, new_n27762_ );
or   ( new_n27771_, new_n27770_, new_n27769_ );
and  ( new_n27772_, new_n27771_, new_n27768_ );
or   ( new_n27773_, new_n755_, new_n24927_ );
or   ( new_n27774_, new_n757_, new_n24543_ );
and  ( new_n27775_, new_n27774_, new_n27773_ );
xor  ( new_n27776_, new_n27775_, new_n523_ );
or   ( new_n27777_, new_n524_, new_n25048_ );
or   ( new_n27778_, new_n526_, new_n24925_ );
and  ( new_n27779_, new_n27778_, new_n27777_ );
xor  ( new_n27780_, new_n27779_, new_n403_ );
or   ( new_n27781_, new_n27780_, new_n27776_ );
and  ( new_n27782_, new_n27780_, new_n27776_ );
or   ( new_n27783_, new_n409_, new_n25486_ );
or   ( new_n27784_, new_n411_, new_n25288_ );
and  ( new_n27785_, new_n27784_, new_n27783_ );
xor  ( new_n27786_, new_n27785_, new_n328_ );
or   ( new_n27787_, new_n27786_, new_n27782_ );
and  ( new_n27788_, new_n27787_, new_n27781_ );
or   ( new_n27789_, new_n27788_, new_n27772_ );
and  ( new_n27790_, new_n27788_, new_n27772_ );
or   ( new_n27791_, new_n337_, new_n26196_ );
or   ( new_n27792_, new_n340_, new_n25813_ );
and  ( new_n27793_, new_n27792_, new_n27791_ );
xor  ( new_n27794_, new_n27793_, new_n332_ );
or   ( new_n27795_, new_n317_, new_n26372_ );
or   ( new_n27796_, new_n320_, new_n26063_ );
and  ( new_n27797_, new_n27796_, new_n27795_ );
xor  ( new_n27798_, new_n27797_, new_n312_ );
nor  ( new_n27799_, new_n27798_, new_n27794_ );
and  ( new_n27800_, new_n27798_, new_n27794_ );
or   ( new_n27801_, new_n283_, new_n26762_ );
or   ( new_n27802_, new_n286_, new_n26620_ );
and  ( new_n27803_, new_n27802_, new_n27801_ );
xor  ( new_n27804_, new_n27803_, new_n278_ );
nor  ( new_n27805_, new_n27804_, new_n27800_ );
nor  ( new_n27806_, new_n27805_, new_n27799_ );
or   ( new_n27807_, new_n27806_, new_n27790_ );
and  ( new_n27808_, new_n27807_, new_n27789_ );
or   ( new_n27809_, new_n6173_, new_n21701_ );
or   ( new_n27810_, new_n6175_, new_n21703_ );
and  ( new_n27811_, new_n27810_, new_n27809_ );
xor  ( new_n27812_, new_n27811_, new_n5597_ );
and  ( new_n27813_, new_n27812_, new_n6638_ );
or   ( new_n27814_, new_n27812_, new_n6638_ );
or   ( new_n27815_, new_n6645_, new_n21694_ );
or   ( new_n27816_, new_n6647_, new_n21696_ );
and  ( new_n27817_, new_n27816_, new_n27815_ );
xor  ( new_n27818_, new_n27817_, new_n6166_ );
and  ( new_n27819_, new_n27818_, new_n27814_ );
or   ( new_n27820_, new_n27819_, new_n27813_ );
or   ( new_n27821_, new_n5604_, new_n21672_ );
or   ( new_n27822_, new_n5606_, new_n21674_ );
and  ( new_n27823_, new_n27822_, new_n27821_ );
xor  ( new_n27824_, new_n27823_, new_n5206_ );
or   ( new_n27825_, new_n5207_, new_n21678_ );
or   ( new_n27826_, new_n5209_, new_n21680_ );
and  ( new_n27827_, new_n27826_, new_n27825_ );
xor  ( new_n27828_, new_n27827_, new_n4708_ );
or   ( new_n27829_, new_n27828_, new_n27824_ );
and  ( new_n27830_, new_n27828_, new_n27824_ );
or   ( new_n27831_, new_n4709_, new_n21685_ );
or   ( new_n27832_, new_n4711_, new_n21687_ );
and  ( new_n27833_, new_n27832_, new_n27831_ );
xor  ( new_n27834_, new_n27833_, new_n4295_ );
or   ( new_n27835_, new_n27834_, new_n27830_ );
and  ( new_n27836_, new_n27835_, new_n27829_ );
or   ( new_n27837_, new_n27836_, new_n27820_ );
and  ( new_n27838_, new_n27836_, new_n27820_ );
or   ( new_n27839_, new_n4302_, new_n21792_ );
or   ( new_n27840_, new_n4304_, new_n21751_ );
and  ( new_n27841_, new_n27840_, new_n27839_ );
xor  ( new_n27842_, new_n27841_, new_n3895_ );
or   ( new_n27843_, new_n3896_, new_n21840_ );
or   ( new_n27844_, new_n3898_, new_n21842_ );
and  ( new_n27845_, new_n27844_, new_n27843_ );
xor  ( new_n27846_, new_n27845_, new_n3460_ );
nor  ( new_n27847_, new_n27846_, new_n27842_ );
and  ( new_n27848_, new_n27846_, new_n27842_ );
or   ( new_n27849_, new_n3461_, new_n22098_ );
or   ( new_n27850_, new_n3463_, new_n21847_ );
and  ( new_n27851_, new_n27850_, new_n27849_ );
xor  ( new_n27852_, new_n27851_, new_n3116_ );
nor  ( new_n27853_, new_n27852_, new_n27848_ );
nor  ( new_n27854_, new_n27853_, new_n27847_ );
or   ( new_n27855_, new_n27854_, new_n27838_ );
and  ( new_n27856_, new_n27855_, new_n27837_ );
or   ( new_n27857_, new_n27856_, new_n27808_ );
and  ( new_n27858_, new_n27856_, new_n27808_ );
or   ( new_n27859_, new_n2122_, new_n22975_ );
or   ( new_n27860_, new_n2124_, new_n22829_ );
and  ( new_n27861_, new_n27860_, new_n27859_ );
xor  ( new_n27862_, new_n27861_, new_n1843_ );
or   ( new_n27863_, new_n1844_, new_n23166_ );
or   ( new_n27864_, new_n1846_, new_n22973_ );
and  ( new_n27865_, new_n27864_, new_n27863_ );
xor  ( new_n27866_, new_n27865_, new_n1586_ );
or   ( new_n27867_, new_n27866_, new_n27862_ );
and  ( new_n27868_, new_n27866_, new_n27862_ );
or   ( new_n27869_, new_n1593_, new_n23370_ );
or   ( new_n27870_, new_n1595_, new_n23252_ );
and  ( new_n27871_, new_n27870_, new_n27869_ );
xor  ( new_n27872_, new_n27871_, new_n1358_ );
or   ( new_n27873_, new_n27872_, new_n27868_ );
and  ( new_n27874_, new_n27873_, new_n27867_ );
or   ( new_n27875_, new_n3117_, new_n22207_ );
or   ( new_n27876_, new_n3119_, new_n22129_ );
and  ( new_n27877_, new_n27876_, new_n27875_ );
xor  ( new_n27878_, new_n27877_, new_n2800_ );
or   ( new_n27879_, new_n2807_, new_n22423_ );
or   ( new_n27880_, new_n2809_, new_n22304_ );
and  ( new_n27881_, new_n27880_, new_n27879_ );
xor  ( new_n27882_, new_n27881_, new_n2424_ );
or   ( new_n27883_, new_n27882_, new_n27878_ );
and  ( new_n27884_, new_n27882_, new_n27878_ );
or   ( new_n27885_, new_n2425_, new_n22641_ );
or   ( new_n27886_, new_n2427_, new_n22590_ );
and  ( new_n27887_, new_n27886_, new_n27885_ );
xor  ( new_n27888_, new_n27887_, new_n2121_ );
or   ( new_n27889_, new_n27888_, new_n27884_ );
and  ( new_n27890_, new_n27889_, new_n27883_ );
nor  ( new_n27891_, new_n27890_, new_n27874_ );
and  ( new_n27892_, new_n27890_, new_n27874_ );
or   ( new_n27893_, new_n1364_, new_n23733_ );
or   ( new_n27894_, new_n1366_, new_n23554_ );
and  ( new_n27895_, new_n27894_, new_n27893_ );
xor  ( new_n27896_, new_n27895_, new_n1129_ );
or   ( new_n27897_, new_n1135_, new_n24006_ );
or   ( new_n27898_, new_n1137_, new_n23895_ );
and  ( new_n27899_, new_n27898_, new_n27897_ );
xor  ( new_n27900_, new_n27899_, new_n896_ );
nor  ( new_n27901_, new_n27900_, new_n27896_ );
and  ( new_n27902_, new_n27900_, new_n27896_ );
or   ( new_n27903_, new_n897_, new_n24418_ );
or   ( new_n27904_, new_n899_, new_n24227_ );
and  ( new_n27905_, new_n27904_, new_n27903_ );
xor  ( new_n27906_, new_n27905_, new_n748_ );
nor  ( new_n27907_, new_n27906_, new_n27902_ );
nor  ( new_n27908_, new_n27907_, new_n27901_ );
nor  ( new_n27909_, new_n27908_, new_n27892_ );
nor  ( new_n27910_, new_n27909_, new_n27891_ );
or   ( new_n27911_, new_n27910_, new_n27858_ );
and  ( new_n27912_, new_n27911_, new_n27857_ );
or   ( new_n27913_, new_n27912_, new_n27758_ );
nand ( new_n27914_, new_n27912_, new_n27758_ );
xnor ( new_n27915_, new_n27670_, new_n27666_ );
xor  ( new_n27916_, new_n27915_, new_n27676_ );
xnor ( new_n27917_, new_n27654_, new_n27650_ );
xor  ( new_n27918_, new_n27917_, new_n27660_ );
or   ( new_n27919_, new_n27918_, new_n27916_ );
and  ( new_n27920_, new_n27918_, new_n27916_ );
xor  ( new_n27921_, new_n27686_, new_n27684_ );
xnor ( new_n27922_, new_n27921_, new_n27692_ );
or   ( new_n27923_, new_n27922_, new_n27920_ );
and  ( new_n27924_, new_n27923_, new_n27919_ );
xnor ( new_n27925_, new_n27616_, new_n27612_ );
xor  ( new_n27926_, new_n27925_, new_n27622_ );
xnor ( new_n27927_, new_n27634_, new_n27630_ );
xor  ( new_n27928_, new_n27927_, new_n27640_ );
or   ( new_n27929_, new_n27928_, new_n27926_ );
and  ( new_n27930_, new_n27928_, new_n27926_ );
xor  ( new_n27931_, new_n27607_, new_n27606_ );
or   ( new_n27932_, new_n27931_, new_n27930_ );
and  ( new_n27933_, new_n27932_, new_n27929_ );
nor  ( new_n27934_, new_n27933_, new_n27924_ );
and  ( new_n27935_, new_n27933_, new_n27924_ );
xnor ( new_n27936_, new_n27573_, new_n27569_ );
xor  ( new_n27937_, new_n27936_, new_n27579_ );
xnor ( new_n27938_, new_n27557_, new_n27553_ );
xor  ( new_n27939_, new_n27938_, new_n27563_ );
nor  ( new_n27940_, new_n27939_, new_n27937_ );
and  ( new_n27941_, new_n27939_, new_n27937_ );
xor  ( new_n27942_, new_n27591_, new_n27587_ );
xnor ( new_n27943_, new_n27942_, new_n27597_ );
nor  ( new_n27944_, new_n27943_, new_n27941_ );
nor  ( new_n27945_, new_n27944_, new_n27940_ );
nor  ( new_n27946_, new_n27945_, new_n27935_ );
nor  ( new_n27947_, new_n27946_, new_n27934_ );
nand ( new_n27948_, new_n27947_, new_n27914_ );
and  ( new_n27949_, new_n27948_, new_n27913_ );
nor  ( new_n27950_, new_n27949_, new_n27748_ );
and  ( new_n27951_, new_n27949_, new_n27748_ );
xnor ( new_n27952_, new_n27581_, new_n27565_ );
xor  ( new_n27953_, new_n27952_, new_n27599_ );
xnor ( new_n27954_, new_n27624_, new_n27608_ );
xor  ( new_n27955_, new_n27954_, new_n27642_ );
nor  ( new_n27956_, new_n27955_, new_n27953_ );
nand ( new_n27957_, new_n27955_, new_n27953_ );
xor  ( new_n27958_, new_n27678_, new_n27662_ );
xor  ( new_n27959_, new_n27958_, new_n27694_ );
and  ( new_n27960_, new_n27959_, new_n27957_ );
or   ( new_n27961_, new_n27960_, new_n27956_ );
xnor ( new_n27962_, new_n27704_, new_n27702_ );
xor  ( new_n27963_, new_n27962_, new_n27708_ );
nor  ( new_n27964_, new_n27963_, new_n27961_ );
and  ( new_n27965_, new_n27963_, new_n27961_ );
xor  ( new_n27966_, new_n27505_, new_n27503_ );
xnor ( new_n27967_, new_n27966_, new_n27509_ );
nor  ( new_n27968_, new_n27967_, new_n27965_ );
nor  ( new_n27969_, new_n27968_, new_n27964_ );
nor  ( new_n27970_, new_n27969_, new_n27951_ );
nor  ( new_n27971_, new_n27970_, new_n27950_ );
or   ( new_n27972_, new_n27971_, new_n27743_ );
and  ( new_n27973_, new_n27972_, new_n27742_ );
or   ( new_n27974_, new_n27973_, new_n27730_ );
and  ( new_n27975_, new_n27973_, new_n27730_ );
xor  ( new_n27976_, new_n27488_, new_n27486_ );
xor  ( new_n27977_, new_n27976_, new_n27715_ );
or   ( new_n27978_, new_n27977_, new_n27975_ );
and  ( new_n27979_, new_n27978_, new_n27974_ );
xor  ( new_n27980_, new_n27719_, new_n27717_ );
xor  ( new_n27981_, new_n27980_, new_n27723_ );
and  ( new_n27982_, new_n27981_, new_n27979_ );
xor  ( new_n27983_, new_n27725_, new_n27477_ );
and  ( new_n27984_, new_n27983_, new_n27982_ );
xor  ( new_n27985_, new_n27734_, new_n27732_ );
xor  ( new_n27986_, new_n27985_, new_n27737_ );
xor  ( new_n27987_, new_n27912_, new_n27758_ );
xor  ( new_n27988_, new_n27987_, new_n27947_ );
xnor ( new_n27989_, new_n27963_, new_n27961_ );
xor  ( new_n27990_, new_n27989_, new_n27967_ );
or   ( new_n27991_, new_n27990_, new_n27988_ );
and  ( new_n27992_, new_n27990_, new_n27988_ );
xnor ( new_n27993_, new_n27747_, new_n27745_ );
or   ( new_n27994_, new_n27993_, new_n27992_ );
and  ( new_n27995_, new_n27994_, new_n27991_ );
nor  ( new_n27996_, new_n27995_, new_n27986_ );
and  ( new_n27997_, new_n27995_, new_n27986_ );
xor  ( new_n27998_, new_n27933_, new_n27924_ );
xnor ( new_n27999_, new_n27998_, new_n27945_ );
xnor ( new_n28000_, new_n27856_, new_n27808_ );
xnor ( new_n28001_, new_n28000_, new_n27910_ );
and  ( new_n28002_, new_n28001_, new_n27999_ );
xnor ( new_n28003_, new_n27882_, new_n27878_ );
xor  ( new_n28004_, new_n28003_, new_n27888_ );
xnor ( new_n28005_, new_n27866_, new_n27862_ );
xor  ( new_n28006_, new_n28005_, new_n27872_ );
or   ( new_n28007_, new_n28006_, new_n28004_ );
and  ( new_n28008_, new_n28006_, new_n28004_ );
xor  ( new_n28009_, new_n27900_, new_n27896_ );
xnor ( new_n28010_, new_n28009_, new_n27906_ );
or   ( new_n28011_, new_n28010_, new_n28008_ );
and  ( new_n28012_, new_n28011_, new_n28007_ );
xnor ( new_n28013_, new_n27828_, new_n27824_ );
xor  ( new_n28014_, new_n28013_, new_n27834_ );
xnor ( new_n28015_, new_n27846_, new_n27842_ );
xor  ( new_n28016_, new_n28015_, new_n27852_ );
or   ( new_n28017_, new_n28016_, new_n28014_ );
and  ( new_n28018_, new_n28016_, new_n28014_ );
xor  ( new_n28019_, new_n27812_, new_n6638_ );
xor  ( new_n28020_, new_n28019_, new_n27818_ );
not  ( new_n28021_, new_n28020_ );
or   ( new_n28022_, new_n28021_, new_n28018_ );
and  ( new_n28023_, new_n28022_, new_n28017_ );
nor  ( new_n28024_, new_n28023_, new_n28012_ );
nand ( new_n28025_, new_n28023_, new_n28012_ );
xnor ( new_n28026_, new_n27767_, new_n27762_ );
xor  ( new_n28027_, new_n28026_, new_n27769_ );
xnor ( new_n28028_, new_n27780_, new_n27776_ );
xor  ( new_n28029_, new_n28028_, new_n27786_ );
nor  ( new_n28030_, new_n28029_, new_n28027_ );
nand ( new_n28031_, new_n28029_, new_n28027_ );
xor  ( new_n28032_, new_n27798_, new_n27794_ );
xor  ( new_n28033_, new_n28032_, new_n27804_ );
and  ( new_n28034_, new_n28033_, new_n28031_ );
or   ( new_n28035_, new_n28034_, new_n28030_ );
and  ( new_n28036_, new_n28035_, new_n28025_ );
or   ( new_n28037_, new_n28036_, new_n28024_ );
or   ( new_n28038_, new_n4302_, new_n21842_ );
or   ( new_n28039_, new_n4304_, new_n21792_ );
and  ( new_n28040_, new_n28039_, new_n28038_ );
xor  ( new_n28041_, new_n28040_, new_n3895_ );
or   ( new_n28042_, new_n3896_, new_n21847_ );
or   ( new_n28043_, new_n3898_, new_n21840_ );
and  ( new_n28044_, new_n28043_, new_n28042_ );
xor  ( new_n28045_, new_n28044_, new_n3460_ );
or   ( new_n28046_, new_n28045_, new_n28041_ );
and  ( new_n28047_, new_n28045_, new_n28041_ );
or   ( new_n28048_, new_n3461_, new_n22129_ );
or   ( new_n28049_, new_n3463_, new_n22098_ );
and  ( new_n28050_, new_n28049_, new_n28048_ );
xor  ( new_n28051_, new_n28050_, new_n3116_ );
or   ( new_n28052_, new_n28051_, new_n28047_ );
and  ( new_n28053_, new_n28052_, new_n28046_ );
or   ( new_n28054_, new_n5604_, new_n21680_ );
or   ( new_n28055_, new_n5606_, new_n21672_ );
and  ( new_n28056_, new_n28055_, new_n28054_ );
xor  ( new_n28057_, new_n28056_, new_n5206_ );
or   ( new_n28058_, new_n5207_, new_n21687_ );
or   ( new_n28059_, new_n5209_, new_n21678_ );
and  ( new_n28060_, new_n28059_, new_n28058_ );
xor  ( new_n28061_, new_n28060_, new_n4708_ );
or   ( new_n28062_, new_n28061_, new_n28057_ );
and  ( new_n28063_, new_n28061_, new_n28057_ );
or   ( new_n28064_, new_n4709_, new_n21751_ );
or   ( new_n28065_, new_n4711_, new_n21685_ );
and  ( new_n28066_, new_n28065_, new_n28064_ );
xor  ( new_n28067_, new_n28066_, new_n4295_ );
or   ( new_n28068_, new_n28067_, new_n28063_ );
and  ( new_n28069_, new_n28068_, new_n28062_ );
or   ( new_n28070_, new_n28069_, new_n28053_ );
and  ( new_n28071_, new_n28069_, new_n28053_ );
or   ( new_n28072_, new_n6645_, new_n21703_ );
or   ( new_n28073_, new_n6647_, new_n21694_ );
and  ( new_n28074_, new_n28073_, new_n28072_ );
xor  ( new_n28075_, new_n28074_, new_n6165_ );
and  ( new_n28076_, new_n6910_, RIbb315f0_129 );
xor  ( new_n28077_, new_n28076_, new_n6638_ );
and  ( new_n28078_, new_n28077_, new_n28075_ );
nor  ( new_n28079_, new_n28077_, new_n28075_ );
or   ( new_n28080_, new_n6173_, new_n21674_ );
or   ( new_n28081_, new_n6175_, new_n21701_ );
and  ( new_n28082_, new_n28081_, new_n28080_ );
xor  ( new_n28083_, new_n28082_, new_n5597_ );
nor  ( new_n28084_, new_n28083_, new_n28079_ );
nor  ( new_n28085_, new_n28084_, new_n28078_ );
or   ( new_n28086_, new_n28085_, new_n28071_ );
and  ( new_n28087_, new_n28086_, new_n28070_ );
or   ( new_n28088_, new_n755_, new_n24925_ );
or   ( new_n28089_, new_n757_, new_n24927_ );
and  ( new_n28090_, new_n28089_, new_n28088_ );
xor  ( new_n28091_, new_n28090_, new_n523_ );
or   ( new_n28092_, new_n524_, new_n25288_ );
or   ( new_n28093_, new_n526_, new_n25048_ );
and  ( new_n28094_, new_n28093_, new_n28092_ );
xor  ( new_n28095_, new_n28094_, new_n403_ );
or   ( new_n28096_, new_n28095_, new_n28091_ );
and  ( new_n28097_, new_n28095_, new_n28091_ );
or   ( new_n28098_, new_n409_, new_n25813_ );
or   ( new_n28099_, new_n411_, new_n25486_ );
and  ( new_n28100_, new_n28099_, new_n28098_ );
xor  ( new_n28101_, new_n28100_, new_n328_ );
or   ( new_n28102_, new_n28101_, new_n28097_ );
and  ( new_n28103_, new_n28102_, new_n28096_ );
or   ( new_n28104_, new_n299_, new_n27602_ );
or   ( new_n28105_, new_n302_, new_n27396_ );
and  ( new_n28106_, new_n28105_, new_n28104_ );
xor  ( new_n28107_, new_n28106_, new_n293_ );
not  ( new_n28108_, RIbb32d60_179 );
or   ( new_n28109_, new_n268_, new_n28108_ );
or   ( new_n28110_, new_n271_, new_n27763_ );
and  ( new_n28111_, new_n28110_, new_n28109_ );
xor  ( new_n28112_, new_n28111_, new_n263_ );
nor  ( new_n28113_, new_n28112_, new_n28107_ );
and  ( new_n28114_, RIbb32dd8_180, RIbb2f610_1 );
and  ( new_n28115_, new_n28112_, new_n28107_ );
nor  ( new_n28116_, new_n28115_, new_n28114_ );
nor  ( new_n28117_, new_n28116_, new_n28113_ );
or   ( new_n28118_, new_n337_, new_n26063_ );
or   ( new_n28119_, new_n340_, new_n26196_ );
and  ( new_n28120_, new_n28119_, new_n28118_ );
xor  ( new_n28121_, new_n28120_, new_n332_ );
or   ( new_n28122_, new_n317_, new_n26620_ );
or   ( new_n28123_, new_n320_, new_n26372_ );
and  ( new_n28124_, new_n28123_, new_n28122_ );
xor  ( new_n28125_, new_n28124_, new_n312_ );
or   ( new_n28126_, new_n28125_, new_n28121_ );
and  ( new_n28127_, new_n28125_, new_n28121_ );
or   ( new_n28128_, new_n283_, new_n27085_ );
or   ( new_n28129_, new_n286_, new_n26762_ );
and  ( new_n28130_, new_n28129_, new_n28128_ );
xor  ( new_n28131_, new_n28130_, new_n278_ );
or   ( new_n28132_, new_n28131_, new_n28127_ );
and  ( new_n28133_, new_n28132_, new_n28126_ );
and  ( new_n28134_, new_n28133_, new_n28117_ );
or   ( new_n28135_, new_n28134_, new_n28103_ );
or   ( new_n28136_, new_n28133_, new_n28117_ );
and  ( new_n28137_, new_n28136_, new_n28135_ );
or   ( new_n28138_, new_n28137_, new_n28087_ );
or   ( new_n28139_, new_n2122_, new_n22973_ );
or   ( new_n28140_, new_n2124_, new_n22975_ );
and  ( new_n28141_, new_n28140_, new_n28139_ );
xor  ( new_n28142_, new_n28141_, new_n1843_ );
or   ( new_n28143_, new_n1844_, new_n23252_ );
or   ( new_n28144_, new_n1846_, new_n23166_ );
and  ( new_n28145_, new_n28144_, new_n28143_ );
xor  ( new_n28146_, new_n28145_, new_n1586_ );
or   ( new_n28147_, new_n28146_, new_n28142_ );
and  ( new_n28148_, new_n28146_, new_n28142_ );
or   ( new_n28149_, new_n1593_, new_n23554_ );
or   ( new_n28150_, new_n1595_, new_n23370_ );
and  ( new_n28151_, new_n28150_, new_n28149_ );
xor  ( new_n28152_, new_n28151_, new_n1358_ );
or   ( new_n28153_, new_n28152_, new_n28148_ );
and  ( new_n28154_, new_n28153_, new_n28147_ );
or   ( new_n28155_, new_n3117_, new_n22304_ );
or   ( new_n28156_, new_n3119_, new_n22207_ );
and  ( new_n28157_, new_n28156_, new_n28155_ );
xor  ( new_n28158_, new_n28157_, new_n2800_ );
or   ( new_n28159_, new_n2807_, new_n22590_ );
or   ( new_n28160_, new_n2809_, new_n22423_ );
and  ( new_n28161_, new_n28160_, new_n28159_ );
xor  ( new_n28162_, new_n28161_, new_n2424_ );
or   ( new_n28163_, new_n28162_, new_n28158_ );
and  ( new_n28164_, new_n28162_, new_n28158_ );
or   ( new_n28165_, new_n2425_, new_n22829_ );
or   ( new_n28166_, new_n2427_, new_n22641_ );
and  ( new_n28167_, new_n28166_, new_n28165_ );
xor  ( new_n28168_, new_n28167_, new_n2121_ );
or   ( new_n28169_, new_n28168_, new_n28164_ );
and  ( new_n28170_, new_n28169_, new_n28163_ );
nor  ( new_n28171_, new_n28170_, new_n28154_ );
and  ( new_n28172_, new_n28170_, new_n28154_ );
or   ( new_n28173_, new_n1364_, new_n23895_ );
or   ( new_n28174_, new_n1366_, new_n23733_ );
and  ( new_n28175_, new_n28174_, new_n28173_ );
xor  ( new_n28176_, new_n28175_, new_n1129_ );
or   ( new_n28177_, new_n1135_, new_n24227_ );
or   ( new_n28178_, new_n1137_, new_n24006_ );
and  ( new_n28179_, new_n28178_, new_n28177_ );
xor  ( new_n28180_, new_n28179_, new_n896_ );
nor  ( new_n28181_, new_n28180_, new_n28176_ );
and  ( new_n28182_, new_n28180_, new_n28176_ );
or   ( new_n28183_, new_n897_, new_n24543_ );
or   ( new_n28184_, new_n899_, new_n24418_ );
and  ( new_n28185_, new_n28184_, new_n28183_ );
xor  ( new_n28186_, new_n28185_, new_n748_ );
nor  ( new_n28187_, new_n28186_, new_n28182_ );
nor  ( new_n28188_, new_n28187_, new_n28181_ );
nor  ( new_n28189_, new_n28188_, new_n28172_ );
nor  ( new_n28190_, new_n28189_, new_n28171_ );
and  ( new_n28191_, new_n28137_, new_n28087_ );
or   ( new_n28192_, new_n28191_, new_n28190_ );
and  ( new_n28193_, new_n28192_, new_n28138_ );
or   ( new_n28194_, new_n28193_, new_n28037_ );
and  ( new_n28195_, new_n28193_, new_n28037_ );
xnor ( new_n28196_, new_n27939_, new_n27937_ );
xor  ( new_n28197_, new_n28196_, new_n27943_ );
xnor ( new_n28198_, new_n27918_, new_n27916_ );
xor  ( new_n28199_, new_n28198_, new_n27922_ );
and  ( new_n28200_, new_n28199_, new_n28197_ );
or   ( new_n28201_, new_n28199_, new_n28197_ );
xor  ( new_n28202_, new_n27928_, new_n27926_ );
xor  ( new_n28203_, new_n28202_, new_n27931_ );
not  ( new_n28204_, new_n28203_ );
and  ( new_n28205_, new_n28204_, new_n28201_ );
or   ( new_n28206_, new_n28205_, new_n28200_ );
or   ( new_n28207_, new_n28206_, new_n28195_ );
and  ( new_n28208_, new_n28207_, new_n28194_ );
and  ( new_n28209_, new_n28208_, new_n28002_ );
nor  ( new_n28210_, new_n28208_, new_n28002_ );
xnor ( new_n28211_, new_n27788_, new_n27772_ );
xor  ( new_n28212_, new_n28211_, new_n27806_ );
xnor ( new_n28213_, new_n27836_, new_n27820_ );
xor  ( new_n28214_, new_n28213_, new_n27854_ );
nor  ( new_n28215_, new_n28214_, new_n28212_ );
nand ( new_n28216_, new_n28214_, new_n28212_ );
xor  ( new_n28217_, new_n27890_, new_n27874_ );
xor  ( new_n28218_, new_n28217_, new_n27908_ );
and  ( new_n28219_, new_n28218_, new_n28216_ );
or   ( new_n28220_, new_n28219_, new_n28215_ );
xor  ( new_n28221_, new_n27955_, new_n27953_ );
xor  ( new_n28222_, new_n28221_, new_n27959_ );
and  ( new_n28223_, new_n28222_, new_n28220_ );
nor  ( new_n28224_, new_n28222_, new_n28220_ );
xor  ( new_n28225_, new_n27752_, new_n27750_ );
xnor ( new_n28226_, new_n28225_, new_n27756_ );
nor  ( new_n28227_, new_n28226_, new_n28224_ );
nor  ( new_n28228_, new_n28227_, new_n28223_ );
nor  ( new_n28229_, new_n28228_, new_n28210_ );
nor  ( new_n28230_, new_n28229_, new_n28209_ );
nor  ( new_n28231_, new_n28230_, new_n27997_ );
or   ( new_n28232_, new_n28231_, new_n27996_ );
xnor ( new_n28233_, new_n27513_, new_n27495_ );
xor  ( new_n28234_, new_n28233_, new_n27712_ );
nor  ( new_n28235_, new_n28234_, new_n28232_ );
nand ( new_n28236_, new_n28234_, new_n28232_ );
xnor ( new_n28237_, new_n27741_, new_n27739_ );
xor  ( new_n28238_, new_n28237_, new_n27971_ );
and  ( new_n28239_, new_n28238_, new_n28236_ );
or   ( new_n28240_, new_n28239_, new_n28235_ );
xnor ( new_n28241_, new_n27973_, new_n27730_ );
xor  ( new_n28242_, new_n28241_, new_n27977_ );
nor  ( new_n28243_, new_n28242_, new_n28240_ );
xor  ( new_n28244_, new_n27981_, new_n27979_ );
and  ( new_n28245_, new_n28244_, new_n28243_ );
xor  ( new_n28246_, new_n27995_, new_n27986_ );
xor  ( new_n28247_, new_n28246_, new_n28230_ );
xnor ( new_n28248_, new_n27949_, new_n27748_ );
xor  ( new_n28249_, new_n28248_, new_n27969_ );
or   ( new_n28250_, new_n28249_, new_n28247_ );
and  ( new_n28251_, new_n28249_, new_n28247_ );
xor  ( new_n28252_, new_n27990_, new_n27988_ );
xor  ( new_n28253_, new_n28252_, new_n27993_ );
xor  ( new_n28254_, new_n28193_, new_n28037_ );
xor  ( new_n28255_, new_n28254_, new_n28206_ );
xnor ( new_n28256_, new_n28222_, new_n28220_ );
xor  ( new_n28257_, new_n28256_, new_n28226_ );
nand ( new_n28258_, new_n28257_, new_n28255_ );
nor  ( new_n28259_, new_n28257_, new_n28255_ );
xnor ( new_n28260_, new_n28001_, new_n27999_ );
or   ( new_n28261_, new_n28260_, new_n28259_ );
and  ( new_n28262_, new_n28261_, new_n28258_ );
nor  ( new_n28263_, new_n28262_, new_n28253_ );
and  ( new_n28264_, new_n28262_, new_n28253_ );
xor  ( new_n28265_, new_n28137_, new_n28087_ );
xnor ( new_n28266_, new_n28265_, new_n28190_ );
xor  ( new_n28267_, new_n28023_, new_n28012_ );
xnor ( new_n28268_, new_n28267_, new_n28035_ );
or   ( new_n28269_, new_n28268_, new_n28266_ );
or   ( new_n28270_, new_n409_, new_n26196_ );
or   ( new_n28271_, new_n411_, new_n25813_ );
and  ( new_n28272_, new_n28271_, new_n28270_ );
xor  ( new_n28273_, new_n28272_, new_n328_ );
or   ( new_n28274_, new_n337_, new_n26372_ );
or   ( new_n28275_, new_n340_, new_n26063_ );
and  ( new_n28276_, new_n28275_, new_n28274_ );
xor  ( new_n28277_, new_n28276_, new_n332_ );
or   ( new_n28278_, new_n28277_, new_n28273_ );
and  ( new_n28279_, new_n28277_, new_n28273_ );
or   ( new_n28280_, new_n317_, new_n26762_ );
or   ( new_n28281_, new_n320_, new_n26620_ );
and  ( new_n28282_, new_n28281_, new_n28280_ );
xor  ( new_n28283_, new_n28282_, new_n312_ );
or   ( new_n28284_, new_n28283_, new_n28279_ );
and  ( new_n28285_, new_n28284_, new_n28278_ );
or   ( new_n28286_, new_n897_, new_n24927_ );
or   ( new_n28287_, new_n899_, new_n24543_ );
and  ( new_n28288_, new_n28287_, new_n28286_ );
xor  ( new_n28289_, new_n28288_, new_n748_ );
or   ( new_n28290_, new_n755_, new_n25048_ );
or   ( new_n28291_, new_n757_, new_n24925_ );
and  ( new_n28292_, new_n28291_, new_n28290_ );
xor  ( new_n28293_, new_n28292_, new_n523_ );
or   ( new_n28294_, new_n28293_, new_n28289_ );
and  ( new_n28295_, new_n28293_, new_n28289_ );
or   ( new_n28296_, new_n524_, new_n25486_ );
or   ( new_n28297_, new_n526_, new_n25288_ );
and  ( new_n28298_, new_n28297_, new_n28296_ );
xor  ( new_n28299_, new_n28298_, new_n403_ );
or   ( new_n28300_, new_n28299_, new_n28295_ );
and  ( new_n28301_, new_n28300_, new_n28294_ );
or   ( new_n28302_, new_n28301_, new_n28285_ );
and  ( new_n28303_, new_n28301_, new_n28285_ );
or   ( new_n28304_, new_n283_, new_n27396_ );
or   ( new_n28305_, new_n286_, new_n27085_ );
and  ( new_n28306_, new_n28305_, new_n28304_ );
xor  ( new_n28307_, new_n28306_, new_n278_ );
or   ( new_n28308_, new_n299_, new_n27763_ );
or   ( new_n28309_, new_n302_, new_n27602_ );
and  ( new_n28310_, new_n28309_, new_n28308_ );
xor  ( new_n28311_, new_n28310_, new_n293_ );
nor  ( new_n28312_, new_n28311_, new_n28307_ );
and  ( new_n28313_, new_n28311_, new_n28307_ );
not  ( new_n28314_, RIbb32dd8_180 );
or   ( new_n28315_, new_n268_, new_n28314_ );
or   ( new_n28316_, new_n271_, new_n28108_ );
and  ( new_n28317_, new_n28316_, new_n28315_ );
xor  ( new_n28318_, new_n28317_, new_n263_ );
nor  ( new_n28319_, new_n28318_, new_n28313_ );
nor  ( new_n28320_, new_n28319_, new_n28312_ );
or   ( new_n28321_, new_n28320_, new_n28303_ );
and  ( new_n28322_, new_n28321_, new_n28302_ );
or   ( new_n28323_, new_n6173_, new_n21672_ );
or   ( new_n28324_, new_n6175_, new_n21674_ );
and  ( new_n28325_, new_n28324_, new_n28323_ );
xor  ( new_n28326_, new_n28325_, new_n5597_ );
or   ( new_n28327_, new_n5604_, new_n21678_ );
or   ( new_n28328_, new_n5606_, new_n21680_ );
and  ( new_n28329_, new_n28328_, new_n28327_ );
xor  ( new_n28330_, new_n28329_, new_n5206_ );
nor  ( new_n28331_, new_n28330_, new_n28326_ );
nand ( new_n28332_, new_n28330_, new_n28326_ );
or   ( new_n28333_, new_n5207_, new_n21685_ );
or   ( new_n28334_, new_n5209_, new_n21687_ );
and  ( new_n28335_, new_n28334_, new_n28333_ );
xor  ( new_n28336_, new_n28335_, new_n4707_ );
and  ( new_n28337_, new_n28336_, new_n28332_ );
or   ( new_n28338_, new_n28337_, new_n28331_ );
or   ( new_n28339_, new_n6645_, new_n21701_ );
or   ( new_n28340_, new_n6647_, new_n21703_ );
and  ( new_n28341_, new_n28340_, new_n28339_ );
xor  ( new_n28342_, new_n28341_, new_n6166_ );
nand ( new_n28343_, new_n28342_, new_n7177_ );
or   ( new_n28344_, new_n28342_, new_n7177_ );
or   ( new_n28345_, new_n7184_, new_n21694_ );
or   ( new_n28346_, new_n7186_, new_n21696_ );
and  ( new_n28347_, new_n28346_, new_n28345_ );
xor  ( new_n28348_, new_n28347_, new_n6638_ );
nand ( new_n28349_, new_n28348_, new_n28344_ );
and  ( new_n28350_, new_n28349_, new_n28343_ );
nand ( new_n28351_, new_n28350_, new_n28338_ );
nor  ( new_n28352_, new_n28350_, new_n28338_ );
or   ( new_n28353_, new_n4709_, new_n21792_ );
or   ( new_n28354_, new_n4711_, new_n21751_ );
and  ( new_n28355_, new_n28354_, new_n28353_ );
xor  ( new_n28356_, new_n28355_, new_n4295_ );
or   ( new_n28357_, new_n4302_, new_n21840_ );
or   ( new_n28358_, new_n4304_, new_n21842_ );
and  ( new_n28359_, new_n28358_, new_n28357_ );
xor  ( new_n28360_, new_n28359_, new_n3895_ );
nor  ( new_n28361_, new_n28360_, new_n28356_ );
and  ( new_n28362_, new_n28360_, new_n28356_ );
or   ( new_n28363_, new_n3896_, new_n22098_ );
or   ( new_n28364_, new_n3898_, new_n21847_ );
and  ( new_n28365_, new_n28364_, new_n28363_ );
xor  ( new_n28366_, new_n28365_, new_n3460_ );
nor  ( new_n28367_, new_n28366_, new_n28362_ );
nor  ( new_n28368_, new_n28367_, new_n28361_ );
or   ( new_n28369_, new_n28368_, new_n28352_ );
and  ( new_n28370_, new_n28369_, new_n28351_ );
nor  ( new_n28371_, new_n28370_, new_n28322_ );
nand ( new_n28372_, new_n28370_, new_n28322_ );
or   ( new_n28373_, new_n3461_, new_n22207_ );
or   ( new_n28374_, new_n3463_, new_n22129_ );
and  ( new_n28375_, new_n28374_, new_n28373_ );
xor  ( new_n28376_, new_n28375_, new_n3116_ );
or   ( new_n28377_, new_n3117_, new_n22423_ );
or   ( new_n28378_, new_n3119_, new_n22304_ );
and  ( new_n28379_, new_n28378_, new_n28377_ );
xor  ( new_n28380_, new_n28379_, new_n2800_ );
or   ( new_n28381_, new_n28380_, new_n28376_ );
and  ( new_n28382_, new_n28380_, new_n28376_ );
or   ( new_n28383_, new_n2807_, new_n22641_ );
or   ( new_n28384_, new_n2809_, new_n22590_ );
and  ( new_n28385_, new_n28384_, new_n28383_ );
xor  ( new_n28386_, new_n28385_, new_n2424_ );
or   ( new_n28387_, new_n28386_, new_n28382_ );
and  ( new_n28388_, new_n28387_, new_n28381_ );
or   ( new_n28389_, new_n2425_, new_n22975_ );
or   ( new_n28390_, new_n2427_, new_n22829_ );
and  ( new_n28391_, new_n28390_, new_n28389_ );
xor  ( new_n28392_, new_n28391_, new_n2121_ );
or   ( new_n28393_, new_n2122_, new_n23166_ );
or   ( new_n28394_, new_n2124_, new_n22973_ );
and  ( new_n28395_, new_n28394_, new_n28393_ );
xor  ( new_n28396_, new_n28395_, new_n1843_ );
or   ( new_n28397_, new_n28396_, new_n28392_ );
and  ( new_n28398_, new_n28396_, new_n28392_ );
or   ( new_n28399_, new_n1844_, new_n23370_ );
or   ( new_n28400_, new_n1846_, new_n23252_ );
and  ( new_n28401_, new_n28400_, new_n28399_ );
xor  ( new_n28402_, new_n28401_, new_n1586_ );
or   ( new_n28403_, new_n28402_, new_n28398_ );
and  ( new_n28404_, new_n28403_, new_n28397_ );
nor  ( new_n28405_, new_n28404_, new_n28388_ );
nand ( new_n28406_, new_n28404_, new_n28388_ );
or   ( new_n28407_, new_n1593_, new_n23733_ );
or   ( new_n28408_, new_n1595_, new_n23554_ );
and  ( new_n28409_, new_n28408_, new_n28407_ );
xor  ( new_n28410_, new_n28409_, new_n1358_ );
or   ( new_n28411_, new_n1364_, new_n24006_ );
or   ( new_n28412_, new_n1366_, new_n23895_ );
and  ( new_n28413_, new_n28412_, new_n28411_ );
xor  ( new_n28414_, new_n28413_, new_n1129_ );
nor  ( new_n28415_, new_n28414_, new_n28410_ );
and  ( new_n28416_, new_n28414_, new_n28410_ );
or   ( new_n28417_, new_n1135_, new_n24418_ );
or   ( new_n28418_, new_n1137_, new_n24227_ );
and  ( new_n28419_, new_n28418_, new_n28417_ );
xor  ( new_n28420_, new_n28419_, new_n896_ );
nor  ( new_n28421_, new_n28420_, new_n28416_ );
or   ( new_n28422_, new_n28421_, new_n28415_ );
and  ( new_n28423_, new_n28422_, new_n28406_ );
or   ( new_n28424_, new_n28423_, new_n28405_ );
and  ( new_n28425_, new_n28424_, new_n28372_ );
or   ( new_n28426_, new_n28425_, new_n28371_ );
xor  ( new_n28427_, new_n28029_, new_n28027_ );
xor  ( new_n28428_, new_n28427_, new_n28033_ );
xnor ( new_n28429_, new_n28006_, new_n28004_ );
xor  ( new_n28430_, new_n28429_, new_n28010_ );
nand ( new_n28431_, new_n28430_, new_n28428_ );
nor  ( new_n28432_, new_n28430_, new_n28428_ );
xor  ( new_n28433_, new_n28016_, new_n28014_ );
xor  ( new_n28434_, new_n28433_, new_n28021_ );
or   ( new_n28435_, new_n28434_, new_n28432_ );
and  ( new_n28436_, new_n28435_, new_n28431_ );
or   ( new_n28437_, new_n28436_, new_n28426_ );
and  ( new_n28438_, new_n28436_, new_n28426_ );
xor  ( new_n28439_, new_n28112_, new_n28107_ );
xnor ( new_n28440_, new_n28439_, new_n28114_ );
xnor ( new_n28441_, new_n28125_, new_n28121_ );
xor  ( new_n28442_, new_n28441_, new_n28131_ );
and  ( new_n28443_, new_n28442_, new_n28440_ );
xnor ( new_n28444_, new_n28146_, new_n28142_ );
xor  ( new_n28445_, new_n28444_, new_n28152_ );
xnor ( new_n28446_, new_n28095_, new_n28091_ );
xor  ( new_n28447_, new_n28446_, new_n28101_ );
or   ( new_n28448_, new_n28447_, new_n28445_ );
and  ( new_n28449_, new_n28447_, new_n28445_ );
xor  ( new_n28450_, new_n28180_, new_n28176_ );
xnor ( new_n28451_, new_n28450_, new_n28186_ );
or   ( new_n28452_, new_n28451_, new_n28449_ );
and  ( new_n28453_, new_n28452_, new_n28448_ );
or   ( new_n28454_, new_n28453_, new_n28443_ );
and  ( new_n28455_, new_n28453_, new_n28443_ );
xnor ( new_n28456_, new_n28061_, new_n28057_ );
xor  ( new_n28457_, new_n28456_, new_n28067_ );
xnor ( new_n28458_, new_n28162_, new_n28158_ );
xor  ( new_n28459_, new_n28458_, new_n28168_ );
nor  ( new_n28460_, new_n28459_, new_n28457_ );
and  ( new_n28461_, new_n28459_, new_n28457_ );
xor  ( new_n28462_, new_n28045_, new_n28041_ );
xnor ( new_n28463_, new_n28462_, new_n28051_ );
nor  ( new_n28464_, new_n28463_, new_n28461_ );
nor  ( new_n28465_, new_n28464_, new_n28460_ );
or   ( new_n28466_, new_n28465_, new_n28455_ );
and  ( new_n28467_, new_n28466_, new_n28454_ );
or   ( new_n28468_, new_n28467_, new_n28438_ );
and  ( new_n28469_, new_n28468_, new_n28437_ );
nor  ( new_n28470_, new_n28469_, new_n28269_ );
and  ( new_n28471_, new_n28469_, new_n28269_ );
xnor ( new_n28472_, new_n28133_, new_n28117_ );
xor  ( new_n28473_, new_n28472_, new_n28103_ );
xnor ( new_n28474_, new_n28069_, new_n28053_ );
xor  ( new_n28475_, new_n28474_, new_n28085_ );
nor  ( new_n28476_, new_n28475_, new_n28473_ );
nand ( new_n28477_, new_n28475_, new_n28473_ );
xor  ( new_n28478_, new_n28170_, new_n28154_ );
xor  ( new_n28479_, new_n28478_, new_n28188_ );
and  ( new_n28480_, new_n28479_, new_n28477_ );
or   ( new_n28481_, new_n28480_, new_n28476_ );
xor  ( new_n28482_, new_n28214_, new_n28212_ );
xor  ( new_n28483_, new_n28482_, new_n28218_ );
and  ( new_n28484_, new_n28483_, new_n28481_ );
nor  ( new_n28485_, new_n28483_, new_n28481_ );
xor  ( new_n28486_, new_n28199_, new_n28197_ );
xor  ( new_n28487_, new_n28486_, new_n28204_ );
not  ( new_n28488_, new_n28487_ );
nor  ( new_n28489_, new_n28488_, new_n28485_ );
nor  ( new_n28490_, new_n28489_, new_n28484_ );
nor  ( new_n28491_, new_n28490_, new_n28471_ );
nor  ( new_n28492_, new_n28491_, new_n28470_ );
nor  ( new_n28493_, new_n28492_, new_n28264_ );
nor  ( new_n28494_, new_n28493_, new_n28263_ );
or   ( new_n28495_, new_n28494_, new_n28251_ );
and  ( new_n28496_, new_n28495_, new_n28250_ );
xor  ( new_n28497_, new_n28234_, new_n28232_ );
xor  ( new_n28498_, new_n28497_, new_n28238_ );
nor  ( new_n28499_, new_n28498_, new_n28496_ );
xor  ( new_n28500_, new_n28242_, new_n28240_ );
and  ( new_n28501_, new_n28500_, new_n28499_ );
xor  ( new_n28502_, new_n28257_, new_n28255_ );
xor  ( new_n28503_, new_n28502_, new_n28260_ );
xor  ( new_n28504_, new_n28436_, new_n28426_ );
xor  ( new_n28505_, new_n28504_, new_n28467_ );
xor  ( new_n28506_, new_n28483_, new_n28481_ );
xor  ( new_n28507_, new_n28506_, new_n28488_ );
or   ( new_n28508_, new_n28507_, new_n28505_ );
and  ( new_n28509_, new_n28507_, new_n28505_ );
xnor ( new_n28510_, new_n28268_, new_n28266_ );
or   ( new_n28511_, new_n28510_, new_n28509_ );
and  ( new_n28512_, new_n28511_, new_n28508_ );
nor  ( new_n28513_, new_n28512_, new_n28503_ );
and  ( new_n28514_, new_n28512_, new_n28503_ );
xor  ( new_n28515_, new_n28453_, new_n28443_ );
xnor ( new_n28516_, new_n28515_, new_n28465_ );
xor  ( new_n28517_, new_n28370_, new_n28322_ );
xnor ( new_n28518_, new_n28517_, new_n28424_ );
and  ( new_n28519_, new_n28518_, new_n28516_ );
xor  ( new_n28520_, new_n28330_, new_n28326_ );
xor  ( new_n28521_, new_n28520_, new_n28336_ );
xnor ( new_n28522_, new_n28380_, new_n28376_ );
xor  ( new_n28523_, new_n28522_, new_n28386_ );
nor  ( new_n28524_, new_n28523_, new_n28521_ );
nand ( new_n28525_, new_n28523_, new_n28521_ );
xor  ( new_n28526_, new_n28360_, new_n28356_ );
xnor ( new_n28527_, new_n28526_, new_n28366_ );
not  ( new_n28528_, new_n28527_ );
and  ( new_n28529_, new_n28528_, new_n28525_ );
or   ( new_n28530_, new_n28529_, new_n28524_ );
not  ( new_n28531_, RIbb32e50_181 );
or   ( new_n28532_, new_n28531_, new_n260_ );
xnor ( new_n28533_, new_n28277_, new_n28273_ );
xor  ( new_n28534_, new_n28533_, new_n28283_ );
nand ( new_n28535_, new_n28534_, new_n28532_ );
or   ( new_n28536_, new_n28534_, new_n28532_ );
xor  ( new_n28537_, new_n28311_, new_n28307_ );
xnor ( new_n28538_, new_n28537_, new_n28318_ );
nand ( new_n28539_, new_n28538_, new_n28536_ );
and  ( new_n28540_, new_n28539_, new_n28535_ );
and  ( new_n28541_, new_n28540_, new_n28530_ );
or   ( new_n28542_, new_n28540_, new_n28530_ );
xnor ( new_n28543_, new_n28293_, new_n28289_ );
xor  ( new_n28544_, new_n28543_, new_n28299_ );
xnor ( new_n28545_, new_n28396_, new_n28392_ );
xor  ( new_n28546_, new_n28545_, new_n28402_ );
nor  ( new_n28547_, new_n28546_, new_n28544_ );
nand ( new_n28548_, new_n28546_, new_n28544_ );
xor  ( new_n28549_, new_n28414_, new_n28410_ );
xor  ( new_n28550_, new_n28549_, new_n28420_ );
and  ( new_n28551_, new_n28550_, new_n28548_ );
or   ( new_n28552_, new_n28551_, new_n28547_ );
and  ( new_n28553_, new_n28552_, new_n28542_ );
or   ( new_n28554_, new_n28553_, new_n28541_ );
or   ( new_n28555_, new_n283_, new_n27602_ );
or   ( new_n28556_, new_n286_, new_n27396_ );
and  ( new_n28557_, new_n28556_, new_n28555_ );
xor  ( new_n28558_, new_n28557_, new_n278_ );
or   ( new_n28559_, new_n299_, new_n28108_ );
or   ( new_n28560_, new_n302_, new_n27763_ );
and  ( new_n28561_, new_n28560_, new_n28559_ );
xor  ( new_n28562_, new_n28561_, new_n293_ );
or   ( new_n28563_, new_n28562_, new_n28558_ );
and  ( new_n28564_, new_n28562_, new_n28558_ );
or   ( new_n28565_, new_n268_, new_n28531_ );
or   ( new_n28566_, new_n271_, new_n28314_ );
and  ( new_n28567_, new_n28566_, new_n28565_ );
xor  ( new_n28568_, new_n28567_, new_n263_ );
or   ( new_n28569_, new_n28568_, new_n28564_ );
and  ( new_n28570_, new_n28569_, new_n28563_ );
or   ( new_n28571_, new_n897_, new_n24925_ );
or   ( new_n28572_, new_n899_, new_n24927_ );
and  ( new_n28573_, new_n28572_, new_n28571_ );
xor  ( new_n28574_, new_n28573_, new_n748_ );
or   ( new_n28575_, new_n755_, new_n25288_ );
or   ( new_n28576_, new_n757_, new_n25048_ );
and  ( new_n28577_, new_n28576_, new_n28575_ );
xor  ( new_n28578_, new_n28577_, new_n523_ );
or   ( new_n28579_, new_n28578_, new_n28574_ );
and  ( new_n28580_, new_n28578_, new_n28574_ );
or   ( new_n28581_, new_n524_, new_n25813_ );
or   ( new_n28582_, new_n526_, new_n25486_ );
and  ( new_n28583_, new_n28582_, new_n28581_ );
xor  ( new_n28584_, new_n28583_, new_n403_ );
or   ( new_n28585_, new_n28584_, new_n28580_ );
and  ( new_n28586_, new_n28585_, new_n28579_ );
or   ( new_n28587_, new_n28586_, new_n28570_ );
and  ( new_n28588_, new_n28586_, new_n28570_ );
or   ( new_n28589_, new_n409_, new_n26063_ );
or   ( new_n28590_, new_n411_, new_n26196_ );
and  ( new_n28591_, new_n28590_, new_n28589_ );
xor  ( new_n28592_, new_n28591_, new_n328_ );
or   ( new_n28593_, new_n337_, new_n26620_ );
or   ( new_n28594_, new_n340_, new_n26372_ );
and  ( new_n28595_, new_n28594_, new_n28593_ );
xor  ( new_n28596_, new_n28595_, new_n332_ );
nor  ( new_n28597_, new_n28596_, new_n28592_ );
and  ( new_n28598_, new_n28596_, new_n28592_ );
or   ( new_n28599_, new_n317_, new_n27085_ );
or   ( new_n28600_, new_n320_, new_n26762_ );
and  ( new_n28601_, new_n28600_, new_n28599_ );
xor  ( new_n28602_, new_n28601_, new_n312_ );
nor  ( new_n28603_, new_n28602_, new_n28598_ );
nor  ( new_n28604_, new_n28603_, new_n28597_ );
or   ( new_n28605_, new_n28604_, new_n28588_ );
and  ( new_n28606_, new_n28605_, new_n28587_ );
or   ( new_n28607_, new_n4709_, new_n21842_ );
or   ( new_n28608_, new_n4711_, new_n21792_ );
and  ( new_n28609_, new_n28608_, new_n28607_ );
xor  ( new_n28610_, new_n28609_, new_n4295_ );
or   ( new_n28611_, new_n4302_, new_n21847_ );
or   ( new_n28612_, new_n4304_, new_n21840_ );
and  ( new_n28613_, new_n28612_, new_n28611_ );
xor  ( new_n28614_, new_n28613_, new_n3895_ );
or   ( new_n28615_, new_n28614_, new_n28610_ );
and  ( new_n28616_, new_n28614_, new_n28610_ );
or   ( new_n28617_, new_n3896_, new_n22129_ );
or   ( new_n28618_, new_n3898_, new_n22098_ );
and  ( new_n28619_, new_n28618_, new_n28617_ );
xor  ( new_n28620_, new_n28619_, new_n3460_ );
or   ( new_n28621_, new_n28620_, new_n28616_ );
and  ( new_n28622_, new_n28621_, new_n28615_ );
or   ( new_n28623_, new_n6173_, new_n21680_ );
or   ( new_n28624_, new_n6175_, new_n21672_ );
and  ( new_n28625_, new_n28624_, new_n28623_ );
xor  ( new_n28626_, new_n28625_, new_n5597_ );
or   ( new_n28627_, new_n5604_, new_n21687_ );
or   ( new_n28628_, new_n5606_, new_n21678_ );
and  ( new_n28629_, new_n28628_, new_n28627_ );
xor  ( new_n28630_, new_n28629_, new_n5206_ );
or   ( new_n28631_, new_n28630_, new_n28626_ );
and  ( new_n28632_, new_n28630_, new_n28626_ );
or   ( new_n28633_, new_n5207_, new_n21751_ );
or   ( new_n28634_, new_n5209_, new_n21685_ );
and  ( new_n28635_, new_n28634_, new_n28633_ );
xor  ( new_n28636_, new_n28635_, new_n4708_ );
or   ( new_n28637_, new_n28636_, new_n28632_ );
and  ( new_n28638_, new_n28637_, new_n28631_ );
or   ( new_n28639_, new_n28638_, new_n28622_ );
and  ( new_n28640_, new_n28638_, new_n28622_ );
or   ( new_n28641_, new_n7184_, new_n21703_ );
or   ( new_n28642_, new_n7186_, new_n21694_ );
and  ( new_n28643_, new_n28642_, new_n28641_ );
xor  ( new_n28644_, new_n28643_, new_n6637_ );
and  ( new_n28645_, new_n7489_, RIbb315f0_129 );
xor  ( new_n28646_, new_n28645_, new_n7177_ );
and  ( new_n28647_, new_n28646_, new_n28644_ );
nor  ( new_n28648_, new_n28646_, new_n28644_ );
or   ( new_n28649_, new_n6645_, new_n21674_ );
or   ( new_n28650_, new_n6647_, new_n21701_ );
and  ( new_n28651_, new_n28650_, new_n28649_ );
xor  ( new_n28652_, new_n28651_, new_n6166_ );
nor  ( new_n28653_, new_n28652_, new_n28648_ );
nor  ( new_n28654_, new_n28653_, new_n28647_ );
or   ( new_n28655_, new_n28654_, new_n28640_ );
and  ( new_n28656_, new_n28655_, new_n28639_ );
or   ( new_n28657_, new_n28656_, new_n28606_ );
or   ( new_n28658_, new_n3461_, new_n22304_ );
or   ( new_n28659_, new_n3463_, new_n22207_ );
and  ( new_n28660_, new_n28659_, new_n28658_ );
xor  ( new_n28661_, new_n28660_, new_n3116_ );
or   ( new_n28662_, new_n3117_, new_n22590_ );
or   ( new_n28663_, new_n3119_, new_n22423_ );
and  ( new_n28664_, new_n28663_, new_n28662_ );
xor  ( new_n28665_, new_n28664_, new_n2800_ );
or   ( new_n28666_, new_n28665_, new_n28661_ );
and  ( new_n28667_, new_n28665_, new_n28661_ );
or   ( new_n28668_, new_n2807_, new_n22829_ );
or   ( new_n28669_, new_n2809_, new_n22641_ );
and  ( new_n28670_, new_n28669_, new_n28668_ );
xor  ( new_n28671_, new_n28670_, new_n2424_ );
or   ( new_n28672_, new_n28671_, new_n28667_ );
and  ( new_n28673_, new_n28672_, new_n28666_ );
or   ( new_n28674_, new_n1593_, new_n23895_ );
or   ( new_n28675_, new_n1595_, new_n23733_ );
and  ( new_n28676_, new_n28675_, new_n28674_ );
xor  ( new_n28677_, new_n28676_, new_n1358_ );
or   ( new_n28678_, new_n1364_, new_n24227_ );
or   ( new_n28679_, new_n1366_, new_n24006_ );
and  ( new_n28680_, new_n28679_, new_n28678_ );
xor  ( new_n28681_, new_n28680_, new_n1129_ );
or   ( new_n28682_, new_n28681_, new_n28677_ );
and  ( new_n28683_, new_n28681_, new_n28677_ );
or   ( new_n28684_, new_n1135_, new_n24543_ );
or   ( new_n28685_, new_n1137_, new_n24418_ );
and  ( new_n28686_, new_n28685_, new_n28684_ );
xor  ( new_n28687_, new_n28686_, new_n896_ );
or   ( new_n28688_, new_n28687_, new_n28683_ );
and  ( new_n28689_, new_n28688_, new_n28682_ );
or   ( new_n28690_, new_n28689_, new_n28673_ );
and  ( new_n28691_, new_n28689_, new_n28673_ );
or   ( new_n28692_, new_n2425_, new_n22973_ );
or   ( new_n28693_, new_n2427_, new_n22975_ );
and  ( new_n28694_, new_n28693_, new_n28692_ );
xor  ( new_n28695_, new_n28694_, new_n2121_ );
or   ( new_n28696_, new_n2122_, new_n23252_ );
or   ( new_n28697_, new_n2124_, new_n23166_ );
and  ( new_n28698_, new_n28697_, new_n28696_ );
xor  ( new_n28699_, new_n28698_, new_n1843_ );
nor  ( new_n28700_, new_n28699_, new_n28695_ );
and  ( new_n28701_, new_n28699_, new_n28695_ );
or   ( new_n28702_, new_n1844_, new_n23554_ );
or   ( new_n28703_, new_n1846_, new_n23370_ );
and  ( new_n28704_, new_n28703_, new_n28702_ );
xor  ( new_n28705_, new_n28704_, new_n1586_ );
nor  ( new_n28706_, new_n28705_, new_n28701_ );
nor  ( new_n28707_, new_n28706_, new_n28700_ );
or   ( new_n28708_, new_n28707_, new_n28691_ );
and  ( new_n28709_, new_n28708_, new_n28690_ );
and  ( new_n28710_, new_n28656_, new_n28606_ );
or   ( new_n28711_, new_n28710_, new_n28709_ );
and  ( new_n28712_, new_n28711_, new_n28657_ );
or   ( new_n28713_, new_n28712_, new_n28554_ );
and  ( new_n28714_, new_n28712_, new_n28554_ );
xor  ( new_n28715_, new_n28077_, new_n28075_ );
xor  ( new_n28716_, new_n28715_, new_n28083_ );
xnor ( new_n28717_, new_n28459_, new_n28457_ );
xor  ( new_n28718_, new_n28717_, new_n28463_ );
and  ( new_n28719_, new_n28718_, new_n28716_ );
or   ( new_n28720_, new_n28718_, new_n28716_ );
xor  ( new_n28721_, new_n28447_, new_n28445_ );
xnor ( new_n28722_, new_n28721_, new_n28451_ );
and  ( new_n28723_, new_n28722_, new_n28720_ );
or   ( new_n28724_, new_n28723_, new_n28719_ );
or   ( new_n28725_, new_n28724_, new_n28714_ );
and  ( new_n28726_, new_n28725_, new_n28713_ );
and  ( new_n28727_, new_n28726_, new_n28519_ );
nor  ( new_n28728_, new_n28726_, new_n28519_ );
xnor ( new_n28729_, new_n28430_, new_n28428_ );
xor  ( new_n28730_, new_n28729_, new_n28434_ );
xor  ( new_n28731_, new_n28475_, new_n28473_ );
xor  ( new_n28732_, new_n28731_, new_n28479_ );
and  ( new_n28733_, new_n28732_, new_n28730_ );
nor  ( new_n28734_, new_n28732_, new_n28730_ );
xor  ( new_n28735_, new_n28404_, new_n28388_ );
xor  ( new_n28736_, new_n28735_, new_n28422_ );
xnor ( new_n28737_, new_n28301_, new_n28285_ );
xor  ( new_n28738_, new_n28737_, new_n28320_ );
nor  ( new_n28739_, new_n28738_, new_n28736_ );
and  ( new_n28740_, new_n28738_, new_n28736_ );
xor  ( new_n28741_, new_n28442_, new_n28440_ );
nor  ( new_n28742_, new_n28741_, new_n28740_ );
nor  ( new_n28743_, new_n28742_, new_n28739_ );
nor  ( new_n28744_, new_n28743_, new_n28734_ );
nor  ( new_n28745_, new_n28744_, new_n28733_ );
nor  ( new_n28746_, new_n28745_, new_n28728_ );
nor  ( new_n28747_, new_n28746_, new_n28727_ );
nor  ( new_n28748_, new_n28747_, new_n28514_ );
or   ( new_n28749_, new_n28748_, new_n28513_ );
xnor ( new_n28750_, new_n28208_, new_n28002_ );
xor  ( new_n28751_, new_n28750_, new_n28228_ );
or   ( new_n28752_, new_n28751_, new_n28749_ );
and  ( new_n28753_, new_n28751_, new_n28749_ );
xor  ( new_n28754_, new_n28262_, new_n28253_ );
xnor ( new_n28755_, new_n28754_, new_n28492_ );
or   ( new_n28756_, new_n28755_, new_n28753_ );
and  ( new_n28757_, new_n28756_, new_n28752_ );
xnor ( new_n28758_, new_n28249_, new_n28247_ );
xor  ( new_n28759_, new_n28758_, new_n28494_ );
and  ( new_n28760_, new_n28759_, new_n28757_ );
xor  ( new_n28761_, new_n28498_, new_n28496_ );
and  ( new_n28762_, new_n28761_, new_n28760_ );
xnor ( new_n28763_, new_n28469_, new_n28269_ );
xor  ( new_n28764_, new_n28763_, new_n28490_ );
xor  ( new_n28765_, new_n28507_, new_n28505_ );
xor  ( new_n28766_, new_n28765_, new_n28510_ );
xor  ( new_n28767_, new_n28712_, new_n28554_ );
xor  ( new_n28768_, new_n28767_, new_n28724_ );
xnor ( new_n28769_, new_n28732_, new_n28730_ );
xor  ( new_n28770_, new_n28769_, new_n28743_ );
nand ( new_n28771_, new_n28770_, new_n28768_ );
nor  ( new_n28772_, new_n28770_, new_n28768_ );
xnor ( new_n28773_, new_n28518_, new_n28516_ );
or   ( new_n28774_, new_n28773_, new_n28772_ );
and  ( new_n28775_, new_n28774_, new_n28771_ );
nand ( new_n28776_, new_n28775_, new_n28766_ );
or   ( new_n28777_, new_n28775_, new_n28766_ );
xor  ( new_n28778_, new_n28656_, new_n28606_ );
xor  ( new_n28779_, new_n28778_, new_n28709_ );
xor  ( new_n28780_, new_n28540_, new_n28530_ );
xor  ( new_n28781_, new_n28780_, new_n28552_ );
nand ( new_n28782_, new_n28781_, new_n28779_ );
nor  ( new_n28783_, new_n28781_, new_n28779_ );
xor  ( new_n28784_, new_n28718_, new_n28716_ );
xnor ( new_n28785_, new_n28784_, new_n28722_ );
or   ( new_n28786_, new_n28785_, new_n28783_ );
and  ( new_n28787_, new_n28786_, new_n28782_ );
xnor ( new_n28788_, new_n28350_, new_n28338_ );
xor  ( new_n28789_, new_n28788_, new_n28368_ );
xnor ( new_n28790_, new_n28586_, new_n28570_ );
xor  ( new_n28791_, new_n28790_, new_n28604_ );
xnor ( new_n28792_, new_n28689_, new_n28673_ );
xor  ( new_n28793_, new_n28792_, new_n28707_ );
or   ( new_n28794_, new_n28793_, new_n28791_ );
and  ( new_n28795_, new_n28793_, new_n28791_ );
xor  ( new_n28796_, new_n28534_, new_n28532_ );
xor  ( new_n28797_, new_n28796_, new_n28538_ );
or   ( new_n28798_, new_n28797_, new_n28795_ );
and  ( new_n28799_, new_n28798_, new_n28794_ );
or   ( new_n28800_, new_n28799_, new_n28789_ );
and  ( new_n28801_, new_n28799_, new_n28789_ );
xor  ( new_n28802_, new_n28738_, new_n28736_ );
xor  ( new_n28803_, new_n28802_, new_n28741_ );
or   ( new_n28804_, new_n28803_, new_n28801_ );
and  ( new_n28805_, new_n28804_, new_n28800_ );
nor  ( new_n28806_, new_n28805_, new_n28787_ );
and  ( new_n28807_, new_n28805_, new_n28787_ );
or   ( new_n28808_, new_n317_, new_n27396_ );
or   ( new_n28809_, new_n320_, new_n27085_ );
and  ( new_n28810_, new_n28809_, new_n28808_ );
xor  ( new_n28811_, new_n28810_, new_n312_ );
or   ( new_n28812_, new_n283_, new_n27763_ );
or   ( new_n28813_, new_n286_, new_n27602_ );
and  ( new_n28814_, new_n28813_, new_n28812_ );
xor  ( new_n28815_, new_n28814_, new_n278_ );
or   ( new_n28816_, new_n28815_, new_n28811_ );
and  ( new_n28817_, new_n28815_, new_n28811_ );
or   ( new_n28818_, new_n299_, new_n28314_ );
or   ( new_n28819_, new_n302_, new_n28108_ );
and  ( new_n28820_, new_n28819_, new_n28818_ );
xor  ( new_n28821_, new_n28820_, new_n293_ );
or   ( new_n28822_, new_n28821_, new_n28817_ );
and  ( new_n28823_, new_n28822_, new_n28816_ );
or   ( new_n28824_, new_n524_, new_n26196_ );
or   ( new_n28825_, new_n526_, new_n25813_ );
and  ( new_n28826_, new_n28825_, new_n28824_ );
xor  ( new_n28827_, new_n28826_, new_n403_ );
or   ( new_n28828_, new_n409_, new_n26372_ );
or   ( new_n28829_, new_n411_, new_n26063_ );
and  ( new_n28830_, new_n28829_, new_n28828_ );
xor  ( new_n28831_, new_n28830_, new_n328_ );
or   ( new_n28832_, new_n28831_, new_n28827_ );
and  ( new_n28833_, new_n28831_, new_n28827_ );
or   ( new_n28834_, new_n337_, new_n26762_ );
or   ( new_n28835_, new_n340_, new_n26620_ );
and  ( new_n28836_, new_n28835_, new_n28834_ );
xor  ( new_n28837_, new_n28836_, new_n332_ );
or   ( new_n28838_, new_n28837_, new_n28833_ );
and  ( new_n28839_, new_n28838_, new_n28832_ );
or   ( new_n28840_, new_n28839_, new_n28823_ );
and  ( new_n28841_, new_n28839_, new_n28823_ );
or   ( new_n28842_, new_n1135_, new_n24927_ );
or   ( new_n28843_, new_n1137_, new_n24543_ );
and  ( new_n28844_, new_n28843_, new_n28842_ );
xor  ( new_n28845_, new_n28844_, new_n896_ );
or   ( new_n28846_, new_n897_, new_n25048_ );
or   ( new_n28847_, new_n899_, new_n24925_ );
and  ( new_n28848_, new_n28847_, new_n28846_ );
xor  ( new_n28849_, new_n28848_, new_n748_ );
nor  ( new_n28850_, new_n28849_, new_n28845_ );
and  ( new_n28851_, new_n28849_, new_n28845_ );
or   ( new_n28852_, new_n755_, new_n25486_ );
or   ( new_n28853_, new_n757_, new_n25288_ );
and  ( new_n28854_, new_n28853_, new_n28852_ );
xor  ( new_n28855_, new_n28854_, new_n523_ );
nor  ( new_n28856_, new_n28855_, new_n28851_ );
nor  ( new_n28857_, new_n28856_, new_n28850_ );
or   ( new_n28858_, new_n28857_, new_n28841_ );
and  ( new_n28859_, new_n28858_, new_n28840_ );
or   ( new_n28860_, new_n5207_, new_n21792_ );
or   ( new_n28861_, new_n5209_, new_n21751_ );
and  ( new_n28862_, new_n28861_, new_n28860_ );
xor  ( new_n28863_, new_n28862_, new_n4708_ );
or   ( new_n28864_, new_n4709_, new_n21840_ );
or   ( new_n28865_, new_n4711_, new_n21842_ );
and  ( new_n28866_, new_n28865_, new_n28864_ );
xor  ( new_n28867_, new_n28866_, new_n4295_ );
nor  ( new_n28868_, new_n28867_, new_n28863_ );
nand ( new_n28869_, new_n28867_, new_n28863_ );
or   ( new_n28870_, new_n4302_, new_n22098_ );
or   ( new_n28871_, new_n4304_, new_n21847_ );
and  ( new_n28872_, new_n28871_, new_n28870_ );
xor  ( new_n28873_, new_n28872_, new_n3895_ );
not  ( new_n28874_, new_n28873_ );
and  ( new_n28875_, new_n28874_, new_n28869_ );
or   ( new_n28876_, new_n28875_, new_n28868_ );
or   ( new_n28877_, new_n7184_, new_n21701_ );
or   ( new_n28878_, new_n7186_, new_n21703_ );
and  ( new_n28879_, new_n28878_, new_n28877_ );
xor  ( new_n28880_, new_n28879_, new_n6638_ );
nand ( new_n28881_, new_n28880_, new_n7725_ );
or   ( new_n28882_, new_n28880_, new_n7725_ );
or   ( new_n28883_, new_n7732_, new_n21694_ );
or   ( new_n28884_, new_n7734_, new_n21696_ );
and  ( new_n28885_, new_n28884_, new_n28883_ );
xor  ( new_n28886_, new_n28885_, new_n7177_ );
nand ( new_n28887_, new_n28886_, new_n28882_ );
and  ( new_n28888_, new_n28887_, new_n28881_ );
nand ( new_n28889_, new_n28888_, new_n28876_ );
nor  ( new_n28890_, new_n28888_, new_n28876_ );
or   ( new_n28891_, new_n6645_, new_n21672_ );
or   ( new_n28892_, new_n6647_, new_n21674_ );
and  ( new_n28893_, new_n28892_, new_n28891_ );
xor  ( new_n28894_, new_n28893_, new_n6166_ );
or   ( new_n28895_, new_n6173_, new_n21678_ );
or   ( new_n28896_, new_n6175_, new_n21680_ );
and  ( new_n28897_, new_n28896_, new_n28895_ );
xor  ( new_n28898_, new_n28897_, new_n5597_ );
nor  ( new_n28899_, new_n28898_, new_n28894_ );
and  ( new_n28900_, new_n28898_, new_n28894_ );
or   ( new_n28901_, new_n5604_, new_n21685_ );
or   ( new_n28902_, new_n5606_, new_n21687_ );
and  ( new_n28903_, new_n28902_, new_n28901_ );
xor  ( new_n28904_, new_n28903_, new_n5206_ );
nor  ( new_n28905_, new_n28904_, new_n28900_ );
nor  ( new_n28906_, new_n28905_, new_n28899_ );
or   ( new_n28907_, new_n28906_, new_n28890_ );
and  ( new_n28908_, new_n28907_, new_n28889_ );
or   ( new_n28909_, new_n28908_, new_n28859_ );
and  ( new_n28910_, new_n28908_, new_n28859_ );
or   ( new_n28911_, new_n3896_, new_n22207_ );
or   ( new_n28912_, new_n3898_, new_n22129_ );
and  ( new_n28913_, new_n28912_, new_n28911_ );
xor  ( new_n28914_, new_n28913_, new_n3460_ );
or   ( new_n28915_, new_n3461_, new_n22423_ );
or   ( new_n28916_, new_n3463_, new_n22304_ );
and  ( new_n28917_, new_n28916_, new_n28915_ );
xor  ( new_n28918_, new_n28917_, new_n3116_ );
or   ( new_n28919_, new_n28918_, new_n28914_ );
and  ( new_n28920_, new_n28918_, new_n28914_ );
or   ( new_n28921_, new_n3117_, new_n22641_ );
or   ( new_n28922_, new_n3119_, new_n22590_ );
and  ( new_n28923_, new_n28922_, new_n28921_ );
xor  ( new_n28924_, new_n28923_, new_n2800_ );
or   ( new_n28925_, new_n28924_, new_n28920_ );
and  ( new_n28926_, new_n28925_, new_n28919_ );
or   ( new_n28927_, new_n1844_, new_n23733_ );
or   ( new_n28928_, new_n1846_, new_n23554_ );
and  ( new_n28929_, new_n28928_, new_n28927_ );
xor  ( new_n28930_, new_n28929_, new_n1586_ );
or   ( new_n28931_, new_n1593_, new_n24006_ );
or   ( new_n28932_, new_n1595_, new_n23895_ );
and  ( new_n28933_, new_n28932_, new_n28931_ );
xor  ( new_n28934_, new_n28933_, new_n1358_ );
or   ( new_n28935_, new_n28934_, new_n28930_ );
and  ( new_n28936_, new_n28934_, new_n28930_ );
or   ( new_n28937_, new_n1364_, new_n24418_ );
or   ( new_n28938_, new_n1366_, new_n24227_ );
and  ( new_n28939_, new_n28938_, new_n28937_ );
xor  ( new_n28940_, new_n28939_, new_n1129_ );
or   ( new_n28941_, new_n28940_, new_n28936_ );
and  ( new_n28942_, new_n28941_, new_n28935_ );
nor  ( new_n28943_, new_n28942_, new_n28926_ );
and  ( new_n28944_, new_n28942_, new_n28926_ );
or   ( new_n28945_, new_n2807_, new_n22975_ );
or   ( new_n28946_, new_n2809_, new_n22829_ );
and  ( new_n28947_, new_n28946_, new_n28945_ );
xor  ( new_n28948_, new_n28947_, new_n2424_ );
or   ( new_n28949_, new_n2425_, new_n23166_ );
or   ( new_n28950_, new_n2427_, new_n22973_ );
and  ( new_n28951_, new_n28950_, new_n28949_ );
xor  ( new_n28952_, new_n28951_, new_n2121_ );
nor  ( new_n28953_, new_n28952_, new_n28948_ );
and  ( new_n28954_, new_n28952_, new_n28948_ );
or   ( new_n28955_, new_n2122_, new_n23370_ );
or   ( new_n28956_, new_n2124_, new_n23252_ );
and  ( new_n28957_, new_n28956_, new_n28955_ );
xor  ( new_n28958_, new_n28957_, new_n1843_ );
nor  ( new_n28959_, new_n28958_, new_n28954_ );
nor  ( new_n28960_, new_n28959_, new_n28953_ );
nor  ( new_n28961_, new_n28960_, new_n28944_ );
nor  ( new_n28962_, new_n28961_, new_n28943_ );
or   ( new_n28963_, new_n28962_, new_n28910_ );
and  ( new_n28964_, new_n28963_, new_n28909_ );
xor  ( new_n28965_, new_n28546_, new_n28544_ );
xor  ( new_n28966_, new_n28965_, new_n28550_ );
xor  ( new_n28967_, new_n28342_, new_n7177_ );
xor  ( new_n28968_, new_n28967_, new_n28348_ );
or   ( new_n28969_, new_n28968_, new_n28966_ );
and  ( new_n28970_, new_n28968_, new_n28966_ );
xor  ( new_n28971_, new_n28523_, new_n28521_ );
xor  ( new_n28972_, new_n28971_, new_n28528_ );
or   ( new_n28973_, new_n28972_, new_n28970_ );
and  ( new_n28974_, new_n28973_, new_n28969_ );
and  ( new_n28975_, new_n28974_, new_n28964_ );
nor  ( new_n28976_, new_n28974_, new_n28964_ );
and  ( new_n28977_, RIbb32ec8_182, RIbb2f610_1 );
not  ( new_n28978_, new_n28977_ );
xnor ( new_n28979_, new_n28562_, new_n28558_ );
xor  ( new_n28980_, new_n28979_, new_n28568_ );
and  ( new_n28981_, new_n28980_, new_n28978_ );
xnor ( new_n28982_, new_n28614_, new_n28610_ );
xor  ( new_n28983_, new_n28982_, new_n28620_ );
xnor ( new_n28984_, new_n28665_, new_n28661_ );
xor  ( new_n28985_, new_n28984_, new_n28671_ );
or   ( new_n28986_, new_n28985_, new_n28983_ );
and  ( new_n28987_, new_n28985_, new_n28983_ );
xor  ( new_n28988_, new_n28699_, new_n28695_ );
xnor ( new_n28989_, new_n28988_, new_n28705_ );
or   ( new_n28990_, new_n28989_, new_n28987_ );
and  ( new_n28991_, new_n28990_, new_n28986_ );
nor  ( new_n28992_, new_n28991_, new_n28981_ );
and  ( new_n28993_, new_n28991_, new_n28981_ );
xnor ( new_n28994_, new_n28578_, new_n28574_ );
xor  ( new_n28995_, new_n28994_, new_n28584_ );
xnor ( new_n28996_, new_n28681_, new_n28677_ );
xor  ( new_n28997_, new_n28996_, new_n28687_ );
nor  ( new_n28998_, new_n28997_, new_n28995_ );
and  ( new_n28999_, new_n28997_, new_n28995_ );
xor  ( new_n29000_, new_n28596_, new_n28592_ );
xnor ( new_n29001_, new_n29000_, new_n28602_ );
nor  ( new_n29002_, new_n29001_, new_n28999_ );
nor  ( new_n29003_, new_n29002_, new_n28998_ );
nor  ( new_n29004_, new_n29003_, new_n28993_ );
nor  ( new_n29005_, new_n29004_, new_n28992_ );
nor  ( new_n29006_, new_n29005_, new_n28976_ );
nor  ( new_n29007_, new_n29006_, new_n28975_ );
nor  ( new_n29008_, new_n29007_, new_n28807_ );
nor  ( new_n29009_, new_n29008_, new_n28806_ );
nand ( new_n29010_, new_n29009_, new_n28777_ );
and  ( new_n29011_, new_n29010_, new_n28776_ );
nor  ( new_n29012_, new_n29011_, new_n28764_ );
nand ( new_n29013_, new_n29011_, new_n28764_ );
xor  ( new_n29014_, new_n28512_, new_n28503_ );
xor  ( new_n29015_, new_n29014_, new_n28747_ );
and  ( new_n29016_, new_n29015_, new_n29013_ );
or   ( new_n29017_, new_n29016_, new_n29012_ );
xnor ( new_n29018_, new_n28751_, new_n28749_ );
xor  ( new_n29019_, new_n29018_, new_n28755_ );
nor  ( new_n29020_, new_n29019_, new_n29017_ );
xor  ( new_n29021_, new_n28759_, new_n28757_ );
and  ( new_n29022_, new_n29021_, new_n29020_ );
xor  ( new_n29023_, new_n29011_, new_n28764_ );
xor  ( new_n29024_, new_n29023_, new_n29015_ );
xor  ( new_n29025_, new_n28726_, new_n28519_ );
xor  ( new_n29026_, new_n29025_, new_n28745_ );
xnor ( new_n29027_, new_n28781_, new_n28779_ );
xor  ( new_n29028_, new_n29027_, new_n28785_ );
xnor ( new_n29029_, new_n28974_, new_n28964_ );
xor  ( new_n29030_, new_n29029_, new_n29005_ );
or   ( new_n29031_, new_n29030_, new_n29028_ );
and  ( new_n29032_, new_n29030_, new_n29028_ );
xor  ( new_n29033_, new_n28799_, new_n28789_ );
xnor ( new_n29034_, new_n29033_, new_n28803_ );
or   ( new_n29035_, new_n29034_, new_n29032_ );
and  ( new_n29036_, new_n29035_, new_n29031_ );
xnor ( new_n29037_, new_n28997_, new_n28995_ );
xor  ( new_n29038_, new_n29037_, new_n29001_ );
xnor ( new_n29039_, new_n28985_, new_n28983_ );
xor  ( new_n29040_, new_n29039_, new_n28989_ );
nor  ( new_n29041_, new_n29040_, new_n29038_ );
nand ( new_n29042_, new_n29040_, new_n29038_ );
xor  ( new_n29043_, new_n28980_, new_n28978_ );
and  ( new_n29044_, new_n29043_, new_n29042_ );
or   ( new_n29045_, new_n29044_, new_n29041_ );
xnor ( new_n29046_, new_n28638_, new_n28622_ );
xor  ( new_n29047_, new_n29046_, new_n28654_ );
nor  ( new_n29048_, new_n29047_, new_n29045_ );
and  ( new_n29049_, new_n29047_, new_n29045_ );
xnor ( new_n29050_, new_n28942_, new_n28926_ );
xor  ( new_n29051_, new_n29050_, new_n28960_ );
xnor ( new_n29052_, new_n28888_, new_n28876_ );
xor  ( new_n29053_, new_n29052_, new_n28906_ );
nor  ( new_n29054_, new_n29053_, new_n29051_ );
and  ( new_n29055_, new_n29053_, new_n29051_ );
xor  ( new_n29056_, new_n28839_, new_n28823_ );
xnor ( new_n29057_, new_n29056_, new_n28857_ );
nor  ( new_n29058_, new_n29057_, new_n29055_ );
nor  ( new_n29059_, new_n29058_, new_n29054_ );
nor  ( new_n29060_, new_n29059_, new_n29049_ );
or   ( new_n29061_, new_n29060_, new_n29048_ );
xor  ( new_n29062_, new_n28898_, new_n28894_ );
xor  ( new_n29063_, new_n29062_, new_n28904_ );
xor  ( new_n29064_, new_n28880_, new_n7725_ );
xor  ( new_n29065_, new_n29064_, new_n28886_ );
nand ( new_n29066_, new_n29065_, new_n29063_ );
nor  ( new_n29067_, new_n29065_, new_n29063_ );
xor  ( new_n29068_, new_n28867_, new_n28863_ );
xor  ( new_n29069_, new_n29068_, new_n28874_ );
or   ( new_n29070_, new_n29069_, new_n29067_ );
and  ( new_n29071_, new_n29070_, new_n29066_ );
xnor ( new_n29072_, new_n28630_, new_n28626_ );
xor  ( new_n29073_, new_n29072_, new_n28636_ );
nor  ( new_n29074_, new_n29073_, new_n29071_ );
and  ( new_n29075_, new_n29073_, new_n29071_ );
xor  ( new_n29076_, new_n28646_, new_n28644_ );
xnor ( new_n29077_, new_n29076_, new_n28652_ );
nor  ( new_n29078_, new_n29077_, new_n29075_ );
or   ( new_n29079_, new_n29078_, new_n29074_ );
or   ( new_n29080_, new_n1844_, new_n23895_ );
or   ( new_n29081_, new_n1846_, new_n23733_ );
and  ( new_n29082_, new_n29081_, new_n29080_ );
xor  ( new_n29083_, new_n29082_, new_n1586_ );
or   ( new_n29084_, new_n1593_, new_n24227_ );
or   ( new_n29085_, new_n1595_, new_n24006_ );
and  ( new_n29086_, new_n29085_, new_n29084_ );
xor  ( new_n29087_, new_n29086_, new_n1358_ );
or   ( new_n29088_, new_n29087_, new_n29083_ );
and  ( new_n29089_, new_n29087_, new_n29083_ );
or   ( new_n29090_, new_n1364_, new_n24543_ );
or   ( new_n29091_, new_n1366_, new_n24418_ );
and  ( new_n29092_, new_n29091_, new_n29090_ );
xor  ( new_n29093_, new_n29092_, new_n1129_ );
or   ( new_n29094_, new_n29093_, new_n29089_ );
and  ( new_n29095_, new_n29094_, new_n29088_ );
or   ( new_n29096_, new_n2807_, new_n22973_ );
or   ( new_n29097_, new_n2809_, new_n22975_ );
and  ( new_n29098_, new_n29097_, new_n29096_ );
xor  ( new_n29099_, new_n29098_, new_n2424_ );
or   ( new_n29100_, new_n2425_, new_n23252_ );
or   ( new_n29101_, new_n2427_, new_n23166_ );
and  ( new_n29102_, new_n29101_, new_n29100_ );
xor  ( new_n29103_, new_n29102_, new_n2121_ );
or   ( new_n29104_, new_n29103_, new_n29099_ );
and  ( new_n29105_, new_n29103_, new_n29099_ );
or   ( new_n29106_, new_n2122_, new_n23554_ );
or   ( new_n29107_, new_n2124_, new_n23370_ );
and  ( new_n29108_, new_n29107_, new_n29106_ );
xor  ( new_n29109_, new_n29108_, new_n1843_ );
or   ( new_n29110_, new_n29109_, new_n29105_ );
and  ( new_n29111_, new_n29110_, new_n29104_ );
or   ( new_n29112_, new_n29111_, new_n29095_ );
and  ( new_n29113_, new_n29111_, new_n29095_ );
or   ( new_n29114_, new_n3896_, new_n22304_ );
or   ( new_n29115_, new_n3898_, new_n22207_ );
and  ( new_n29116_, new_n29115_, new_n29114_ );
xor  ( new_n29117_, new_n29116_, new_n3460_ );
or   ( new_n29118_, new_n3461_, new_n22590_ );
or   ( new_n29119_, new_n3463_, new_n22423_ );
and  ( new_n29120_, new_n29119_, new_n29118_ );
xor  ( new_n29121_, new_n29120_, new_n3116_ );
nor  ( new_n29122_, new_n29121_, new_n29117_ );
and  ( new_n29123_, new_n29121_, new_n29117_ );
or   ( new_n29124_, new_n3117_, new_n22829_ );
or   ( new_n29125_, new_n3119_, new_n22641_ );
and  ( new_n29126_, new_n29125_, new_n29124_ );
xor  ( new_n29127_, new_n29126_, new_n2800_ );
nor  ( new_n29128_, new_n29127_, new_n29123_ );
nor  ( new_n29129_, new_n29128_, new_n29122_ );
or   ( new_n29130_, new_n29129_, new_n29113_ );
and  ( new_n29131_, new_n29130_, new_n29112_ );
or   ( new_n29132_, new_n1135_, new_n24925_ );
or   ( new_n29133_, new_n1137_, new_n24927_ );
and  ( new_n29134_, new_n29133_, new_n29132_ );
xor  ( new_n29135_, new_n29134_, new_n896_ );
or   ( new_n29136_, new_n897_, new_n25288_ );
or   ( new_n29137_, new_n899_, new_n25048_ );
and  ( new_n29138_, new_n29137_, new_n29136_ );
xor  ( new_n29139_, new_n29138_, new_n748_ );
or   ( new_n29140_, new_n29139_, new_n29135_ );
and  ( new_n29141_, new_n29139_, new_n29135_ );
or   ( new_n29142_, new_n755_, new_n25813_ );
or   ( new_n29143_, new_n757_, new_n25486_ );
and  ( new_n29144_, new_n29143_, new_n29142_ );
xor  ( new_n29145_, new_n29144_, new_n523_ );
or   ( new_n29146_, new_n29145_, new_n29141_ );
and  ( new_n29147_, new_n29146_, new_n29140_ );
or   ( new_n29148_, new_n524_, new_n26063_ );
or   ( new_n29149_, new_n526_, new_n26196_ );
and  ( new_n29150_, new_n29149_, new_n29148_ );
xor  ( new_n29151_, new_n29150_, new_n403_ );
or   ( new_n29152_, new_n409_, new_n26620_ );
or   ( new_n29153_, new_n411_, new_n26372_ );
and  ( new_n29154_, new_n29153_, new_n29152_ );
xor  ( new_n29155_, new_n29154_, new_n328_ );
or   ( new_n29156_, new_n29155_, new_n29151_ );
and  ( new_n29157_, new_n29155_, new_n29151_ );
or   ( new_n29158_, new_n337_, new_n27085_ );
or   ( new_n29159_, new_n340_, new_n26762_ );
and  ( new_n29160_, new_n29159_, new_n29158_ );
xor  ( new_n29161_, new_n29160_, new_n332_ );
or   ( new_n29162_, new_n29161_, new_n29157_ );
and  ( new_n29163_, new_n29162_, new_n29156_ );
or   ( new_n29164_, new_n29163_, new_n29147_ );
and  ( new_n29165_, new_n29163_, new_n29147_ );
or   ( new_n29166_, new_n317_, new_n27602_ );
or   ( new_n29167_, new_n320_, new_n27396_ );
and  ( new_n29168_, new_n29167_, new_n29166_ );
xor  ( new_n29169_, new_n29168_, new_n312_ );
or   ( new_n29170_, new_n283_, new_n28108_ );
or   ( new_n29171_, new_n286_, new_n27763_ );
and  ( new_n29172_, new_n29171_, new_n29170_ );
xor  ( new_n29173_, new_n29172_, new_n278_ );
nor  ( new_n29174_, new_n29173_, new_n29169_ );
and  ( new_n29175_, new_n29173_, new_n29169_ );
or   ( new_n29176_, new_n299_, new_n28531_ );
or   ( new_n29177_, new_n302_, new_n28314_ );
and  ( new_n29178_, new_n29177_, new_n29176_ );
xor  ( new_n29179_, new_n29178_, new_n293_ );
nor  ( new_n29180_, new_n29179_, new_n29175_ );
nor  ( new_n29181_, new_n29180_, new_n29174_ );
or   ( new_n29182_, new_n29181_, new_n29165_ );
and  ( new_n29183_, new_n29182_, new_n29164_ );
or   ( new_n29184_, new_n29183_, new_n29131_ );
or   ( new_n29185_, new_n7732_, new_n21703_ );
or   ( new_n29186_, new_n7734_, new_n21694_ );
and  ( new_n29187_, new_n29186_, new_n29185_ );
xor  ( new_n29188_, new_n29187_, new_n7176_ );
and  ( new_n29189_, new_n8042_, RIbb315f0_129 );
xor  ( new_n29190_, new_n29189_, new_n7725_ );
nand ( new_n29191_, new_n29190_, new_n29188_ );
nor  ( new_n29192_, new_n29190_, new_n29188_ );
or   ( new_n29193_, new_n7184_, new_n21674_ );
or   ( new_n29194_, new_n7186_, new_n21701_ );
and  ( new_n29195_, new_n29194_, new_n29193_ );
xor  ( new_n29196_, new_n29195_, new_n6638_ );
or   ( new_n29197_, new_n29196_, new_n29192_ );
and  ( new_n29198_, new_n29197_, new_n29191_ );
or   ( new_n29199_, new_n5207_, new_n21842_ );
or   ( new_n29200_, new_n5209_, new_n21792_ );
and  ( new_n29201_, new_n29200_, new_n29199_ );
xor  ( new_n29202_, new_n29201_, new_n4708_ );
or   ( new_n29203_, new_n4709_, new_n21847_ );
or   ( new_n29204_, new_n4711_, new_n21840_ );
and  ( new_n29205_, new_n29204_, new_n29203_ );
xor  ( new_n29206_, new_n29205_, new_n4295_ );
or   ( new_n29207_, new_n29206_, new_n29202_ );
and  ( new_n29208_, new_n29206_, new_n29202_ );
or   ( new_n29209_, new_n4302_, new_n22129_ );
or   ( new_n29210_, new_n4304_, new_n22098_ );
and  ( new_n29211_, new_n29210_, new_n29209_ );
xor  ( new_n29212_, new_n29211_, new_n3895_ );
or   ( new_n29213_, new_n29212_, new_n29208_ );
and  ( new_n29214_, new_n29213_, new_n29207_ );
nor  ( new_n29215_, new_n29214_, new_n29198_ );
and  ( new_n29216_, new_n29214_, new_n29198_ );
or   ( new_n29217_, new_n6645_, new_n21680_ );
or   ( new_n29218_, new_n6647_, new_n21672_ );
and  ( new_n29219_, new_n29218_, new_n29217_ );
xor  ( new_n29220_, new_n29219_, new_n6166_ );
or   ( new_n29221_, new_n6173_, new_n21687_ );
or   ( new_n29222_, new_n6175_, new_n21678_ );
and  ( new_n29223_, new_n29222_, new_n29221_ );
xor  ( new_n29224_, new_n29223_, new_n5597_ );
nor  ( new_n29225_, new_n29224_, new_n29220_ );
and  ( new_n29226_, new_n29224_, new_n29220_ );
or   ( new_n29227_, new_n5604_, new_n21751_ );
or   ( new_n29228_, new_n5606_, new_n21685_ );
and  ( new_n29229_, new_n29228_, new_n29227_ );
xor  ( new_n29230_, new_n29229_, new_n5206_ );
nor  ( new_n29231_, new_n29230_, new_n29226_ );
nor  ( new_n29232_, new_n29231_, new_n29225_ );
nor  ( new_n29233_, new_n29232_, new_n29216_ );
nor  ( new_n29234_, new_n29233_, new_n29215_ );
and  ( new_n29235_, new_n29183_, new_n29131_ );
or   ( new_n29236_, new_n29235_, new_n29234_ );
and  ( new_n29237_, new_n29236_, new_n29184_ );
or   ( new_n29238_, new_n29237_, new_n29079_ );
xnor ( new_n29239_, new_n28831_, new_n28827_ );
xor  ( new_n29240_, new_n29239_, new_n28837_ );
xnor ( new_n29241_, new_n28815_, new_n28811_ );
xor  ( new_n29242_, new_n29241_, new_n28821_ );
or   ( new_n29243_, new_n29242_, new_n29240_ );
and  ( new_n29244_, new_n29242_, new_n29240_ );
xor  ( new_n29245_, new_n28849_, new_n28845_ );
xnor ( new_n29246_, new_n29245_, new_n28855_ );
or   ( new_n29247_, new_n29246_, new_n29244_ );
and  ( new_n29248_, new_n29247_, new_n29243_ );
xnor ( new_n29249_, new_n28934_, new_n28930_ );
xor  ( new_n29250_, new_n29249_, new_n28940_ );
xnor ( new_n29251_, new_n28918_, new_n28914_ );
xor  ( new_n29252_, new_n29251_, new_n28924_ );
or   ( new_n29253_, new_n29252_, new_n29250_ );
and  ( new_n29254_, new_n29252_, new_n29250_ );
xor  ( new_n29255_, new_n28952_, new_n28948_ );
xnor ( new_n29256_, new_n29255_, new_n28958_ );
or   ( new_n29257_, new_n29256_, new_n29254_ );
and  ( new_n29258_, new_n29257_, new_n29253_ );
nor  ( new_n29259_, new_n29258_, new_n29248_ );
nand ( new_n29260_, new_n29258_, new_n29248_ );
not  ( new_n29261_, RIbb32f40_183 );
or   ( new_n29262_, new_n268_, new_n29261_ );
not  ( new_n29263_, RIbb32ec8_182 );
or   ( new_n29264_, new_n271_, new_n29263_ );
and  ( new_n29265_, new_n29264_, new_n29262_ );
xor  ( new_n29266_, new_n29265_, new_n263_ );
and  ( new_n29267_, RIbb32fb8_184, RIbb2f610_1 );
or   ( new_n29268_, new_n29267_, new_n29266_ );
or   ( new_n29269_, new_n268_, new_n29263_ );
or   ( new_n29270_, new_n271_, new_n28531_ );
and  ( new_n29271_, new_n29270_, new_n29269_ );
xor  ( new_n29272_, new_n29271_, new_n263_ );
nor  ( new_n29273_, new_n29272_, new_n29268_ );
and  ( new_n29274_, new_n29272_, new_n29268_ );
and  ( new_n29275_, RIbb32f40_183, RIbb2f610_1 );
nor  ( new_n29276_, new_n29275_, new_n29274_ );
nor  ( new_n29277_, new_n29276_, new_n29273_ );
and  ( new_n29278_, new_n29277_, new_n29260_ );
or   ( new_n29279_, new_n29278_, new_n29259_ );
and  ( new_n29280_, new_n29237_, new_n29079_ );
or   ( new_n29281_, new_n29280_, new_n29279_ );
and  ( new_n29282_, new_n29281_, new_n29238_ );
or   ( new_n29283_, new_n29282_, new_n29061_ );
nand ( new_n29284_, new_n29282_, new_n29061_ );
xnor ( new_n29285_, new_n28991_, new_n28981_ );
xor  ( new_n29286_, new_n29285_, new_n29003_ );
xnor ( new_n29287_, new_n28793_, new_n28791_ );
xor  ( new_n29288_, new_n29287_, new_n28797_ );
and  ( new_n29289_, new_n29288_, new_n29286_ );
nor  ( new_n29290_, new_n29288_, new_n29286_ );
xor  ( new_n29291_, new_n28968_, new_n28966_ );
xnor ( new_n29292_, new_n29291_, new_n28972_ );
nor  ( new_n29293_, new_n29292_, new_n29290_ );
nor  ( new_n29294_, new_n29293_, new_n29289_ );
nand ( new_n29295_, new_n29294_, new_n29284_ );
and  ( new_n29296_, new_n29295_, new_n29283_ );
nand ( new_n29297_, new_n29296_, new_n29036_ );
nor  ( new_n29298_, new_n29296_, new_n29036_ );
xor  ( new_n29299_, new_n28770_, new_n28768_ );
xor  ( new_n29300_, new_n29299_, new_n28773_ );
or   ( new_n29301_, new_n29300_, new_n29298_ );
and  ( new_n29302_, new_n29301_, new_n29297_ );
or   ( new_n29303_, new_n29302_, new_n29026_ );
and  ( new_n29304_, new_n29302_, new_n29026_ );
xor  ( new_n29305_, new_n28775_, new_n28766_ );
xor  ( new_n29306_, new_n29305_, new_n29009_ );
or   ( new_n29307_, new_n29306_, new_n29304_ );
and  ( new_n29308_, new_n29307_, new_n29303_ );
nor  ( new_n29309_, new_n29308_, new_n29024_ );
xor  ( new_n29310_, new_n29019_, new_n29017_ );
and  ( new_n29311_, new_n29310_, new_n29309_ );
xnor ( new_n29312_, new_n29302_, new_n29026_ );
xor  ( new_n29313_, new_n29312_, new_n29306_ );
or   ( new_n29314_, new_n1364_, new_n24927_ );
or   ( new_n29315_, new_n1366_, new_n24543_ );
and  ( new_n29316_, new_n29315_, new_n29314_ );
xor  ( new_n29317_, new_n29316_, new_n1129_ );
or   ( new_n29318_, new_n1135_, new_n25048_ );
or   ( new_n29319_, new_n1137_, new_n24925_ );
and  ( new_n29320_, new_n29319_, new_n29318_ );
xor  ( new_n29321_, new_n29320_, new_n896_ );
or   ( new_n29322_, new_n29321_, new_n29317_ );
and  ( new_n29323_, new_n29321_, new_n29317_ );
or   ( new_n29324_, new_n897_, new_n25486_ );
or   ( new_n29325_, new_n899_, new_n25288_ );
and  ( new_n29326_, new_n29325_, new_n29324_ );
xor  ( new_n29327_, new_n29326_, new_n748_ );
or   ( new_n29328_, new_n29327_, new_n29323_ );
and  ( new_n29329_, new_n29328_, new_n29322_ );
or   ( new_n29330_, new_n755_, new_n26196_ );
or   ( new_n29331_, new_n757_, new_n25813_ );
and  ( new_n29332_, new_n29331_, new_n29330_ );
xor  ( new_n29333_, new_n29332_, new_n523_ );
or   ( new_n29334_, new_n524_, new_n26372_ );
or   ( new_n29335_, new_n526_, new_n26063_ );
and  ( new_n29336_, new_n29335_, new_n29334_ );
xor  ( new_n29337_, new_n29336_, new_n403_ );
or   ( new_n29338_, new_n29337_, new_n29333_ );
and  ( new_n29339_, new_n29337_, new_n29333_ );
or   ( new_n29340_, new_n409_, new_n26762_ );
or   ( new_n29341_, new_n411_, new_n26620_ );
and  ( new_n29342_, new_n29341_, new_n29340_ );
xor  ( new_n29343_, new_n29342_, new_n328_ );
or   ( new_n29344_, new_n29343_, new_n29339_ );
and  ( new_n29345_, new_n29344_, new_n29338_ );
or   ( new_n29346_, new_n29345_, new_n29329_ );
and  ( new_n29347_, new_n29345_, new_n29329_ );
or   ( new_n29348_, new_n337_, new_n27396_ );
or   ( new_n29349_, new_n340_, new_n27085_ );
and  ( new_n29350_, new_n29349_, new_n29348_ );
xor  ( new_n29351_, new_n29350_, new_n332_ );
or   ( new_n29352_, new_n317_, new_n27763_ );
or   ( new_n29353_, new_n320_, new_n27602_ );
and  ( new_n29354_, new_n29353_, new_n29352_ );
xor  ( new_n29355_, new_n29354_, new_n312_ );
or   ( new_n29356_, new_n29355_, new_n29351_ );
and  ( new_n29357_, new_n29355_, new_n29351_ );
or   ( new_n29358_, new_n283_, new_n28314_ );
or   ( new_n29359_, new_n286_, new_n28108_ );
and  ( new_n29360_, new_n29359_, new_n29358_ );
xor  ( new_n29361_, new_n29360_, new_n278_ );
or   ( new_n29362_, new_n29361_, new_n29357_ );
and  ( new_n29363_, new_n29362_, new_n29356_ );
or   ( new_n29364_, new_n29363_, new_n29347_ );
and  ( new_n29365_, new_n29364_, new_n29346_ );
or   ( new_n29366_, new_n7184_, new_n21672_ );
or   ( new_n29367_, new_n7186_, new_n21674_ );
and  ( new_n29368_, new_n29367_, new_n29366_ );
xor  ( new_n29369_, new_n29368_, new_n6638_ );
or   ( new_n29370_, new_n6645_, new_n21678_ );
or   ( new_n29371_, new_n6647_, new_n21680_ );
and  ( new_n29372_, new_n29371_, new_n29370_ );
xor  ( new_n29373_, new_n29372_, new_n6166_ );
nor  ( new_n29374_, new_n29373_, new_n29369_ );
nand ( new_n29375_, new_n29373_, new_n29369_ );
or   ( new_n29376_, new_n6173_, new_n21685_ );
or   ( new_n29377_, new_n6175_, new_n21687_ );
and  ( new_n29378_, new_n29377_, new_n29376_ );
xor  ( new_n29379_, new_n29378_, new_n5596_ );
and  ( new_n29380_, new_n29379_, new_n29375_ );
or   ( new_n29381_, new_n29380_, new_n29374_ );
or   ( new_n29382_, new_n7732_, new_n21701_ );
or   ( new_n29383_, new_n7734_, new_n21703_ );
and  ( new_n29384_, new_n29383_, new_n29382_ );
xor  ( new_n29385_, new_n29384_, new_n7177_ );
nand ( new_n29386_, new_n29385_, new_n8257_ );
or   ( new_n29387_, new_n29385_, new_n8257_ );
or   ( new_n29388_, new_n8264_, new_n21694_ );
or   ( new_n29389_, new_n8266_, new_n21696_ );
and  ( new_n29390_, new_n29389_, new_n29388_ );
xor  ( new_n29391_, new_n29390_, new_n7725_ );
nand ( new_n29392_, new_n29391_, new_n29387_ );
and  ( new_n29393_, new_n29392_, new_n29386_ );
nand ( new_n29394_, new_n29393_, new_n29381_ );
nor  ( new_n29395_, new_n29393_, new_n29381_ );
or   ( new_n29396_, new_n5604_, new_n21792_ );
or   ( new_n29397_, new_n5606_, new_n21751_ );
and  ( new_n29398_, new_n29397_, new_n29396_ );
xor  ( new_n29399_, new_n29398_, new_n5206_ );
or   ( new_n29400_, new_n5207_, new_n21840_ );
or   ( new_n29401_, new_n5209_, new_n21842_ );
and  ( new_n29402_, new_n29401_, new_n29400_ );
xor  ( new_n29403_, new_n29402_, new_n4708_ );
nor  ( new_n29404_, new_n29403_, new_n29399_ );
and  ( new_n29405_, new_n29403_, new_n29399_ );
or   ( new_n29406_, new_n4709_, new_n22098_ );
or   ( new_n29407_, new_n4711_, new_n21847_ );
and  ( new_n29408_, new_n29407_, new_n29406_ );
xor  ( new_n29409_, new_n29408_, new_n4295_ );
nor  ( new_n29410_, new_n29409_, new_n29405_ );
nor  ( new_n29411_, new_n29410_, new_n29404_ );
or   ( new_n29412_, new_n29411_, new_n29395_ );
and  ( new_n29413_, new_n29412_, new_n29394_ );
nor  ( new_n29414_, new_n29413_, new_n29365_ );
and  ( new_n29415_, new_n29413_, new_n29365_ );
or   ( new_n29416_, new_n3117_, new_n22975_ );
or   ( new_n29417_, new_n3119_, new_n22829_ );
and  ( new_n29418_, new_n29417_, new_n29416_ );
xor  ( new_n29419_, new_n29418_, new_n2800_ );
or   ( new_n29420_, new_n2807_, new_n23166_ );
or   ( new_n29421_, new_n2809_, new_n22973_ );
and  ( new_n29422_, new_n29421_, new_n29420_ );
xor  ( new_n29423_, new_n29422_, new_n2424_ );
or   ( new_n29424_, new_n29423_, new_n29419_ );
and  ( new_n29425_, new_n29423_, new_n29419_ );
or   ( new_n29426_, new_n2425_, new_n23370_ );
or   ( new_n29427_, new_n2427_, new_n23252_ );
and  ( new_n29428_, new_n29427_, new_n29426_ );
xor  ( new_n29429_, new_n29428_, new_n2121_ );
or   ( new_n29430_, new_n29429_, new_n29425_ );
and  ( new_n29431_, new_n29430_, new_n29424_ );
or   ( new_n29432_, new_n2122_, new_n23733_ );
or   ( new_n29433_, new_n2124_, new_n23554_ );
and  ( new_n29434_, new_n29433_, new_n29432_ );
xor  ( new_n29435_, new_n29434_, new_n1843_ );
or   ( new_n29436_, new_n1844_, new_n24006_ );
or   ( new_n29437_, new_n1846_, new_n23895_ );
and  ( new_n29438_, new_n29437_, new_n29436_ );
xor  ( new_n29439_, new_n29438_, new_n1586_ );
or   ( new_n29440_, new_n29439_, new_n29435_ );
and  ( new_n29441_, new_n29439_, new_n29435_ );
or   ( new_n29442_, new_n1593_, new_n24418_ );
or   ( new_n29443_, new_n1595_, new_n24227_ );
and  ( new_n29444_, new_n29443_, new_n29442_ );
xor  ( new_n29445_, new_n29444_, new_n1358_ );
or   ( new_n29446_, new_n29445_, new_n29441_ );
and  ( new_n29447_, new_n29446_, new_n29440_ );
nor  ( new_n29448_, new_n29447_, new_n29431_ );
and  ( new_n29449_, new_n29447_, new_n29431_ );
or   ( new_n29450_, new_n4302_, new_n22207_ );
or   ( new_n29451_, new_n4304_, new_n22129_ );
and  ( new_n29452_, new_n29451_, new_n29450_ );
xor  ( new_n29453_, new_n29452_, new_n3895_ );
or   ( new_n29454_, new_n3896_, new_n22423_ );
or   ( new_n29455_, new_n3898_, new_n22304_ );
and  ( new_n29456_, new_n29455_, new_n29454_ );
xor  ( new_n29457_, new_n29456_, new_n3460_ );
nor  ( new_n29458_, new_n29457_, new_n29453_ );
and  ( new_n29459_, new_n29457_, new_n29453_ );
or   ( new_n29460_, new_n3461_, new_n22641_ );
or   ( new_n29461_, new_n3463_, new_n22590_ );
and  ( new_n29462_, new_n29461_, new_n29460_ );
xor  ( new_n29463_, new_n29462_, new_n3116_ );
nor  ( new_n29464_, new_n29463_, new_n29459_ );
nor  ( new_n29465_, new_n29464_, new_n29458_ );
nor  ( new_n29466_, new_n29465_, new_n29449_ );
nor  ( new_n29467_, new_n29466_, new_n29448_ );
nor  ( new_n29468_, new_n29467_, new_n29415_ );
or   ( new_n29469_, new_n29468_, new_n29414_ );
or   ( new_n29470_, new_n299_, new_n29263_ );
or   ( new_n29471_, new_n302_, new_n28531_ );
and  ( new_n29472_, new_n29471_, new_n29470_ );
xor  ( new_n29473_, new_n29472_, new_n293_ );
not  ( new_n29474_, RIbb32fb8_184 );
or   ( new_n29475_, new_n268_, new_n29474_ );
or   ( new_n29476_, new_n271_, new_n29261_ );
and  ( new_n29477_, new_n29476_, new_n29475_ );
xor  ( new_n29478_, new_n29477_, new_n263_ );
nor  ( new_n29479_, new_n29478_, new_n29473_ );
and  ( new_n29480_, RIbb33030_185, RIbb2f610_1 );
not  ( new_n29481_, new_n29480_ );
nand ( new_n29482_, new_n29478_, new_n29473_ );
and  ( new_n29483_, new_n29482_, new_n29481_ );
or   ( new_n29484_, new_n29483_, new_n29479_ );
xnor ( new_n29485_, new_n29173_, new_n29169_ );
xor  ( new_n29486_, new_n29485_, new_n29179_ );
or   ( new_n29487_, new_n29486_, new_n29484_ );
and  ( new_n29488_, new_n29486_, new_n29484_ );
xor  ( new_n29489_, new_n29267_, new_n29266_ );
or   ( new_n29490_, new_n29489_, new_n29488_ );
and  ( new_n29491_, new_n29490_, new_n29487_ );
xnor ( new_n29492_, new_n29103_, new_n29099_ );
xor  ( new_n29493_, new_n29492_, new_n29109_ );
xnor ( new_n29494_, new_n29206_, new_n29202_ );
xor  ( new_n29495_, new_n29494_, new_n29212_ );
or   ( new_n29496_, new_n29495_, new_n29493_ );
and  ( new_n29497_, new_n29495_, new_n29493_ );
xor  ( new_n29498_, new_n29121_, new_n29117_ );
xnor ( new_n29499_, new_n29498_, new_n29127_ );
or   ( new_n29500_, new_n29499_, new_n29497_ );
and  ( new_n29501_, new_n29500_, new_n29496_ );
or   ( new_n29502_, new_n29501_, new_n29491_ );
and  ( new_n29503_, new_n29501_, new_n29491_ );
xnor ( new_n29504_, new_n29087_, new_n29083_ );
xor  ( new_n29505_, new_n29504_, new_n29093_ );
xnor ( new_n29506_, new_n29155_, new_n29151_ );
xor  ( new_n29507_, new_n29506_, new_n29161_ );
nor  ( new_n29508_, new_n29507_, new_n29505_ );
and  ( new_n29509_, new_n29507_, new_n29505_ );
xor  ( new_n29510_, new_n29139_, new_n29135_ );
xnor ( new_n29511_, new_n29510_, new_n29145_ );
nor  ( new_n29512_, new_n29511_, new_n29509_ );
nor  ( new_n29513_, new_n29512_, new_n29508_ );
or   ( new_n29514_, new_n29513_, new_n29503_ );
and  ( new_n29515_, new_n29514_, new_n29502_ );
and  ( new_n29516_, new_n29515_, new_n29469_ );
or   ( new_n29517_, new_n29515_, new_n29469_ );
xnor ( new_n29518_, new_n29242_, new_n29240_ );
xor  ( new_n29519_, new_n29518_, new_n29246_ );
xnor ( new_n29520_, new_n29252_, new_n29250_ );
xor  ( new_n29521_, new_n29520_, new_n29256_ );
nor  ( new_n29522_, new_n29521_, new_n29519_ );
nand ( new_n29523_, new_n29521_, new_n29519_ );
xor  ( new_n29524_, new_n29065_, new_n29063_ );
xnor ( new_n29525_, new_n29524_, new_n29069_ );
not  ( new_n29526_, new_n29525_ );
and  ( new_n29527_, new_n29526_, new_n29523_ );
or   ( new_n29528_, new_n29527_, new_n29522_ );
and  ( new_n29529_, new_n29528_, new_n29517_ );
or   ( new_n29530_, new_n29529_, new_n29516_ );
xnor ( new_n29531_, new_n29258_, new_n29248_ );
xor  ( new_n29532_, new_n29531_, new_n29277_ );
xnor ( new_n29533_, new_n29183_, new_n29131_ );
xor  ( new_n29534_, new_n29533_, new_n29234_ );
or   ( new_n29535_, new_n29534_, new_n29532_ );
and  ( new_n29536_, new_n29534_, new_n29532_ );
xor  ( new_n29537_, new_n29073_, new_n29071_ );
xor  ( new_n29538_, new_n29537_, new_n29077_ );
or   ( new_n29539_, new_n29538_, new_n29536_ );
and  ( new_n29540_, new_n29539_, new_n29535_ );
or   ( new_n29541_, new_n29540_, new_n29530_ );
and  ( new_n29542_, new_n29540_, new_n29530_ );
xnor ( new_n29543_, new_n29040_, new_n29038_ );
xor  ( new_n29544_, new_n29543_, new_n29043_ );
xnor ( new_n29545_, new_n29053_, new_n29051_ );
xor  ( new_n29546_, new_n29545_, new_n29057_ );
and  ( new_n29547_, new_n29546_, new_n29544_ );
nor  ( new_n29548_, new_n29546_, new_n29544_ );
xnor ( new_n29549_, new_n29111_, new_n29095_ );
xor  ( new_n29550_, new_n29549_, new_n29129_ );
xnor ( new_n29551_, new_n29163_, new_n29147_ );
xor  ( new_n29552_, new_n29551_, new_n29181_ );
nor  ( new_n29553_, new_n29552_, new_n29550_ );
and  ( new_n29554_, new_n29552_, new_n29550_ );
xor  ( new_n29555_, new_n29272_, new_n29268_ );
xnor ( new_n29556_, new_n29555_, new_n29275_ );
nor  ( new_n29557_, new_n29556_, new_n29554_ );
nor  ( new_n29558_, new_n29557_, new_n29553_ );
nor  ( new_n29559_, new_n29558_, new_n29548_ );
nor  ( new_n29560_, new_n29559_, new_n29547_ );
or   ( new_n29561_, new_n29560_, new_n29542_ );
and  ( new_n29562_, new_n29561_, new_n29541_ );
xor  ( new_n29563_, new_n29047_, new_n29045_ );
xor  ( new_n29564_, new_n29563_, new_n29059_ );
xnor ( new_n29565_, new_n28908_, new_n28859_ );
xor  ( new_n29566_, new_n29565_, new_n28962_ );
or   ( new_n29567_, new_n29566_, new_n29564_ );
and  ( new_n29568_, new_n29566_, new_n29564_ );
xor  ( new_n29569_, new_n29288_, new_n29286_ );
xor  ( new_n29570_, new_n29569_, new_n29292_ );
or   ( new_n29571_, new_n29570_, new_n29568_ );
and  ( new_n29572_, new_n29571_, new_n29567_ );
or   ( new_n29573_, new_n29572_, new_n29562_ );
and  ( new_n29574_, new_n29572_, new_n29562_ );
xor  ( new_n29575_, new_n29030_, new_n29028_ );
xnor ( new_n29576_, new_n29575_, new_n29034_ );
or   ( new_n29577_, new_n29576_, new_n29574_ );
and  ( new_n29578_, new_n29577_, new_n29573_ );
xor  ( new_n29579_, new_n29296_, new_n29036_ );
xor  ( new_n29580_, new_n29579_, new_n29300_ );
nand ( new_n29581_, new_n29580_, new_n29578_ );
nor  ( new_n29582_, new_n29580_, new_n29578_ );
xor  ( new_n29583_, new_n28805_, new_n28787_ );
xnor ( new_n29584_, new_n29583_, new_n29007_ );
or   ( new_n29585_, new_n29584_, new_n29582_ );
and  ( new_n29586_, new_n29585_, new_n29581_ );
and  ( new_n29587_, new_n29586_, new_n29313_ );
xor  ( new_n29588_, new_n29308_, new_n29024_ );
and  ( new_n29589_, new_n29588_, new_n29587_ );
xor  ( new_n29590_, new_n29540_, new_n29530_ );
xnor ( new_n29591_, new_n29590_, new_n29560_ );
xor  ( new_n29592_, new_n29566_, new_n29564_ );
xnor ( new_n29593_, new_n29592_, new_n29570_ );
and  ( new_n29594_, new_n29593_, new_n29591_ );
xor  ( new_n29595_, new_n29237_, new_n29079_ );
xor  ( new_n29596_, new_n29595_, new_n29279_ );
xnor ( new_n29597_, new_n29214_, new_n29198_ );
xor  ( new_n29598_, new_n29597_, new_n29232_ );
xor  ( new_n29599_, new_n29345_, new_n29329_ );
xor  ( new_n29600_, new_n29599_, new_n29363_ );
xnor ( new_n29601_, new_n29507_, new_n29505_ );
xor  ( new_n29602_, new_n29601_, new_n29511_ );
nand ( new_n29603_, new_n29602_, new_n29600_ );
nor  ( new_n29604_, new_n29602_, new_n29600_ );
xor  ( new_n29605_, new_n29486_, new_n29484_ );
xor  ( new_n29606_, new_n29605_, new_n29489_ );
or   ( new_n29607_, new_n29606_, new_n29604_ );
and  ( new_n29608_, new_n29607_, new_n29603_ );
nor  ( new_n29609_, new_n29608_, new_n29598_ );
nand ( new_n29610_, new_n29608_, new_n29598_ );
xor  ( new_n29611_, new_n29552_, new_n29550_ );
xnor ( new_n29612_, new_n29611_, new_n29556_ );
and  ( new_n29613_, new_n29612_, new_n29610_ );
or   ( new_n29614_, new_n29613_, new_n29609_ );
or   ( new_n29615_, new_n299_, new_n29261_ );
or   ( new_n29616_, new_n302_, new_n29263_ );
and  ( new_n29617_, new_n29616_, new_n29615_ );
xor  ( new_n29618_, new_n29617_, new_n293_ );
not  ( new_n29619_, RIbb33030_185 );
or   ( new_n29620_, new_n268_, new_n29619_ );
or   ( new_n29621_, new_n271_, new_n29474_ );
and  ( new_n29622_, new_n29621_, new_n29620_ );
xor  ( new_n29623_, new_n29622_, new_n263_ );
nor  ( new_n29624_, new_n29623_, new_n29618_ );
and  ( new_n29625_, RIbb330a8_186, RIbb2f610_1 );
not  ( new_n29626_, new_n29625_ );
nand ( new_n29627_, new_n29623_, new_n29618_ );
and  ( new_n29628_, new_n29627_, new_n29626_ );
or   ( new_n29629_, new_n29628_, new_n29624_ );
xnor ( new_n29630_, new_n29355_, new_n29351_ );
xor  ( new_n29631_, new_n29630_, new_n29361_ );
and  ( new_n29632_, new_n29631_, new_n29629_ );
or   ( new_n29633_, new_n29631_, new_n29629_ );
xor  ( new_n29634_, new_n29478_, new_n29473_ );
xor  ( new_n29635_, new_n29634_, new_n29481_ );
and  ( new_n29636_, new_n29635_, new_n29633_ );
or   ( new_n29637_, new_n29636_, new_n29632_ );
xnor ( new_n29638_, new_n29403_, new_n29399_ );
xor  ( new_n29639_, new_n29638_, new_n29409_ );
xnor ( new_n29640_, new_n29423_, new_n29419_ );
xor  ( new_n29641_, new_n29640_, new_n29429_ );
or   ( new_n29642_, new_n29641_, new_n29639_ );
and  ( new_n29643_, new_n29641_, new_n29639_ );
xor  ( new_n29644_, new_n29457_, new_n29453_ );
xnor ( new_n29645_, new_n29644_, new_n29463_ );
or   ( new_n29646_, new_n29645_, new_n29643_ );
and  ( new_n29647_, new_n29646_, new_n29642_ );
nor  ( new_n29648_, new_n29647_, new_n29637_ );
nand ( new_n29649_, new_n29647_, new_n29637_ );
xnor ( new_n29650_, new_n29439_, new_n29435_ );
xor  ( new_n29651_, new_n29650_, new_n29445_ );
xnor ( new_n29652_, new_n29337_, new_n29333_ );
xor  ( new_n29653_, new_n29652_, new_n29343_ );
nor  ( new_n29654_, new_n29653_, new_n29651_ );
nand ( new_n29655_, new_n29653_, new_n29651_ );
xor  ( new_n29656_, new_n29321_, new_n29317_ );
xor  ( new_n29657_, new_n29656_, new_n29327_ );
and  ( new_n29658_, new_n29657_, new_n29655_ );
or   ( new_n29659_, new_n29658_, new_n29654_ );
and  ( new_n29660_, new_n29659_, new_n29649_ );
or   ( new_n29661_, new_n29660_, new_n29648_ );
or   ( new_n29662_, new_n4302_, new_n22304_ );
or   ( new_n29663_, new_n4304_, new_n22207_ );
and  ( new_n29664_, new_n29663_, new_n29662_ );
xor  ( new_n29665_, new_n29664_, new_n3895_ );
or   ( new_n29666_, new_n3896_, new_n22590_ );
or   ( new_n29667_, new_n3898_, new_n22423_ );
and  ( new_n29668_, new_n29667_, new_n29666_ );
xor  ( new_n29669_, new_n29668_, new_n3460_ );
or   ( new_n29670_, new_n29669_, new_n29665_ );
and  ( new_n29671_, new_n29669_, new_n29665_ );
or   ( new_n29672_, new_n3461_, new_n22829_ );
or   ( new_n29673_, new_n3463_, new_n22641_ );
and  ( new_n29674_, new_n29673_, new_n29672_ );
xor  ( new_n29675_, new_n29674_, new_n3116_ );
or   ( new_n29676_, new_n29675_, new_n29671_ );
and  ( new_n29677_, new_n29676_, new_n29670_ );
or   ( new_n29678_, new_n2122_, new_n23895_ );
or   ( new_n29679_, new_n2124_, new_n23733_ );
and  ( new_n29680_, new_n29679_, new_n29678_ );
xor  ( new_n29681_, new_n29680_, new_n1843_ );
or   ( new_n29682_, new_n1844_, new_n24227_ );
or   ( new_n29683_, new_n1846_, new_n24006_ );
and  ( new_n29684_, new_n29683_, new_n29682_ );
xor  ( new_n29685_, new_n29684_, new_n1586_ );
or   ( new_n29686_, new_n29685_, new_n29681_ );
and  ( new_n29687_, new_n29685_, new_n29681_ );
or   ( new_n29688_, new_n1593_, new_n24543_ );
or   ( new_n29689_, new_n1595_, new_n24418_ );
and  ( new_n29690_, new_n29689_, new_n29688_ );
xor  ( new_n29691_, new_n29690_, new_n1358_ );
or   ( new_n29692_, new_n29691_, new_n29687_ );
and  ( new_n29693_, new_n29692_, new_n29686_ );
or   ( new_n29694_, new_n29693_, new_n29677_ );
and  ( new_n29695_, new_n29693_, new_n29677_ );
or   ( new_n29696_, new_n3117_, new_n22973_ );
or   ( new_n29697_, new_n3119_, new_n22975_ );
and  ( new_n29698_, new_n29697_, new_n29696_ );
xor  ( new_n29699_, new_n29698_, new_n2800_ );
or   ( new_n29700_, new_n2807_, new_n23252_ );
or   ( new_n29701_, new_n2809_, new_n23166_ );
and  ( new_n29702_, new_n29701_, new_n29700_ );
xor  ( new_n29703_, new_n29702_, new_n2424_ );
nor  ( new_n29704_, new_n29703_, new_n29699_ );
and  ( new_n29705_, new_n29703_, new_n29699_ );
or   ( new_n29706_, new_n2425_, new_n23554_ );
or   ( new_n29707_, new_n2427_, new_n23370_ );
and  ( new_n29708_, new_n29707_, new_n29706_ );
xor  ( new_n29709_, new_n29708_, new_n2121_ );
nor  ( new_n29710_, new_n29709_, new_n29705_ );
nor  ( new_n29711_, new_n29710_, new_n29704_ );
or   ( new_n29712_, new_n29711_, new_n29695_ );
and  ( new_n29713_, new_n29712_, new_n29694_ );
or   ( new_n29714_, new_n755_, new_n26063_ );
or   ( new_n29715_, new_n757_, new_n26196_ );
and  ( new_n29716_, new_n29715_, new_n29714_ );
xor  ( new_n29717_, new_n29716_, new_n523_ );
or   ( new_n29718_, new_n524_, new_n26620_ );
or   ( new_n29719_, new_n526_, new_n26372_ );
and  ( new_n29720_, new_n29719_, new_n29718_ );
xor  ( new_n29721_, new_n29720_, new_n403_ );
or   ( new_n29722_, new_n29721_, new_n29717_ );
and  ( new_n29723_, new_n29721_, new_n29717_ );
or   ( new_n29724_, new_n409_, new_n27085_ );
or   ( new_n29725_, new_n411_, new_n26762_ );
and  ( new_n29726_, new_n29725_, new_n29724_ );
xor  ( new_n29727_, new_n29726_, new_n328_ );
or   ( new_n29728_, new_n29727_, new_n29723_ );
and  ( new_n29729_, new_n29728_, new_n29722_ );
or   ( new_n29730_, new_n337_, new_n27602_ );
or   ( new_n29731_, new_n340_, new_n27396_ );
and  ( new_n29732_, new_n29731_, new_n29730_ );
xor  ( new_n29733_, new_n29732_, new_n332_ );
or   ( new_n29734_, new_n317_, new_n28108_ );
or   ( new_n29735_, new_n320_, new_n27763_ );
and  ( new_n29736_, new_n29735_, new_n29734_ );
xor  ( new_n29737_, new_n29736_, new_n312_ );
or   ( new_n29738_, new_n29737_, new_n29733_ );
and  ( new_n29739_, new_n29737_, new_n29733_ );
or   ( new_n29740_, new_n283_, new_n28531_ );
or   ( new_n29741_, new_n286_, new_n28314_ );
and  ( new_n29742_, new_n29741_, new_n29740_ );
xor  ( new_n29743_, new_n29742_, new_n278_ );
or   ( new_n29744_, new_n29743_, new_n29739_ );
and  ( new_n29745_, new_n29744_, new_n29738_ );
or   ( new_n29746_, new_n29745_, new_n29729_ );
and  ( new_n29747_, new_n29745_, new_n29729_ );
or   ( new_n29748_, new_n1364_, new_n24925_ );
or   ( new_n29749_, new_n1366_, new_n24927_ );
and  ( new_n29750_, new_n29749_, new_n29748_ );
xor  ( new_n29751_, new_n29750_, new_n1129_ );
or   ( new_n29752_, new_n1135_, new_n25288_ );
or   ( new_n29753_, new_n1137_, new_n25048_ );
and  ( new_n29754_, new_n29753_, new_n29752_ );
xor  ( new_n29755_, new_n29754_, new_n896_ );
nor  ( new_n29756_, new_n29755_, new_n29751_ );
and  ( new_n29757_, new_n29755_, new_n29751_ );
or   ( new_n29758_, new_n897_, new_n25813_ );
or   ( new_n29759_, new_n899_, new_n25486_ );
and  ( new_n29760_, new_n29759_, new_n29758_ );
xor  ( new_n29761_, new_n29760_, new_n748_ );
nor  ( new_n29762_, new_n29761_, new_n29757_ );
nor  ( new_n29763_, new_n29762_, new_n29756_ );
or   ( new_n29764_, new_n29763_, new_n29747_ );
and  ( new_n29765_, new_n29764_, new_n29746_ );
or   ( new_n29766_, new_n29765_, new_n29713_ );
or   ( new_n29767_, new_n5604_, new_n21842_ );
or   ( new_n29768_, new_n5606_, new_n21792_ );
and  ( new_n29769_, new_n29768_, new_n29767_ );
xor  ( new_n29770_, new_n29769_, new_n5206_ );
or   ( new_n29771_, new_n5207_, new_n21847_ );
or   ( new_n29772_, new_n5209_, new_n21840_ );
and  ( new_n29773_, new_n29772_, new_n29771_ );
xor  ( new_n29774_, new_n29773_, new_n4708_ );
or   ( new_n29775_, new_n29774_, new_n29770_ );
and  ( new_n29776_, new_n29774_, new_n29770_ );
or   ( new_n29777_, new_n4709_, new_n22129_ );
or   ( new_n29778_, new_n4711_, new_n22098_ );
and  ( new_n29779_, new_n29778_, new_n29777_ );
xor  ( new_n29780_, new_n29779_, new_n4295_ );
or   ( new_n29781_, new_n29780_, new_n29776_ );
and  ( new_n29782_, new_n29781_, new_n29775_ );
or   ( new_n29783_, new_n8264_, new_n21703_ );
or   ( new_n29784_, new_n8266_, new_n21694_ );
and  ( new_n29785_, new_n29784_, new_n29783_ );
xor  ( new_n29786_, new_n29785_, new_n7724_ );
and  ( new_n29787_, new_n8651_, RIbb315f0_129 );
xor  ( new_n29788_, new_n29787_, new_n8257_ );
nand ( new_n29789_, new_n29788_, new_n29786_ );
nor  ( new_n29790_, new_n29788_, new_n29786_ );
or   ( new_n29791_, new_n7732_, new_n21674_ );
or   ( new_n29792_, new_n7734_, new_n21701_ );
and  ( new_n29793_, new_n29792_, new_n29791_ );
xor  ( new_n29794_, new_n29793_, new_n7177_ );
or   ( new_n29795_, new_n29794_, new_n29790_ );
and  ( new_n29796_, new_n29795_, new_n29789_ );
or   ( new_n29797_, new_n29796_, new_n29782_ );
and  ( new_n29798_, new_n29796_, new_n29782_ );
or   ( new_n29799_, new_n7184_, new_n21680_ );
or   ( new_n29800_, new_n7186_, new_n21672_ );
and  ( new_n29801_, new_n29800_, new_n29799_ );
xor  ( new_n29802_, new_n29801_, new_n6638_ );
or   ( new_n29803_, new_n6645_, new_n21687_ );
or   ( new_n29804_, new_n6647_, new_n21678_ );
and  ( new_n29805_, new_n29804_, new_n29803_ );
xor  ( new_n29806_, new_n29805_, new_n6166_ );
nor  ( new_n29807_, new_n29806_, new_n29802_ );
and  ( new_n29808_, new_n29806_, new_n29802_ );
or   ( new_n29809_, new_n6173_, new_n21751_ );
or   ( new_n29810_, new_n6175_, new_n21685_ );
and  ( new_n29811_, new_n29810_, new_n29809_ );
xor  ( new_n29812_, new_n29811_, new_n5597_ );
nor  ( new_n29813_, new_n29812_, new_n29808_ );
nor  ( new_n29814_, new_n29813_, new_n29807_ );
or   ( new_n29815_, new_n29814_, new_n29798_ );
and  ( new_n29816_, new_n29815_, new_n29797_ );
and  ( new_n29817_, new_n29765_, new_n29713_ );
or   ( new_n29818_, new_n29817_, new_n29816_ );
and  ( new_n29819_, new_n29818_, new_n29766_ );
or   ( new_n29820_, new_n29819_, new_n29661_ );
nand ( new_n29821_, new_n29819_, new_n29661_ );
xnor ( new_n29822_, new_n29190_, new_n29188_ );
xor  ( new_n29823_, new_n29822_, new_n29196_ );
xnor ( new_n29824_, new_n29224_, new_n29220_ );
xor  ( new_n29825_, new_n29824_, new_n29230_ );
nor  ( new_n29826_, new_n29825_, new_n29823_ );
and  ( new_n29827_, new_n29825_, new_n29823_ );
xor  ( new_n29828_, new_n29495_, new_n29493_ );
xnor ( new_n29829_, new_n29828_, new_n29499_ );
not  ( new_n29830_, new_n29829_ );
nor  ( new_n29831_, new_n29830_, new_n29827_ );
nor  ( new_n29832_, new_n29831_, new_n29826_ );
nand ( new_n29833_, new_n29832_, new_n29821_ );
and  ( new_n29834_, new_n29833_, new_n29820_ );
or   ( new_n29835_, new_n29834_, new_n29614_ );
nand ( new_n29836_, new_n29834_, new_n29614_ );
xor  ( new_n29837_, new_n29413_, new_n29365_ );
xor  ( new_n29838_, new_n29837_, new_n29467_ );
xnor ( new_n29839_, new_n29501_, new_n29491_ );
xor  ( new_n29840_, new_n29839_, new_n29513_ );
and  ( new_n29841_, new_n29840_, new_n29838_ );
nor  ( new_n29842_, new_n29840_, new_n29838_ );
xor  ( new_n29843_, new_n29521_, new_n29519_ );
xor  ( new_n29844_, new_n29843_, new_n29526_ );
nor  ( new_n29845_, new_n29844_, new_n29842_ );
nor  ( new_n29846_, new_n29845_, new_n29841_ );
nand ( new_n29847_, new_n29846_, new_n29836_ );
and  ( new_n29848_, new_n29847_, new_n29835_ );
or   ( new_n29849_, new_n29848_, new_n29596_ );
nand ( new_n29850_, new_n29848_, new_n29596_ );
xor  ( new_n29851_, new_n29515_, new_n29469_ );
xor  ( new_n29852_, new_n29851_, new_n29528_ );
xor  ( new_n29853_, new_n29534_, new_n29532_ );
xor  ( new_n29854_, new_n29853_, new_n29538_ );
nor  ( new_n29855_, new_n29854_, new_n29852_ );
and  ( new_n29856_, new_n29854_, new_n29852_ );
xor  ( new_n29857_, new_n29546_, new_n29544_ );
xnor ( new_n29858_, new_n29857_, new_n29558_ );
not  ( new_n29859_, new_n29858_ );
nor  ( new_n29860_, new_n29859_, new_n29856_ );
nor  ( new_n29861_, new_n29860_, new_n29855_ );
nand ( new_n29862_, new_n29861_, new_n29850_ );
and  ( new_n29863_, new_n29862_, new_n29849_ );
and  ( new_n29864_, new_n29863_, new_n29594_ );
nor  ( new_n29865_, new_n29863_, new_n29594_ );
xor  ( new_n29866_, new_n29282_, new_n29061_ );
xor  ( new_n29867_, new_n29866_, new_n29294_ );
nor  ( new_n29868_, new_n29867_, new_n29865_ );
nor  ( new_n29869_, new_n29868_, new_n29864_ );
xnor ( new_n29870_, new_n29580_, new_n29578_ );
xor  ( new_n29871_, new_n29870_, new_n29584_ );
nor  ( new_n29872_, new_n29871_, new_n29869_ );
xor  ( new_n29873_, new_n29586_, new_n29313_ );
and  ( new_n29874_, new_n29873_, new_n29872_ );
xnor ( new_n29875_, new_n29871_, new_n29869_ );
xor  ( new_n29876_, new_n29863_, new_n29594_ );
xor  ( new_n29877_, new_n29876_, new_n29867_ );
xor  ( new_n29878_, new_n29854_, new_n29852_ );
xor  ( new_n29879_, new_n29878_, new_n29859_ );
xor  ( new_n29880_, new_n29819_, new_n29661_ );
xor  ( new_n29881_, new_n29880_, new_n29832_ );
xnor ( new_n29882_, new_n29608_, new_n29598_ );
xor  ( new_n29883_, new_n29882_, new_n29612_ );
or   ( new_n29884_, new_n29883_, new_n29881_ );
nand ( new_n29885_, new_n29883_, new_n29881_ );
xor  ( new_n29886_, new_n29840_, new_n29838_ );
xnor ( new_n29887_, new_n29886_, new_n29844_ );
nand ( new_n29888_, new_n29887_, new_n29885_ );
and  ( new_n29889_, new_n29888_, new_n29884_ );
or   ( new_n29890_, new_n29889_, new_n29879_ );
and  ( new_n29891_, new_n29889_, new_n29879_ );
xnor ( new_n29892_, new_n29641_, new_n29639_ );
xor  ( new_n29893_, new_n29892_, new_n29645_ );
xor  ( new_n29894_, new_n29653_, new_n29651_ );
xor  ( new_n29895_, new_n29894_, new_n29657_ );
nor  ( new_n29896_, new_n29895_, new_n29893_ );
and  ( new_n29897_, new_n29895_, new_n29893_ );
xor  ( new_n29898_, new_n29631_, new_n29629_ );
xnor ( new_n29899_, new_n29898_, new_n29635_ );
nor  ( new_n29900_, new_n29899_, new_n29897_ );
or   ( new_n29901_, new_n29900_, new_n29896_ );
xnor ( new_n29902_, new_n29447_, new_n29431_ );
xor  ( new_n29903_, new_n29902_, new_n29465_ );
or   ( new_n29904_, new_n29903_, new_n29901_ );
and  ( new_n29905_, new_n29903_, new_n29901_ );
xnor ( new_n29906_, new_n29693_, new_n29677_ );
xor  ( new_n29907_, new_n29906_, new_n29711_ );
xnor ( new_n29908_, new_n29745_, new_n29729_ );
xor  ( new_n29909_, new_n29908_, new_n29763_ );
nor  ( new_n29910_, new_n29909_, new_n29907_ );
and  ( new_n29911_, new_n29909_, new_n29907_ );
xor  ( new_n29912_, new_n29796_, new_n29782_ );
xnor ( new_n29913_, new_n29912_, new_n29814_ );
nor  ( new_n29914_, new_n29913_, new_n29911_ );
nor  ( new_n29915_, new_n29914_, new_n29910_ );
or   ( new_n29916_, new_n29915_, new_n29905_ );
and  ( new_n29917_, new_n29916_, new_n29904_ );
xnor ( new_n29918_, new_n29393_, new_n29381_ );
xor  ( new_n29919_, new_n29918_, new_n29411_ );
xor  ( new_n29920_, new_n29825_, new_n29823_ );
xor  ( new_n29921_, new_n29920_, new_n29830_ );
or   ( new_n29922_, new_n29921_, new_n29919_ );
and  ( new_n29923_, new_n29921_, new_n29919_ );
xor  ( new_n29924_, new_n29602_, new_n29600_ );
xnor ( new_n29925_, new_n29924_, new_n29606_ );
not  ( new_n29926_, new_n29925_ );
or   ( new_n29927_, new_n29926_, new_n29923_ );
and  ( new_n29928_, new_n29927_, new_n29922_ );
nor  ( new_n29929_, new_n29928_, new_n29917_ );
and  ( new_n29930_, new_n29928_, new_n29917_ );
xor  ( new_n29931_, new_n29373_, new_n29369_ );
xor  ( new_n29932_, new_n29931_, new_n29379_ );
xnor ( new_n29933_, new_n29788_, new_n29786_ );
xor  ( new_n29934_, new_n29933_, new_n29794_ );
xnor ( new_n29935_, new_n29774_, new_n29770_ );
xor  ( new_n29936_, new_n29935_, new_n29780_ );
or   ( new_n29937_, new_n29936_, new_n29934_ );
and  ( new_n29938_, new_n29936_, new_n29934_ );
xnor ( new_n29939_, new_n29806_, new_n29802_ );
xor  ( new_n29940_, new_n29939_, new_n29812_ );
or   ( new_n29941_, new_n29940_, new_n29938_ );
and  ( new_n29942_, new_n29941_, new_n29937_ );
nor  ( new_n29943_, new_n29942_, new_n29932_ );
nand ( new_n29944_, new_n29942_, new_n29932_ );
xor  ( new_n29945_, new_n29385_, new_n8257_ );
xor  ( new_n29946_, new_n29945_, new_n29391_ );
and  ( new_n29947_, new_n29946_, new_n29944_ );
or   ( new_n29948_, new_n29947_, new_n29943_ );
or   ( new_n29949_, new_n2425_, new_n23733_ );
or   ( new_n29950_, new_n2427_, new_n23554_ );
and  ( new_n29951_, new_n29950_, new_n29949_ );
xor  ( new_n29952_, new_n29951_, new_n2121_ );
or   ( new_n29953_, new_n2122_, new_n24006_ );
or   ( new_n29954_, new_n2124_, new_n23895_ );
and  ( new_n29955_, new_n29954_, new_n29953_ );
xor  ( new_n29956_, new_n29955_, new_n1843_ );
or   ( new_n29957_, new_n29956_, new_n29952_ );
and  ( new_n29958_, new_n29956_, new_n29952_ );
or   ( new_n29959_, new_n1844_, new_n24418_ );
or   ( new_n29960_, new_n1846_, new_n24227_ );
and  ( new_n29961_, new_n29960_, new_n29959_ );
xor  ( new_n29962_, new_n29961_, new_n1586_ );
or   ( new_n29963_, new_n29962_, new_n29958_ );
and  ( new_n29964_, new_n29963_, new_n29957_ );
or   ( new_n29965_, new_n3461_, new_n22975_ );
or   ( new_n29966_, new_n3463_, new_n22829_ );
and  ( new_n29967_, new_n29966_, new_n29965_ );
xor  ( new_n29968_, new_n29967_, new_n3116_ );
or   ( new_n29969_, new_n3117_, new_n23166_ );
or   ( new_n29970_, new_n3119_, new_n22973_ );
and  ( new_n29971_, new_n29970_, new_n29969_ );
xor  ( new_n29972_, new_n29971_, new_n2800_ );
or   ( new_n29973_, new_n29972_, new_n29968_ );
and  ( new_n29974_, new_n29972_, new_n29968_ );
or   ( new_n29975_, new_n2807_, new_n23370_ );
or   ( new_n29976_, new_n2809_, new_n23252_ );
and  ( new_n29977_, new_n29976_, new_n29975_ );
xor  ( new_n29978_, new_n29977_, new_n2424_ );
or   ( new_n29979_, new_n29978_, new_n29974_ );
and  ( new_n29980_, new_n29979_, new_n29973_ );
or   ( new_n29981_, new_n29980_, new_n29964_ );
and  ( new_n29982_, new_n29980_, new_n29964_ );
or   ( new_n29983_, new_n4709_, new_n22207_ );
or   ( new_n29984_, new_n4711_, new_n22129_ );
and  ( new_n29985_, new_n29984_, new_n29983_ );
xor  ( new_n29986_, new_n29985_, new_n4295_ );
or   ( new_n29987_, new_n4302_, new_n22423_ );
or   ( new_n29988_, new_n4304_, new_n22304_ );
and  ( new_n29989_, new_n29988_, new_n29987_ );
xor  ( new_n29990_, new_n29989_, new_n3895_ );
nor  ( new_n29991_, new_n29990_, new_n29986_ );
and  ( new_n29992_, new_n29990_, new_n29986_ );
or   ( new_n29993_, new_n3896_, new_n22641_ );
or   ( new_n29994_, new_n3898_, new_n22590_ );
and  ( new_n29995_, new_n29994_, new_n29993_ );
xor  ( new_n29996_, new_n29995_, new_n3460_ );
nor  ( new_n29997_, new_n29996_, new_n29992_ );
nor  ( new_n29998_, new_n29997_, new_n29991_ );
or   ( new_n29999_, new_n29998_, new_n29982_ );
and  ( new_n30000_, new_n29999_, new_n29981_ );
or   ( new_n30001_, new_n8874_, new_n21694_ );
or   ( new_n30002_, new_n8876_, new_n21696_ );
and  ( new_n30003_, new_n30002_, new_n30001_ );
xor  ( new_n30004_, new_n30003_, new_n8257_ );
and  ( new_n30005_, new_n30004_, new_n8873_ );
or   ( new_n30006_, new_n30004_, new_n8873_ );
or   ( new_n30007_, new_n8264_, new_n21701_ );
or   ( new_n30008_, new_n8266_, new_n21703_ );
and  ( new_n30009_, new_n30008_, new_n30007_ );
xor  ( new_n30010_, new_n30009_, new_n7725_ );
and  ( new_n30011_, new_n30010_, new_n30006_ );
or   ( new_n30012_, new_n30011_, new_n30005_ );
or   ( new_n30013_, new_n6173_, new_n21792_ );
or   ( new_n30014_, new_n6175_, new_n21751_ );
and  ( new_n30015_, new_n30014_, new_n30013_ );
xor  ( new_n30016_, new_n30015_, new_n5597_ );
or   ( new_n30017_, new_n5604_, new_n21840_ );
or   ( new_n30018_, new_n5606_, new_n21842_ );
and  ( new_n30019_, new_n30018_, new_n30017_ );
xor  ( new_n30020_, new_n30019_, new_n5206_ );
or   ( new_n30021_, new_n30020_, new_n30016_ );
and  ( new_n30022_, new_n30020_, new_n30016_ );
or   ( new_n30023_, new_n5207_, new_n22098_ );
or   ( new_n30024_, new_n5209_, new_n21847_ );
and  ( new_n30025_, new_n30024_, new_n30023_ );
xor  ( new_n30026_, new_n30025_, new_n4708_ );
or   ( new_n30027_, new_n30026_, new_n30022_ );
and  ( new_n30028_, new_n30027_, new_n30021_ );
or   ( new_n30029_, new_n30028_, new_n30012_ );
and  ( new_n30030_, new_n30028_, new_n30012_ );
or   ( new_n30031_, new_n7732_, new_n21672_ );
or   ( new_n30032_, new_n7734_, new_n21674_ );
and  ( new_n30033_, new_n30032_, new_n30031_ );
xor  ( new_n30034_, new_n30033_, new_n7177_ );
or   ( new_n30035_, new_n7184_, new_n21678_ );
or   ( new_n30036_, new_n7186_, new_n21680_ );
and  ( new_n30037_, new_n30036_, new_n30035_ );
xor  ( new_n30038_, new_n30037_, new_n6638_ );
nor  ( new_n30039_, new_n30038_, new_n30034_ );
and  ( new_n30040_, new_n30038_, new_n30034_ );
or   ( new_n30041_, new_n6645_, new_n21685_ );
or   ( new_n30042_, new_n6647_, new_n21687_ );
and  ( new_n30043_, new_n30042_, new_n30041_ );
xor  ( new_n30044_, new_n30043_, new_n6166_ );
nor  ( new_n30045_, new_n30044_, new_n30040_ );
nor  ( new_n30046_, new_n30045_, new_n30039_ );
or   ( new_n30047_, new_n30046_, new_n30030_ );
and  ( new_n30048_, new_n30047_, new_n30029_ );
or   ( new_n30049_, new_n30048_, new_n30000_ );
or   ( new_n30050_, new_n897_, new_n26196_ );
or   ( new_n30051_, new_n899_, new_n25813_ );
and  ( new_n30052_, new_n30051_, new_n30050_ );
xor  ( new_n30053_, new_n30052_, new_n748_ );
or   ( new_n30054_, new_n755_, new_n26372_ );
or   ( new_n30055_, new_n757_, new_n26063_ );
and  ( new_n30056_, new_n30055_, new_n30054_ );
xor  ( new_n30057_, new_n30056_, new_n523_ );
or   ( new_n30058_, new_n30057_, new_n30053_ );
and  ( new_n30059_, new_n30057_, new_n30053_ );
or   ( new_n30060_, new_n524_, new_n26762_ );
or   ( new_n30061_, new_n526_, new_n26620_ );
and  ( new_n30062_, new_n30061_, new_n30060_ );
xor  ( new_n30063_, new_n30062_, new_n403_ );
or   ( new_n30064_, new_n30063_, new_n30059_ );
and  ( new_n30065_, new_n30064_, new_n30058_ );
or   ( new_n30066_, new_n409_, new_n27396_ );
or   ( new_n30067_, new_n411_, new_n27085_ );
and  ( new_n30068_, new_n30067_, new_n30066_ );
xor  ( new_n30069_, new_n30068_, new_n328_ );
or   ( new_n30070_, new_n337_, new_n27763_ );
or   ( new_n30071_, new_n340_, new_n27602_ );
and  ( new_n30072_, new_n30071_, new_n30070_ );
xor  ( new_n30073_, new_n30072_, new_n332_ );
or   ( new_n30074_, new_n30073_, new_n30069_ );
and  ( new_n30075_, new_n30073_, new_n30069_ );
or   ( new_n30076_, new_n317_, new_n28314_ );
or   ( new_n30077_, new_n320_, new_n28108_ );
and  ( new_n30078_, new_n30077_, new_n30076_ );
xor  ( new_n30079_, new_n30078_, new_n312_ );
or   ( new_n30080_, new_n30079_, new_n30075_ );
and  ( new_n30081_, new_n30080_, new_n30074_ );
nor  ( new_n30082_, new_n30081_, new_n30065_ );
and  ( new_n30083_, new_n30081_, new_n30065_ );
or   ( new_n30084_, new_n1593_, new_n24927_ );
or   ( new_n30085_, new_n1595_, new_n24543_ );
and  ( new_n30086_, new_n30085_, new_n30084_ );
xor  ( new_n30087_, new_n30086_, new_n1358_ );
or   ( new_n30088_, new_n1364_, new_n25048_ );
or   ( new_n30089_, new_n1366_, new_n24925_ );
and  ( new_n30090_, new_n30089_, new_n30088_ );
xor  ( new_n30091_, new_n30090_, new_n1129_ );
nor  ( new_n30092_, new_n30091_, new_n30087_ );
and  ( new_n30093_, new_n30091_, new_n30087_ );
or   ( new_n30094_, new_n1135_, new_n25486_ );
or   ( new_n30095_, new_n1137_, new_n25288_ );
and  ( new_n30096_, new_n30095_, new_n30094_ );
xor  ( new_n30097_, new_n30096_, new_n896_ );
nor  ( new_n30098_, new_n30097_, new_n30093_ );
nor  ( new_n30099_, new_n30098_, new_n30092_ );
nor  ( new_n30100_, new_n30099_, new_n30083_ );
nor  ( new_n30101_, new_n30100_, new_n30082_ );
and  ( new_n30102_, new_n30048_, new_n30000_ );
or   ( new_n30103_, new_n30102_, new_n30101_ );
and  ( new_n30104_, new_n30103_, new_n30049_ );
and  ( new_n30105_, new_n30104_, new_n29948_ );
nor  ( new_n30106_, new_n30104_, new_n29948_ );
xor  ( new_n30107_, new_n29623_, new_n29618_ );
xor  ( new_n30108_, new_n30107_, new_n29626_ );
not  ( new_n30109_, new_n30108_ );
or   ( new_n30110_, new_n283_, new_n29263_ );
or   ( new_n30111_, new_n286_, new_n28531_ );
and  ( new_n30112_, new_n30111_, new_n30110_ );
xor  ( new_n30113_, new_n30112_, new_n278_ );
or   ( new_n30114_, new_n299_, new_n29474_ );
or   ( new_n30115_, new_n302_, new_n29261_ );
and  ( new_n30116_, new_n30115_, new_n30114_ );
xor  ( new_n30117_, new_n30116_, new_n293_ );
or   ( new_n30118_, new_n30117_, new_n30113_ );
and  ( new_n30119_, new_n30117_, new_n30113_ );
not  ( new_n30120_, RIbb330a8_186 );
or   ( new_n30121_, new_n268_, new_n30120_ );
or   ( new_n30122_, new_n271_, new_n29619_ );
and  ( new_n30123_, new_n30122_, new_n30121_ );
xor  ( new_n30124_, new_n30123_, new_n263_ );
or   ( new_n30125_, new_n30124_, new_n30119_ );
and  ( new_n30126_, new_n30125_, new_n30118_ );
nor  ( new_n30127_, new_n30126_, new_n30109_ );
xnor ( new_n30128_, new_n29685_, new_n29681_ );
xor  ( new_n30129_, new_n30128_, new_n29691_ );
xnor ( new_n30130_, new_n29669_, new_n29665_ );
xor  ( new_n30131_, new_n30130_, new_n29675_ );
or   ( new_n30132_, new_n30131_, new_n30129_ );
and  ( new_n30133_, new_n30131_, new_n30129_ );
xor  ( new_n30134_, new_n29703_, new_n29699_ );
xnor ( new_n30135_, new_n30134_, new_n29709_ );
or   ( new_n30136_, new_n30135_, new_n30133_ );
and  ( new_n30137_, new_n30136_, new_n30132_ );
nor  ( new_n30138_, new_n30137_, new_n30127_ );
and  ( new_n30139_, new_n30137_, new_n30127_ );
xnor ( new_n30140_, new_n29737_, new_n29733_ );
xor  ( new_n30141_, new_n30140_, new_n29743_ );
xnor ( new_n30142_, new_n29721_, new_n29717_ );
xor  ( new_n30143_, new_n30142_, new_n29727_ );
nor  ( new_n30144_, new_n30143_, new_n30141_ );
and  ( new_n30145_, new_n30143_, new_n30141_ );
xor  ( new_n30146_, new_n29755_, new_n29751_ );
xnor ( new_n30147_, new_n30146_, new_n29761_ );
nor  ( new_n30148_, new_n30147_, new_n30145_ );
nor  ( new_n30149_, new_n30148_, new_n30144_ );
nor  ( new_n30150_, new_n30149_, new_n30139_ );
nor  ( new_n30151_, new_n30150_, new_n30138_ );
nor  ( new_n30152_, new_n30151_, new_n30106_ );
nor  ( new_n30153_, new_n30152_, new_n30105_ );
nor  ( new_n30154_, new_n30153_, new_n29930_ );
nor  ( new_n30155_, new_n30154_, new_n29929_ );
or   ( new_n30156_, new_n30155_, new_n29891_ );
and  ( new_n30157_, new_n30156_, new_n29890_ );
xor  ( new_n30158_, new_n29848_, new_n29596_ );
xor  ( new_n30159_, new_n30158_, new_n29861_ );
or   ( new_n30160_, new_n30159_, new_n30157_ );
and  ( new_n30161_, new_n30159_, new_n30157_ );
xnor ( new_n30162_, new_n29593_, new_n29591_ );
or   ( new_n30163_, new_n30162_, new_n30161_ );
and  ( new_n30164_, new_n30163_, new_n30160_ );
or   ( new_n30165_, new_n30164_, new_n29877_ );
nand ( new_n30166_, new_n30164_, new_n29877_ );
xor  ( new_n30167_, new_n29572_, new_n29562_ );
xnor ( new_n30168_, new_n30167_, new_n29576_ );
nand ( new_n30169_, new_n30168_, new_n30166_ );
and  ( new_n30170_, new_n30169_, new_n30165_ );
nor  ( new_n30171_, new_n30170_, new_n29875_ );
xor  ( new_n30172_, new_n30159_, new_n30157_ );
xor  ( new_n30173_, new_n30172_, new_n30162_ );
xor  ( new_n30174_, new_n29883_, new_n29881_ );
xor  ( new_n30175_, new_n30174_, new_n29887_ );
xor  ( new_n30176_, new_n29895_, new_n29893_ );
xor  ( new_n30177_, new_n30176_, new_n29899_ );
xnor ( new_n30178_, new_n29909_, new_n29907_ );
xor  ( new_n30179_, new_n30178_, new_n29913_ );
and  ( new_n30180_, new_n30179_, new_n30177_ );
or   ( new_n30181_, new_n30179_, new_n30177_ );
xor  ( new_n30182_, new_n30081_, new_n30065_ );
xor  ( new_n30183_, new_n30182_, new_n30099_ );
xnor ( new_n30184_, new_n30143_, new_n30141_ );
xor  ( new_n30185_, new_n30184_, new_n30147_ );
and  ( new_n30186_, new_n30185_, new_n30183_ );
nor  ( new_n30187_, new_n30185_, new_n30183_ );
xor  ( new_n30188_, new_n30126_, new_n30109_ );
nor  ( new_n30189_, new_n30188_, new_n30187_ );
nor  ( new_n30190_, new_n30189_, new_n30186_ );
not  ( new_n30191_, new_n30190_ );
and  ( new_n30192_, new_n30191_, new_n30181_ );
or   ( new_n30193_, new_n30192_, new_n30180_ );
xnor ( new_n30194_, new_n30117_, new_n30113_ );
xor  ( new_n30195_, new_n30194_, new_n30124_ );
xnor ( new_n30196_, new_n30073_, new_n30069_ );
xor  ( new_n30197_, new_n30196_, new_n30079_ );
or   ( new_n30198_, new_n30197_, new_n30195_ );
and  ( new_n30199_, new_n30197_, new_n30195_ );
xor  ( new_n30200_, new_n30057_, new_n30053_ );
xnor ( new_n30201_, new_n30200_, new_n30063_ );
or   ( new_n30202_, new_n30201_, new_n30199_ );
and  ( new_n30203_, new_n30202_, new_n30198_ );
xnor ( new_n30204_, new_n30091_, new_n30087_ );
xor  ( new_n30205_, new_n30204_, new_n30097_ );
xnor ( new_n30206_, new_n29972_, new_n29968_ );
xor  ( new_n30207_, new_n30206_, new_n29978_ );
or   ( new_n30208_, new_n30207_, new_n30205_ );
and  ( new_n30209_, new_n30207_, new_n30205_ );
xor  ( new_n30210_, new_n29956_, new_n29952_ );
xnor ( new_n30211_, new_n30210_, new_n29962_ );
or   ( new_n30212_, new_n30211_, new_n30209_ );
and  ( new_n30213_, new_n30212_, new_n30208_ );
nor  ( new_n30214_, new_n30213_, new_n30203_ );
nand ( new_n30215_, new_n30213_, new_n30203_ );
and  ( new_n30216_, RIbb33198_188, RIbb2f610_1 );
or   ( new_n30217_, new_n283_, new_n29261_ );
or   ( new_n30218_, new_n286_, new_n29263_ );
and  ( new_n30219_, new_n30218_, new_n30217_ );
xor  ( new_n30220_, new_n30219_, new_n278_ );
or   ( new_n30221_, new_n299_, new_n29619_ );
or   ( new_n30222_, new_n302_, new_n29474_ );
and  ( new_n30223_, new_n30222_, new_n30221_ );
xor  ( new_n30224_, new_n30223_, new_n293_ );
or   ( new_n30225_, new_n30224_, new_n30220_ );
and  ( new_n30226_, new_n30224_, new_n30220_ );
not  ( new_n30227_, RIbb33120_187 );
or   ( new_n30228_, new_n268_, new_n30227_ );
or   ( new_n30229_, new_n271_, new_n30120_ );
and  ( new_n30230_, new_n30229_, new_n30228_ );
xor  ( new_n30231_, new_n30230_, new_n263_ );
or   ( new_n30232_, new_n30231_, new_n30226_ );
and  ( new_n30233_, new_n30232_, new_n30225_ );
nor  ( new_n30234_, new_n30233_, new_n30216_ );
and  ( new_n30235_, new_n30233_, new_n30216_ );
and  ( new_n30236_, RIbb33120_187, RIbb2f610_1 );
nor  ( new_n30237_, new_n30236_, new_n30235_ );
nor  ( new_n30238_, new_n30237_, new_n30234_ );
and  ( new_n30239_, new_n30238_, new_n30215_ );
or   ( new_n30240_, new_n30239_, new_n30214_ );
or   ( new_n30241_, new_n1593_, new_n24925_ );
or   ( new_n30242_, new_n1595_, new_n24927_ );
and  ( new_n30243_, new_n30242_, new_n30241_ );
xor  ( new_n30244_, new_n30243_, new_n1358_ );
or   ( new_n30245_, new_n1364_, new_n25288_ );
or   ( new_n30246_, new_n1366_, new_n25048_ );
and  ( new_n30247_, new_n30246_, new_n30245_ );
xor  ( new_n30248_, new_n30247_, new_n1129_ );
or   ( new_n30249_, new_n30248_, new_n30244_ );
and  ( new_n30250_, new_n30248_, new_n30244_ );
or   ( new_n30251_, new_n1135_, new_n25813_ );
or   ( new_n30252_, new_n1137_, new_n25486_ );
and  ( new_n30253_, new_n30252_, new_n30251_ );
xor  ( new_n30254_, new_n30253_, new_n896_ );
or   ( new_n30255_, new_n30254_, new_n30250_ );
and  ( new_n30256_, new_n30255_, new_n30249_ );
or   ( new_n30257_, new_n897_, new_n26063_ );
or   ( new_n30258_, new_n899_, new_n26196_ );
and  ( new_n30259_, new_n30258_, new_n30257_ );
xor  ( new_n30260_, new_n30259_, new_n748_ );
or   ( new_n30261_, new_n755_, new_n26620_ );
or   ( new_n30262_, new_n757_, new_n26372_ );
and  ( new_n30263_, new_n30262_, new_n30261_ );
xor  ( new_n30264_, new_n30263_, new_n523_ );
or   ( new_n30265_, new_n30264_, new_n30260_ );
and  ( new_n30266_, new_n30264_, new_n30260_ );
or   ( new_n30267_, new_n524_, new_n27085_ );
or   ( new_n30268_, new_n526_, new_n26762_ );
and  ( new_n30269_, new_n30268_, new_n30267_ );
xor  ( new_n30270_, new_n30269_, new_n403_ );
or   ( new_n30271_, new_n30270_, new_n30266_ );
and  ( new_n30272_, new_n30271_, new_n30265_ );
or   ( new_n30273_, new_n30272_, new_n30256_ );
and  ( new_n30274_, new_n30272_, new_n30256_ );
or   ( new_n30275_, new_n409_, new_n27602_ );
or   ( new_n30276_, new_n411_, new_n27396_ );
and  ( new_n30277_, new_n30276_, new_n30275_ );
xor  ( new_n30278_, new_n30277_, new_n328_ );
or   ( new_n30279_, new_n337_, new_n28108_ );
or   ( new_n30280_, new_n340_, new_n27763_ );
and  ( new_n30281_, new_n30280_, new_n30279_ );
xor  ( new_n30282_, new_n30281_, new_n332_ );
nor  ( new_n30283_, new_n30282_, new_n30278_ );
and  ( new_n30284_, new_n30282_, new_n30278_ );
or   ( new_n30285_, new_n317_, new_n28531_ );
or   ( new_n30286_, new_n320_, new_n28314_ );
and  ( new_n30287_, new_n30286_, new_n30285_ );
xor  ( new_n30288_, new_n30287_, new_n312_ );
nor  ( new_n30289_, new_n30288_, new_n30284_ );
nor  ( new_n30290_, new_n30289_, new_n30283_ );
or   ( new_n30291_, new_n30290_, new_n30274_ );
and  ( new_n30292_, new_n30291_, new_n30273_ );
or   ( new_n30293_, new_n6173_, new_n21842_ );
or   ( new_n30294_, new_n6175_, new_n21792_ );
and  ( new_n30295_, new_n30294_, new_n30293_ );
xor  ( new_n30296_, new_n30295_, new_n5597_ );
or   ( new_n30297_, new_n5604_, new_n21847_ );
or   ( new_n30298_, new_n5606_, new_n21840_ );
and  ( new_n30299_, new_n30298_, new_n30297_ );
xor  ( new_n30300_, new_n30299_, new_n5206_ );
or   ( new_n30301_, new_n30300_, new_n30296_ );
and  ( new_n30302_, new_n30300_, new_n30296_ );
or   ( new_n30303_, new_n5207_, new_n22129_ );
or   ( new_n30304_, new_n5209_, new_n22098_ );
and  ( new_n30305_, new_n30304_, new_n30303_ );
xor  ( new_n30306_, new_n30305_, new_n4708_ );
or   ( new_n30307_, new_n30306_, new_n30302_ );
and  ( new_n30308_, new_n30307_, new_n30301_ );
or   ( new_n30309_, new_n8874_, new_n21703_ );
or   ( new_n30310_, new_n8876_, new_n21694_ );
and  ( new_n30311_, new_n30310_, new_n30309_ );
xor  ( new_n30312_, new_n30311_, new_n8256_ );
and  ( new_n30313_, new_n9187_, RIbb315f0_129 );
xor  ( new_n30314_, new_n30313_, new_n8873_ );
nand ( new_n30315_, new_n30314_, new_n30312_ );
nor  ( new_n30316_, new_n30314_, new_n30312_ );
or   ( new_n30317_, new_n8264_, new_n21674_ );
or   ( new_n30318_, new_n8266_, new_n21701_ );
and  ( new_n30319_, new_n30318_, new_n30317_ );
xor  ( new_n30320_, new_n30319_, new_n7725_ );
or   ( new_n30321_, new_n30320_, new_n30316_ );
and  ( new_n30322_, new_n30321_, new_n30315_ );
or   ( new_n30323_, new_n30322_, new_n30308_ );
and  ( new_n30324_, new_n30322_, new_n30308_ );
or   ( new_n30325_, new_n7732_, new_n21680_ );
or   ( new_n30326_, new_n7734_, new_n21672_ );
and  ( new_n30327_, new_n30326_, new_n30325_ );
xor  ( new_n30328_, new_n30327_, new_n7177_ );
or   ( new_n30329_, new_n7184_, new_n21687_ );
or   ( new_n30330_, new_n7186_, new_n21678_ );
and  ( new_n30331_, new_n30330_, new_n30329_ );
xor  ( new_n30332_, new_n30331_, new_n6638_ );
nor  ( new_n30333_, new_n30332_, new_n30328_ );
and  ( new_n30334_, new_n30332_, new_n30328_ );
or   ( new_n30335_, new_n6645_, new_n21751_ );
or   ( new_n30336_, new_n6647_, new_n21685_ );
and  ( new_n30337_, new_n30336_, new_n30335_ );
xor  ( new_n30338_, new_n30337_, new_n6166_ );
nor  ( new_n30339_, new_n30338_, new_n30334_ );
nor  ( new_n30340_, new_n30339_, new_n30333_ );
or   ( new_n30341_, new_n30340_, new_n30324_ );
and  ( new_n30342_, new_n30341_, new_n30323_ );
or   ( new_n30343_, new_n30342_, new_n30292_ );
or   ( new_n30344_, new_n2425_, new_n23895_ );
or   ( new_n30345_, new_n2427_, new_n23733_ );
and  ( new_n30346_, new_n30345_, new_n30344_ );
xor  ( new_n30347_, new_n30346_, new_n2121_ );
or   ( new_n30348_, new_n2122_, new_n24227_ );
or   ( new_n30349_, new_n2124_, new_n24006_ );
and  ( new_n30350_, new_n30349_, new_n30348_ );
xor  ( new_n30351_, new_n30350_, new_n1843_ );
or   ( new_n30352_, new_n30351_, new_n30347_ );
and  ( new_n30353_, new_n30351_, new_n30347_ );
or   ( new_n30354_, new_n1844_, new_n24543_ );
or   ( new_n30355_, new_n1846_, new_n24418_ );
and  ( new_n30356_, new_n30355_, new_n30354_ );
xor  ( new_n30357_, new_n30356_, new_n1586_ );
or   ( new_n30358_, new_n30357_, new_n30353_ );
and  ( new_n30359_, new_n30358_, new_n30352_ );
or   ( new_n30360_, new_n4709_, new_n22304_ );
or   ( new_n30361_, new_n4711_, new_n22207_ );
and  ( new_n30362_, new_n30361_, new_n30360_ );
xor  ( new_n30363_, new_n30362_, new_n4295_ );
or   ( new_n30364_, new_n4302_, new_n22590_ );
or   ( new_n30365_, new_n4304_, new_n22423_ );
and  ( new_n30366_, new_n30365_, new_n30364_ );
xor  ( new_n30367_, new_n30366_, new_n3895_ );
or   ( new_n30368_, new_n30367_, new_n30363_ );
and  ( new_n30369_, new_n30367_, new_n30363_ );
or   ( new_n30370_, new_n3896_, new_n22829_ );
or   ( new_n30371_, new_n3898_, new_n22641_ );
and  ( new_n30372_, new_n30371_, new_n30370_ );
xor  ( new_n30373_, new_n30372_, new_n3460_ );
or   ( new_n30374_, new_n30373_, new_n30369_ );
and  ( new_n30375_, new_n30374_, new_n30368_ );
nor  ( new_n30376_, new_n30375_, new_n30359_ );
and  ( new_n30377_, new_n30375_, new_n30359_ );
or   ( new_n30378_, new_n3461_, new_n22973_ );
or   ( new_n30379_, new_n3463_, new_n22975_ );
and  ( new_n30380_, new_n30379_, new_n30378_ );
xor  ( new_n30381_, new_n30380_, new_n3116_ );
or   ( new_n30382_, new_n3117_, new_n23252_ );
or   ( new_n30383_, new_n3119_, new_n23166_ );
and  ( new_n30384_, new_n30383_, new_n30382_ );
xor  ( new_n30385_, new_n30384_, new_n2800_ );
nor  ( new_n30386_, new_n30385_, new_n30381_ );
and  ( new_n30387_, new_n30385_, new_n30381_ );
or   ( new_n30388_, new_n2807_, new_n23554_ );
or   ( new_n30389_, new_n2809_, new_n23370_ );
and  ( new_n30390_, new_n30389_, new_n30388_ );
xor  ( new_n30391_, new_n30390_, new_n2424_ );
nor  ( new_n30392_, new_n30391_, new_n30387_ );
nor  ( new_n30393_, new_n30392_, new_n30386_ );
nor  ( new_n30394_, new_n30393_, new_n30377_ );
nor  ( new_n30395_, new_n30394_, new_n30376_ );
and  ( new_n30396_, new_n30342_, new_n30292_ );
or   ( new_n30397_, new_n30396_, new_n30395_ );
and  ( new_n30398_, new_n30397_, new_n30343_ );
or   ( new_n30399_, new_n30398_, new_n30240_ );
and  ( new_n30400_, new_n30398_, new_n30240_ );
xor  ( new_n30401_, new_n29936_, new_n29934_ );
xor  ( new_n30402_, new_n30401_, new_n29940_ );
xnor ( new_n30403_, new_n30020_, new_n30016_ );
xor  ( new_n30404_, new_n30403_, new_n30026_ );
xnor ( new_n30405_, new_n30038_, new_n30034_ );
xor  ( new_n30406_, new_n30405_, new_n30044_ );
or   ( new_n30407_, new_n30406_, new_n30404_ );
and  ( new_n30408_, new_n30406_, new_n30404_ );
xor  ( new_n30409_, new_n29990_, new_n29986_ );
xnor ( new_n30410_, new_n30409_, new_n29996_ );
or   ( new_n30411_, new_n30410_, new_n30408_ );
and  ( new_n30412_, new_n30411_, new_n30407_ );
nor  ( new_n30413_, new_n30412_, new_n30402_ );
nand ( new_n30414_, new_n30412_, new_n30402_ );
xor  ( new_n30415_, new_n30131_, new_n30129_ );
xnor ( new_n30416_, new_n30415_, new_n30135_ );
and  ( new_n30417_, new_n30416_, new_n30414_ );
or   ( new_n30418_, new_n30417_, new_n30413_ );
or   ( new_n30419_, new_n30418_, new_n30400_ );
and  ( new_n30420_, new_n30419_, new_n30399_ );
or   ( new_n30421_, new_n30420_, new_n30193_ );
nand ( new_n30422_, new_n30420_, new_n30193_ );
xor  ( new_n30423_, new_n30137_, new_n30127_ );
xor  ( new_n30424_, new_n30423_, new_n30149_ );
xnor ( new_n30425_, new_n30048_, new_n30000_ );
xor  ( new_n30426_, new_n30425_, new_n30101_ );
nor  ( new_n30427_, new_n30426_, new_n30424_ );
and  ( new_n30428_, new_n30426_, new_n30424_ );
xor  ( new_n30429_, new_n29942_, new_n29932_ );
xnor ( new_n30430_, new_n30429_, new_n29946_ );
nor  ( new_n30431_, new_n30430_, new_n30428_ );
nor  ( new_n30432_, new_n30431_, new_n30427_ );
nand ( new_n30433_, new_n30432_, new_n30422_ );
and  ( new_n30434_, new_n30433_, new_n30421_ );
nor  ( new_n30435_, new_n30434_, new_n30175_ );
nand ( new_n30436_, new_n30434_, new_n30175_ );
xor  ( new_n30437_, new_n29765_, new_n29713_ );
xor  ( new_n30438_, new_n30437_, new_n29816_ );
xor  ( new_n30439_, new_n29647_, new_n29637_ );
xor  ( new_n30440_, new_n30439_, new_n29659_ );
and  ( new_n30441_, new_n30440_, new_n30438_ );
nor  ( new_n30442_, new_n30440_, new_n30438_ );
xor  ( new_n30443_, new_n29921_, new_n29919_ );
xor  ( new_n30444_, new_n30443_, new_n29926_ );
nor  ( new_n30445_, new_n30444_, new_n30442_ );
nor  ( new_n30446_, new_n30445_, new_n30441_ );
and  ( new_n30447_, new_n30446_, new_n30436_ );
or   ( new_n30448_, new_n30447_, new_n30435_ );
xor  ( new_n30449_, new_n29834_, new_n29614_ );
xor  ( new_n30450_, new_n30449_, new_n29846_ );
or   ( new_n30451_, new_n30450_, new_n30448_ );
and  ( new_n30452_, new_n30450_, new_n30448_ );
xor  ( new_n30453_, new_n29889_, new_n29879_ );
xor  ( new_n30454_, new_n30453_, new_n30155_ );
or   ( new_n30455_, new_n30454_, new_n30452_ );
and  ( new_n30456_, new_n30455_, new_n30451_ );
nor  ( new_n30457_, new_n30456_, new_n30173_ );
xor  ( new_n30458_, new_n30164_, new_n29877_ );
xor  ( new_n30459_, new_n30458_, new_n30168_ );
and  ( new_n30460_, new_n30459_, new_n30457_ );
xor  ( new_n30461_, new_n30450_, new_n30448_ );
xnor ( new_n30462_, new_n30461_, new_n30454_ );
xnor ( new_n30463_, new_n29903_, new_n29901_ );
xor  ( new_n30464_, new_n30463_, new_n29915_ );
xnor ( new_n30465_, new_n29980_, new_n29964_ );
xor  ( new_n30466_, new_n30465_, new_n29998_ );
xor  ( new_n30467_, new_n30233_, new_n30216_ );
xor  ( new_n30468_, new_n30467_, new_n30236_ );
xnor ( new_n30469_, new_n30197_, new_n30195_ );
xor  ( new_n30470_, new_n30469_, new_n30201_ );
nand ( new_n30471_, new_n30470_, new_n30468_ );
or   ( new_n30472_, new_n30470_, new_n30468_ );
xor  ( new_n30473_, new_n30207_, new_n30205_ );
xnor ( new_n30474_, new_n30473_, new_n30211_ );
nand ( new_n30475_, new_n30474_, new_n30472_ );
and  ( new_n30476_, new_n30475_, new_n30471_ );
nor  ( new_n30477_, new_n30476_, new_n30466_ );
and  ( new_n30478_, new_n30476_, new_n30466_ );
xnor ( new_n30479_, new_n30272_, new_n30256_ );
xor  ( new_n30480_, new_n30479_, new_n30290_ );
xnor ( new_n30481_, new_n30322_, new_n30308_ );
xor  ( new_n30482_, new_n30481_, new_n30340_ );
nor  ( new_n30483_, new_n30482_, new_n30480_ );
and  ( new_n30484_, new_n30482_, new_n30480_ );
xor  ( new_n30485_, new_n30375_, new_n30359_ );
xnor ( new_n30486_, new_n30485_, new_n30393_ );
nor  ( new_n30487_, new_n30486_, new_n30484_ );
nor  ( new_n30488_, new_n30487_, new_n30483_ );
nor  ( new_n30489_, new_n30488_, new_n30478_ );
or   ( new_n30490_, new_n30489_, new_n30477_ );
or   ( new_n30491_, new_n1135_, new_n26196_ );
or   ( new_n30492_, new_n1137_, new_n25813_ );
and  ( new_n30493_, new_n30492_, new_n30491_ );
xor  ( new_n30494_, new_n30493_, new_n896_ );
or   ( new_n30495_, new_n897_, new_n26372_ );
or   ( new_n30496_, new_n899_, new_n26063_ );
and  ( new_n30497_, new_n30496_, new_n30495_ );
xor  ( new_n30498_, new_n30497_, new_n748_ );
or   ( new_n30499_, new_n30498_, new_n30494_ );
and  ( new_n30500_, new_n30498_, new_n30494_ );
or   ( new_n30501_, new_n755_, new_n26762_ );
or   ( new_n30502_, new_n757_, new_n26620_ );
and  ( new_n30503_, new_n30502_, new_n30501_ );
xor  ( new_n30504_, new_n30503_, new_n523_ );
or   ( new_n30505_, new_n30504_, new_n30500_ );
and  ( new_n30506_, new_n30505_, new_n30499_ );
or   ( new_n30507_, new_n524_, new_n27396_ );
or   ( new_n30508_, new_n526_, new_n27085_ );
and  ( new_n30509_, new_n30508_, new_n30507_ );
xor  ( new_n30510_, new_n30509_, new_n403_ );
or   ( new_n30511_, new_n409_, new_n27763_ );
or   ( new_n30512_, new_n411_, new_n27602_ );
and  ( new_n30513_, new_n30512_, new_n30511_ );
xor  ( new_n30514_, new_n30513_, new_n328_ );
or   ( new_n30515_, new_n30514_, new_n30510_ );
and  ( new_n30516_, new_n30514_, new_n30510_ );
or   ( new_n30517_, new_n337_, new_n28314_ );
or   ( new_n30518_, new_n340_, new_n28108_ );
and  ( new_n30519_, new_n30518_, new_n30517_ );
xor  ( new_n30520_, new_n30519_, new_n332_ );
or   ( new_n30521_, new_n30520_, new_n30516_ );
and  ( new_n30522_, new_n30521_, new_n30515_ );
or   ( new_n30523_, new_n30522_, new_n30506_ );
and  ( new_n30524_, new_n30522_, new_n30506_ );
or   ( new_n30525_, new_n1844_, new_n24927_ );
or   ( new_n30526_, new_n1846_, new_n24543_ );
and  ( new_n30527_, new_n30526_, new_n30525_ );
xor  ( new_n30528_, new_n30527_, new_n1586_ );
or   ( new_n30529_, new_n1593_, new_n25048_ );
or   ( new_n30530_, new_n1595_, new_n24925_ );
and  ( new_n30531_, new_n30530_, new_n30529_ );
xor  ( new_n30532_, new_n30531_, new_n1358_ );
nor  ( new_n30533_, new_n30532_, new_n30528_ );
and  ( new_n30534_, new_n30532_, new_n30528_ );
or   ( new_n30535_, new_n1364_, new_n25486_ );
or   ( new_n30536_, new_n1366_, new_n25288_ );
and  ( new_n30537_, new_n30536_, new_n30535_ );
xor  ( new_n30538_, new_n30537_, new_n1129_ );
nor  ( new_n30539_, new_n30538_, new_n30534_ );
nor  ( new_n30540_, new_n30539_, new_n30533_ );
or   ( new_n30541_, new_n30540_, new_n30524_ );
and  ( new_n30542_, new_n30541_, new_n30523_ );
or   ( new_n30543_, new_n9422_, new_n21694_ );
or   ( new_n30544_, new_n9424_, new_n21696_ );
and  ( new_n30545_, new_n30544_, new_n30543_ );
xor  ( new_n30546_, new_n30545_, new_n8873_ );
and  ( new_n30547_, new_n30546_, new_n9421_ );
or   ( new_n30548_, new_n30546_, new_n9421_ );
or   ( new_n30549_, new_n8874_, new_n21701_ );
or   ( new_n30550_, new_n8876_, new_n21703_ );
and  ( new_n30551_, new_n30550_, new_n30549_ );
xor  ( new_n30552_, new_n30551_, new_n8257_ );
and  ( new_n30553_, new_n30552_, new_n30548_ );
or   ( new_n30554_, new_n30553_, new_n30547_ );
or   ( new_n30555_, new_n6645_, new_n21792_ );
or   ( new_n30556_, new_n6647_, new_n21751_ );
and  ( new_n30557_, new_n30556_, new_n30555_ );
xor  ( new_n30558_, new_n30557_, new_n6166_ );
or   ( new_n30559_, new_n6173_, new_n21840_ );
or   ( new_n30560_, new_n6175_, new_n21842_ );
and  ( new_n30561_, new_n30560_, new_n30559_ );
xor  ( new_n30562_, new_n30561_, new_n5597_ );
or   ( new_n30563_, new_n30562_, new_n30558_ );
and  ( new_n30564_, new_n30562_, new_n30558_ );
or   ( new_n30565_, new_n5604_, new_n22098_ );
or   ( new_n30566_, new_n5606_, new_n21847_ );
and  ( new_n30567_, new_n30566_, new_n30565_ );
xor  ( new_n30568_, new_n30567_, new_n5206_ );
or   ( new_n30569_, new_n30568_, new_n30564_ );
and  ( new_n30570_, new_n30569_, new_n30563_ );
or   ( new_n30571_, new_n30570_, new_n30554_ );
and  ( new_n30572_, new_n30570_, new_n30554_ );
or   ( new_n30573_, new_n8264_, new_n21672_ );
or   ( new_n30574_, new_n8266_, new_n21674_ );
and  ( new_n30575_, new_n30574_, new_n30573_ );
xor  ( new_n30576_, new_n30575_, new_n7725_ );
or   ( new_n30577_, new_n7732_, new_n21678_ );
or   ( new_n30578_, new_n7734_, new_n21680_ );
and  ( new_n30579_, new_n30578_, new_n30577_ );
xor  ( new_n30580_, new_n30579_, new_n7177_ );
nor  ( new_n30581_, new_n30580_, new_n30576_ );
and  ( new_n30582_, new_n30580_, new_n30576_ );
or   ( new_n30583_, new_n7184_, new_n21685_ );
or   ( new_n30584_, new_n7186_, new_n21687_ );
and  ( new_n30585_, new_n30584_, new_n30583_ );
xor  ( new_n30586_, new_n30585_, new_n6638_ );
nor  ( new_n30587_, new_n30586_, new_n30582_ );
nor  ( new_n30588_, new_n30587_, new_n30581_ );
or   ( new_n30589_, new_n30588_, new_n30572_ );
and  ( new_n30590_, new_n30589_, new_n30571_ );
nor  ( new_n30591_, new_n30590_, new_n30542_ );
nand ( new_n30592_, new_n30590_, new_n30542_ );
or   ( new_n30593_, new_n3896_, new_n22975_ );
or   ( new_n30594_, new_n3898_, new_n22829_ );
and  ( new_n30595_, new_n30594_, new_n30593_ );
xor  ( new_n30596_, new_n30595_, new_n3460_ );
or   ( new_n30597_, new_n3461_, new_n23166_ );
or   ( new_n30598_, new_n3463_, new_n22973_ );
and  ( new_n30599_, new_n30598_, new_n30597_ );
xor  ( new_n30600_, new_n30599_, new_n3116_ );
or   ( new_n30601_, new_n30600_, new_n30596_ );
and  ( new_n30602_, new_n30600_, new_n30596_ );
or   ( new_n30603_, new_n3117_, new_n23370_ );
or   ( new_n30604_, new_n3119_, new_n23252_ );
and  ( new_n30605_, new_n30604_, new_n30603_ );
xor  ( new_n30606_, new_n30605_, new_n2800_ );
or   ( new_n30607_, new_n30606_, new_n30602_ );
and  ( new_n30608_, new_n30607_, new_n30601_ );
or   ( new_n30609_, new_n2807_, new_n23733_ );
or   ( new_n30610_, new_n2809_, new_n23554_ );
and  ( new_n30611_, new_n30610_, new_n30609_ );
xor  ( new_n30612_, new_n30611_, new_n2424_ );
or   ( new_n30613_, new_n2425_, new_n24006_ );
or   ( new_n30614_, new_n2427_, new_n23895_ );
and  ( new_n30615_, new_n30614_, new_n30613_ );
xor  ( new_n30616_, new_n30615_, new_n2121_ );
or   ( new_n30617_, new_n30616_, new_n30612_ );
and  ( new_n30618_, new_n30616_, new_n30612_ );
or   ( new_n30619_, new_n2122_, new_n24418_ );
or   ( new_n30620_, new_n2124_, new_n24227_ );
and  ( new_n30621_, new_n30620_, new_n30619_ );
xor  ( new_n30622_, new_n30621_, new_n1843_ );
or   ( new_n30623_, new_n30622_, new_n30618_ );
and  ( new_n30624_, new_n30623_, new_n30617_ );
nor  ( new_n30625_, new_n30624_, new_n30608_ );
nand ( new_n30626_, new_n30624_, new_n30608_ );
or   ( new_n30627_, new_n5207_, new_n22207_ );
or   ( new_n30628_, new_n5209_, new_n22129_ );
and  ( new_n30629_, new_n30628_, new_n30627_ );
xor  ( new_n30630_, new_n30629_, new_n4708_ );
or   ( new_n30631_, new_n4709_, new_n22423_ );
or   ( new_n30632_, new_n4711_, new_n22304_ );
and  ( new_n30633_, new_n30632_, new_n30631_ );
xor  ( new_n30634_, new_n30633_, new_n4295_ );
nor  ( new_n30635_, new_n30634_, new_n30630_ );
and  ( new_n30636_, new_n30634_, new_n30630_ );
or   ( new_n30637_, new_n4302_, new_n22641_ );
or   ( new_n30638_, new_n4304_, new_n22590_ );
and  ( new_n30639_, new_n30638_, new_n30637_ );
xor  ( new_n30640_, new_n30639_, new_n3895_ );
nor  ( new_n30641_, new_n30640_, new_n30636_ );
nor  ( new_n30642_, new_n30641_, new_n30635_ );
not  ( new_n30643_, new_n30642_ );
and  ( new_n30644_, new_n30643_, new_n30626_ );
or   ( new_n30645_, new_n30644_, new_n30625_ );
and  ( new_n30646_, new_n30645_, new_n30592_ );
or   ( new_n30647_, new_n30646_, new_n30591_ );
not  ( new_n30648_, new_n30216_ );
or   ( new_n30649_, new_n317_, new_n29263_ );
or   ( new_n30650_, new_n320_, new_n28531_ );
and  ( new_n30651_, new_n30650_, new_n30649_ );
xor  ( new_n30652_, new_n30651_, new_n312_ );
or   ( new_n30653_, new_n283_, new_n29474_ );
or   ( new_n30654_, new_n286_, new_n29261_ );
and  ( new_n30655_, new_n30654_, new_n30653_ );
xor  ( new_n30656_, new_n30655_, new_n278_ );
or   ( new_n30657_, new_n30656_, new_n30652_ );
and  ( new_n30658_, new_n30656_, new_n30652_ );
or   ( new_n30659_, new_n299_, new_n30120_ );
or   ( new_n30660_, new_n302_, new_n29619_ );
and  ( new_n30661_, new_n30660_, new_n30659_ );
xor  ( new_n30662_, new_n30661_, new_n293_ );
or   ( new_n30663_, new_n30662_, new_n30658_ );
and  ( new_n30664_, new_n30663_, new_n30657_ );
nor  ( new_n30665_, new_n30664_, new_n30648_ );
nand ( new_n30666_, new_n30664_, new_n30648_ );
xor  ( new_n30667_, new_n30224_, new_n30220_ );
xnor ( new_n30668_, new_n30667_, new_n30231_ );
and  ( new_n30669_, new_n30668_, new_n30666_ );
or   ( new_n30670_, new_n30669_, new_n30665_ );
xnor ( new_n30671_, new_n30367_, new_n30363_ );
xor  ( new_n30672_, new_n30671_, new_n30373_ );
xnor ( new_n30673_, new_n30351_, new_n30347_ );
xor  ( new_n30674_, new_n30673_, new_n30357_ );
or   ( new_n30675_, new_n30674_, new_n30672_ );
and  ( new_n30676_, new_n30674_, new_n30672_ );
xor  ( new_n30677_, new_n30385_, new_n30381_ );
xnor ( new_n30678_, new_n30677_, new_n30391_ );
or   ( new_n30679_, new_n30678_, new_n30676_ );
and  ( new_n30680_, new_n30679_, new_n30675_ );
or   ( new_n30681_, new_n30680_, new_n30670_ );
and  ( new_n30682_, new_n30680_, new_n30670_ );
xnor ( new_n30683_, new_n30264_, new_n30260_ );
xor  ( new_n30684_, new_n30683_, new_n30270_ );
xnor ( new_n30685_, new_n30248_, new_n30244_ );
xor  ( new_n30686_, new_n30685_, new_n30254_ );
nor  ( new_n30687_, new_n30686_, new_n30684_ );
and  ( new_n30688_, new_n30686_, new_n30684_ );
xor  ( new_n30689_, new_n30282_, new_n30278_ );
xnor ( new_n30690_, new_n30689_, new_n30288_ );
nor  ( new_n30691_, new_n30690_, new_n30688_ );
nor  ( new_n30692_, new_n30691_, new_n30687_ );
or   ( new_n30693_, new_n30692_, new_n30682_ );
and  ( new_n30694_, new_n30693_, new_n30681_ );
nand ( new_n30695_, new_n30694_, new_n30647_ );
or   ( new_n30696_, new_n30694_, new_n30647_ );
xor  ( new_n30697_, new_n30004_, new_n8872_ );
xor  ( new_n30698_, new_n30697_, new_n30010_ );
xnor ( new_n30699_, new_n30314_, new_n30312_ );
xor  ( new_n30700_, new_n30699_, new_n30320_ );
xnor ( new_n30701_, new_n30300_, new_n30296_ );
xor  ( new_n30702_, new_n30701_, new_n30306_ );
or   ( new_n30703_, new_n30702_, new_n30700_ );
and  ( new_n30704_, new_n30702_, new_n30700_ );
xor  ( new_n30705_, new_n30332_, new_n30328_ );
xnor ( new_n30706_, new_n30705_, new_n30338_ );
or   ( new_n30707_, new_n30706_, new_n30704_ );
and  ( new_n30708_, new_n30707_, new_n30703_ );
nor  ( new_n30709_, new_n30708_, new_n30698_ );
and  ( new_n30710_, new_n30708_, new_n30698_ );
xor  ( new_n30711_, new_n30406_, new_n30404_ );
xnor ( new_n30712_, new_n30711_, new_n30410_ );
not  ( new_n30713_, new_n30712_ );
nor  ( new_n30714_, new_n30713_, new_n30710_ );
nor  ( new_n30715_, new_n30714_, new_n30709_ );
nand ( new_n30716_, new_n30715_, new_n30696_ );
and  ( new_n30717_, new_n30716_, new_n30695_ );
or   ( new_n30718_, new_n30717_, new_n30490_ );
nand ( new_n30719_, new_n30717_, new_n30490_ );
xnor ( new_n30720_, new_n30028_, new_n30012_ );
xor  ( new_n30721_, new_n30720_, new_n30046_ );
xnor ( new_n30722_, new_n30412_, new_n30402_ );
xor  ( new_n30723_, new_n30722_, new_n30416_ );
nor  ( new_n30724_, new_n30723_, new_n30721_ );
and  ( new_n30725_, new_n30723_, new_n30721_ );
xor  ( new_n30726_, new_n30185_, new_n30183_ );
xnor ( new_n30727_, new_n30726_, new_n30188_ );
not  ( new_n30728_, new_n30727_ );
nor  ( new_n30729_, new_n30728_, new_n30725_ );
nor  ( new_n30730_, new_n30729_, new_n30724_ );
nand ( new_n30731_, new_n30730_, new_n30719_ );
and  ( new_n30732_, new_n30731_, new_n30718_ );
nor  ( new_n30733_, new_n30732_, new_n30464_ );
nand ( new_n30734_, new_n30732_, new_n30464_ );
xor  ( new_n30735_, new_n30398_, new_n30240_ );
xor  ( new_n30736_, new_n30735_, new_n30418_ );
xnor ( new_n30737_, new_n30426_, new_n30424_ );
xor  ( new_n30738_, new_n30737_, new_n30430_ );
nand ( new_n30739_, new_n30738_, new_n30736_ );
or   ( new_n30740_, new_n30738_, new_n30736_ );
xor  ( new_n30741_, new_n30179_, new_n30177_ );
xor  ( new_n30742_, new_n30741_, new_n30191_ );
nand ( new_n30743_, new_n30742_, new_n30740_ );
and  ( new_n30744_, new_n30743_, new_n30739_ );
and  ( new_n30745_, new_n30744_, new_n30734_ );
or   ( new_n30746_, new_n30745_, new_n30733_ );
xor  ( new_n30747_, new_n30104_, new_n29948_ );
xor  ( new_n30748_, new_n30747_, new_n30151_ );
xor  ( new_n30749_, new_n30420_, new_n30193_ );
xor  ( new_n30750_, new_n30749_, new_n30432_ );
or   ( new_n30751_, new_n30750_, new_n30748_ );
and  ( new_n30752_, new_n30750_, new_n30748_ );
xor  ( new_n30753_, new_n30440_, new_n30438_ );
xnor ( new_n30754_, new_n30753_, new_n30444_ );
not  ( new_n30755_, new_n30754_ );
or   ( new_n30756_, new_n30755_, new_n30752_ );
and  ( new_n30757_, new_n30756_, new_n30751_ );
or   ( new_n30758_, new_n30757_, new_n30746_ );
and  ( new_n30759_, new_n30757_, new_n30746_ );
xor  ( new_n30760_, new_n29928_, new_n29917_ );
xor  ( new_n30761_, new_n30760_, new_n30153_ );
or   ( new_n30762_, new_n30761_, new_n30759_ );
nand ( new_n30763_, new_n30762_, new_n30758_ );
and  ( new_n30764_, new_n30763_, new_n30462_ );
xor  ( new_n30765_, new_n30456_, new_n30173_ );
and  ( new_n30766_, new_n30765_, new_n30764_ );
xnor ( new_n30767_, new_n30763_, new_n30462_ );
xor  ( new_n30768_, new_n30757_, new_n30746_ );
xor  ( new_n30769_, new_n30768_, new_n30761_ );
xor  ( new_n30770_, new_n30738_, new_n30736_ );
xor  ( new_n30771_, new_n30770_, new_n30742_ );
xor  ( new_n30772_, new_n30482_, new_n30480_ );
xor  ( new_n30773_, new_n30772_, new_n30486_ );
xnor ( new_n30774_, new_n30674_, new_n30672_ );
xor  ( new_n30775_, new_n30774_, new_n30678_ );
xnor ( new_n30776_, new_n30686_, new_n30684_ );
xor  ( new_n30777_, new_n30776_, new_n30690_ );
nand ( new_n30778_, new_n30777_, new_n30775_ );
nor  ( new_n30779_, new_n30777_, new_n30775_ );
xor  ( new_n30780_, new_n30664_, new_n30648_ );
xor  ( new_n30781_, new_n30780_, new_n30668_ );
or   ( new_n30782_, new_n30781_, new_n30779_ );
and  ( new_n30783_, new_n30782_, new_n30778_ );
nor  ( new_n30784_, new_n30783_, new_n30773_ );
and  ( new_n30785_, new_n30783_, new_n30773_ );
xnor ( new_n30786_, new_n30522_, new_n30506_ );
xor  ( new_n30787_, new_n30786_, new_n30540_ );
xnor ( new_n30788_, new_n30570_, new_n30554_ );
xor  ( new_n30789_, new_n30788_, new_n30588_ );
nor  ( new_n30790_, new_n30789_, new_n30787_ );
and  ( new_n30791_, new_n30789_, new_n30787_ );
xor  ( new_n30792_, new_n30624_, new_n30608_ );
xor  ( new_n30793_, new_n30792_, new_n30643_ );
nor  ( new_n30794_, new_n30793_, new_n30791_ );
nor  ( new_n30795_, new_n30794_, new_n30790_ );
nor  ( new_n30796_, new_n30795_, new_n30785_ );
or   ( new_n30797_, new_n30796_, new_n30784_ );
not  ( new_n30798_, RIbb33210_189 );
or   ( new_n30799_, new_n268_, new_n30798_ );
not  ( new_n30800_, RIbb33198_188 );
or   ( new_n30801_, new_n271_, new_n30800_ );
and  ( new_n30802_, new_n30801_, new_n30799_ );
xor  ( new_n30803_, new_n30802_, new_n263_ );
and  ( new_n30804_, RIbb33288_190, RIbb2f610_1 );
or   ( new_n30805_, new_n30804_, new_n30803_ );
or   ( new_n30806_, new_n317_, new_n29261_ );
or   ( new_n30807_, new_n320_, new_n29263_ );
and  ( new_n30808_, new_n30807_, new_n30806_ );
xor  ( new_n30809_, new_n30808_, new_n312_ );
or   ( new_n30810_, new_n283_, new_n29619_ );
or   ( new_n30811_, new_n286_, new_n29474_ );
and  ( new_n30812_, new_n30811_, new_n30810_ );
xor  ( new_n30813_, new_n30812_, new_n278_ );
or   ( new_n30814_, new_n30813_, new_n30809_ );
and  ( new_n30815_, new_n30813_, new_n30809_ );
or   ( new_n30816_, new_n299_, new_n30227_ );
or   ( new_n30817_, new_n302_, new_n30120_ );
and  ( new_n30818_, new_n30817_, new_n30816_ );
xor  ( new_n30819_, new_n30818_, new_n293_ );
or   ( new_n30820_, new_n30819_, new_n30815_ );
and  ( new_n30821_, new_n30820_, new_n30814_ );
and  ( new_n30822_, new_n30821_, new_n30805_ );
or   ( new_n30823_, new_n30821_, new_n30805_ );
or   ( new_n30824_, new_n268_, new_n30800_ );
or   ( new_n30825_, new_n271_, new_n30227_ );
and  ( new_n30826_, new_n30825_, new_n30824_ );
xor  ( new_n30827_, new_n30826_, new_n263_ );
and  ( new_n30828_, new_n30827_, new_n30823_ );
or   ( new_n30829_, new_n30828_, new_n30822_ );
or   ( new_n30830_, new_n30798_, new_n260_ );
xnor ( new_n30831_, new_n30514_, new_n30510_ );
xor  ( new_n30832_, new_n30831_, new_n30520_ );
nand ( new_n30833_, new_n30832_, new_n30830_ );
or   ( new_n30834_, new_n30832_, new_n30830_ );
xor  ( new_n30835_, new_n30656_, new_n30652_ );
xnor ( new_n30836_, new_n30835_, new_n30662_ );
nand ( new_n30837_, new_n30836_, new_n30834_ );
and  ( new_n30838_, new_n30837_, new_n30833_ );
and  ( new_n30839_, new_n30838_, new_n30829_ );
nor  ( new_n30840_, new_n30838_, new_n30829_ );
xnor ( new_n30841_, new_n30616_, new_n30612_ );
xor  ( new_n30842_, new_n30841_, new_n30622_ );
xnor ( new_n30843_, new_n30498_, new_n30494_ );
xor  ( new_n30844_, new_n30843_, new_n30504_ );
nor  ( new_n30845_, new_n30844_, new_n30842_ );
and  ( new_n30846_, new_n30844_, new_n30842_ );
xor  ( new_n30847_, new_n30532_, new_n30528_ );
xnor ( new_n30848_, new_n30847_, new_n30538_ );
nor  ( new_n30849_, new_n30848_, new_n30846_ );
nor  ( new_n30850_, new_n30849_, new_n30845_ );
nor  ( new_n30851_, new_n30850_, new_n30840_ );
or   ( new_n30852_, new_n30851_, new_n30839_ );
or   ( new_n30853_, new_n9422_, new_n21703_ );
or   ( new_n30854_, new_n9424_, new_n21694_ );
and  ( new_n30855_, new_n30854_, new_n30853_ );
xor  ( new_n30856_, new_n30855_, new_n8872_ );
and  ( new_n30857_, new_n9740_, RIbb315f0_129 );
xor  ( new_n30858_, new_n30857_, new_n9421_ );
nand ( new_n30859_, new_n30858_, new_n30856_ );
nor  ( new_n30860_, new_n30858_, new_n30856_ );
or   ( new_n30861_, new_n8874_, new_n21674_ );
or   ( new_n30862_, new_n8876_, new_n21701_ );
and  ( new_n30863_, new_n30862_, new_n30861_ );
xor  ( new_n30864_, new_n30863_, new_n8257_ );
or   ( new_n30865_, new_n30864_, new_n30860_ );
and  ( new_n30866_, new_n30865_, new_n30859_ );
or   ( new_n30867_, new_n6645_, new_n21842_ );
or   ( new_n30868_, new_n6647_, new_n21792_ );
and  ( new_n30869_, new_n30868_, new_n30867_ );
xor  ( new_n30870_, new_n30869_, new_n6166_ );
or   ( new_n30871_, new_n6173_, new_n21847_ );
or   ( new_n30872_, new_n6175_, new_n21840_ );
and  ( new_n30873_, new_n30872_, new_n30871_ );
xor  ( new_n30874_, new_n30873_, new_n5597_ );
or   ( new_n30875_, new_n30874_, new_n30870_ );
and  ( new_n30876_, new_n30874_, new_n30870_ );
or   ( new_n30877_, new_n5604_, new_n22129_ );
or   ( new_n30878_, new_n5606_, new_n22098_ );
and  ( new_n30879_, new_n30878_, new_n30877_ );
xor  ( new_n30880_, new_n30879_, new_n5206_ );
or   ( new_n30881_, new_n30880_, new_n30876_ );
and  ( new_n30882_, new_n30881_, new_n30875_ );
or   ( new_n30883_, new_n30882_, new_n30866_ );
and  ( new_n30884_, new_n30882_, new_n30866_ );
or   ( new_n30885_, new_n8264_, new_n21680_ );
or   ( new_n30886_, new_n8266_, new_n21672_ );
and  ( new_n30887_, new_n30886_, new_n30885_ );
xor  ( new_n30888_, new_n30887_, new_n7725_ );
or   ( new_n30889_, new_n7732_, new_n21687_ );
or   ( new_n30890_, new_n7734_, new_n21678_ );
and  ( new_n30891_, new_n30890_, new_n30889_ );
xor  ( new_n30892_, new_n30891_, new_n7177_ );
nor  ( new_n30893_, new_n30892_, new_n30888_ );
and  ( new_n30894_, new_n30892_, new_n30888_ );
or   ( new_n30895_, new_n7184_, new_n21751_ );
or   ( new_n30896_, new_n7186_, new_n21685_ );
and  ( new_n30897_, new_n30896_, new_n30895_ );
xor  ( new_n30898_, new_n30897_, new_n6638_ );
nor  ( new_n30899_, new_n30898_, new_n30894_ );
nor  ( new_n30900_, new_n30899_, new_n30893_ );
or   ( new_n30901_, new_n30900_, new_n30884_ );
and  ( new_n30902_, new_n30901_, new_n30883_ );
or   ( new_n30903_, new_n1844_, new_n24925_ );
or   ( new_n30904_, new_n1846_, new_n24927_ );
and  ( new_n30905_, new_n30904_, new_n30903_ );
xor  ( new_n30906_, new_n30905_, new_n1586_ );
or   ( new_n30907_, new_n1593_, new_n25288_ );
or   ( new_n30908_, new_n1595_, new_n25048_ );
and  ( new_n30909_, new_n30908_, new_n30907_ );
xor  ( new_n30910_, new_n30909_, new_n1358_ );
or   ( new_n30911_, new_n30910_, new_n30906_ );
and  ( new_n30912_, new_n30910_, new_n30906_ );
or   ( new_n30913_, new_n1364_, new_n25813_ );
or   ( new_n30914_, new_n1366_, new_n25486_ );
and  ( new_n30915_, new_n30914_, new_n30913_ );
xor  ( new_n30916_, new_n30915_, new_n1129_ );
or   ( new_n30917_, new_n30916_, new_n30912_ );
and  ( new_n30918_, new_n30917_, new_n30911_ );
or   ( new_n30919_, new_n524_, new_n27602_ );
or   ( new_n30920_, new_n526_, new_n27396_ );
and  ( new_n30921_, new_n30920_, new_n30919_ );
xor  ( new_n30922_, new_n30921_, new_n403_ );
or   ( new_n30923_, new_n409_, new_n28108_ );
or   ( new_n30924_, new_n411_, new_n27763_ );
and  ( new_n30925_, new_n30924_, new_n30923_ );
xor  ( new_n30926_, new_n30925_, new_n328_ );
or   ( new_n30927_, new_n30926_, new_n30922_ );
and  ( new_n30928_, new_n30926_, new_n30922_ );
or   ( new_n30929_, new_n337_, new_n28531_ );
or   ( new_n30930_, new_n340_, new_n28314_ );
and  ( new_n30931_, new_n30930_, new_n30929_ );
xor  ( new_n30932_, new_n30931_, new_n332_ );
or   ( new_n30933_, new_n30932_, new_n30928_ );
and  ( new_n30934_, new_n30933_, new_n30927_ );
or   ( new_n30935_, new_n30934_, new_n30918_ );
and  ( new_n30936_, new_n30934_, new_n30918_ );
or   ( new_n30937_, new_n1135_, new_n26063_ );
or   ( new_n30938_, new_n1137_, new_n26196_ );
and  ( new_n30939_, new_n30938_, new_n30937_ );
xor  ( new_n30940_, new_n30939_, new_n896_ );
or   ( new_n30941_, new_n897_, new_n26620_ );
or   ( new_n30942_, new_n899_, new_n26372_ );
and  ( new_n30943_, new_n30942_, new_n30941_ );
xor  ( new_n30944_, new_n30943_, new_n748_ );
nor  ( new_n30945_, new_n30944_, new_n30940_ );
and  ( new_n30946_, new_n30944_, new_n30940_ );
or   ( new_n30947_, new_n755_, new_n27085_ );
or   ( new_n30948_, new_n757_, new_n26762_ );
and  ( new_n30949_, new_n30948_, new_n30947_ );
xor  ( new_n30950_, new_n30949_, new_n523_ );
nor  ( new_n30951_, new_n30950_, new_n30946_ );
nor  ( new_n30952_, new_n30951_, new_n30945_ );
or   ( new_n30953_, new_n30952_, new_n30936_ );
and  ( new_n30954_, new_n30953_, new_n30935_ );
or   ( new_n30955_, new_n30954_, new_n30902_ );
or   ( new_n30956_, new_n2807_, new_n23895_ );
or   ( new_n30957_, new_n2809_, new_n23733_ );
and  ( new_n30958_, new_n30957_, new_n30956_ );
xor  ( new_n30959_, new_n30958_, new_n2424_ );
or   ( new_n30960_, new_n2425_, new_n24227_ );
or   ( new_n30961_, new_n2427_, new_n24006_ );
and  ( new_n30962_, new_n30961_, new_n30960_ );
xor  ( new_n30963_, new_n30962_, new_n2121_ );
or   ( new_n30964_, new_n30963_, new_n30959_ );
and  ( new_n30965_, new_n30963_, new_n30959_ );
or   ( new_n30966_, new_n2122_, new_n24543_ );
or   ( new_n30967_, new_n2124_, new_n24418_ );
and  ( new_n30968_, new_n30967_, new_n30966_ );
xor  ( new_n30969_, new_n30968_, new_n1843_ );
or   ( new_n30970_, new_n30969_, new_n30965_ );
and  ( new_n30971_, new_n30970_, new_n30964_ );
or   ( new_n30972_, new_n5207_, new_n22304_ );
or   ( new_n30973_, new_n5209_, new_n22207_ );
and  ( new_n30974_, new_n30973_, new_n30972_ );
xor  ( new_n30975_, new_n30974_, new_n4708_ );
or   ( new_n30976_, new_n4709_, new_n22590_ );
or   ( new_n30977_, new_n4711_, new_n22423_ );
and  ( new_n30978_, new_n30977_, new_n30976_ );
xor  ( new_n30979_, new_n30978_, new_n4295_ );
or   ( new_n30980_, new_n30979_, new_n30975_ );
and  ( new_n30981_, new_n30979_, new_n30975_ );
or   ( new_n30982_, new_n4302_, new_n22829_ );
or   ( new_n30983_, new_n4304_, new_n22641_ );
and  ( new_n30984_, new_n30983_, new_n30982_ );
xor  ( new_n30985_, new_n30984_, new_n3895_ );
or   ( new_n30986_, new_n30985_, new_n30981_ );
and  ( new_n30987_, new_n30986_, new_n30980_ );
or   ( new_n30988_, new_n30987_, new_n30971_ );
and  ( new_n30989_, new_n30987_, new_n30971_ );
or   ( new_n30990_, new_n3896_, new_n22973_ );
or   ( new_n30991_, new_n3898_, new_n22975_ );
and  ( new_n30992_, new_n30991_, new_n30990_ );
xor  ( new_n30993_, new_n30992_, new_n3460_ );
or   ( new_n30994_, new_n3461_, new_n23252_ );
or   ( new_n30995_, new_n3463_, new_n23166_ );
and  ( new_n30996_, new_n30995_, new_n30994_ );
xor  ( new_n30997_, new_n30996_, new_n3116_ );
nor  ( new_n30998_, new_n30997_, new_n30993_ );
and  ( new_n30999_, new_n30997_, new_n30993_ );
or   ( new_n31000_, new_n3117_, new_n23554_ );
or   ( new_n31001_, new_n3119_, new_n23370_ );
and  ( new_n31002_, new_n31001_, new_n31000_ );
xor  ( new_n31003_, new_n31002_, new_n2800_ );
nor  ( new_n31004_, new_n31003_, new_n30999_ );
nor  ( new_n31005_, new_n31004_, new_n30998_ );
or   ( new_n31006_, new_n31005_, new_n30989_ );
and  ( new_n31007_, new_n31006_, new_n30988_ );
and  ( new_n31008_, new_n30954_, new_n30902_ );
or   ( new_n31009_, new_n31008_, new_n31007_ );
and  ( new_n31010_, new_n31009_, new_n30955_ );
or   ( new_n31011_, new_n31010_, new_n30852_ );
nand ( new_n31012_, new_n31010_, new_n30852_ );
xor  ( new_n31013_, new_n30580_, new_n30576_ );
xnor ( new_n31014_, new_n31013_, new_n30586_ );
not  ( new_n31015_, new_n31014_ );
xor  ( new_n31016_, new_n30546_, new_n9421_ );
xor  ( new_n31017_, new_n31016_, new_n30552_ );
nand ( new_n31018_, new_n31017_, new_n31015_ );
xnor ( new_n31019_, new_n30562_, new_n30558_ );
xor  ( new_n31020_, new_n31019_, new_n30568_ );
xnor ( new_n31021_, new_n30600_, new_n30596_ );
xor  ( new_n31022_, new_n31021_, new_n30606_ );
or   ( new_n31023_, new_n31022_, new_n31020_ );
and  ( new_n31024_, new_n31022_, new_n31020_ );
xnor ( new_n31025_, new_n30634_, new_n30630_ );
xor  ( new_n31026_, new_n31025_, new_n30640_ );
or   ( new_n31027_, new_n31026_, new_n31024_ );
and  ( new_n31028_, new_n31027_, new_n31023_ );
nor  ( new_n31029_, new_n31028_, new_n31018_ );
and  ( new_n31030_, new_n31028_, new_n31018_ );
xor  ( new_n31031_, new_n30702_, new_n30700_ );
xnor ( new_n31032_, new_n31031_, new_n30706_ );
not  ( new_n31033_, new_n31032_ );
nor  ( new_n31034_, new_n31033_, new_n31030_ );
nor  ( new_n31035_, new_n31034_, new_n31029_ );
nand ( new_n31036_, new_n31035_, new_n31012_ );
and  ( new_n31037_, new_n31036_, new_n31011_ );
or   ( new_n31038_, new_n31037_, new_n30797_ );
nand ( new_n31039_, new_n31037_, new_n30797_ );
xor  ( new_n31040_, new_n30470_, new_n30468_ );
xor  ( new_n31041_, new_n31040_, new_n30474_ );
xnor ( new_n31042_, new_n30680_, new_n30670_ );
xor  ( new_n31043_, new_n31042_, new_n30692_ );
and  ( new_n31044_, new_n31043_, new_n31041_ );
nor  ( new_n31045_, new_n31043_, new_n31041_ );
xor  ( new_n31046_, new_n30708_, new_n30698_ );
xor  ( new_n31047_, new_n31046_, new_n30713_ );
nor  ( new_n31048_, new_n31047_, new_n31045_ );
nor  ( new_n31049_, new_n31048_, new_n31044_ );
nand ( new_n31050_, new_n31049_, new_n31039_ );
and  ( new_n31051_, new_n31050_, new_n31038_ );
nor  ( new_n31052_, new_n31051_, new_n30771_ );
nand ( new_n31053_, new_n31051_, new_n30771_ );
xnor ( new_n31054_, new_n30213_, new_n30203_ );
xor  ( new_n31055_, new_n31054_, new_n30238_ );
xnor ( new_n31056_, new_n30342_, new_n30292_ );
xor  ( new_n31057_, new_n31056_, new_n30395_ );
or   ( new_n31058_, new_n31057_, new_n31055_ );
and  ( new_n31059_, new_n31057_, new_n31055_ );
xor  ( new_n31060_, new_n30723_, new_n30721_ );
xor  ( new_n31061_, new_n31060_, new_n30728_ );
or   ( new_n31062_, new_n31061_, new_n31059_ );
and  ( new_n31063_, new_n31062_, new_n31058_ );
and  ( new_n31064_, new_n31063_, new_n31053_ );
or   ( new_n31065_, new_n31064_, new_n31052_ );
xor  ( new_n31066_, new_n30732_, new_n30464_ );
xor  ( new_n31067_, new_n31066_, new_n30744_ );
or   ( new_n31068_, new_n31067_, new_n31065_ );
and  ( new_n31069_, new_n31067_, new_n31065_ );
xor  ( new_n31070_, new_n30750_, new_n30748_ );
xor  ( new_n31071_, new_n31070_, new_n30755_ );
or   ( new_n31072_, new_n31071_, new_n31069_ );
and  ( new_n31073_, new_n31072_, new_n31068_ );
or   ( new_n31074_, new_n31073_, new_n30769_ );
and  ( new_n31075_, new_n31073_, new_n30769_ );
xor  ( new_n31076_, new_n30434_, new_n30175_ );
xor  ( new_n31077_, new_n31076_, new_n30446_ );
or   ( new_n31078_, new_n31077_, new_n31075_ );
and  ( new_n31079_, new_n31078_, new_n31074_ );
nor  ( new_n31080_, new_n31079_, new_n30767_ );
xor  ( new_n31081_, new_n30476_, new_n30466_ );
xor  ( new_n31082_, new_n31081_, new_n30488_ );
xor  ( new_n31083_, new_n30783_, new_n30773_ );
xor  ( new_n31084_, new_n31083_, new_n30795_ );
xor  ( new_n31085_, new_n30590_, new_n30542_ );
xor  ( new_n31086_, new_n31085_, new_n30645_ );
or   ( new_n31087_, new_n31086_, new_n31084_ );
and  ( new_n31088_, new_n31086_, new_n31084_ );
xor  ( new_n31089_, new_n31043_, new_n31041_ );
xnor ( new_n31090_, new_n31089_, new_n31047_ );
not  ( new_n31091_, new_n31090_ );
or   ( new_n31092_, new_n31091_, new_n31088_ );
and  ( new_n31093_, new_n31092_, new_n31087_ );
or   ( new_n31094_, new_n31093_, new_n31082_ );
and  ( new_n31095_, new_n31093_, new_n31082_ );
xnor ( new_n31096_, new_n30821_, new_n30805_ );
xor  ( new_n31097_, new_n31096_, new_n30827_ );
xor  ( new_n31098_, new_n30832_, new_n30830_ );
xor  ( new_n31099_, new_n31098_, new_n30836_ );
nor  ( new_n31100_, new_n31099_, new_n31097_ );
nand ( new_n31101_, new_n31099_, new_n31097_ );
xnor ( new_n31102_, new_n30844_, new_n30842_ );
xor  ( new_n31103_, new_n31102_, new_n30848_ );
and  ( new_n31104_, new_n31103_, new_n31101_ );
or   ( new_n31105_, new_n31104_, new_n31100_ );
xnor ( new_n31106_, new_n30789_, new_n30787_ );
xor  ( new_n31107_, new_n31106_, new_n30793_ );
nand ( new_n31108_, new_n31107_, new_n31105_ );
nor  ( new_n31109_, new_n31107_, new_n31105_ );
xnor ( new_n31110_, new_n30882_, new_n30866_ );
xor  ( new_n31111_, new_n31110_, new_n30900_ );
xnor ( new_n31112_, new_n30934_, new_n30918_ );
xor  ( new_n31113_, new_n31112_, new_n30952_ );
nor  ( new_n31114_, new_n31113_, new_n31111_ );
and  ( new_n31115_, new_n31113_, new_n31111_ );
xor  ( new_n31116_, new_n30987_, new_n30971_ );
xnor ( new_n31117_, new_n31116_, new_n31005_ );
nor  ( new_n31118_, new_n31117_, new_n31115_ );
nor  ( new_n31119_, new_n31118_, new_n31114_ );
or   ( new_n31120_, new_n31119_, new_n31109_ );
and  ( new_n31121_, new_n31120_, new_n31108_ );
xor  ( new_n31122_, new_n30838_, new_n30829_ );
xor  ( new_n31123_, new_n31122_, new_n30850_ );
xor  ( new_n31124_, new_n31028_, new_n31018_ );
xor  ( new_n31125_, new_n31124_, new_n31033_ );
or   ( new_n31126_, new_n31125_, new_n31123_ );
and  ( new_n31127_, new_n31125_, new_n31123_ );
xor  ( new_n31128_, new_n30777_, new_n30775_ );
xnor ( new_n31129_, new_n31128_, new_n30781_ );
not  ( new_n31130_, new_n31129_ );
or   ( new_n31131_, new_n31130_, new_n31127_ );
and  ( new_n31132_, new_n31131_, new_n31126_ );
or   ( new_n31133_, new_n31132_, new_n31121_ );
and  ( new_n31134_, new_n31132_, new_n31121_ );
xor  ( new_n31135_, new_n31022_, new_n31020_ );
xor  ( new_n31136_, new_n31135_, new_n31026_ );
xnor ( new_n31137_, new_n30979_, new_n30975_ );
xor  ( new_n31138_, new_n31137_, new_n30985_ );
xnor ( new_n31139_, new_n30874_, new_n30870_ );
xor  ( new_n31140_, new_n31139_, new_n30880_ );
or   ( new_n31141_, new_n31140_, new_n31138_ );
and  ( new_n31142_, new_n31140_, new_n31138_ );
xor  ( new_n31143_, new_n30892_, new_n30888_ );
xnor ( new_n31144_, new_n31143_, new_n30898_ );
or   ( new_n31145_, new_n31144_, new_n31142_ );
and  ( new_n31146_, new_n31145_, new_n31141_ );
nor  ( new_n31147_, new_n31146_, new_n31136_ );
nand ( new_n31148_, new_n31146_, new_n31136_ );
xor  ( new_n31149_, new_n31017_, new_n31015_ );
and  ( new_n31150_, new_n31149_, new_n31148_ );
or   ( new_n31151_, new_n31150_, new_n31147_ );
or   ( new_n31152_, new_n8874_, new_n21672_ );
or   ( new_n31153_, new_n8876_, new_n21674_ );
and  ( new_n31154_, new_n31153_, new_n31152_ );
xor  ( new_n31155_, new_n31154_, new_n8257_ );
or   ( new_n31156_, new_n8264_, new_n21678_ );
or   ( new_n31157_, new_n8266_, new_n21680_ );
and  ( new_n31158_, new_n31157_, new_n31156_ );
xor  ( new_n31159_, new_n31158_, new_n7725_ );
or   ( new_n31160_, new_n31159_, new_n31155_ );
and  ( new_n31161_, new_n31159_, new_n31155_ );
or   ( new_n31162_, new_n7732_, new_n21685_ );
or   ( new_n31163_, new_n7734_, new_n21687_ );
and  ( new_n31164_, new_n31163_, new_n31162_ );
xor  ( new_n31165_, new_n31164_, new_n7177_ );
or   ( new_n31166_, new_n31165_, new_n31161_ );
and  ( new_n31167_, new_n31166_, new_n31160_ );
or   ( new_n31168_, new_n9422_, new_n21701_ );
or   ( new_n31169_, new_n9424_, new_n21703_ );
and  ( new_n31170_, new_n31169_, new_n31168_ );
xor  ( new_n31171_, new_n31170_, new_n8873_ );
or   ( new_n31172_, new_n31171_, new_n10052_ );
and  ( new_n31173_, new_n31171_, new_n10052_ );
or   ( new_n31174_, new_n10059_, new_n21694_ );
or   ( new_n31175_, new_n10061_, new_n21696_ );
and  ( new_n31176_, new_n31175_, new_n31174_ );
xor  ( new_n31177_, new_n31176_, new_n9421_ );
or   ( new_n31178_, new_n31177_, new_n31173_ );
and  ( new_n31179_, new_n31178_, new_n31172_ );
or   ( new_n31180_, new_n31179_, new_n31167_ );
and  ( new_n31181_, new_n31179_, new_n31167_ );
or   ( new_n31182_, new_n7184_, new_n21792_ );
or   ( new_n31183_, new_n7186_, new_n21751_ );
and  ( new_n31184_, new_n31183_, new_n31182_ );
xor  ( new_n31185_, new_n31184_, new_n6638_ );
or   ( new_n31186_, new_n6645_, new_n21840_ );
or   ( new_n31187_, new_n6647_, new_n21842_ );
and  ( new_n31188_, new_n31187_, new_n31186_ );
xor  ( new_n31189_, new_n31188_, new_n6166_ );
nor  ( new_n31190_, new_n31189_, new_n31185_ );
and  ( new_n31191_, new_n31189_, new_n31185_ );
or   ( new_n31192_, new_n6173_, new_n22098_ );
or   ( new_n31193_, new_n6175_, new_n21847_ );
and  ( new_n31194_, new_n31193_, new_n31192_ );
xor  ( new_n31195_, new_n31194_, new_n5597_ );
nor  ( new_n31196_, new_n31195_, new_n31191_ );
nor  ( new_n31197_, new_n31196_, new_n31190_ );
or   ( new_n31198_, new_n31197_, new_n31181_ );
and  ( new_n31199_, new_n31198_, new_n31180_ );
or   ( new_n31200_, new_n2122_, new_n24927_ );
or   ( new_n31201_, new_n2124_, new_n24543_ );
and  ( new_n31202_, new_n31201_, new_n31200_ );
xor  ( new_n31203_, new_n31202_, new_n1843_ );
or   ( new_n31204_, new_n1844_, new_n25048_ );
or   ( new_n31205_, new_n1846_, new_n24925_ );
and  ( new_n31206_, new_n31205_, new_n31204_ );
xor  ( new_n31207_, new_n31206_, new_n1586_ );
or   ( new_n31208_, new_n31207_, new_n31203_ );
and  ( new_n31209_, new_n31207_, new_n31203_ );
or   ( new_n31210_, new_n1593_, new_n25486_ );
or   ( new_n31211_, new_n1595_, new_n25288_ );
and  ( new_n31212_, new_n31211_, new_n31210_ );
xor  ( new_n31213_, new_n31212_, new_n1358_ );
or   ( new_n31214_, new_n31213_, new_n31209_ );
and  ( new_n31215_, new_n31214_, new_n31208_ );
or   ( new_n31216_, new_n1364_, new_n26196_ );
or   ( new_n31217_, new_n1366_, new_n25813_ );
and  ( new_n31218_, new_n31217_, new_n31216_ );
xor  ( new_n31219_, new_n31218_, new_n1129_ );
or   ( new_n31220_, new_n1135_, new_n26372_ );
or   ( new_n31221_, new_n1137_, new_n26063_ );
and  ( new_n31222_, new_n31221_, new_n31220_ );
xor  ( new_n31223_, new_n31222_, new_n896_ );
or   ( new_n31224_, new_n31223_, new_n31219_ );
and  ( new_n31225_, new_n31223_, new_n31219_ );
or   ( new_n31226_, new_n897_, new_n26762_ );
or   ( new_n31227_, new_n899_, new_n26620_ );
and  ( new_n31228_, new_n31227_, new_n31226_ );
xor  ( new_n31229_, new_n31228_, new_n748_ );
or   ( new_n31230_, new_n31229_, new_n31225_ );
and  ( new_n31231_, new_n31230_, new_n31224_ );
or   ( new_n31232_, new_n31231_, new_n31215_ );
and  ( new_n31233_, new_n31231_, new_n31215_ );
or   ( new_n31234_, new_n755_, new_n27396_ );
or   ( new_n31235_, new_n757_, new_n27085_ );
and  ( new_n31236_, new_n31235_, new_n31234_ );
xor  ( new_n31237_, new_n31236_, new_n523_ );
or   ( new_n31238_, new_n524_, new_n27763_ );
or   ( new_n31239_, new_n526_, new_n27602_ );
and  ( new_n31240_, new_n31239_, new_n31238_ );
xor  ( new_n31241_, new_n31240_, new_n403_ );
nor  ( new_n31242_, new_n31241_, new_n31237_ );
and  ( new_n31243_, new_n31241_, new_n31237_ );
or   ( new_n31244_, new_n409_, new_n28314_ );
or   ( new_n31245_, new_n411_, new_n28108_ );
and  ( new_n31246_, new_n31245_, new_n31244_ );
xor  ( new_n31247_, new_n31246_, new_n328_ );
nor  ( new_n31248_, new_n31247_, new_n31243_ );
nor  ( new_n31249_, new_n31248_, new_n31242_ );
or   ( new_n31250_, new_n31249_, new_n31233_ );
and  ( new_n31251_, new_n31250_, new_n31232_ );
or   ( new_n31252_, new_n31251_, new_n31199_ );
or   ( new_n31253_, new_n3117_, new_n23733_ );
or   ( new_n31254_, new_n3119_, new_n23554_ );
and  ( new_n31255_, new_n31254_, new_n31253_ );
xor  ( new_n31256_, new_n31255_, new_n2800_ );
or   ( new_n31257_, new_n2807_, new_n24006_ );
or   ( new_n31258_, new_n2809_, new_n23895_ );
and  ( new_n31259_, new_n31258_, new_n31257_ );
xor  ( new_n31260_, new_n31259_, new_n2424_ );
or   ( new_n31261_, new_n31260_, new_n31256_ );
and  ( new_n31262_, new_n31260_, new_n31256_ );
or   ( new_n31263_, new_n2425_, new_n24418_ );
or   ( new_n31264_, new_n2427_, new_n24227_ );
and  ( new_n31265_, new_n31264_, new_n31263_ );
xor  ( new_n31266_, new_n31265_, new_n2121_ );
or   ( new_n31267_, new_n31266_, new_n31262_ );
and  ( new_n31268_, new_n31267_, new_n31261_ );
or   ( new_n31269_, new_n4302_, new_n22975_ );
or   ( new_n31270_, new_n4304_, new_n22829_ );
and  ( new_n31271_, new_n31270_, new_n31269_ );
xor  ( new_n31272_, new_n31271_, new_n3895_ );
or   ( new_n31273_, new_n3896_, new_n23166_ );
or   ( new_n31274_, new_n3898_, new_n22973_ );
and  ( new_n31275_, new_n31274_, new_n31273_ );
xor  ( new_n31276_, new_n31275_, new_n3460_ );
or   ( new_n31277_, new_n31276_, new_n31272_ );
and  ( new_n31278_, new_n31276_, new_n31272_ );
or   ( new_n31279_, new_n3461_, new_n23370_ );
or   ( new_n31280_, new_n3463_, new_n23252_ );
and  ( new_n31281_, new_n31280_, new_n31279_ );
xor  ( new_n31282_, new_n31281_, new_n3116_ );
or   ( new_n31283_, new_n31282_, new_n31278_ );
and  ( new_n31284_, new_n31283_, new_n31277_ );
nor  ( new_n31285_, new_n31284_, new_n31268_ );
and  ( new_n31286_, new_n31284_, new_n31268_ );
or   ( new_n31287_, new_n5604_, new_n22207_ );
or   ( new_n31288_, new_n5606_, new_n22129_ );
and  ( new_n31289_, new_n31288_, new_n31287_ );
xor  ( new_n31290_, new_n31289_, new_n5206_ );
or   ( new_n31291_, new_n5207_, new_n22423_ );
or   ( new_n31292_, new_n5209_, new_n22304_ );
and  ( new_n31293_, new_n31292_, new_n31291_ );
xor  ( new_n31294_, new_n31293_, new_n4708_ );
nor  ( new_n31295_, new_n31294_, new_n31290_ );
and  ( new_n31296_, new_n31294_, new_n31290_ );
or   ( new_n31297_, new_n4709_, new_n22641_ );
or   ( new_n31298_, new_n4711_, new_n22590_ );
and  ( new_n31299_, new_n31298_, new_n31297_ );
xor  ( new_n31300_, new_n31299_, new_n4295_ );
nor  ( new_n31301_, new_n31300_, new_n31296_ );
nor  ( new_n31302_, new_n31301_, new_n31295_ );
nor  ( new_n31303_, new_n31302_, new_n31286_ );
nor  ( new_n31304_, new_n31303_, new_n31285_ );
and  ( new_n31305_, new_n31251_, new_n31199_ );
or   ( new_n31306_, new_n31305_, new_n31304_ );
and  ( new_n31307_, new_n31306_, new_n31252_ );
and  ( new_n31308_, new_n31307_, new_n31151_ );
nor  ( new_n31309_, new_n31307_, new_n31151_ );
xnor ( new_n31310_, new_n30804_, new_n30803_ );
or   ( new_n31311_, new_n337_, new_n29263_ );
or   ( new_n31312_, new_n340_, new_n28531_ );
and  ( new_n31313_, new_n31312_, new_n31311_ );
xor  ( new_n31314_, new_n31313_, new_n332_ );
or   ( new_n31315_, new_n317_, new_n29474_ );
or   ( new_n31316_, new_n320_, new_n29261_ );
and  ( new_n31317_, new_n31316_, new_n31315_ );
xor  ( new_n31318_, new_n31317_, new_n312_ );
or   ( new_n31319_, new_n31318_, new_n31314_ );
and  ( new_n31320_, new_n31318_, new_n31314_ );
or   ( new_n31321_, new_n283_, new_n30120_ );
or   ( new_n31322_, new_n286_, new_n29619_ );
and  ( new_n31323_, new_n31322_, new_n31321_ );
xor  ( new_n31324_, new_n31323_, new_n278_ );
or   ( new_n31325_, new_n31324_, new_n31320_ );
and  ( new_n31326_, new_n31325_, new_n31319_ );
nor  ( new_n31327_, new_n31326_, new_n31310_ );
and  ( new_n31328_, new_n31326_, new_n31310_ );
or   ( new_n31329_, new_n299_, new_n30800_ );
or   ( new_n31330_, new_n302_, new_n30227_ );
and  ( new_n31331_, new_n31330_, new_n31329_ );
xor  ( new_n31332_, new_n31331_, new_n293_ );
not  ( new_n31333_, RIbb33288_190 );
or   ( new_n31334_, new_n268_, new_n31333_ );
or   ( new_n31335_, new_n271_, new_n30798_ );
and  ( new_n31336_, new_n31335_, new_n31334_ );
xor  ( new_n31337_, new_n31336_, new_n263_ );
nor  ( new_n31338_, new_n31337_, new_n31332_ );
and  ( new_n31339_, RIbb33300_191, RIbb2f610_1 );
and  ( new_n31340_, new_n31337_, new_n31332_ );
nor  ( new_n31341_, new_n31340_, new_n31339_ );
nor  ( new_n31342_, new_n31341_, new_n31338_ );
nor  ( new_n31343_, new_n31342_, new_n31328_ );
or   ( new_n31344_, new_n31343_, new_n31327_ );
xnor ( new_n31345_, new_n30963_, new_n30959_ );
xor  ( new_n31346_, new_n31345_, new_n30969_ );
xnor ( new_n31347_, new_n30997_, new_n30993_ );
xor  ( new_n31348_, new_n31347_, new_n31003_ );
or   ( new_n31349_, new_n31348_, new_n31346_ );
and  ( new_n31350_, new_n31348_, new_n31346_ );
xor  ( new_n31351_, new_n30910_, new_n30906_ );
xnor ( new_n31352_, new_n31351_, new_n30916_ );
or   ( new_n31353_, new_n31352_, new_n31350_ );
and  ( new_n31354_, new_n31353_, new_n31349_ );
nor  ( new_n31355_, new_n31354_, new_n31344_ );
and  ( new_n31356_, new_n31354_, new_n31344_ );
xnor ( new_n31357_, new_n30926_, new_n30922_ );
xor  ( new_n31358_, new_n31357_, new_n30932_ );
xnor ( new_n31359_, new_n30813_, new_n30809_ );
xor  ( new_n31360_, new_n31359_, new_n30819_ );
nor  ( new_n31361_, new_n31360_, new_n31358_ );
and  ( new_n31362_, new_n31360_, new_n31358_ );
xor  ( new_n31363_, new_n30944_, new_n30940_ );
xnor ( new_n31364_, new_n31363_, new_n30950_ );
nor  ( new_n31365_, new_n31364_, new_n31362_ );
nor  ( new_n31366_, new_n31365_, new_n31361_ );
nor  ( new_n31367_, new_n31366_, new_n31356_ );
nor  ( new_n31368_, new_n31367_, new_n31355_ );
nor  ( new_n31369_, new_n31368_, new_n31309_ );
nor  ( new_n31370_, new_n31369_, new_n31308_ );
or   ( new_n31371_, new_n31370_, new_n31134_ );
and  ( new_n31372_, new_n31371_, new_n31133_ );
or   ( new_n31373_, new_n31372_, new_n31095_ );
and  ( new_n31374_, new_n31373_, new_n31094_ );
xor  ( new_n31375_, new_n30694_, new_n30647_ );
xor  ( new_n31376_, new_n31375_, new_n30715_ );
xor  ( new_n31377_, new_n31037_, new_n30797_ );
xor  ( new_n31378_, new_n31377_, new_n31049_ );
or   ( new_n31379_, new_n31378_, new_n31376_ );
and  ( new_n31380_, new_n31378_, new_n31376_ );
xor  ( new_n31381_, new_n31057_, new_n31055_ );
xnor ( new_n31382_, new_n31381_, new_n31061_ );
not  ( new_n31383_, new_n31382_ );
or   ( new_n31384_, new_n31383_, new_n31380_ );
and  ( new_n31385_, new_n31384_, new_n31379_ );
nor  ( new_n31386_, new_n31385_, new_n31374_ );
and  ( new_n31387_, new_n31385_, new_n31374_ );
xor  ( new_n31388_, new_n30717_, new_n30490_ );
xor  ( new_n31389_, new_n31388_, new_n30730_ );
nor  ( new_n31390_, new_n31389_, new_n31387_ );
nor  ( new_n31391_, new_n31390_, new_n31386_ );
xnor ( new_n31392_, new_n31067_, new_n31065_ );
xnor ( new_n31393_, new_n31392_, new_n31071_ );
nor  ( new_n31394_, new_n31393_, new_n31391_ );
xnor ( new_n31395_, new_n31073_, new_n30769_ );
xor  ( new_n31396_, new_n31395_, new_n31077_ );
and  ( new_n31397_, new_n31396_, new_n31394_ );
xnor ( new_n31398_, new_n31393_, new_n31391_ );
xor  ( new_n31399_, new_n31385_, new_n31374_ );
xor  ( new_n31400_, new_n31399_, new_n31389_ );
xor  ( new_n31401_, new_n31010_, new_n30852_ );
xor  ( new_n31402_, new_n31401_, new_n31035_ );
xor  ( new_n31403_, new_n30954_, new_n30902_ );
xor  ( new_n31404_, new_n31403_, new_n31007_ );
xnor ( new_n31405_, new_n31107_, new_n31105_ );
xor  ( new_n31406_, new_n31405_, new_n31119_ );
nand ( new_n31407_, new_n31406_, new_n31404_ );
nor  ( new_n31408_, new_n31406_, new_n31404_ );
xor  ( new_n31409_, new_n31125_, new_n31123_ );
xor  ( new_n31410_, new_n31409_, new_n31130_ );
or   ( new_n31411_, new_n31410_, new_n31408_ );
and  ( new_n31412_, new_n31411_, new_n31407_ );
or   ( new_n31413_, new_n31412_, new_n31402_ );
and  ( new_n31414_, new_n31412_, new_n31402_ );
xor  ( new_n31415_, new_n31099_, new_n31097_ );
xor  ( new_n31416_, new_n31415_, new_n31103_ );
xnor ( new_n31417_, new_n31354_, new_n31344_ );
xor  ( new_n31418_, new_n31417_, new_n31366_ );
or   ( new_n31419_, new_n31418_, new_n31416_ );
and  ( new_n31420_, new_n31418_, new_n31416_ );
xor  ( new_n31421_, new_n31146_, new_n31136_ );
xor  ( new_n31422_, new_n31421_, new_n31149_ );
or   ( new_n31423_, new_n31422_, new_n31420_ );
and  ( new_n31424_, new_n31423_, new_n31419_ );
xnor ( new_n31425_, new_n31140_, new_n31138_ );
xor  ( new_n31426_, new_n31425_, new_n31144_ );
xnor ( new_n31427_, new_n31348_, new_n31346_ );
xor  ( new_n31428_, new_n31427_, new_n31352_ );
or   ( new_n31429_, new_n31428_, new_n31426_ );
and  ( new_n31430_, new_n31428_, new_n31426_ );
xor  ( new_n31431_, new_n31360_, new_n31358_ );
xnor ( new_n31432_, new_n31431_, new_n31364_ );
or   ( new_n31433_, new_n31432_, new_n31430_ );
and  ( new_n31434_, new_n31433_, new_n31429_ );
xnor ( new_n31435_, new_n31113_, new_n31111_ );
xor  ( new_n31436_, new_n31435_, new_n31117_ );
or   ( new_n31437_, new_n31436_, new_n31434_ );
nand ( new_n31438_, new_n31436_, new_n31434_ );
xnor ( new_n31439_, new_n31231_, new_n31215_ );
xor  ( new_n31440_, new_n31439_, new_n31249_ );
xnor ( new_n31441_, new_n31284_, new_n31268_ );
xor  ( new_n31442_, new_n31441_, new_n31302_ );
nor  ( new_n31443_, new_n31442_, new_n31440_ );
and  ( new_n31444_, new_n31442_, new_n31440_ );
xor  ( new_n31445_, new_n31326_, new_n31310_ );
xor  ( new_n31446_, new_n31445_, new_n31342_ );
not  ( new_n31447_, new_n31446_ );
nor  ( new_n31448_, new_n31447_, new_n31444_ );
nor  ( new_n31449_, new_n31448_, new_n31443_ );
nand ( new_n31450_, new_n31449_, new_n31438_ );
and  ( new_n31451_, new_n31450_, new_n31437_ );
and  ( new_n31452_, new_n31451_, new_n31424_ );
nor  ( new_n31453_, new_n31451_, new_n31424_ );
xor  ( new_n31454_, new_n31159_, new_n31155_ );
xnor ( new_n31455_, new_n31454_, new_n31165_ );
xor  ( new_n31456_, new_n31171_, RIbb2d900_63 );
xor  ( new_n31457_, new_n31456_, new_n31177_ );
or   ( new_n31458_, new_n31457_, new_n31455_ );
xnor ( new_n31459_, new_n31276_, new_n31272_ );
xor  ( new_n31460_, new_n31459_, new_n31282_ );
xnor ( new_n31461_, new_n31189_, new_n31185_ );
xor  ( new_n31462_, new_n31461_, new_n31195_ );
or   ( new_n31463_, new_n31462_, new_n31460_ );
and  ( new_n31464_, new_n31462_, new_n31460_ );
xnor ( new_n31465_, new_n31294_, new_n31290_ );
xor  ( new_n31466_, new_n31465_, new_n31300_ );
or   ( new_n31467_, new_n31466_, new_n31464_ );
and  ( new_n31468_, new_n31467_, new_n31463_ );
nor  ( new_n31469_, new_n31468_, new_n31458_ );
and  ( new_n31470_, new_n31468_, new_n31458_ );
xor  ( new_n31471_, new_n30858_, new_n30856_ );
xnor ( new_n31472_, new_n31471_, new_n30864_ );
nor  ( new_n31473_, new_n31472_, new_n31470_ );
or   ( new_n31474_, new_n31473_, new_n31469_ );
or   ( new_n31475_, new_n897_, new_n27085_ );
or   ( new_n31476_, new_n899_, new_n26762_ );
and  ( new_n31477_, new_n31476_, new_n31475_ );
xor  ( new_n31478_, new_n31477_, new_n748_ );
or   ( new_n31479_, new_n755_, new_n27602_ );
or   ( new_n31480_, new_n757_, new_n27396_ );
and  ( new_n31481_, new_n31480_, new_n31479_ );
xor  ( new_n31482_, new_n31481_, new_n523_ );
or   ( new_n31483_, new_n31482_, new_n31478_ );
and  ( new_n31484_, new_n31482_, new_n31478_ );
or   ( new_n31485_, new_n524_, new_n28108_ );
or   ( new_n31486_, new_n526_, new_n27763_ );
and  ( new_n31487_, new_n31486_, new_n31485_ );
xor  ( new_n31488_, new_n31487_, new_n403_ );
or   ( new_n31489_, new_n31488_, new_n31484_ );
and  ( new_n31490_, new_n31489_, new_n31483_ );
or   ( new_n31491_, new_n1593_, new_n25813_ );
or   ( new_n31492_, new_n1595_, new_n25486_ );
and  ( new_n31493_, new_n31492_, new_n31491_ );
xor  ( new_n31494_, new_n31493_, new_n1358_ );
or   ( new_n31495_, new_n1364_, new_n26063_ );
or   ( new_n31496_, new_n1366_, new_n26196_ );
and  ( new_n31497_, new_n31496_, new_n31495_ );
xor  ( new_n31498_, new_n31497_, new_n1129_ );
or   ( new_n31499_, new_n31498_, new_n31494_ );
and  ( new_n31500_, new_n31498_, new_n31494_ );
or   ( new_n31501_, new_n1135_, new_n26620_ );
or   ( new_n31502_, new_n1137_, new_n26372_ );
and  ( new_n31503_, new_n31502_, new_n31501_ );
xor  ( new_n31504_, new_n31503_, new_n896_ );
or   ( new_n31505_, new_n31504_, new_n31500_ );
and  ( new_n31506_, new_n31505_, new_n31499_ );
or   ( new_n31507_, new_n31506_, new_n31490_ );
and  ( new_n31508_, new_n31506_, new_n31490_ );
or   ( new_n31509_, new_n2425_, new_n24543_ );
or   ( new_n31510_, new_n2427_, new_n24418_ );
and  ( new_n31511_, new_n31510_, new_n31509_ );
xor  ( new_n31512_, new_n31511_, new_n2121_ );
or   ( new_n31513_, new_n2122_, new_n24925_ );
or   ( new_n31514_, new_n2124_, new_n24927_ );
and  ( new_n31515_, new_n31514_, new_n31513_ );
xor  ( new_n31516_, new_n31515_, new_n1843_ );
nor  ( new_n31517_, new_n31516_, new_n31512_ );
and  ( new_n31518_, new_n31516_, new_n31512_ );
or   ( new_n31519_, new_n1844_, new_n25288_ );
or   ( new_n31520_, new_n1846_, new_n25048_ );
and  ( new_n31521_, new_n31520_, new_n31519_ );
xor  ( new_n31522_, new_n31521_, new_n1586_ );
nor  ( new_n31523_, new_n31522_, new_n31518_ );
nor  ( new_n31524_, new_n31523_, new_n31517_ );
or   ( new_n31525_, new_n31524_, new_n31508_ );
and  ( new_n31526_, new_n31525_, new_n31507_ );
or   ( new_n31527_, new_n3461_, new_n23554_ );
or   ( new_n31528_, new_n3463_, new_n23370_ );
and  ( new_n31529_, new_n31528_, new_n31527_ );
xor  ( new_n31530_, new_n31529_, new_n3116_ );
or   ( new_n31531_, new_n3117_, new_n23895_ );
or   ( new_n31532_, new_n3119_, new_n23733_ );
and  ( new_n31533_, new_n31532_, new_n31531_ );
xor  ( new_n31534_, new_n31533_, new_n2800_ );
or   ( new_n31535_, new_n31534_, new_n31530_ );
and  ( new_n31536_, new_n31534_, new_n31530_ );
or   ( new_n31537_, new_n2807_, new_n24227_ );
or   ( new_n31538_, new_n2809_, new_n24006_ );
and  ( new_n31539_, new_n31538_, new_n31537_ );
xor  ( new_n31540_, new_n31539_, new_n2424_ );
or   ( new_n31541_, new_n31540_, new_n31536_ );
and  ( new_n31542_, new_n31541_, new_n31535_ );
or   ( new_n31543_, new_n4709_, new_n22829_ );
or   ( new_n31544_, new_n4711_, new_n22641_ );
and  ( new_n31545_, new_n31544_, new_n31543_ );
xor  ( new_n31546_, new_n31545_, new_n4295_ );
or   ( new_n31547_, new_n4302_, new_n22973_ );
or   ( new_n31548_, new_n4304_, new_n22975_ );
and  ( new_n31549_, new_n31548_, new_n31547_ );
xor  ( new_n31550_, new_n31549_, new_n3895_ );
or   ( new_n31551_, new_n31550_, new_n31546_ );
and  ( new_n31552_, new_n31550_, new_n31546_ );
or   ( new_n31553_, new_n3896_, new_n23252_ );
or   ( new_n31554_, new_n3898_, new_n23166_ );
and  ( new_n31555_, new_n31554_, new_n31553_ );
xor  ( new_n31556_, new_n31555_, new_n3460_ );
or   ( new_n31557_, new_n31556_, new_n31552_ );
and  ( new_n31558_, new_n31557_, new_n31551_ );
or   ( new_n31559_, new_n31558_, new_n31542_ );
and  ( new_n31560_, new_n31558_, new_n31542_ );
or   ( new_n31561_, new_n6173_, new_n22129_ );
or   ( new_n31562_, new_n6175_, new_n22098_ );
and  ( new_n31563_, new_n31562_, new_n31561_ );
xor  ( new_n31564_, new_n31563_, new_n5597_ );
or   ( new_n31565_, new_n5604_, new_n22304_ );
or   ( new_n31566_, new_n5606_, new_n22207_ );
and  ( new_n31567_, new_n31566_, new_n31565_ );
xor  ( new_n31568_, new_n31567_, new_n5206_ );
nor  ( new_n31569_, new_n31568_, new_n31564_ );
and  ( new_n31570_, new_n31568_, new_n31564_ );
or   ( new_n31571_, new_n5207_, new_n22590_ );
or   ( new_n31572_, new_n5209_, new_n22423_ );
and  ( new_n31573_, new_n31572_, new_n31571_ );
xor  ( new_n31574_, new_n31573_, new_n4708_ );
nor  ( new_n31575_, new_n31574_, new_n31570_ );
nor  ( new_n31576_, new_n31575_, new_n31569_ );
or   ( new_n31577_, new_n31576_, new_n31560_ );
and  ( new_n31578_, new_n31577_, new_n31559_ );
or   ( new_n31579_, new_n31578_, new_n31526_ );
and  ( new_n31580_, new_n31578_, new_n31526_ );
or   ( new_n31581_, new_n9422_, new_n21674_ );
or   ( new_n31582_, new_n9424_, new_n21701_ );
and  ( new_n31583_, new_n31582_, new_n31581_ );
xor  ( new_n31584_, new_n31583_, new_n8873_ );
or   ( new_n31585_, new_n8874_, new_n21680_ );
or   ( new_n31586_, new_n8876_, new_n21672_ );
and  ( new_n31587_, new_n31586_, new_n31585_ );
xor  ( new_n31588_, new_n31587_, new_n8257_ );
nor  ( new_n31589_, new_n31588_, new_n31584_ );
and  ( new_n31590_, new_n31588_, new_n31584_ );
or   ( new_n31591_, new_n8264_, new_n21687_ );
or   ( new_n31592_, new_n8266_, new_n21678_ );
and  ( new_n31593_, new_n31592_, new_n31591_ );
xor  ( new_n31594_, new_n31593_, new_n7725_ );
nor  ( new_n31595_, new_n31594_, new_n31590_ );
nor  ( new_n31596_, new_n31595_, new_n31589_ );
or   ( new_n31597_, new_n10059_, new_n21703_ );
or   ( new_n31598_, new_n10061_, new_n21694_ );
and  ( new_n31599_, new_n31598_, new_n31597_ );
xor  ( new_n31600_, new_n31599_, new_n9421_ );
or   ( new_n31601_, new_n21696_, RIbb2d888_64 );
and  ( new_n31602_, new_n31601_, RIbb2d900_63 );
and  ( new_n31603_, new_n31602_, new_n31600_ );
or   ( new_n31604_, new_n7732_, new_n21751_ );
or   ( new_n31605_, new_n7734_, new_n21685_ );
and  ( new_n31606_, new_n31605_, new_n31604_ );
xor  ( new_n31607_, new_n31606_, new_n7177_ );
or   ( new_n31608_, new_n7184_, new_n21842_ );
or   ( new_n31609_, new_n7186_, new_n21792_ );
and  ( new_n31610_, new_n31609_, new_n31608_ );
xor  ( new_n31611_, new_n31610_, new_n6638_ );
nor  ( new_n31612_, new_n31611_, new_n31607_ );
and  ( new_n31613_, new_n31611_, new_n31607_ );
or   ( new_n31614_, new_n6645_, new_n21847_ );
or   ( new_n31615_, new_n6647_, new_n21840_ );
and  ( new_n31616_, new_n31615_, new_n31614_ );
xor  ( new_n31617_, new_n31616_, new_n6166_ );
nor  ( new_n31618_, new_n31617_, new_n31613_ );
nor  ( new_n31619_, new_n31618_, new_n31612_ );
and  ( new_n31620_, new_n31619_, new_n31603_ );
nor  ( new_n31621_, new_n31620_, new_n31596_ );
nor  ( new_n31622_, new_n31619_, new_n31603_ );
nor  ( new_n31623_, new_n31622_, new_n31621_ );
or   ( new_n31624_, new_n31623_, new_n31580_ );
and  ( new_n31625_, new_n31624_, new_n31579_ );
and  ( new_n31626_, new_n31625_, new_n31474_ );
nor  ( new_n31627_, new_n31625_, new_n31474_ );
or   ( new_n31628_, new_n409_, new_n28531_ );
or   ( new_n31629_, new_n411_, new_n28314_ );
and  ( new_n31630_, new_n31629_, new_n31628_ );
xor  ( new_n31631_, new_n31630_, new_n328_ );
or   ( new_n31632_, new_n337_, new_n29261_ );
or   ( new_n31633_, new_n340_, new_n29263_ );
and  ( new_n31634_, new_n31633_, new_n31632_ );
xor  ( new_n31635_, new_n31634_, new_n332_ );
or   ( new_n31636_, new_n31635_, new_n31631_ );
and  ( new_n31637_, new_n31635_, new_n31631_ );
or   ( new_n31638_, new_n317_, new_n29619_ );
or   ( new_n31639_, new_n320_, new_n29474_ );
and  ( new_n31640_, new_n31639_, new_n31638_ );
xor  ( new_n31641_, new_n31640_, new_n312_ );
or   ( new_n31642_, new_n31641_, new_n31637_ );
and  ( new_n31643_, new_n31642_, new_n31636_ );
or   ( new_n31644_, new_n283_, new_n30227_ );
or   ( new_n31645_, new_n286_, new_n30120_ );
and  ( new_n31646_, new_n31645_, new_n31644_ );
xor  ( new_n31647_, new_n31646_, new_n278_ );
or   ( new_n31648_, new_n299_, new_n30798_ );
or   ( new_n31649_, new_n302_, new_n30800_ );
and  ( new_n31650_, new_n31649_, new_n31648_ );
xor  ( new_n31651_, new_n31650_, new_n293_ );
or   ( new_n31652_, new_n31651_, new_n31647_ );
and  ( new_n31653_, new_n31651_, new_n31647_ );
not  ( new_n31654_, RIbb33300_191 );
or   ( new_n31655_, new_n268_, new_n31654_ );
or   ( new_n31656_, new_n271_, new_n31333_ );
and  ( new_n31657_, new_n31656_, new_n31655_ );
xor  ( new_n31658_, new_n31657_, new_n263_ );
or   ( new_n31659_, new_n31658_, new_n31653_ );
and  ( new_n31660_, new_n31659_, new_n31652_ );
nor  ( new_n31661_, new_n31660_, new_n31643_ );
xnor ( new_n31662_, new_n31318_, new_n31314_ );
xor  ( new_n31663_, new_n31662_, new_n31324_ );
xnor ( new_n31664_, new_n31337_, new_n31332_ );
xor  ( new_n31665_, new_n31664_, new_n31339_ );
or   ( new_n31666_, new_n31665_, new_n31663_ );
and  ( new_n31667_, new_n31665_, new_n31663_ );
xor  ( new_n31668_, new_n31241_, new_n31237_ );
xnor ( new_n31669_, new_n31668_, new_n31247_ );
or   ( new_n31670_, new_n31669_, new_n31667_ );
and  ( new_n31671_, new_n31670_, new_n31666_ );
nor  ( new_n31672_, new_n31671_, new_n31661_ );
and  ( new_n31673_, new_n31671_, new_n31661_ );
xnor ( new_n31674_, new_n31223_, new_n31219_ );
xor  ( new_n31675_, new_n31674_, new_n31229_ );
xnor ( new_n31676_, new_n31207_, new_n31203_ );
xor  ( new_n31677_, new_n31676_, new_n31213_ );
nor  ( new_n31678_, new_n31677_, new_n31675_ );
and  ( new_n31679_, new_n31677_, new_n31675_ );
xor  ( new_n31680_, new_n31260_, new_n31256_ );
xnor ( new_n31681_, new_n31680_, new_n31266_ );
nor  ( new_n31682_, new_n31681_, new_n31679_ );
nor  ( new_n31683_, new_n31682_, new_n31678_ );
nor  ( new_n31684_, new_n31683_, new_n31673_ );
nor  ( new_n31685_, new_n31684_, new_n31672_ );
nor  ( new_n31686_, new_n31685_, new_n31627_ );
nor  ( new_n31687_, new_n31686_, new_n31626_ );
nor  ( new_n31688_, new_n31687_, new_n31453_ );
nor  ( new_n31689_, new_n31688_, new_n31452_ );
or   ( new_n31690_, new_n31689_, new_n31414_ );
and  ( new_n31691_, new_n31690_, new_n31413_ );
xor  ( new_n31692_, new_n31093_, new_n31082_ );
xor  ( new_n31693_, new_n31692_, new_n31372_ );
or   ( new_n31694_, new_n31693_, new_n31691_ );
and  ( new_n31695_, new_n31693_, new_n31691_ );
xor  ( new_n31696_, new_n31378_, new_n31376_ );
xor  ( new_n31697_, new_n31696_, new_n31383_ );
or   ( new_n31698_, new_n31697_, new_n31695_ );
and  ( new_n31699_, new_n31698_, new_n31694_ );
or   ( new_n31700_, new_n31699_, new_n31400_ );
and  ( new_n31701_, new_n31699_, new_n31400_ );
xor  ( new_n31702_, new_n31051_, new_n30771_ );
xor  ( new_n31703_, new_n31702_, new_n31063_ );
or   ( new_n31704_, new_n31703_, new_n31701_ );
and  ( new_n31705_, new_n31704_, new_n31700_ );
nor  ( new_n31706_, new_n31705_, new_n31398_ );
xor  ( new_n31707_, new_n31699_, new_n31400_ );
xor  ( new_n31708_, new_n31707_, new_n31703_ );
xor  ( new_n31709_, new_n31132_, new_n31121_ );
xnor ( new_n31710_, new_n31709_, new_n31370_ );
xnor ( new_n31711_, new_n31412_, new_n31402_ );
xor  ( new_n31712_, new_n31711_, new_n31689_ );
nand ( new_n31713_, new_n31712_, new_n31710_ );
xor  ( new_n31714_, new_n31451_, new_n31424_ );
xnor ( new_n31715_, new_n31714_, new_n31687_ );
xnor ( new_n31716_, new_n31406_, new_n31404_ );
xor  ( new_n31717_, new_n31716_, new_n31410_ );
and  ( new_n31718_, new_n31717_, new_n31715_ );
xor  ( new_n31719_, new_n31307_, new_n31151_ );
xor  ( new_n31720_, new_n31719_, new_n31368_ );
xnor ( new_n31721_, new_n31251_, new_n31199_ );
xor  ( new_n31722_, new_n31721_, new_n31304_ );
xor  ( new_n31723_, new_n31436_, new_n31434_ );
xor  ( new_n31724_, new_n31723_, new_n31449_ );
or   ( new_n31725_, new_n31724_, new_n31722_ );
and  ( new_n31726_, new_n31724_, new_n31722_ );
xnor ( new_n31727_, new_n31418_, new_n31416_ );
xor  ( new_n31728_, new_n31727_, new_n31422_ );
or   ( new_n31729_, new_n31728_, new_n31726_ );
and  ( new_n31730_, new_n31729_, new_n31725_ );
nand ( new_n31731_, new_n31730_, new_n31720_ );
or   ( new_n31732_, new_n31730_, new_n31720_ );
xnor ( new_n31733_, new_n31677_, new_n31675_ );
xor  ( new_n31734_, new_n31733_, new_n31681_ );
xnor ( new_n31735_, new_n31665_, new_n31663_ );
xor  ( new_n31736_, new_n31735_, new_n31669_ );
nor  ( new_n31737_, new_n31736_, new_n31734_ );
nand ( new_n31738_, new_n31736_, new_n31734_ );
xor  ( new_n31739_, new_n31660_, new_n31643_ );
and  ( new_n31740_, new_n31739_, new_n31738_ );
or   ( new_n31741_, new_n31740_, new_n31737_ );
xnor ( new_n31742_, new_n31179_, new_n31167_ );
xor  ( new_n31743_, new_n31742_, new_n31197_ );
or   ( new_n31744_, new_n31743_, new_n31741_ );
and  ( new_n31745_, new_n31743_, new_n31741_ );
xnor ( new_n31746_, new_n31506_, new_n31490_ );
xor  ( new_n31747_, new_n31746_, new_n31524_ );
xnor ( new_n31748_, new_n31558_, new_n31542_ );
xor  ( new_n31749_, new_n31748_, new_n31576_ );
nor  ( new_n31750_, new_n31749_, new_n31747_ );
and  ( new_n31751_, new_n31749_, new_n31747_ );
xnor ( new_n31752_, new_n31619_, new_n31603_ );
xnor ( new_n31753_, new_n31752_, new_n31596_ );
not  ( new_n31754_, new_n31753_ );
nor  ( new_n31755_, new_n31754_, new_n31751_ );
nor  ( new_n31756_, new_n31755_, new_n31750_ );
or   ( new_n31757_, new_n31756_, new_n31745_ );
and  ( new_n31758_, new_n31757_, new_n31744_ );
xor  ( new_n31759_, new_n31468_, new_n31458_ );
xor  ( new_n31760_, new_n31759_, new_n31472_ );
xnor ( new_n31761_, new_n31428_, new_n31426_ );
xor  ( new_n31762_, new_n31761_, new_n31432_ );
or   ( new_n31763_, new_n31762_, new_n31760_ );
and  ( new_n31764_, new_n31762_, new_n31760_ );
xor  ( new_n31765_, new_n31442_, new_n31440_ );
xor  ( new_n31766_, new_n31765_, new_n31447_ );
or   ( new_n31767_, new_n31766_, new_n31764_ );
and  ( new_n31768_, new_n31767_, new_n31763_ );
nor  ( new_n31769_, new_n31768_, new_n31758_ );
and  ( new_n31770_, new_n31768_, new_n31758_ );
xor  ( new_n31771_, new_n31462_, new_n31460_ );
xor  ( new_n31772_, new_n31771_, new_n31466_ );
xnor ( new_n31773_, new_n31588_, new_n31584_ );
xor  ( new_n31774_, new_n31773_, new_n31594_ );
xnor ( new_n31775_, new_n31611_, new_n31607_ );
xor  ( new_n31776_, new_n31775_, new_n31617_ );
or   ( new_n31777_, new_n31776_, new_n31774_ );
and  ( new_n31778_, new_n31776_, new_n31774_ );
xor  ( new_n31779_, new_n31568_, new_n31564_ );
xnor ( new_n31780_, new_n31779_, new_n31574_ );
or   ( new_n31781_, new_n31780_, new_n31778_ );
and  ( new_n31782_, new_n31781_, new_n31777_ );
nor  ( new_n31783_, new_n31782_, new_n31772_ );
nand ( new_n31784_, new_n31782_, new_n31772_ );
xor  ( new_n31785_, new_n31457_, new_n31455_ );
and  ( new_n31786_, new_n31785_, new_n31784_ );
or   ( new_n31787_, new_n31786_, new_n31783_ );
or   ( new_n31788_, new_n5604_, new_n22423_ );
or   ( new_n31789_, new_n5606_, new_n22304_ );
and  ( new_n31790_, new_n31789_, new_n31788_ );
xor  ( new_n31791_, new_n31790_, new_n5206_ );
or   ( new_n31792_, new_n5207_, new_n22641_ );
or   ( new_n31793_, new_n5209_, new_n22590_ );
and  ( new_n31794_, new_n31793_, new_n31792_ );
xor  ( new_n31795_, new_n31794_, new_n4708_ );
or   ( new_n31796_, new_n31795_, new_n31791_ );
and  ( new_n31797_, new_n31795_, new_n31791_ );
or   ( new_n31798_, new_n4709_, new_n22975_ );
or   ( new_n31799_, new_n4711_, new_n22829_ );
and  ( new_n31800_, new_n31799_, new_n31798_ );
xor  ( new_n31801_, new_n31800_, new_n4295_ );
or   ( new_n31802_, new_n31801_, new_n31797_ );
and  ( new_n31803_, new_n31802_, new_n31796_ );
or   ( new_n31804_, new_n4302_, new_n23166_ );
or   ( new_n31805_, new_n4304_, new_n22973_ );
and  ( new_n31806_, new_n31805_, new_n31804_ );
xor  ( new_n31807_, new_n31806_, new_n3895_ );
or   ( new_n31808_, new_n3896_, new_n23370_ );
or   ( new_n31809_, new_n3898_, new_n23252_ );
and  ( new_n31810_, new_n31809_, new_n31808_ );
xor  ( new_n31811_, new_n31810_, new_n3460_ );
or   ( new_n31812_, new_n31811_, new_n31807_ );
and  ( new_n31813_, new_n31811_, new_n31807_ );
or   ( new_n31814_, new_n3461_, new_n23733_ );
or   ( new_n31815_, new_n3463_, new_n23554_ );
and  ( new_n31816_, new_n31815_, new_n31814_ );
xor  ( new_n31817_, new_n31816_, new_n3116_ );
or   ( new_n31818_, new_n31817_, new_n31813_ );
and  ( new_n31819_, new_n31818_, new_n31812_ );
or   ( new_n31820_, new_n31819_, new_n31803_ );
and  ( new_n31821_, new_n31819_, new_n31803_ );
or   ( new_n31822_, new_n3117_, new_n24006_ );
or   ( new_n31823_, new_n3119_, new_n23895_ );
and  ( new_n31824_, new_n31823_, new_n31822_ );
xor  ( new_n31825_, new_n31824_, new_n2800_ );
or   ( new_n31826_, new_n2807_, new_n24418_ );
or   ( new_n31827_, new_n2809_, new_n24227_ );
and  ( new_n31828_, new_n31827_, new_n31826_ );
xor  ( new_n31829_, new_n31828_, new_n2424_ );
nor  ( new_n31830_, new_n31829_, new_n31825_ );
and  ( new_n31831_, new_n31829_, new_n31825_ );
or   ( new_n31832_, new_n2425_, new_n24927_ );
or   ( new_n31833_, new_n2427_, new_n24543_ );
and  ( new_n31834_, new_n31833_, new_n31832_ );
xor  ( new_n31835_, new_n31834_, new_n2121_ );
nor  ( new_n31836_, new_n31835_, new_n31831_ );
nor  ( new_n31837_, new_n31836_, new_n31830_ );
or   ( new_n31838_, new_n31837_, new_n31821_ );
and  ( new_n31839_, new_n31838_, new_n31820_ );
or   ( new_n31840_, new_n8874_, new_n21678_ );
or   ( new_n31841_, new_n8876_, new_n21680_ );
and  ( new_n31842_, new_n31841_, new_n31840_ );
xor  ( new_n31843_, new_n31842_, new_n8257_ );
or   ( new_n31844_, new_n8264_, new_n21685_ );
or   ( new_n31845_, new_n8266_, new_n21687_ );
and  ( new_n31846_, new_n31845_, new_n31844_ );
xor  ( new_n31847_, new_n31846_, new_n7725_ );
or   ( new_n31848_, new_n31847_, new_n31843_ );
and  ( new_n31849_, new_n31847_, new_n31843_ );
or   ( new_n31850_, new_n7732_, new_n21792_ );
or   ( new_n31851_, new_n7734_, new_n21751_ );
and  ( new_n31852_, new_n31851_, new_n31850_ );
xor  ( new_n31853_, new_n31852_, new_n7177_ );
or   ( new_n31854_, new_n31853_, new_n31849_ );
and  ( new_n31855_, new_n31854_, new_n31848_ );
or   ( new_n31856_, new_n7184_, new_n21840_ );
or   ( new_n31857_, new_n7186_, new_n21842_ );
and  ( new_n31858_, new_n31857_, new_n31856_ );
xor  ( new_n31859_, new_n31858_, new_n6638_ );
or   ( new_n31860_, new_n6645_, new_n22098_ );
or   ( new_n31861_, new_n6647_, new_n21847_ );
and  ( new_n31862_, new_n31861_, new_n31860_ );
xor  ( new_n31863_, new_n31862_, new_n6166_ );
or   ( new_n31864_, new_n31863_, new_n31859_ );
and  ( new_n31865_, new_n31863_, new_n31859_ );
or   ( new_n31866_, new_n6173_, new_n22207_ );
or   ( new_n31867_, new_n6175_, new_n22129_ );
and  ( new_n31868_, new_n31867_, new_n31866_ );
xor  ( new_n31869_, new_n31868_, new_n5597_ );
or   ( new_n31870_, new_n31869_, new_n31865_ );
and  ( new_n31871_, new_n31870_, new_n31864_ );
or   ( new_n31872_, new_n31871_, new_n31855_ );
and  ( new_n31873_, new_n31871_, new_n31855_ );
or   ( new_n31874_, new_n10059_, new_n21701_ );
or   ( new_n31875_, new_n10061_, new_n21703_ );
and  ( new_n31876_, new_n31875_, new_n31874_ );
xor  ( new_n31877_, new_n31876_, new_n9421_ );
and  ( new_n31878_, RIbb315f0_129, RIbb2d888_64 );
or   ( new_n31879_, new_n21694_, RIbb2d888_64 );
and  ( new_n31880_, new_n31879_, RIbb2d900_63 );
or   ( new_n31881_, new_n31880_, new_n31878_ );
or   ( new_n31882_, new_n10770_, new_n21696_ );
and  ( new_n31883_, new_n31882_, new_n31881_ );
nor  ( new_n31884_, new_n31883_, new_n31877_ );
and  ( new_n31885_, new_n31883_, new_n31877_ );
or   ( new_n31886_, new_n9422_, new_n21672_ );
or   ( new_n31887_, new_n9424_, new_n21674_ );
and  ( new_n31888_, new_n31887_, new_n31886_ );
xor  ( new_n31889_, new_n31888_, new_n8873_ );
nor  ( new_n31890_, new_n31889_, new_n31885_ );
nor  ( new_n31891_, new_n31890_, new_n31884_ );
or   ( new_n31892_, new_n31891_, new_n31873_ );
and  ( new_n31893_, new_n31892_, new_n31872_ );
or   ( new_n31894_, new_n31893_, new_n31839_ );
or   ( new_n31895_, new_n2122_, new_n25048_ );
or   ( new_n31896_, new_n2124_, new_n24925_ );
and  ( new_n31897_, new_n31896_, new_n31895_ );
xor  ( new_n31898_, new_n31897_, new_n1843_ );
or   ( new_n31899_, new_n1844_, new_n25486_ );
or   ( new_n31900_, new_n1846_, new_n25288_ );
and  ( new_n31901_, new_n31900_, new_n31899_ );
xor  ( new_n31902_, new_n31901_, new_n1586_ );
or   ( new_n31903_, new_n31902_, new_n31898_ );
and  ( new_n31904_, new_n31902_, new_n31898_ );
or   ( new_n31905_, new_n1593_, new_n26196_ );
or   ( new_n31906_, new_n1595_, new_n25813_ );
and  ( new_n31907_, new_n31906_, new_n31905_ );
xor  ( new_n31908_, new_n31907_, new_n1358_ );
or   ( new_n31909_, new_n31908_, new_n31904_ );
and  ( new_n31910_, new_n31909_, new_n31903_ );
or   ( new_n31911_, new_n1364_, new_n26372_ );
or   ( new_n31912_, new_n1366_, new_n26063_ );
and  ( new_n31913_, new_n31912_, new_n31911_ );
xor  ( new_n31914_, new_n31913_, new_n1129_ );
or   ( new_n31915_, new_n1135_, new_n26762_ );
or   ( new_n31916_, new_n1137_, new_n26620_ );
and  ( new_n31917_, new_n31916_, new_n31915_ );
xor  ( new_n31918_, new_n31917_, new_n896_ );
or   ( new_n31919_, new_n31918_, new_n31914_ );
and  ( new_n31920_, new_n31918_, new_n31914_ );
or   ( new_n31921_, new_n897_, new_n27396_ );
or   ( new_n31922_, new_n899_, new_n27085_ );
and  ( new_n31923_, new_n31922_, new_n31921_ );
xor  ( new_n31924_, new_n31923_, new_n748_ );
or   ( new_n31925_, new_n31924_, new_n31920_ );
and  ( new_n31926_, new_n31925_, new_n31919_ );
or   ( new_n31927_, new_n31926_, new_n31910_ );
and  ( new_n31928_, new_n31926_, new_n31910_ );
or   ( new_n31929_, new_n755_, new_n27763_ );
or   ( new_n31930_, new_n757_, new_n27602_ );
and  ( new_n31931_, new_n31930_, new_n31929_ );
xor  ( new_n31932_, new_n31931_, new_n523_ );
or   ( new_n31933_, new_n524_, new_n28314_ );
or   ( new_n31934_, new_n526_, new_n28108_ );
and  ( new_n31935_, new_n31934_, new_n31933_ );
xor  ( new_n31936_, new_n31935_, new_n403_ );
nor  ( new_n31937_, new_n31936_, new_n31932_ );
and  ( new_n31938_, new_n31936_, new_n31932_ );
or   ( new_n31939_, new_n409_, new_n29263_ );
or   ( new_n31940_, new_n411_, new_n28531_ );
and  ( new_n31941_, new_n31940_, new_n31939_ );
xor  ( new_n31942_, new_n31941_, new_n328_ );
nor  ( new_n31943_, new_n31942_, new_n31938_ );
nor  ( new_n31944_, new_n31943_, new_n31937_ );
or   ( new_n31945_, new_n31944_, new_n31928_ );
and  ( new_n31946_, new_n31945_, new_n31927_ );
and  ( new_n31947_, new_n31893_, new_n31839_ );
or   ( new_n31948_, new_n31947_, new_n31946_ );
and  ( new_n31949_, new_n31948_, new_n31894_ );
and  ( new_n31950_, new_n31949_, new_n31787_ );
nor  ( new_n31951_, new_n31949_, new_n31787_ );
not  ( new_n31952_, RIbb33378_192 );
or   ( new_n31953_, new_n31952_, new_n260_ );
xnor ( new_n31954_, new_n31651_, new_n31647_ );
xor  ( new_n31955_, new_n31954_, new_n31658_ );
or   ( new_n31956_, new_n31955_, new_n31953_ );
and  ( new_n31957_, new_n31955_, new_n31953_ );
or   ( new_n31958_, new_n337_, new_n29474_ );
or   ( new_n31959_, new_n340_, new_n29261_ );
and  ( new_n31960_, new_n31959_, new_n31958_ );
xor  ( new_n31961_, new_n31960_, new_n332_ );
or   ( new_n31962_, new_n317_, new_n30120_ );
or   ( new_n31963_, new_n320_, new_n29619_ );
and  ( new_n31964_, new_n31963_, new_n31962_ );
xor  ( new_n31965_, new_n31964_, new_n312_ );
nor  ( new_n31966_, new_n31965_, new_n31961_ );
and  ( new_n31967_, new_n31965_, new_n31961_ );
or   ( new_n31968_, new_n283_, new_n30800_ );
or   ( new_n31969_, new_n286_, new_n30227_ );
and  ( new_n31970_, new_n31969_, new_n31968_ );
xor  ( new_n31971_, new_n31970_, new_n278_ );
nor  ( new_n31972_, new_n31971_, new_n31967_ );
nor  ( new_n31973_, new_n31972_, new_n31966_ );
not  ( new_n31974_, new_n31973_ );
or   ( new_n31975_, new_n31974_, new_n31957_ );
and  ( new_n31976_, new_n31975_, new_n31956_ );
xnor ( new_n31977_, new_n31550_, new_n31546_ );
xor  ( new_n31978_, new_n31977_, new_n31556_ );
xnor ( new_n31979_, new_n31534_, new_n31530_ );
xor  ( new_n31980_, new_n31979_, new_n31540_ );
or   ( new_n31981_, new_n31980_, new_n31978_ );
and  ( new_n31982_, new_n31980_, new_n31978_ );
xnor ( new_n31983_, new_n31516_, new_n31512_ );
xor  ( new_n31984_, new_n31983_, new_n31522_ );
or   ( new_n31985_, new_n31984_, new_n31982_ );
and  ( new_n31986_, new_n31985_, new_n31981_ );
nor  ( new_n31987_, new_n31986_, new_n31976_ );
and  ( new_n31988_, new_n31986_, new_n31976_ );
xnor ( new_n31989_, new_n31498_, new_n31494_ );
xor  ( new_n31990_, new_n31989_, new_n31504_ );
xnor ( new_n31991_, new_n31635_, new_n31631_ );
xor  ( new_n31992_, new_n31991_, new_n31641_ );
nor  ( new_n31993_, new_n31992_, new_n31990_ );
and  ( new_n31994_, new_n31992_, new_n31990_ );
xor  ( new_n31995_, new_n31482_, new_n31478_ );
xnor ( new_n31996_, new_n31995_, new_n31488_ );
nor  ( new_n31997_, new_n31996_, new_n31994_ );
nor  ( new_n31998_, new_n31997_, new_n31993_ );
nor  ( new_n31999_, new_n31998_, new_n31988_ );
nor  ( new_n32000_, new_n31999_, new_n31987_ );
nor  ( new_n32001_, new_n32000_, new_n31951_ );
nor  ( new_n32002_, new_n32001_, new_n31950_ );
nor  ( new_n32003_, new_n32002_, new_n31770_ );
nor  ( new_n32004_, new_n32003_, new_n31769_ );
nand ( new_n32005_, new_n32004_, new_n31732_ );
and  ( new_n32006_, new_n32005_, new_n31731_ );
nand ( new_n32007_, new_n32006_, new_n31718_ );
nor  ( new_n32008_, new_n32006_, new_n31718_ );
xor  ( new_n32009_, new_n31086_, new_n31084_ );
xor  ( new_n32010_, new_n32009_, new_n31091_ );
or   ( new_n32011_, new_n32010_, new_n32008_ );
and  ( new_n32012_, new_n32011_, new_n32007_ );
or   ( new_n32013_, new_n32012_, new_n31713_ );
nand ( new_n32014_, new_n32012_, new_n31713_ );
xor  ( new_n32015_, new_n31693_, new_n31691_ );
xnor ( new_n32016_, new_n32015_, new_n31697_ );
nand ( new_n32017_, new_n32016_, new_n32014_ );
and  ( new_n32018_, new_n32017_, new_n32013_ );
nor  ( new_n32019_, new_n32018_, new_n31708_ );
xor  ( new_n32020_, new_n32012_, new_n31713_ );
xor  ( new_n32021_, new_n32020_, new_n32016_ );
xnor ( new_n32022_, new_n31776_, new_n31774_ );
xor  ( new_n32023_, new_n32022_, new_n31780_ );
xnor ( new_n32024_, new_n31992_, new_n31990_ );
xor  ( new_n32025_, new_n32024_, new_n31996_ );
nor  ( new_n32026_, new_n32025_, new_n32023_ );
nand ( new_n32027_, new_n32025_, new_n32023_ );
xor  ( new_n32028_, new_n31980_, new_n31978_ );
xor  ( new_n32029_, new_n32028_, new_n31984_ );
and  ( new_n32030_, new_n32029_, new_n32027_ );
or   ( new_n32031_, new_n32030_, new_n32026_ );
xor  ( new_n32032_, new_n31749_, new_n31747_ );
xor  ( new_n32033_, new_n32032_, new_n31754_ );
nor  ( new_n32034_, new_n32033_, new_n32031_ );
nand ( new_n32035_, new_n32033_, new_n32031_ );
xnor ( new_n32036_, new_n31819_, new_n31803_ );
xor  ( new_n32037_, new_n32036_, new_n31837_ );
xnor ( new_n32038_, new_n31926_, new_n31910_ );
xor  ( new_n32039_, new_n32038_, new_n31944_ );
nor  ( new_n32040_, new_n32039_, new_n32037_ );
and  ( new_n32041_, new_n32039_, new_n32037_ );
xor  ( new_n32042_, new_n31955_, new_n31953_ );
xor  ( new_n32043_, new_n32042_, new_n31974_ );
nor  ( new_n32044_, new_n32043_, new_n32041_ );
or   ( new_n32045_, new_n32044_, new_n32040_ );
and  ( new_n32046_, new_n32045_, new_n32035_ );
or   ( new_n32047_, new_n32046_, new_n32034_ );
xor  ( new_n32048_, new_n31847_, new_n31843_ );
xnor ( new_n32049_, new_n32048_, new_n31853_ );
xnor ( new_n32050_, new_n31883_, new_n31877_ );
xor  ( new_n32051_, new_n32050_, new_n31889_ );
or   ( new_n32052_, new_n32051_, new_n32049_ );
xnor ( new_n32053_, new_n31811_, new_n31807_ );
xor  ( new_n32054_, new_n32053_, new_n31817_ );
xnor ( new_n32055_, new_n31795_, new_n31791_ );
xor  ( new_n32056_, new_n32055_, new_n31801_ );
or   ( new_n32057_, new_n32056_, new_n32054_ );
and  ( new_n32058_, new_n32056_, new_n32054_ );
xnor ( new_n32059_, new_n31863_, new_n31859_ );
xor  ( new_n32060_, new_n32059_, new_n31869_ );
or   ( new_n32061_, new_n32060_, new_n32058_ );
and  ( new_n32062_, new_n32061_, new_n32057_ );
nor  ( new_n32063_, new_n32062_, new_n32052_ );
nand ( new_n32064_, new_n32062_, new_n32052_ );
xor  ( new_n32065_, new_n31602_, new_n31600_ );
and  ( new_n32066_, new_n32065_, new_n32064_ );
or   ( new_n32067_, new_n32066_, new_n32063_ );
xnor ( new_n32068_, new_n31918_, new_n31914_ );
xor  ( new_n32069_, new_n32068_, new_n31924_ );
xnor ( new_n32070_, new_n31902_, new_n31898_ );
xor  ( new_n32071_, new_n32070_, new_n31908_ );
nor  ( new_n32072_, new_n32071_, new_n32069_ );
and  ( new_n32073_, new_n32071_, new_n32069_ );
xor  ( new_n32074_, new_n31829_, new_n31825_ );
xnor ( new_n32075_, new_n32074_, new_n31835_ );
nor  ( new_n32076_, new_n32075_, new_n32073_ );
or   ( new_n32077_, new_n32076_, new_n32072_ );
or   ( new_n32078_, new_n299_, new_n31333_ );
or   ( new_n32079_, new_n302_, new_n30798_ );
and  ( new_n32080_, new_n32079_, new_n32078_ );
xor  ( new_n32081_, new_n32080_, new_n293_ );
or   ( new_n32082_, new_n283_, new_n30798_ );
or   ( new_n32083_, new_n286_, new_n30800_ );
and  ( new_n32084_, new_n32083_, new_n32082_ );
xor  ( new_n32085_, new_n32084_, new_n278_ );
or   ( new_n32086_, new_n299_, new_n31654_ );
or   ( new_n32087_, new_n302_, new_n31333_ );
and  ( new_n32088_, new_n32087_, new_n32086_ );
xor  ( new_n32089_, new_n32088_, new_n293_ );
or   ( new_n32090_, new_n32089_, new_n32085_ );
and  ( new_n32091_, new_n32089_, new_n32085_ );
and  ( new_n32092_, new_n265_, RIbb33378_192 );
nor  ( new_n32093_, new_n32092_, new_n262_ );
and  ( new_n32094_, new_n32092_, RIbb2f610_1 );
nor  ( new_n32095_, new_n32094_, new_n32093_ );
or   ( new_n32096_, new_n32095_, new_n32091_ );
and  ( new_n32097_, new_n32096_, new_n32090_ );
or   ( new_n32098_, new_n32097_, new_n32081_ );
and  ( new_n32099_, new_n32097_, new_n32081_ );
or   ( new_n32100_, new_n409_, new_n29261_ );
or   ( new_n32101_, new_n411_, new_n29263_ );
and  ( new_n32102_, new_n32101_, new_n32100_ );
xor  ( new_n32103_, new_n32102_, new_n328_ );
or   ( new_n32104_, new_n337_, new_n29619_ );
or   ( new_n32105_, new_n340_, new_n29474_ );
and  ( new_n32106_, new_n32105_, new_n32104_ );
xor  ( new_n32107_, new_n32106_, new_n332_ );
nor  ( new_n32108_, new_n32107_, new_n32103_ );
and  ( new_n32109_, new_n32107_, new_n32103_ );
or   ( new_n32110_, new_n317_, new_n30227_ );
or   ( new_n32111_, new_n320_, new_n30120_ );
and  ( new_n32112_, new_n32111_, new_n32110_ );
xor  ( new_n32113_, new_n32112_, new_n312_ );
nor  ( new_n32114_, new_n32113_, new_n32109_ );
nor  ( new_n32115_, new_n32114_, new_n32108_ );
or   ( new_n32116_, new_n32115_, new_n32099_ );
and  ( new_n32117_, new_n32116_, new_n32098_ );
or   ( new_n32118_, new_n32117_, new_n32077_ );
and  ( new_n32119_, new_n32117_, new_n32077_ );
or   ( new_n32120_, new_n268_, new_n31952_ );
or   ( new_n32121_, new_n271_, new_n31654_ );
and  ( new_n32122_, new_n32121_, new_n32120_ );
xor  ( new_n32123_, new_n32122_, new_n262_ );
xnor ( new_n32124_, new_n31936_, new_n31932_ );
xor  ( new_n32125_, new_n32124_, new_n31942_ );
and  ( new_n32126_, new_n32125_, new_n32123_ );
nor  ( new_n32127_, new_n32125_, new_n32123_ );
xor  ( new_n32128_, new_n31965_, new_n31961_ );
xnor ( new_n32129_, new_n32128_, new_n31971_ );
not  ( new_n32130_, new_n32129_ );
nor  ( new_n32131_, new_n32130_, new_n32127_ );
nor  ( new_n32132_, new_n32131_, new_n32126_ );
or   ( new_n32133_, new_n32132_, new_n32119_ );
and  ( new_n32134_, new_n32133_, new_n32118_ );
or   ( new_n32135_, new_n32134_, new_n32067_ );
and  ( new_n32136_, new_n32134_, new_n32067_ );
or   ( new_n32137_, new_n2425_, new_n24925_ );
or   ( new_n32138_, new_n2427_, new_n24927_ );
and  ( new_n32139_, new_n32138_, new_n32137_ );
xor  ( new_n32140_, new_n32139_, new_n2121_ );
or   ( new_n32141_, new_n2122_, new_n25288_ );
or   ( new_n32142_, new_n2124_, new_n25048_ );
and  ( new_n32143_, new_n32142_, new_n32141_ );
xor  ( new_n32144_, new_n32143_, new_n1843_ );
or   ( new_n32145_, new_n32144_, new_n32140_ );
and  ( new_n32146_, new_n32144_, new_n32140_ );
or   ( new_n32147_, new_n1844_, new_n25813_ );
or   ( new_n32148_, new_n1846_, new_n25486_ );
and  ( new_n32149_, new_n32148_, new_n32147_ );
xor  ( new_n32150_, new_n32149_, new_n1586_ );
or   ( new_n32151_, new_n32150_, new_n32146_ );
and  ( new_n32152_, new_n32151_, new_n32145_ );
or   ( new_n32153_, new_n1593_, new_n26063_ );
or   ( new_n32154_, new_n1595_, new_n26196_ );
and  ( new_n32155_, new_n32154_, new_n32153_ );
xor  ( new_n32156_, new_n32155_, new_n1358_ );
or   ( new_n32157_, new_n1364_, new_n26620_ );
or   ( new_n32158_, new_n1366_, new_n26372_ );
and  ( new_n32159_, new_n32158_, new_n32157_ );
xor  ( new_n32160_, new_n32159_, new_n1129_ );
or   ( new_n32161_, new_n32160_, new_n32156_ );
and  ( new_n32162_, new_n32160_, new_n32156_ );
or   ( new_n32163_, new_n1135_, new_n27085_ );
or   ( new_n32164_, new_n1137_, new_n26762_ );
and  ( new_n32165_, new_n32164_, new_n32163_ );
xor  ( new_n32166_, new_n32165_, new_n896_ );
or   ( new_n32167_, new_n32166_, new_n32162_ );
and  ( new_n32168_, new_n32167_, new_n32161_ );
or   ( new_n32169_, new_n32168_, new_n32152_ );
and  ( new_n32170_, new_n32168_, new_n32152_ );
or   ( new_n32171_, new_n897_, new_n27602_ );
or   ( new_n32172_, new_n899_, new_n27396_ );
and  ( new_n32173_, new_n32172_, new_n32171_ );
xor  ( new_n32174_, new_n32173_, new_n748_ );
or   ( new_n32175_, new_n755_, new_n28108_ );
or   ( new_n32176_, new_n757_, new_n27763_ );
and  ( new_n32177_, new_n32176_, new_n32175_ );
xor  ( new_n32178_, new_n32177_, new_n523_ );
or   ( new_n32179_, new_n32178_, new_n32174_ );
and  ( new_n32180_, new_n32178_, new_n32174_ );
or   ( new_n32181_, new_n524_, new_n28531_ );
or   ( new_n32182_, new_n526_, new_n28314_ );
and  ( new_n32183_, new_n32182_, new_n32181_ );
xor  ( new_n32184_, new_n32183_, new_n403_ );
or   ( new_n32185_, new_n32184_, new_n32180_ );
and  ( new_n32186_, new_n32185_, new_n32179_ );
or   ( new_n32187_, new_n32186_, new_n32170_ );
and  ( new_n32188_, new_n32187_, new_n32169_ );
or   ( new_n32189_, new_n7732_, new_n21842_ );
or   ( new_n32190_, new_n7734_, new_n21792_ );
and  ( new_n32191_, new_n32190_, new_n32189_ );
xor  ( new_n32192_, new_n32191_, new_n7177_ );
or   ( new_n32193_, new_n7184_, new_n21847_ );
or   ( new_n32194_, new_n7186_, new_n21840_ );
and  ( new_n32195_, new_n32194_, new_n32193_ );
xor  ( new_n32196_, new_n32195_, new_n6638_ );
nor  ( new_n32197_, new_n32196_, new_n32192_ );
and  ( new_n32198_, new_n32196_, new_n32192_ );
or   ( new_n32199_, new_n6645_, new_n22129_ );
or   ( new_n32200_, new_n6647_, new_n22098_ );
and  ( new_n32201_, new_n32200_, new_n32199_ );
xor  ( new_n32202_, new_n32201_, new_n6166_ );
nor  ( new_n32203_, new_n32202_, new_n32198_ );
nor  ( new_n32204_, new_n32203_, new_n32197_ );
or   ( new_n32205_, new_n10059_, new_n21674_ );
or   ( new_n32206_, new_n10061_, new_n21701_ );
and  ( new_n32207_, new_n32206_, new_n32205_ );
xor  ( new_n32208_, new_n32207_, new_n9421_ );
and  ( new_n32209_, RIbb31668_130, RIbb2d888_64 );
or   ( new_n32210_, new_n21703_, RIbb2d888_64 );
and  ( new_n32211_, new_n32210_, RIbb2d900_63 );
or   ( new_n32212_, new_n32211_, new_n32209_ );
or   ( new_n32213_, new_n10770_, new_n21694_ );
and  ( new_n32214_, new_n32213_, new_n32212_ );
nor  ( new_n32215_, new_n32214_, new_n32208_ );
and  ( new_n32216_, new_n32214_, new_n32208_ );
nor  ( new_n32217_, new_n32216_, new_n262_ );
nor  ( new_n32218_, new_n32217_, new_n32215_ );
or   ( new_n32219_, new_n9422_, new_n21680_ );
or   ( new_n32220_, new_n9424_, new_n21672_ );
and  ( new_n32221_, new_n32220_, new_n32219_ );
xor  ( new_n32222_, new_n32221_, new_n8873_ );
or   ( new_n32223_, new_n8874_, new_n21687_ );
or   ( new_n32224_, new_n8876_, new_n21678_ );
and  ( new_n32225_, new_n32224_, new_n32223_ );
xor  ( new_n32226_, new_n32225_, new_n8257_ );
or   ( new_n32227_, new_n32226_, new_n32222_ );
and  ( new_n32228_, new_n32226_, new_n32222_ );
or   ( new_n32229_, new_n8264_, new_n21751_ );
or   ( new_n32230_, new_n8266_, new_n21685_ );
and  ( new_n32231_, new_n32230_, new_n32229_ );
xor  ( new_n32232_, new_n32231_, new_n7725_ );
or   ( new_n32233_, new_n32232_, new_n32228_ );
and  ( new_n32234_, new_n32233_, new_n32227_ );
and  ( new_n32235_, new_n32234_, new_n32218_ );
or   ( new_n32236_, new_n32235_, new_n32204_ );
or   ( new_n32237_, new_n32234_, new_n32218_ );
and  ( new_n32238_, new_n32237_, new_n32236_ );
nor  ( new_n32239_, new_n32238_, new_n32188_ );
or   ( new_n32240_, new_n6173_, new_n22304_ );
or   ( new_n32241_, new_n6175_, new_n22207_ );
and  ( new_n32242_, new_n32241_, new_n32240_ );
xor  ( new_n32243_, new_n32242_, new_n5597_ );
or   ( new_n32244_, new_n5604_, new_n22590_ );
or   ( new_n32245_, new_n5606_, new_n22423_ );
and  ( new_n32246_, new_n32245_, new_n32244_ );
xor  ( new_n32247_, new_n32246_, new_n5206_ );
or   ( new_n32248_, new_n32247_, new_n32243_ );
and  ( new_n32249_, new_n32247_, new_n32243_ );
or   ( new_n32250_, new_n5207_, new_n22829_ );
or   ( new_n32251_, new_n5209_, new_n22641_ );
and  ( new_n32252_, new_n32251_, new_n32250_ );
xor  ( new_n32253_, new_n32252_, new_n4708_ );
or   ( new_n32254_, new_n32253_, new_n32249_ );
and  ( new_n32255_, new_n32254_, new_n32248_ );
or   ( new_n32256_, new_n4709_, new_n22973_ );
or   ( new_n32257_, new_n4711_, new_n22975_ );
and  ( new_n32258_, new_n32257_, new_n32256_ );
xor  ( new_n32259_, new_n32258_, new_n4295_ );
or   ( new_n32260_, new_n4302_, new_n23252_ );
or   ( new_n32261_, new_n4304_, new_n23166_ );
and  ( new_n32262_, new_n32261_, new_n32260_ );
xor  ( new_n32263_, new_n32262_, new_n3895_ );
or   ( new_n32264_, new_n32263_, new_n32259_ );
and  ( new_n32265_, new_n32263_, new_n32259_ );
or   ( new_n32266_, new_n3896_, new_n23554_ );
or   ( new_n32267_, new_n3898_, new_n23370_ );
and  ( new_n32268_, new_n32267_, new_n32266_ );
xor  ( new_n32269_, new_n32268_, new_n3460_ );
or   ( new_n32270_, new_n32269_, new_n32265_ );
and  ( new_n32271_, new_n32270_, new_n32264_ );
nor  ( new_n32272_, new_n32271_, new_n32255_ );
and  ( new_n32273_, new_n32271_, new_n32255_ );
or   ( new_n32274_, new_n3461_, new_n23895_ );
or   ( new_n32275_, new_n3463_, new_n23733_ );
and  ( new_n32276_, new_n32275_, new_n32274_ );
xor  ( new_n32277_, new_n32276_, new_n3116_ );
or   ( new_n32278_, new_n3117_, new_n24227_ );
or   ( new_n32279_, new_n3119_, new_n24006_ );
and  ( new_n32280_, new_n32279_, new_n32278_ );
xor  ( new_n32281_, new_n32280_, new_n2800_ );
nor  ( new_n32282_, new_n32281_, new_n32277_ );
and  ( new_n32283_, new_n32281_, new_n32277_ );
or   ( new_n32284_, new_n2807_, new_n24543_ );
or   ( new_n32285_, new_n2809_, new_n24418_ );
and  ( new_n32286_, new_n32285_, new_n32284_ );
xor  ( new_n32287_, new_n32286_, new_n2424_ );
nor  ( new_n32288_, new_n32287_, new_n32283_ );
nor  ( new_n32289_, new_n32288_, new_n32282_ );
nor  ( new_n32290_, new_n32289_, new_n32273_ );
nor  ( new_n32291_, new_n32290_, new_n32272_ );
and  ( new_n32292_, new_n32238_, new_n32188_ );
nor  ( new_n32293_, new_n32292_, new_n32291_ );
nor  ( new_n32294_, new_n32293_, new_n32239_ );
or   ( new_n32295_, new_n32294_, new_n32136_ );
and  ( new_n32296_, new_n32295_, new_n32135_ );
nor  ( new_n32297_, new_n32296_, new_n32047_ );
nand ( new_n32298_, new_n32296_, new_n32047_ );
xor  ( new_n32299_, new_n31986_, new_n31976_ );
xor  ( new_n32300_, new_n32299_, new_n31998_ );
xor  ( new_n32301_, new_n31736_, new_n31734_ );
xor  ( new_n32302_, new_n32301_, new_n31739_ );
or   ( new_n32303_, new_n32302_, new_n32300_ );
nand ( new_n32304_, new_n32302_, new_n32300_ );
xor  ( new_n32305_, new_n31782_, new_n31772_ );
xor  ( new_n32306_, new_n32305_, new_n31785_ );
nand ( new_n32307_, new_n32306_, new_n32304_ );
and  ( new_n32308_, new_n32307_, new_n32303_ );
and  ( new_n32309_, new_n32308_, new_n32298_ );
or   ( new_n32310_, new_n32309_, new_n32297_ );
xor  ( new_n32311_, new_n31671_, new_n31661_ );
xor  ( new_n32312_, new_n32311_, new_n31683_ );
xnor ( new_n32313_, new_n31578_, new_n31526_ );
xor  ( new_n32314_, new_n32313_, new_n31623_ );
or   ( new_n32315_, new_n32314_, new_n32312_ );
and  ( new_n32316_, new_n32314_, new_n32312_ );
xor  ( new_n32317_, new_n31762_, new_n31760_ );
xnor ( new_n32318_, new_n32317_, new_n31766_ );
not  ( new_n32319_, new_n32318_ );
or   ( new_n32320_, new_n32319_, new_n32316_ );
and  ( new_n32321_, new_n32320_, new_n32315_ );
or   ( new_n32322_, new_n32321_, new_n32310_ );
nand ( new_n32323_, new_n32321_, new_n32310_ );
xor  ( new_n32324_, new_n31625_, new_n31474_ );
xnor ( new_n32325_, new_n32324_, new_n31685_ );
nand ( new_n32326_, new_n32325_, new_n32323_ );
and  ( new_n32327_, new_n32326_, new_n32322_ );
xor  ( new_n32328_, new_n31730_, new_n31720_ );
xor  ( new_n32329_, new_n32328_, new_n32004_ );
nor  ( new_n32330_, new_n32329_, new_n32327_ );
nand ( new_n32331_, new_n32329_, new_n32327_ );
xor  ( new_n32332_, new_n31717_, new_n31715_ );
and  ( new_n32333_, new_n32332_, new_n32331_ );
or   ( new_n32334_, new_n32333_, new_n32330_ );
xnor ( new_n32335_, new_n32006_, new_n31718_ );
xor  ( new_n32336_, new_n32335_, new_n32010_ );
or   ( new_n32337_, new_n32336_, new_n32334_ );
and  ( new_n32338_, new_n32336_, new_n32334_ );
xor  ( new_n32339_, new_n31712_, new_n31710_ );
or   ( new_n32340_, new_n32339_, new_n32338_ );
and  ( new_n32341_, new_n32340_, new_n32337_ );
and  ( new_n32342_, new_n32341_, new_n32021_ );
xnor ( new_n32343_, new_n32336_, new_n32334_ );
xor  ( new_n32344_, new_n32343_, new_n32339_ );
xor  ( new_n32345_, new_n31768_, new_n31758_ );
xnor ( new_n32346_, new_n32345_, new_n32002_ );
xor  ( new_n32347_, new_n32321_, new_n32310_ );
xor  ( new_n32348_, new_n32347_, new_n32325_ );
nand ( new_n32349_, new_n32348_, new_n32346_ );
xor  ( new_n32350_, new_n31949_, new_n31787_ );
xor  ( new_n32351_, new_n32350_, new_n32000_ );
xor  ( new_n32352_, new_n32296_, new_n32047_ );
xor  ( new_n32353_, new_n32352_, new_n32308_ );
nor  ( new_n32354_, new_n32353_, new_n32351_ );
and  ( new_n32355_, new_n32353_, new_n32351_ );
xor  ( new_n32356_, new_n32314_, new_n32312_ );
xor  ( new_n32357_, new_n32356_, new_n32319_ );
nor  ( new_n32358_, new_n32357_, new_n32355_ );
or   ( new_n32359_, new_n32358_, new_n32354_ );
xor  ( new_n32360_, new_n31893_, new_n31839_ );
xor  ( new_n32361_, new_n32360_, new_n31946_ );
xor  ( new_n32362_, new_n32033_, new_n32031_ );
xor  ( new_n32363_, new_n32362_, new_n32045_ );
or   ( new_n32364_, new_n32363_, new_n32361_ );
and  ( new_n32365_, new_n32363_, new_n32361_ );
xor  ( new_n32366_, new_n32302_, new_n32300_ );
xor  ( new_n32367_, new_n32366_, new_n32306_ );
or   ( new_n32368_, new_n32367_, new_n32365_ );
and  ( new_n32369_, new_n32368_, new_n32364_ );
xor  ( new_n32370_, new_n32071_, new_n32069_ );
xor  ( new_n32371_, new_n32370_, new_n32075_ );
xnor ( new_n32372_, new_n32097_, new_n32081_ );
xor  ( new_n32373_, new_n32372_, new_n32115_ );
or   ( new_n32374_, new_n32373_, new_n32371_ );
and  ( new_n32375_, new_n32373_, new_n32371_ );
xor  ( new_n32376_, new_n32125_, new_n32123_ );
xor  ( new_n32377_, new_n32376_, new_n32129_ );
or   ( new_n32378_, new_n32377_, new_n32375_ );
and  ( new_n32379_, new_n32378_, new_n32374_ );
xor  ( new_n32380_, new_n32168_, new_n32152_ );
xor  ( new_n32381_, new_n32380_, new_n32186_ );
xor  ( new_n32382_, new_n32234_, new_n32218_ );
xor  ( new_n32383_, new_n32382_, new_n32204_ );
nand ( new_n32384_, new_n32383_, new_n32381_ );
nor  ( new_n32385_, new_n32383_, new_n32381_ );
xor  ( new_n32386_, new_n32271_, new_n32255_ );
xnor ( new_n32387_, new_n32386_, new_n32289_ );
or   ( new_n32388_, new_n32387_, new_n32385_ );
and  ( new_n32389_, new_n32388_, new_n32384_ );
nor  ( new_n32390_, new_n32389_, new_n32379_ );
and  ( new_n32391_, new_n32389_, new_n32379_ );
xor  ( new_n32392_, new_n31871_, new_n31855_ );
xnor ( new_n32393_, new_n32392_, new_n31891_ );
nor  ( new_n32394_, new_n32393_, new_n32391_ );
or   ( new_n32395_, new_n32394_, new_n32390_ );
xnor ( new_n32396_, new_n32263_, new_n32259_ );
xor  ( new_n32397_, new_n32396_, new_n32269_ );
xnor ( new_n32398_, new_n32247_, new_n32243_ );
xor  ( new_n32399_, new_n32398_, new_n32253_ );
nor  ( new_n32400_, new_n32399_, new_n32397_ );
nand ( new_n32401_, new_n32399_, new_n32397_ );
xor  ( new_n32402_, new_n32281_, new_n32277_ );
xnor ( new_n32403_, new_n32402_, new_n32287_ );
not  ( new_n32404_, new_n32403_ );
and  ( new_n32405_, new_n32404_, new_n32401_ );
or   ( new_n32406_, new_n32405_, new_n32400_ );
xor  ( new_n32407_, new_n32107_, new_n32103_ );
xor  ( new_n32408_, new_n32407_, new_n32113_ );
or   ( new_n32409_, new_n337_, new_n30120_ );
or   ( new_n32410_, new_n340_, new_n29619_ );
and  ( new_n32411_, new_n32410_, new_n32409_ );
xor  ( new_n32412_, new_n32411_, new_n332_ );
or   ( new_n32413_, new_n317_, new_n30800_ );
or   ( new_n32414_, new_n320_, new_n30227_ );
and  ( new_n32415_, new_n32414_, new_n32413_ );
xor  ( new_n32416_, new_n32415_, new_n312_ );
or   ( new_n32417_, new_n32416_, new_n32412_ );
and  ( new_n32418_, new_n32416_, new_n32412_ );
or   ( new_n32419_, new_n283_, new_n31333_ );
or   ( new_n32420_, new_n286_, new_n30798_ );
and  ( new_n32421_, new_n32420_, new_n32419_ );
xor  ( new_n32422_, new_n32421_, new_n278_ );
or   ( new_n32423_, new_n32422_, new_n32418_ );
and  ( new_n32424_, new_n32423_, new_n32417_ );
or   ( new_n32425_, new_n32424_, new_n32408_ );
nand ( new_n32426_, new_n32424_, new_n32408_ );
xor  ( new_n32427_, new_n32089_, new_n32085_ );
xnor ( new_n32428_, new_n32427_, new_n32095_ );
nand ( new_n32429_, new_n32428_, new_n32426_ );
and  ( new_n32430_, new_n32429_, new_n32425_ );
and  ( new_n32431_, new_n32430_, new_n32406_ );
or   ( new_n32432_, new_n32430_, new_n32406_ );
xnor ( new_n32433_, new_n32160_, new_n32156_ );
xor  ( new_n32434_, new_n32433_, new_n32166_ );
xnor ( new_n32435_, new_n32144_, new_n32140_ );
xor  ( new_n32436_, new_n32435_, new_n32150_ );
nor  ( new_n32437_, new_n32436_, new_n32434_ );
nand ( new_n32438_, new_n32436_, new_n32434_ );
xor  ( new_n32439_, new_n32178_, new_n32174_ );
xnor ( new_n32440_, new_n32439_, new_n32184_ );
not  ( new_n32441_, new_n32440_ );
and  ( new_n32442_, new_n32441_, new_n32438_ );
or   ( new_n32443_, new_n32442_, new_n32437_ );
and  ( new_n32444_, new_n32443_, new_n32432_ );
or   ( new_n32445_, new_n32444_, new_n32431_ );
or   ( new_n32446_, new_n10059_, new_n21672_ );
or   ( new_n32447_, new_n10061_, new_n21674_ );
and  ( new_n32448_, new_n32447_, new_n32446_ );
xor  ( new_n32449_, new_n32448_, new_n9421_ );
and  ( new_n32450_, RIbb316e0_131, RIbb2d888_64 );
or   ( new_n32451_, new_n21701_, RIbb2d888_64 );
and  ( new_n32452_, new_n32451_, RIbb2d900_63 );
or   ( new_n32453_, new_n32452_, new_n32450_ );
or   ( new_n32454_, new_n10770_, new_n21703_ );
and  ( new_n32455_, new_n32454_, new_n32453_ );
or   ( new_n32456_, new_n32455_, new_n32449_ );
and  ( new_n32457_, new_n32455_, new_n32449_ );
or   ( new_n32458_, new_n9422_, new_n21678_ );
or   ( new_n32459_, new_n9424_, new_n21680_ );
and  ( new_n32460_, new_n32459_, new_n32458_ );
xor  ( new_n32461_, new_n32460_, new_n8873_ );
or   ( new_n32462_, new_n32461_, new_n32457_ );
and  ( new_n32463_, new_n32462_, new_n32456_ );
or   ( new_n32464_, new_n8874_, new_n21685_ );
or   ( new_n32465_, new_n8876_, new_n21687_ );
and  ( new_n32466_, new_n32465_, new_n32464_ );
xor  ( new_n32467_, new_n32466_, new_n8257_ );
or   ( new_n32468_, new_n8264_, new_n21792_ );
or   ( new_n32469_, new_n8266_, new_n21751_ );
and  ( new_n32470_, new_n32469_, new_n32468_ );
xor  ( new_n32471_, new_n32470_, new_n7725_ );
or   ( new_n32472_, new_n32471_, new_n32467_ );
and  ( new_n32473_, new_n32471_, new_n32467_ );
or   ( new_n32474_, new_n7732_, new_n21840_ );
or   ( new_n32475_, new_n7734_, new_n21842_ );
and  ( new_n32476_, new_n32475_, new_n32474_ );
xor  ( new_n32477_, new_n32476_, new_n7177_ );
or   ( new_n32478_, new_n32477_, new_n32473_ );
and  ( new_n32479_, new_n32478_, new_n32472_ );
or   ( new_n32480_, new_n32479_, new_n32463_ );
and  ( new_n32481_, new_n32479_, new_n32463_ );
or   ( new_n32482_, new_n7184_, new_n22098_ );
or   ( new_n32483_, new_n7186_, new_n21847_ );
and  ( new_n32484_, new_n32483_, new_n32482_ );
xor  ( new_n32485_, new_n32484_, new_n6638_ );
or   ( new_n32486_, new_n6645_, new_n22207_ );
or   ( new_n32487_, new_n6647_, new_n22129_ );
and  ( new_n32488_, new_n32487_, new_n32486_ );
xor  ( new_n32489_, new_n32488_, new_n6166_ );
nor  ( new_n32490_, new_n32489_, new_n32485_ );
and  ( new_n32491_, new_n32489_, new_n32485_ );
or   ( new_n32492_, new_n6173_, new_n22423_ );
or   ( new_n32493_, new_n6175_, new_n22304_ );
and  ( new_n32494_, new_n32493_, new_n32492_ );
xor  ( new_n32495_, new_n32494_, new_n5597_ );
nor  ( new_n32496_, new_n32495_, new_n32491_ );
nor  ( new_n32497_, new_n32496_, new_n32490_ );
or   ( new_n32498_, new_n32497_, new_n32481_ );
and  ( new_n32499_, new_n32498_, new_n32480_ );
or   ( new_n32500_, new_n755_, new_n28314_ );
or   ( new_n32501_, new_n757_, new_n28108_ );
and  ( new_n32502_, new_n32501_, new_n32500_ );
xor  ( new_n32503_, new_n32502_, new_n523_ );
or   ( new_n32504_, new_n524_, new_n29263_ );
or   ( new_n32505_, new_n526_, new_n28531_ );
and  ( new_n32506_, new_n32505_, new_n32504_ );
xor  ( new_n32507_, new_n32506_, new_n403_ );
or   ( new_n32508_, new_n32507_, new_n32503_ );
and  ( new_n32509_, new_n32507_, new_n32503_ );
or   ( new_n32510_, new_n409_, new_n29474_ );
or   ( new_n32511_, new_n411_, new_n29261_ );
and  ( new_n32512_, new_n32511_, new_n32510_ );
xor  ( new_n32513_, new_n32512_, new_n328_ );
or   ( new_n32514_, new_n32513_, new_n32509_ );
and  ( new_n32515_, new_n32514_, new_n32508_ );
or   ( new_n32516_, new_n1364_, new_n26762_ );
or   ( new_n32517_, new_n1366_, new_n26620_ );
and  ( new_n32518_, new_n32517_, new_n32516_ );
xor  ( new_n32519_, new_n32518_, new_n1129_ );
or   ( new_n32520_, new_n1135_, new_n27396_ );
or   ( new_n32521_, new_n1137_, new_n27085_ );
and  ( new_n32522_, new_n32521_, new_n32520_ );
xor  ( new_n32523_, new_n32522_, new_n896_ );
or   ( new_n32524_, new_n32523_, new_n32519_ );
and  ( new_n32525_, new_n32523_, new_n32519_ );
or   ( new_n32526_, new_n897_, new_n27763_ );
or   ( new_n32527_, new_n899_, new_n27602_ );
and  ( new_n32528_, new_n32527_, new_n32526_ );
xor  ( new_n32529_, new_n32528_, new_n748_ );
or   ( new_n32530_, new_n32529_, new_n32525_ );
and  ( new_n32531_, new_n32530_, new_n32524_ );
or   ( new_n32532_, new_n32531_, new_n32515_ );
and  ( new_n32533_, new_n32531_, new_n32515_ );
or   ( new_n32534_, new_n2122_, new_n25486_ );
or   ( new_n32535_, new_n2124_, new_n25288_ );
and  ( new_n32536_, new_n32535_, new_n32534_ );
xor  ( new_n32537_, new_n32536_, new_n1843_ );
or   ( new_n32538_, new_n1844_, new_n26196_ );
or   ( new_n32539_, new_n1846_, new_n25813_ );
and  ( new_n32540_, new_n32539_, new_n32538_ );
xor  ( new_n32541_, new_n32540_, new_n1586_ );
nor  ( new_n32542_, new_n32541_, new_n32537_ );
and  ( new_n32543_, new_n32541_, new_n32537_ );
or   ( new_n32544_, new_n1593_, new_n26372_ );
or   ( new_n32545_, new_n1595_, new_n26063_ );
and  ( new_n32546_, new_n32545_, new_n32544_ );
xor  ( new_n32547_, new_n32546_, new_n1358_ );
nor  ( new_n32548_, new_n32547_, new_n32543_ );
nor  ( new_n32549_, new_n32548_, new_n32542_ );
or   ( new_n32550_, new_n32549_, new_n32533_ );
and  ( new_n32551_, new_n32550_, new_n32532_ );
or   ( new_n32552_, new_n32551_, new_n32499_ );
or   ( new_n32553_, new_n3117_, new_n24418_ );
or   ( new_n32554_, new_n3119_, new_n24227_ );
and  ( new_n32555_, new_n32554_, new_n32553_ );
xor  ( new_n32556_, new_n32555_, new_n2800_ );
or   ( new_n32557_, new_n2807_, new_n24927_ );
or   ( new_n32558_, new_n2809_, new_n24543_ );
and  ( new_n32559_, new_n32558_, new_n32557_ );
xor  ( new_n32560_, new_n32559_, new_n2424_ );
or   ( new_n32561_, new_n32560_, new_n32556_ );
and  ( new_n32562_, new_n32560_, new_n32556_ );
or   ( new_n32563_, new_n2425_, new_n25048_ );
or   ( new_n32564_, new_n2427_, new_n24925_ );
and  ( new_n32565_, new_n32564_, new_n32563_ );
xor  ( new_n32566_, new_n32565_, new_n2121_ );
or   ( new_n32567_, new_n32566_, new_n32562_ );
and  ( new_n32568_, new_n32567_, new_n32561_ );
or   ( new_n32569_, new_n5604_, new_n22641_ );
or   ( new_n32570_, new_n5606_, new_n22590_ );
and  ( new_n32571_, new_n32570_, new_n32569_ );
xor  ( new_n32572_, new_n32571_, new_n5206_ );
or   ( new_n32573_, new_n5207_, new_n22975_ );
or   ( new_n32574_, new_n5209_, new_n22829_ );
and  ( new_n32575_, new_n32574_, new_n32573_ );
xor  ( new_n32576_, new_n32575_, new_n4708_ );
or   ( new_n32577_, new_n32576_, new_n32572_ );
and  ( new_n32578_, new_n32576_, new_n32572_ );
or   ( new_n32579_, new_n4709_, new_n23166_ );
or   ( new_n32580_, new_n4711_, new_n22973_ );
and  ( new_n32581_, new_n32580_, new_n32579_ );
xor  ( new_n32582_, new_n32581_, new_n4295_ );
or   ( new_n32583_, new_n32582_, new_n32578_ );
and  ( new_n32584_, new_n32583_, new_n32577_ );
or   ( new_n32585_, new_n32584_, new_n32568_ );
and  ( new_n32586_, new_n32584_, new_n32568_ );
or   ( new_n32587_, new_n4302_, new_n23370_ );
or   ( new_n32588_, new_n4304_, new_n23252_ );
and  ( new_n32589_, new_n32588_, new_n32587_ );
xor  ( new_n32590_, new_n32589_, new_n3895_ );
or   ( new_n32591_, new_n3896_, new_n23733_ );
or   ( new_n32592_, new_n3898_, new_n23554_ );
and  ( new_n32593_, new_n32592_, new_n32591_ );
xor  ( new_n32594_, new_n32593_, new_n3460_ );
nor  ( new_n32595_, new_n32594_, new_n32590_ );
and  ( new_n32596_, new_n32594_, new_n32590_ );
or   ( new_n32597_, new_n3461_, new_n24006_ );
or   ( new_n32598_, new_n3463_, new_n23895_ );
and  ( new_n32599_, new_n32598_, new_n32597_ );
xor  ( new_n32600_, new_n32599_, new_n3116_ );
nor  ( new_n32601_, new_n32600_, new_n32596_ );
nor  ( new_n32602_, new_n32601_, new_n32595_ );
or   ( new_n32603_, new_n32602_, new_n32586_ );
and  ( new_n32604_, new_n32603_, new_n32585_ );
and  ( new_n32605_, new_n32551_, new_n32499_ );
or   ( new_n32606_, new_n32605_, new_n32604_ );
and  ( new_n32607_, new_n32606_, new_n32552_ );
or   ( new_n32608_, new_n32607_, new_n32445_ );
and  ( new_n32609_, new_n32607_, new_n32445_ );
xor  ( new_n32610_, new_n32056_, new_n32054_ );
xor  ( new_n32611_, new_n32610_, new_n32060_ );
xnor ( new_n32612_, new_n32196_, new_n32192_ );
xor  ( new_n32613_, new_n32612_, new_n32202_ );
xor  ( new_n32614_, new_n32214_, new_n32208_ );
xor  ( new_n32615_, new_n32614_, new_n263_ );
or   ( new_n32616_, new_n32615_, new_n32613_ );
and  ( new_n32617_, new_n32615_, new_n32613_ );
xnor ( new_n32618_, new_n32226_, new_n32222_ );
xor  ( new_n32619_, new_n32618_, new_n32232_ );
or   ( new_n32620_, new_n32619_, new_n32617_ );
and  ( new_n32621_, new_n32620_, new_n32616_ );
nor  ( new_n32622_, new_n32621_, new_n32611_ );
nand ( new_n32623_, new_n32621_, new_n32611_ );
xor  ( new_n32624_, new_n32051_, new_n32049_ );
and  ( new_n32625_, new_n32624_, new_n32623_ );
or   ( new_n32626_, new_n32625_, new_n32622_ );
or   ( new_n32627_, new_n32626_, new_n32609_ );
and  ( new_n32628_, new_n32627_, new_n32608_ );
or   ( new_n32629_, new_n32628_, new_n32395_ );
nand ( new_n32630_, new_n32628_, new_n32395_ );
xor  ( new_n32631_, new_n32039_, new_n32037_ );
xor  ( new_n32632_, new_n32631_, new_n32043_ );
xor  ( new_n32633_, new_n32025_, new_n32023_ );
xor  ( new_n32634_, new_n32633_, new_n32029_ );
nor  ( new_n32635_, new_n32634_, new_n32632_ );
and  ( new_n32636_, new_n32634_, new_n32632_ );
xor  ( new_n32637_, new_n32062_, new_n32052_ );
xor  ( new_n32638_, new_n32637_, new_n32065_ );
not  ( new_n32639_, new_n32638_ );
nor  ( new_n32640_, new_n32639_, new_n32636_ );
nor  ( new_n32641_, new_n32640_, new_n32635_ );
nand ( new_n32642_, new_n32641_, new_n32630_ );
and  ( new_n32643_, new_n32642_, new_n32629_ );
or   ( new_n32644_, new_n32643_, new_n32369_ );
and  ( new_n32645_, new_n32643_, new_n32369_ );
xor  ( new_n32646_, new_n31743_, new_n31741_ );
xnor ( new_n32647_, new_n32646_, new_n31756_ );
or   ( new_n32648_, new_n32647_, new_n32645_ );
and  ( new_n32649_, new_n32648_, new_n32644_ );
nand ( new_n32650_, new_n32649_, new_n32359_ );
nor  ( new_n32651_, new_n32649_, new_n32359_ );
xor  ( new_n32652_, new_n31724_, new_n31722_ );
xor  ( new_n32653_, new_n32652_, new_n31728_ );
or   ( new_n32654_, new_n32653_, new_n32651_ );
and  ( new_n32655_, new_n32654_, new_n32650_ );
or   ( new_n32656_, new_n32655_, new_n32349_ );
and  ( new_n32657_, new_n32655_, new_n32349_ );
xnor ( new_n32658_, new_n32329_, new_n32327_ );
xor  ( new_n32659_, new_n32658_, new_n32332_ );
or   ( new_n32660_, new_n32659_, new_n32657_ );
and  ( new_n32661_, new_n32660_, new_n32656_ );
nor  ( new_n32662_, new_n32661_, new_n32344_ );
xor  ( new_n32663_, new_n32655_, new_n32349_ );
xor  ( new_n32664_, new_n32663_, new_n32659_ );
xor  ( new_n32665_, new_n32649_, new_n32359_ );
xor  ( new_n32666_, new_n32665_, new_n32653_ );
xnor ( new_n32667_, new_n32643_, new_n32369_ );
xor  ( new_n32668_, new_n32667_, new_n32647_ );
xor  ( new_n32669_, new_n32634_, new_n32632_ );
xor  ( new_n32670_, new_n32669_, new_n32639_ );
xnor ( new_n32671_, new_n32117_, new_n32077_ );
xor  ( new_n32672_, new_n32671_, new_n32132_ );
or   ( new_n32673_, new_n32672_, new_n32670_ );
and  ( new_n32674_, new_n32672_, new_n32670_ );
xor  ( new_n32675_, new_n32238_, new_n32188_ );
xnor ( new_n32676_, new_n32675_, new_n32291_ );
or   ( new_n32677_, new_n32676_, new_n32674_ );
and  ( new_n32678_, new_n32677_, new_n32673_ );
xor  ( new_n32679_, new_n32551_, new_n32499_ );
xor  ( new_n32680_, new_n32679_, new_n32604_ );
xor  ( new_n32681_, new_n32430_, new_n32406_ );
xor  ( new_n32682_, new_n32681_, new_n32443_ );
nor  ( new_n32683_, new_n32682_, new_n32680_ );
nand ( new_n32684_, new_n32682_, new_n32680_ );
xnor ( new_n32685_, new_n32621_, new_n32611_ );
xor  ( new_n32686_, new_n32685_, new_n32624_ );
and  ( new_n32687_, new_n32686_, new_n32684_ );
or   ( new_n32688_, new_n32687_, new_n32683_ );
xnor ( new_n32689_, new_n32383_, new_n32381_ );
xor  ( new_n32690_, new_n32689_, new_n32387_ );
xnor ( new_n32691_, new_n32373_, new_n32371_ );
xor  ( new_n32692_, new_n32691_, new_n32377_ );
nand ( new_n32693_, new_n32692_, new_n32690_ );
nor  ( new_n32694_, new_n32692_, new_n32690_ );
xnor ( new_n32695_, new_n32531_, new_n32515_ );
xor  ( new_n32696_, new_n32695_, new_n32549_ );
xor  ( new_n32697_, new_n32424_, new_n32408_ );
xor  ( new_n32698_, new_n32697_, new_n32428_ );
nor  ( new_n32699_, new_n32698_, new_n32696_ );
and  ( new_n32700_, new_n32698_, new_n32696_ );
xor  ( new_n32701_, new_n32436_, new_n32434_ );
xor  ( new_n32702_, new_n32701_, new_n32441_ );
not  ( new_n32703_, new_n32702_ );
nor  ( new_n32704_, new_n32703_, new_n32700_ );
nor  ( new_n32705_, new_n32704_, new_n32699_ );
or   ( new_n32706_, new_n32705_, new_n32694_ );
and  ( new_n32707_, new_n32706_, new_n32693_ );
or   ( new_n32708_, new_n32707_, new_n32688_ );
and  ( new_n32709_, new_n32707_, new_n32688_ );
or   ( new_n32710_, new_n283_, new_n31654_ );
or   ( new_n32711_, new_n286_, new_n31333_ );
and  ( new_n32712_, new_n32711_, new_n32710_ );
xor  ( new_n32713_, new_n32712_, new_n278_ );
and  ( new_n32714_, new_n295_, RIbb33378_192 );
or   ( new_n32715_, new_n32714_, new_n292_ );
nand ( new_n32716_, new_n32714_, RIbb2f520_3 );
and  ( new_n32717_, new_n32716_, new_n32715_ );
and  ( new_n32718_, new_n32717_, new_n32713_ );
or   ( new_n32719_, new_n299_, new_n31952_ );
or   ( new_n32720_, new_n302_, new_n31654_ );
and  ( new_n32721_, new_n32720_, new_n32719_ );
xor  ( new_n32722_, new_n32721_, new_n293_ );
nor  ( new_n32723_, new_n32722_, new_n32718_ );
nand ( new_n32724_, new_n32722_, new_n32718_ );
or   ( new_n32725_, new_n409_, new_n29619_ );
or   ( new_n32726_, new_n411_, new_n29474_ );
and  ( new_n32727_, new_n32726_, new_n32725_ );
xor  ( new_n32728_, new_n32727_, new_n328_ );
or   ( new_n32729_, new_n337_, new_n30227_ );
or   ( new_n32730_, new_n340_, new_n30120_ );
and  ( new_n32731_, new_n32730_, new_n32729_ );
xor  ( new_n32732_, new_n32731_, new_n332_ );
nor  ( new_n32733_, new_n32732_, new_n32728_ );
and  ( new_n32734_, new_n32732_, new_n32728_ );
or   ( new_n32735_, new_n317_, new_n30798_ );
or   ( new_n32736_, new_n320_, new_n30800_ );
and  ( new_n32737_, new_n32736_, new_n32735_ );
xor  ( new_n32738_, new_n32737_, new_n312_ );
nor  ( new_n32739_, new_n32738_, new_n32734_ );
or   ( new_n32740_, new_n32739_, new_n32733_ );
and  ( new_n32741_, new_n32740_, new_n32724_ );
or   ( new_n32742_, new_n32741_, new_n32723_ );
xnor ( new_n32743_, new_n32541_, new_n32537_ );
xor  ( new_n32744_, new_n32743_, new_n32547_ );
xnor ( new_n32745_, new_n32560_, new_n32556_ );
xor  ( new_n32746_, new_n32745_, new_n32566_ );
or   ( new_n32747_, new_n32746_, new_n32744_ );
and  ( new_n32748_, new_n32746_, new_n32744_ );
xor  ( new_n32749_, new_n32594_, new_n32590_ );
xnor ( new_n32750_, new_n32749_, new_n32600_ );
or   ( new_n32751_, new_n32750_, new_n32748_ );
and  ( new_n32752_, new_n32751_, new_n32747_ );
nor  ( new_n32753_, new_n32752_, new_n32742_ );
nand ( new_n32754_, new_n32752_, new_n32742_ );
xnor ( new_n32755_, new_n32523_, new_n32519_ );
xor  ( new_n32756_, new_n32755_, new_n32529_ );
xnor ( new_n32757_, new_n32507_, new_n32503_ );
xor  ( new_n32758_, new_n32757_, new_n32513_ );
nor  ( new_n32759_, new_n32758_, new_n32756_ );
and  ( new_n32760_, new_n32758_, new_n32756_ );
xor  ( new_n32761_, new_n32416_, new_n32412_ );
xnor ( new_n32762_, new_n32761_, new_n32422_ );
nor  ( new_n32763_, new_n32762_, new_n32760_ );
or   ( new_n32764_, new_n32763_, new_n32759_ );
and  ( new_n32765_, new_n32764_, new_n32754_ );
or   ( new_n32766_, new_n32765_, new_n32753_ );
or   ( new_n32767_, new_n2425_, new_n25288_ );
or   ( new_n32768_, new_n2427_, new_n25048_ );
and  ( new_n32769_, new_n32768_, new_n32767_ );
xor  ( new_n32770_, new_n32769_, new_n2121_ );
or   ( new_n32771_, new_n2122_, new_n25813_ );
or   ( new_n32772_, new_n2124_, new_n25486_ );
and  ( new_n32773_, new_n32772_, new_n32771_ );
xor  ( new_n32774_, new_n32773_, new_n1843_ );
or   ( new_n32775_, new_n32774_, new_n32770_ );
and  ( new_n32776_, new_n32774_, new_n32770_ );
or   ( new_n32777_, new_n1844_, new_n26063_ );
or   ( new_n32778_, new_n1846_, new_n26196_ );
and  ( new_n32779_, new_n32778_, new_n32777_ );
xor  ( new_n32780_, new_n32779_, new_n1586_ );
or   ( new_n32781_, new_n32780_, new_n32776_ );
and  ( new_n32782_, new_n32781_, new_n32775_ );
or   ( new_n32783_, new_n897_, new_n28108_ );
or   ( new_n32784_, new_n899_, new_n27763_ );
and  ( new_n32785_, new_n32784_, new_n32783_ );
xor  ( new_n32786_, new_n32785_, new_n748_ );
or   ( new_n32787_, new_n755_, new_n28531_ );
or   ( new_n32788_, new_n757_, new_n28314_ );
and  ( new_n32789_, new_n32788_, new_n32787_ );
xor  ( new_n32790_, new_n32789_, new_n523_ );
or   ( new_n32791_, new_n32790_, new_n32786_ );
and  ( new_n32792_, new_n32790_, new_n32786_ );
or   ( new_n32793_, new_n524_, new_n29261_ );
or   ( new_n32794_, new_n526_, new_n29263_ );
and  ( new_n32795_, new_n32794_, new_n32793_ );
xor  ( new_n32796_, new_n32795_, new_n403_ );
or   ( new_n32797_, new_n32796_, new_n32792_ );
and  ( new_n32798_, new_n32797_, new_n32791_ );
or   ( new_n32799_, new_n32798_, new_n32782_ );
and  ( new_n32800_, new_n32798_, new_n32782_ );
or   ( new_n32801_, new_n1593_, new_n26620_ );
or   ( new_n32802_, new_n1595_, new_n26372_ );
and  ( new_n32803_, new_n32802_, new_n32801_ );
xor  ( new_n32804_, new_n32803_, new_n1358_ );
or   ( new_n32805_, new_n1364_, new_n27085_ );
or   ( new_n32806_, new_n1366_, new_n26762_ );
and  ( new_n32807_, new_n32806_, new_n32805_ );
xor  ( new_n32808_, new_n32807_, new_n1129_ );
or   ( new_n32809_, new_n32808_, new_n32804_ );
and  ( new_n32810_, new_n32808_, new_n32804_ );
or   ( new_n32811_, new_n1135_, new_n27602_ );
or   ( new_n32812_, new_n1137_, new_n27396_ );
and  ( new_n32813_, new_n32812_, new_n32811_ );
xor  ( new_n32814_, new_n32813_, new_n896_ );
or   ( new_n32815_, new_n32814_, new_n32810_ );
and  ( new_n32816_, new_n32815_, new_n32809_ );
or   ( new_n32817_, new_n32816_, new_n32800_ );
and  ( new_n32818_, new_n32817_, new_n32799_ );
or   ( new_n32819_, new_n7732_, new_n21847_ );
or   ( new_n32820_, new_n7734_, new_n21840_ );
and  ( new_n32821_, new_n32820_, new_n32819_ );
xor  ( new_n32822_, new_n32821_, new_n7177_ );
or   ( new_n32823_, new_n7184_, new_n22129_ );
or   ( new_n32824_, new_n7186_, new_n22098_ );
and  ( new_n32825_, new_n32824_, new_n32823_ );
xor  ( new_n32826_, new_n32825_, new_n6638_ );
nor  ( new_n32827_, new_n32826_, new_n32822_ );
and  ( new_n32828_, new_n32826_, new_n32822_ );
or   ( new_n32829_, new_n6645_, new_n22304_ );
or   ( new_n32830_, new_n6647_, new_n22207_ );
and  ( new_n32831_, new_n32830_, new_n32829_ );
xor  ( new_n32832_, new_n32831_, new_n6166_ );
nor  ( new_n32833_, new_n32832_, new_n32828_ );
nor  ( new_n32834_, new_n32833_, new_n32827_ );
or   ( new_n32835_, new_n10059_, new_n21680_ );
or   ( new_n32836_, new_n10061_, new_n21672_ );
and  ( new_n32837_, new_n32836_, new_n32835_ );
xor  ( new_n32838_, new_n32837_, new_n9421_ );
and  ( new_n32839_, RIbb31758_132, RIbb2d888_64 );
or   ( new_n32840_, new_n21674_, RIbb2d888_64 );
and  ( new_n32841_, new_n32840_, RIbb2d900_63 );
or   ( new_n32842_, new_n32841_, new_n32839_ );
or   ( new_n32843_, new_n10770_, new_n21701_ );
and  ( new_n32844_, new_n32843_, new_n32842_ );
nor  ( new_n32845_, new_n32844_, new_n32838_ );
and  ( new_n32846_, new_n32844_, new_n32838_ );
nor  ( new_n32847_, new_n32846_, new_n292_ );
nor  ( new_n32848_, new_n32847_, new_n32845_ );
or   ( new_n32849_, new_n9422_, new_n21687_ );
or   ( new_n32850_, new_n9424_, new_n21678_ );
and  ( new_n32851_, new_n32850_, new_n32849_ );
xor  ( new_n32852_, new_n32851_, new_n8873_ );
or   ( new_n32853_, new_n8874_, new_n21751_ );
or   ( new_n32854_, new_n8876_, new_n21685_ );
and  ( new_n32855_, new_n32854_, new_n32853_ );
xor  ( new_n32856_, new_n32855_, new_n8257_ );
or   ( new_n32857_, new_n32856_, new_n32852_ );
and  ( new_n32858_, new_n32856_, new_n32852_ );
or   ( new_n32859_, new_n8264_, new_n21842_ );
or   ( new_n32860_, new_n8266_, new_n21792_ );
and  ( new_n32861_, new_n32860_, new_n32859_ );
xor  ( new_n32862_, new_n32861_, new_n7725_ );
or   ( new_n32863_, new_n32862_, new_n32858_ );
and  ( new_n32864_, new_n32863_, new_n32857_ );
and  ( new_n32865_, new_n32864_, new_n32848_ );
or   ( new_n32866_, new_n32865_, new_n32834_ );
or   ( new_n32867_, new_n32864_, new_n32848_ );
and  ( new_n32868_, new_n32867_, new_n32866_ );
or   ( new_n32869_, new_n32868_, new_n32818_ );
or   ( new_n32870_, new_n4709_, new_n23252_ );
or   ( new_n32871_, new_n4711_, new_n23166_ );
and  ( new_n32872_, new_n32871_, new_n32870_ );
xor  ( new_n32873_, new_n32872_, new_n4295_ );
or   ( new_n32874_, new_n4302_, new_n23554_ );
or   ( new_n32875_, new_n4304_, new_n23370_ );
and  ( new_n32876_, new_n32875_, new_n32874_ );
xor  ( new_n32877_, new_n32876_, new_n3895_ );
or   ( new_n32878_, new_n32877_, new_n32873_ );
and  ( new_n32879_, new_n32877_, new_n32873_ );
or   ( new_n32880_, new_n3896_, new_n23895_ );
or   ( new_n32881_, new_n3898_, new_n23733_ );
and  ( new_n32882_, new_n32881_, new_n32880_ );
xor  ( new_n32883_, new_n32882_, new_n3460_ );
or   ( new_n32884_, new_n32883_, new_n32879_ );
and  ( new_n32885_, new_n32884_, new_n32878_ );
or   ( new_n32886_, new_n6173_, new_n22590_ );
or   ( new_n32887_, new_n6175_, new_n22423_ );
and  ( new_n32888_, new_n32887_, new_n32886_ );
xor  ( new_n32889_, new_n32888_, new_n5597_ );
or   ( new_n32890_, new_n5604_, new_n22829_ );
or   ( new_n32891_, new_n5606_, new_n22641_ );
and  ( new_n32892_, new_n32891_, new_n32890_ );
xor  ( new_n32893_, new_n32892_, new_n5206_ );
or   ( new_n32894_, new_n32893_, new_n32889_ );
and  ( new_n32895_, new_n32893_, new_n32889_ );
or   ( new_n32896_, new_n5207_, new_n22973_ );
or   ( new_n32897_, new_n5209_, new_n22975_ );
and  ( new_n32898_, new_n32897_, new_n32896_ );
xor  ( new_n32899_, new_n32898_, new_n4708_ );
or   ( new_n32900_, new_n32899_, new_n32895_ );
and  ( new_n32901_, new_n32900_, new_n32894_ );
or   ( new_n32902_, new_n32901_, new_n32885_ );
and  ( new_n32903_, new_n32901_, new_n32885_ );
or   ( new_n32904_, new_n3461_, new_n24227_ );
or   ( new_n32905_, new_n3463_, new_n24006_ );
and  ( new_n32906_, new_n32905_, new_n32904_ );
xor  ( new_n32907_, new_n32906_, new_n3116_ );
or   ( new_n32908_, new_n3117_, new_n24543_ );
or   ( new_n32909_, new_n3119_, new_n24418_ );
and  ( new_n32910_, new_n32909_, new_n32908_ );
xor  ( new_n32911_, new_n32910_, new_n2800_ );
nor  ( new_n32912_, new_n32911_, new_n32907_ );
and  ( new_n32913_, new_n32911_, new_n32907_ );
or   ( new_n32914_, new_n2807_, new_n24925_ );
or   ( new_n32915_, new_n2809_, new_n24927_ );
and  ( new_n32916_, new_n32915_, new_n32914_ );
xor  ( new_n32917_, new_n32916_, new_n2424_ );
nor  ( new_n32918_, new_n32917_, new_n32913_ );
nor  ( new_n32919_, new_n32918_, new_n32912_ );
or   ( new_n32920_, new_n32919_, new_n32903_ );
and  ( new_n32921_, new_n32920_, new_n32902_ );
and  ( new_n32922_, new_n32868_, new_n32818_ );
or   ( new_n32923_, new_n32922_, new_n32921_ );
and  ( new_n32924_, new_n32923_, new_n32869_ );
and  ( new_n32925_, new_n32924_, new_n32766_ );
nor  ( new_n32926_, new_n32924_, new_n32766_ );
xor  ( new_n32927_, new_n32615_, new_n32613_ );
xor  ( new_n32928_, new_n32927_, new_n32619_ );
xnor ( new_n32929_, new_n32471_, new_n32467_ );
xor  ( new_n32930_, new_n32929_, new_n32477_ );
xnor ( new_n32931_, new_n32576_, new_n32572_ );
xor  ( new_n32932_, new_n32931_, new_n32582_ );
or   ( new_n32933_, new_n32932_, new_n32930_ );
and  ( new_n32934_, new_n32932_, new_n32930_ );
xor  ( new_n32935_, new_n32489_, new_n32485_ );
xnor ( new_n32936_, new_n32935_, new_n32495_ );
or   ( new_n32937_, new_n32936_, new_n32934_ );
and  ( new_n32938_, new_n32937_, new_n32933_ );
nor  ( new_n32939_, new_n32938_, new_n32928_ );
and  ( new_n32940_, new_n32938_, new_n32928_ );
xor  ( new_n32941_, new_n32399_, new_n32397_ );
xor  ( new_n32942_, new_n32941_, new_n32404_ );
not  ( new_n32943_, new_n32942_ );
nor  ( new_n32944_, new_n32943_, new_n32940_ );
nor  ( new_n32945_, new_n32944_, new_n32939_ );
nor  ( new_n32946_, new_n32945_, new_n32926_ );
nor  ( new_n32947_, new_n32946_, new_n32925_ );
or   ( new_n32948_, new_n32947_, new_n32709_ );
and  ( new_n32949_, new_n32948_, new_n32708_ );
or   ( new_n32950_, new_n32949_, new_n32678_ );
and  ( new_n32951_, new_n32949_, new_n32678_ );
xor  ( new_n32952_, new_n32134_, new_n32067_ );
xnor ( new_n32953_, new_n32952_, new_n32294_ );
or   ( new_n32954_, new_n32953_, new_n32951_ );
and  ( new_n32955_, new_n32954_, new_n32950_ );
or   ( new_n32956_, new_n32955_, new_n32668_ );
and  ( new_n32957_, new_n32955_, new_n32668_ );
xor  ( new_n32958_, new_n32353_, new_n32351_ );
xor  ( new_n32959_, new_n32958_, new_n32357_ );
or   ( new_n32960_, new_n32959_, new_n32957_ );
and  ( new_n32961_, new_n32960_, new_n32956_ );
or   ( new_n32962_, new_n32961_, new_n32666_ );
and  ( new_n32963_, new_n32961_, new_n32666_ );
xnor ( new_n32964_, new_n32348_, new_n32346_ );
or   ( new_n32965_, new_n32964_, new_n32963_ );
and  ( new_n32966_, new_n32965_, new_n32962_ );
nor  ( new_n32967_, new_n32966_, new_n32664_ );
xor  ( new_n32968_, new_n32961_, new_n32666_ );
xor  ( new_n32969_, new_n32968_, new_n32964_ );
xor  ( new_n32970_, new_n32628_, new_n32395_ );
xor  ( new_n32971_, new_n32970_, new_n32641_ );
not  ( new_n32972_, new_n32971_ );
xnor ( new_n32973_, new_n32949_, new_n32678_ );
xor  ( new_n32974_, new_n32973_, new_n32953_ );
nand ( new_n32975_, new_n32974_, new_n32972_ );
xnor ( new_n32976_, new_n32363_, new_n32361_ );
xor  ( new_n32977_, new_n32976_, new_n32367_ );
xor  ( new_n32978_, new_n32607_, new_n32445_ );
xor  ( new_n32979_, new_n32978_, new_n32626_ );
xnor ( new_n32980_, new_n32707_, new_n32688_ );
xor  ( new_n32981_, new_n32980_, new_n32947_ );
nand ( new_n32982_, new_n32981_, new_n32979_ );
or   ( new_n32983_, new_n32981_, new_n32979_ );
xor  ( new_n32984_, new_n32672_, new_n32670_ );
xnor ( new_n32985_, new_n32984_, new_n32676_ );
nand ( new_n32986_, new_n32985_, new_n32983_ );
and  ( new_n32987_, new_n32986_, new_n32982_ );
or   ( new_n32988_, new_n32987_, new_n32977_ );
and  ( new_n32989_, new_n32987_, new_n32977_ );
xor  ( new_n32990_, new_n32389_, new_n32379_ );
xor  ( new_n32991_, new_n32990_, new_n32393_ );
xnor ( new_n32992_, new_n32692_, new_n32690_ );
xor  ( new_n32993_, new_n32992_, new_n32705_ );
xnor ( new_n32994_, new_n32924_, new_n32766_ );
xor  ( new_n32995_, new_n32994_, new_n32945_ );
nand ( new_n32996_, new_n32995_, new_n32993_ );
nor  ( new_n32997_, new_n32995_, new_n32993_ );
xor  ( new_n32998_, new_n32682_, new_n32680_ );
xor  ( new_n32999_, new_n32998_, new_n32686_ );
or   ( new_n33000_, new_n32999_, new_n32997_ );
and  ( new_n33001_, new_n33000_, new_n32996_ );
or   ( new_n33002_, new_n33001_, new_n32991_ );
and  ( new_n33003_, new_n33001_, new_n32991_ );
xor  ( new_n33004_, new_n32798_, new_n32782_ );
xor  ( new_n33005_, new_n33004_, new_n32816_ );
xor  ( new_n33006_, new_n32864_, new_n32848_ );
xor  ( new_n33007_, new_n33006_, new_n32834_ );
and  ( new_n33008_, new_n33007_, new_n33005_ );
nor  ( new_n33009_, new_n33007_, new_n33005_ );
xor  ( new_n33010_, new_n32901_, new_n32885_ );
xnor ( new_n33011_, new_n33010_, new_n32919_ );
nor  ( new_n33012_, new_n33011_, new_n33009_ );
or   ( new_n33013_, new_n33012_, new_n33008_ );
xor  ( new_n33014_, new_n32758_, new_n32756_ );
xor  ( new_n33015_, new_n33014_, new_n32762_ );
xor  ( new_n33016_, new_n32722_, new_n32718_ );
xor  ( new_n33017_, new_n33016_, new_n32740_ );
nand ( new_n33018_, new_n33017_, new_n33015_ );
nor  ( new_n33019_, new_n33017_, new_n33015_ );
xor  ( new_n33020_, new_n32746_, new_n32744_ );
xnor ( new_n33021_, new_n33020_, new_n32750_ );
or   ( new_n33022_, new_n33021_, new_n33019_ );
and  ( new_n33023_, new_n33022_, new_n33018_ );
nand ( new_n33024_, new_n33023_, new_n33013_ );
nor  ( new_n33025_, new_n33023_, new_n33013_ );
xor  ( new_n33026_, new_n32584_, new_n32568_ );
xnor ( new_n33027_, new_n33026_, new_n32602_ );
or   ( new_n33028_, new_n33027_, new_n33025_ );
and  ( new_n33029_, new_n33028_, new_n33024_ );
xnor ( new_n33030_, new_n32479_, new_n32463_ );
xor  ( new_n33031_, new_n33030_, new_n32497_ );
xor  ( new_n33032_, new_n32698_, new_n32696_ );
xor  ( new_n33033_, new_n33032_, new_n32703_ );
or   ( new_n33034_, new_n33033_, new_n33031_ );
and  ( new_n33035_, new_n33033_, new_n33031_ );
xor  ( new_n33036_, new_n32938_, new_n32928_ );
xor  ( new_n33037_, new_n33036_, new_n32943_ );
or   ( new_n33038_, new_n33037_, new_n33035_ );
and  ( new_n33039_, new_n33038_, new_n33034_ );
or   ( new_n33040_, new_n33039_, new_n33029_ );
and  ( new_n33041_, new_n33039_, new_n33029_ );
xnor ( new_n33042_, new_n32455_, new_n32449_ );
xor  ( new_n33043_, new_n33042_, new_n32461_ );
xnor ( new_n33044_, new_n32826_, new_n32822_ );
xor  ( new_n33045_, new_n33044_, new_n32832_ );
xnor ( new_n33046_, new_n32856_, new_n32852_ );
xor  ( new_n33047_, new_n33046_, new_n32862_ );
or   ( new_n33048_, new_n33047_, new_n33045_ );
and  ( new_n33049_, new_n33047_, new_n33045_ );
xor  ( new_n33050_, new_n32844_, new_n32838_ );
xor  ( new_n33051_, new_n33050_, new_n293_ );
or   ( new_n33052_, new_n33051_, new_n33049_ );
and  ( new_n33053_, new_n33052_, new_n33048_ );
nor  ( new_n33054_, new_n33053_, new_n33043_ );
nand ( new_n33055_, new_n33053_, new_n33043_ );
xor  ( new_n33056_, new_n32932_, new_n32930_ );
xnor ( new_n33057_, new_n33056_, new_n32936_ );
and  ( new_n33058_, new_n33057_, new_n33055_ );
or   ( new_n33059_, new_n33058_, new_n33054_ );
or   ( new_n33060_, new_n5604_, new_n22975_ );
or   ( new_n33061_, new_n5606_, new_n22829_ );
and  ( new_n33062_, new_n33061_, new_n33060_ );
xor  ( new_n33063_, new_n33062_, new_n5206_ );
or   ( new_n33064_, new_n5207_, new_n23166_ );
or   ( new_n33065_, new_n5209_, new_n22973_ );
and  ( new_n33066_, new_n33065_, new_n33064_ );
xor  ( new_n33067_, new_n33066_, new_n4708_ );
or   ( new_n33068_, new_n33067_, new_n33063_ );
and  ( new_n33069_, new_n33067_, new_n33063_ );
or   ( new_n33070_, new_n4709_, new_n23370_ );
or   ( new_n33071_, new_n4711_, new_n23252_ );
and  ( new_n33072_, new_n33071_, new_n33070_ );
xor  ( new_n33073_, new_n33072_, new_n4295_ );
or   ( new_n33074_, new_n33073_, new_n33069_ );
and  ( new_n33075_, new_n33074_, new_n33068_ );
or   ( new_n33076_, new_n3117_, new_n24927_ );
or   ( new_n33077_, new_n3119_, new_n24543_ );
and  ( new_n33078_, new_n33077_, new_n33076_ );
xor  ( new_n33079_, new_n33078_, new_n2800_ );
or   ( new_n33080_, new_n2807_, new_n25048_ );
or   ( new_n33081_, new_n2809_, new_n24925_ );
and  ( new_n33082_, new_n33081_, new_n33080_ );
xor  ( new_n33083_, new_n33082_, new_n2424_ );
or   ( new_n33084_, new_n33083_, new_n33079_ );
and  ( new_n33085_, new_n33083_, new_n33079_ );
or   ( new_n33086_, new_n2425_, new_n25486_ );
or   ( new_n33087_, new_n2427_, new_n25288_ );
and  ( new_n33088_, new_n33087_, new_n33086_ );
xor  ( new_n33089_, new_n33088_, new_n2121_ );
or   ( new_n33090_, new_n33089_, new_n33085_ );
and  ( new_n33091_, new_n33090_, new_n33084_ );
or   ( new_n33092_, new_n33091_, new_n33075_ );
and  ( new_n33093_, new_n33091_, new_n33075_ );
or   ( new_n33094_, new_n4302_, new_n23733_ );
or   ( new_n33095_, new_n4304_, new_n23554_ );
and  ( new_n33096_, new_n33095_, new_n33094_ );
xor  ( new_n33097_, new_n33096_, new_n3895_ );
or   ( new_n33098_, new_n3896_, new_n24006_ );
or   ( new_n33099_, new_n3898_, new_n23895_ );
and  ( new_n33100_, new_n33099_, new_n33098_ );
xor  ( new_n33101_, new_n33100_, new_n3460_ );
nor  ( new_n33102_, new_n33101_, new_n33097_ );
and  ( new_n33103_, new_n33101_, new_n33097_ );
or   ( new_n33104_, new_n3461_, new_n24418_ );
or   ( new_n33105_, new_n3463_, new_n24227_ );
and  ( new_n33106_, new_n33105_, new_n33104_ );
xor  ( new_n33107_, new_n33106_, new_n3116_ );
nor  ( new_n33108_, new_n33107_, new_n33103_ );
nor  ( new_n33109_, new_n33108_, new_n33102_ );
or   ( new_n33110_, new_n33109_, new_n33093_ );
and  ( new_n33111_, new_n33110_, new_n33092_ );
or   ( new_n33112_, new_n10059_, new_n21678_ );
or   ( new_n33113_, new_n10061_, new_n21680_ );
and  ( new_n33114_, new_n33113_, new_n33112_ );
xor  ( new_n33115_, new_n33114_, new_n9421_ );
and  ( new_n33116_, RIbb317d0_133, RIbb2d888_64 );
or   ( new_n33117_, new_n21672_, RIbb2d888_64 );
and  ( new_n33118_, new_n33117_, RIbb2d900_63 );
or   ( new_n33119_, new_n33118_, new_n33116_ );
or   ( new_n33120_, new_n10770_, new_n21674_ );
and  ( new_n33121_, new_n33120_, new_n33119_ );
or   ( new_n33122_, new_n33121_, new_n33115_ );
and  ( new_n33123_, new_n33121_, new_n33115_ );
or   ( new_n33124_, new_n9422_, new_n21685_ );
or   ( new_n33125_, new_n9424_, new_n21687_ );
and  ( new_n33126_, new_n33125_, new_n33124_ );
xor  ( new_n33127_, new_n33126_, new_n8873_ );
or   ( new_n33128_, new_n33127_, new_n33123_ );
and  ( new_n33129_, new_n33128_, new_n33122_ );
or   ( new_n33130_, new_n7184_, new_n22207_ );
or   ( new_n33131_, new_n7186_, new_n22129_ );
and  ( new_n33132_, new_n33131_, new_n33130_ );
xor  ( new_n33133_, new_n33132_, new_n6638_ );
or   ( new_n33134_, new_n6645_, new_n22423_ );
or   ( new_n33135_, new_n6647_, new_n22304_ );
and  ( new_n33136_, new_n33135_, new_n33134_ );
xor  ( new_n33137_, new_n33136_, new_n6166_ );
or   ( new_n33138_, new_n33137_, new_n33133_ );
and  ( new_n33139_, new_n33137_, new_n33133_ );
or   ( new_n33140_, new_n6173_, new_n22641_ );
or   ( new_n33141_, new_n6175_, new_n22590_ );
and  ( new_n33142_, new_n33141_, new_n33140_ );
xor  ( new_n33143_, new_n33142_, new_n5597_ );
or   ( new_n33144_, new_n33143_, new_n33139_ );
and  ( new_n33145_, new_n33144_, new_n33138_ );
or   ( new_n33146_, new_n33145_, new_n33129_ );
and  ( new_n33147_, new_n33145_, new_n33129_ );
or   ( new_n33148_, new_n8874_, new_n21792_ );
or   ( new_n33149_, new_n8876_, new_n21751_ );
and  ( new_n33150_, new_n33149_, new_n33148_ );
xor  ( new_n33151_, new_n33150_, new_n8257_ );
or   ( new_n33152_, new_n8264_, new_n21840_ );
or   ( new_n33153_, new_n8266_, new_n21842_ );
and  ( new_n33154_, new_n33153_, new_n33152_ );
xor  ( new_n33155_, new_n33154_, new_n7725_ );
nor  ( new_n33156_, new_n33155_, new_n33151_ );
and  ( new_n33157_, new_n33155_, new_n33151_ );
or   ( new_n33158_, new_n7732_, new_n22098_ );
or   ( new_n33159_, new_n7734_, new_n21847_ );
and  ( new_n33160_, new_n33159_, new_n33158_ );
xor  ( new_n33161_, new_n33160_, new_n7177_ );
nor  ( new_n33162_, new_n33161_, new_n33157_ );
nor  ( new_n33163_, new_n33162_, new_n33156_ );
or   ( new_n33164_, new_n33163_, new_n33147_ );
and  ( new_n33165_, new_n33164_, new_n33146_ );
or   ( new_n33166_, new_n33165_, new_n33111_ );
or   ( new_n33167_, new_n755_, new_n29263_ );
or   ( new_n33168_, new_n757_, new_n28531_ );
and  ( new_n33169_, new_n33168_, new_n33167_ );
xor  ( new_n33170_, new_n33169_, new_n523_ );
or   ( new_n33171_, new_n524_, new_n29474_ );
or   ( new_n33172_, new_n526_, new_n29261_ );
and  ( new_n33173_, new_n33172_, new_n33171_ );
xor  ( new_n33174_, new_n33173_, new_n403_ );
or   ( new_n33175_, new_n33174_, new_n33170_ );
and  ( new_n33176_, new_n33174_, new_n33170_ );
or   ( new_n33177_, new_n409_, new_n30120_ );
or   ( new_n33178_, new_n411_, new_n29619_ );
and  ( new_n33179_, new_n33178_, new_n33177_ );
xor  ( new_n33180_, new_n33179_, new_n328_ );
or   ( new_n33181_, new_n33180_, new_n33176_ );
and  ( new_n33182_, new_n33181_, new_n33175_ );
or   ( new_n33183_, new_n2122_, new_n26196_ );
or   ( new_n33184_, new_n2124_, new_n25813_ );
and  ( new_n33185_, new_n33184_, new_n33183_ );
xor  ( new_n33186_, new_n33185_, new_n1843_ );
or   ( new_n33187_, new_n1844_, new_n26372_ );
or   ( new_n33188_, new_n1846_, new_n26063_ );
and  ( new_n33189_, new_n33188_, new_n33187_ );
xor  ( new_n33190_, new_n33189_, new_n1586_ );
or   ( new_n33191_, new_n33190_, new_n33186_ );
and  ( new_n33192_, new_n33190_, new_n33186_ );
or   ( new_n33193_, new_n1593_, new_n26762_ );
or   ( new_n33194_, new_n1595_, new_n26620_ );
and  ( new_n33195_, new_n33194_, new_n33193_ );
xor  ( new_n33196_, new_n33195_, new_n1358_ );
or   ( new_n33197_, new_n33196_, new_n33192_ );
and  ( new_n33198_, new_n33197_, new_n33191_ );
or   ( new_n33199_, new_n33198_, new_n33182_ );
and  ( new_n33200_, new_n33198_, new_n33182_ );
or   ( new_n33201_, new_n1364_, new_n27396_ );
or   ( new_n33202_, new_n1366_, new_n27085_ );
and  ( new_n33203_, new_n33202_, new_n33201_ );
xor  ( new_n33204_, new_n33203_, new_n1129_ );
or   ( new_n33205_, new_n1135_, new_n27763_ );
or   ( new_n33206_, new_n1137_, new_n27602_ );
and  ( new_n33207_, new_n33206_, new_n33205_ );
xor  ( new_n33208_, new_n33207_, new_n896_ );
nor  ( new_n33209_, new_n33208_, new_n33204_ );
and  ( new_n33210_, new_n33208_, new_n33204_ );
or   ( new_n33211_, new_n897_, new_n28314_ );
or   ( new_n33212_, new_n899_, new_n28108_ );
and  ( new_n33213_, new_n33212_, new_n33211_ );
xor  ( new_n33214_, new_n33213_, new_n748_ );
nor  ( new_n33215_, new_n33214_, new_n33210_ );
nor  ( new_n33216_, new_n33215_, new_n33209_ );
or   ( new_n33217_, new_n33216_, new_n33200_ );
and  ( new_n33218_, new_n33217_, new_n33199_ );
and  ( new_n33219_, new_n33165_, new_n33111_ );
or   ( new_n33220_, new_n33219_, new_n33218_ );
and  ( new_n33221_, new_n33220_, new_n33166_ );
nand ( new_n33222_, new_n33221_, new_n33059_ );
nor  ( new_n33223_, new_n33221_, new_n33059_ );
xor  ( new_n33224_, new_n32732_, new_n32728_ );
xor  ( new_n33225_, new_n33224_, new_n32738_ );
or   ( new_n33226_, new_n337_, new_n30800_ );
or   ( new_n33227_, new_n340_, new_n30227_ );
and  ( new_n33228_, new_n33227_, new_n33226_ );
xor  ( new_n33229_, new_n33228_, new_n332_ );
or   ( new_n33230_, new_n317_, new_n31333_ );
or   ( new_n33231_, new_n320_, new_n30798_ );
and  ( new_n33232_, new_n33231_, new_n33230_ );
xor  ( new_n33233_, new_n33232_, new_n312_ );
or   ( new_n33234_, new_n33233_, new_n33229_ );
and  ( new_n33235_, new_n33233_, new_n33229_ );
or   ( new_n33236_, new_n283_, new_n31952_ );
or   ( new_n33237_, new_n286_, new_n31654_ );
and  ( new_n33238_, new_n33237_, new_n33236_ );
xor  ( new_n33239_, new_n33238_, new_n278_ );
or   ( new_n33240_, new_n33239_, new_n33235_ );
and  ( new_n33241_, new_n33240_, new_n33234_ );
nor  ( new_n33242_, new_n33241_, new_n33225_ );
nand ( new_n33243_, new_n33241_, new_n33225_ );
xor  ( new_n33244_, new_n32717_, new_n32713_ );
not  ( new_n33245_, new_n33244_ );
and  ( new_n33246_, new_n33245_, new_n33243_ );
or   ( new_n33247_, new_n33246_, new_n33242_ );
xnor ( new_n33248_, new_n32790_, new_n32786_ );
xor  ( new_n33249_, new_n33248_, new_n32796_ );
xnor ( new_n33250_, new_n32774_, new_n32770_ );
xor  ( new_n33251_, new_n33250_, new_n32780_ );
or   ( new_n33252_, new_n33251_, new_n33249_ );
and  ( new_n33253_, new_n33251_, new_n33249_ );
xor  ( new_n33254_, new_n32808_, new_n32804_ );
xnor ( new_n33255_, new_n33254_, new_n32814_ );
or   ( new_n33256_, new_n33255_, new_n33253_ );
and  ( new_n33257_, new_n33256_, new_n33252_ );
or   ( new_n33258_, new_n33257_, new_n33247_ );
and  ( new_n33259_, new_n33257_, new_n33247_ );
xnor ( new_n33260_, new_n32893_, new_n32889_ );
xor  ( new_n33261_, new_n33260_, new_n32899_ );
xnor ( new_n33262_, new_n32877_, new_n32873_ );
xor  ( new_n33263_, new_n33262_, new_n32883_ );
nor  ( new_n33264_, new_n33263_, new_n33261_ );
and  ( new_n33265_, new_n33263_, new_n33261_ );
xor  ( new_n33266_, new_n32911_, new_n32907_ );
xnor ( new_n33267_, new_n33266_, new_n32917_ );
nor  ( new_n33268_, new_n33267_, new_n33265_ );
nor  ( new_n33269_, new_n33268_, new_n33264_ );
or   ( new_n33270_, new_n33269_, new_n33259_ );
and  ( new_n33271_, new_n33270_, new_n33258_ );
or   ( new_n33272_, new_n33271_, new_n33223_ );
and  ( new_n33273_, new_n33272_, new_n33222_ );
or   ( new_n33274_, new_n33273_, new_n33041_ );
and  ( new_n33275_, new_n33274_, new_n33040_ );
or   ( new_n33276_, new_n33275_, new_n33003_ );
and  ( new_n33277_, new_n33276_, new_n33002_ );
or   ( new_n33278_, new_n33277_, new_n32989_ );
and  ( new_n33279_, new_n33278_, new_n32988_ );
or   ( new_n33280_, new_n33279_, new_n32975_ );
and  ( new_n33281_, new_n33279_, new_n32975_ );
xor  ( new_n33282_, new_n32955_, new_n32668_ );
xor  ( new_n33283_, new_n33282_, new_n32959_ );
or   ( new_n33284_, new_n33283_, new_n33281_ );
and  ( new_n33285_, new_n33284_, new_n33280_ );
nor  ( new_n33286_, new_n33285_, new_n32969_ );
xor  ( new_n33287_, new_n33279_, new_n32975_ );
xor  ( new_n33288_, new_n33287_, new_n33283_ );
xor  ( new_n33289_, new_n32987_, new_n32977_ );
xor  ( new_n33290_, new_n33289_, new_n33277_ );
xor  ( new_n33291_, new_n32995_, new_n32993_ );
xor  ( new_n33292_, new_n33291_, new_n32999_ );
xor  ( new_n33293_, new_n32868_, new_n32818_ );
xor  ( new_n33294_, new_n33293_, new_n32921_ );
xor  ( new_n33295_, new_n32752_, new_n32742_ );
xor  ( new_n33296_, new_n33295_, new_n32764_ );
nand ( new_n33297_, new_n33296_, new_n33294_ );
nor  ( new_n33298_, new_n33296_, new_n33294_ );
xor  ( new_n33299_, new_n33033_, new_n33031_ );
xor  ( new_n33300_, new_n33299_, new_n33037_ );
or   ( new_n33301_, new_n33300_, new_n33298_ );
and  ( new_n33302_, new_n33301_, new_n33297_ );
or   ( new_n33303_, new_n33302_, new_n33292_ );
and  ( new_n33304_, new_n33302_, new_n33292_ );
xor  ( new_n33305_, new_n33007_, new_n33005_ );
xor  ( new_n33306_, new_n33305_, new_n33011_ );
xnor ( new_n33307_, new_n33017_, new_n33015_ );
xor  ( new_n33308_, new_n33307_, new_n33021_ );
or   ( new_n33309_, new_n33308_, new_n33306_ );
and  ( new_n33310_, new_n33308_, new_n33306_ );
xnor ( new_n33311_, new_n33091_, new_n33075_ );
xor  ( new_n33312_, new_n33311_, new_n33109_ );
xnor ( new_n33313_, new_n33198_, new_n33182_ );
xor  ( new_n33314_, new_n33313_, new_n33216_ );
nor  ( new_n33315_, new_n33314_, new_n33312_ );
and  ( new_n33316_, new_n33314_, new_n33312_ );
xor  ( new_n33317_, new_n33241_, new_n33225_ );
xor  ( new_n33318_, new_n33317_, new_n33245_ );
nor  ( new_n33319_, new_n33318_, new_n33316_ );
nor  ( new_n33320_, new_n33319_, new_n33315_ );
or   ( new_n33321_, new_n33320_, new_n33310_ );
and  ( new_n33322_, new_n33321_, new_n33309_ );
xor  ( new_n33323_, new_n33165_, new_n33111_ );
xor  ( new_n33324_, new_n33323_, new_n33218_ );
xnor ( new_n33325_, new_n33257_, new_n33247_ );
xor  ( new_n33326_, new_n33325_, new_n33269_ );
nand ( new_n33327_, new_n33326_, new_n33324_ );
nor  ( new_n33328_, new_n33326_, new_n33324_ );
xnor ( new_n33329_, new_n33053_, new_n33043_ );
xor  ( new_n33330_, new_n33329_, new_n33057_ );
or   ( new_n33331_, new_n33330_, new_n33328_ );
and  ( new_n33332_, new_n33331_, new_n33327_ );
and  ( new_n33333_, new_n33332_, new_n33322_ );
nor  ( new_n33334_, new_n33332_, new_n33322_ );
xnor ( new_n33335_, new_n33047_, new_n33045_ );
xor  ( new_n33336_, new_n33335_, new_n33051_ );
xnor ( new_n33337_, new_n33251_, new_n33249_ );
xor  ( new_n33338_, new_n33337_, new_n33255_ );
or   ( new_n33339_, new_n33338_, new_n33336_ );
and  ( new_n33340_, new_n33338_, new_n33336_ );
xnor ( new_n33341_, new_n33263_, new_n33261_ );
xor  ( new_n33342_, new_n33341_, new_n33267_ );
or   ( new_n33343_, new_n33342_, new_n33340_ );
and  ( new_n33344_, new_n33343_, new_n33339_ );
or   ( new_n33345_, new_n4709_, new_n23554_ );
or   ( new_n33346_, new_n4711_, new_n23370_ );
and  ( new_n33347_, new_n33346_, new_n33345_ );
xor  ( new_n33348_, new_n33347_, new_n4295_ );
or   ( new_n33349_, new_n4302_, new_n23895_ );
or   ( new_n33350_, new_n4304_, new_n23733_ );
and  ( new_n33351_, new_n33350_, new_n33349_ );
xor  ( new_n33352_, new_n33351_, new_n3895_ );
or   ( new_n33353_, new_n33352_, new_n33348_ );
and  ( new_n33354_, new_n33352_, new_n33348_ );
or   ( new_n33355_, new_n3896_, new_n24227_ );
or   ( new_n33356_, new_n3898_, new_n24006_ );
and  ( new_n33357_, new_n33356_, new_n33355_ );
xor  ( new_n33358_, new_n33357_, new_n3460_ );
or   ( new_n33359_, new_n33358_, new_n33354_ );
and  ( new_n33360_, new_n33359_, new_n33353_ );
or   ( new_n33361_, new_n3461_, new_n24543_ );
or   ( new_n33362_, new_n3463_, new_n24418_ );
and  ( new_n33363_, new_n33362_, new_n33361_ );
xor  ( new_n33364_, new_n33363_, new_n3116_ );
or   ( new_n33365_, new_n3117_, new_n24925_ );
or   ( new_n33366_, new_n3119_, new_n24927_ );
and  ( new_n33367_, new_n33366_, new_n33365_ );
xor  ( new_n33368_, new_n33367_, new_n2800_ );
or   ( new_n33369_, new_n33368_, new_n33364_ );
and  ( new_n33370_, new_n33368_, new_n33364_ );
or   ( new_n33371_, new_n2807_, new_n25288_ );
or   ( new_n33372_, new_n2809_, new_n25048_ );
and  ( new_n33373_, new_n33372_, new_n33371_ );
xor  ( new_n33374_, new_n33373_, new_n2424_ );
or   ( new_n33375_, new_n33374_, new_n33370_ );
and  ( new_n33376_, new_n33375_, new_n33369_ );
or   ( new_n33377_, new_n33376_, new_n33360_ );
and  ( new_n33378_, new_n33376_, new_n33360_ );
or   ( new_n33379_, new_n6173_, new_n22829_ );
or   ( new_n33380_, new_n6175_, new_n22641_ );
and  ( new_n33381_, new_n33380_, new_n33379_ );
xor  ( new_n33382_, new_n33381_, new_n5597_ );
or   ( new_n33383_, new_n5604_, new_n22973_ );
or   ( new_n33384_, new_n5606_, new_n22975_ );
and  ( new_n33385_, new_n33384_, new_n33383_ );
xor  ( new_n33386_, new_n33385_, new_n5206_ );
nor  ( new_n33387_, new_n33386_, new_n33382_ );
and  ( new_n33388_, new_n33386_, new_n33382_ );
or   ( new_n33389_, new_n5207_, new_n23252_ );
or   ( new_n33390_, new_n5209_, new_n23166_ );
and  ( new_n33391_, new_n33390_, new_n33389_ );
xor  ( new_n33392_, new_n33391_, new_n4708_ );
nor  ( new_n33393_, new_n33392_, new_n33388_ );
nor  ( new_n33394_, new_n33393_, new_n33387_ );
or   ( new_n33395_, new_n33394_, new_n33378_ );
and  ( new_n33396_, new_n33395_, new_n33377_ );
or   ( new_n33397_, new_n7732_, new_n22129_ );
or   ( new_n33398_, new_n7734_, new_n22098_ );
and  ( new_n33399_, new_n33398_, new_n33397_ );
xor  ( new_n33400_, new_n33399_, new_n7177_ );
or   ( new_n33401_, new_n7184_, new_n22304_ );
or   ( new_n33402_, new_n7186_, new_n22207_ );
and  ( new_n33403_, new_n33402_, new_n33401_ );
xor  ( new_n33404_, new_n33403_, new_n6638_ );
or   ( new_n33405_, new_n33404_, new_n33400_ );
and  ( new_n33406_, new_n33404_, new_n33400_ );
or   ( new_n33407_, new_n6645_, new_n22590_ );
or   ( new_n33408_, new_n6647_, new_n22423_ );
and  ( new_n33409_, new_n33408_, new_n33407_ );
xor  ( new_n33410_, new_n33409_, new_n6166_ );
or   ( new_n33411_, new_n33410_, new_n33406_ );
and  ( new_n33412_, new_n33411_, new_n33405_ );
or   ( new_n33413_, new_n10059_, new_n21687_ );
or   ( new_n33414_, new_n10061_, new_n21678_ );
and  ( new_n33415_, new_n33414_, new_n33413_ );
xor  ( new_n33416_, new_n33415_, new_n9421_ );
and  ( new_n33417_, RIbb31848_134, RIbb2d888_64 );
or   ( new_n33418_, new_n21680_, RIbb2d888_64 );
and  ( new_n33419_, new_n33418_, RIbb2d900_63 );
or   ( new_n33420_, new_n33419_, new_n33417_ );
or   ( new_n33421_, new_n10770_, new_n21672_ );
and  ( new_n33422_, new_n33421_, new_n33420_ );
nor  ( new_n33423_, new_n33422_, new_n33416_ );
and  ( new_n33424_, new_n33422_, new_n33416_ );
nor  ( new_n33425_, new_n33424_, new_n277_ );
nor  ( new_n33426_, new_n33425_, new_n33423_ );
or   ( new_n33427_, new_n9422_, new_n21751_ );
or   ( new_n33428_, new_n9424_, new_n21685_ );
and  ( new_n33429_, new_n33428_, new_n33427_ );
xor  ( new_n33430_, new_n33429_, new_n8873_ );
or   ( new_n33431_, new_n8874_, new_n21842_ );
or   ( new_n33432_, new_n8876_, new_n21792_ );
and  ( new_n33433_, new_n33432_, new_n33431_ );
xor  ( new_n33434_, new_n33433_, new_n8257_ );
or   ( new_n33435_, new_n33434_, new_n33430_ );
and  ( new_n33436_, new_n33434_, new_n33430_ );
or   ( new_n33437_, new_n8264_, new_n21847_ );
or   ( new_n33438_, new_n8266_, new_n21840_ );
and  ( new_n33439_, new_n33438_, new_n33437_ );
xor  ( new_n33440_, new_n33439_, new_n7725_ );
or   ( new_n33441_, new_n33440_, new_n33436_ );
and  ( new_n33442_, new_n33441_, new_n33435_ );
and  ( new_n33443_, new_n33442_, new_n33426_ );
or   ( new_n33444_, new_n33443_, new_n33412_ );
or   ( new_n33445_, new_n33442_, new_n33426_ );
and  ( new_n33446_, new_n33445_, new_n33444_ );
or   ( new_n33447_, new_n33446_, new_n33396_ );
or   ( new_n33448_, new_n1593_, new_n27085_ );
or   ( new_n33449_, new_n1595_, new_n26762_ );
and  ( new_n33450_, new_n33449_, new_n33448_ );
xor  ( new_n33451_, new_n33450_, new_n1358_ );
or   ( new_n33452_, new_n1364_, new_n27602_ );
or   ( new_n33453_, new_n1366_, new_n27396_ );
and  ( new_n33454_, new_n33453_, new_n33452_ );
xor  ( new_n33455_, new_n33454_, new_n1129_ );
or   ( new_n33456_, new_n33455_, new_n33451_ );
and  ( new_n33457_, new_n33455_, new_n33451_ );
or   ( new_n33458_, new_n1135_, new_n28108_ );
or   ( new_n33459_, new_n1137_, new_n27763_ );
and  ( new_n33460_, new_n33459_, new_n33458_ );
xor  ( new_n33461_, new_n33460_, new_n896_ );
or   ( new_n33462_, new_n33461_, new_n33457_ );
and  ( new_n33463_, new_n33462_, new_n33456_ );
or   ( new_n33464_, new_n2425_, new_n25813_ );
or   ( new_n33465_, new_n2427_, new_n25486_ );
and  ( new_n33466_, new_n33465_, new_n33464_ );
xor  ( new_n33467_, new_n33466_, new_n2121_ );
or   ( new_n33468_, new_n2122_, new_n26063_ );
or   ( new_n33469_, new_n2124_, new_n26196_ );
and  ( new_n33470_, new_n33469_, new_n33468_ );
xor  ( new_n33471_, new_n33470_, new_n1843_ );
or   ( new_n33472_, new_n33471_, new_n33467_ );
and  ( new_n33473_, new_n33471_, new_n33467_ );
or   ( new_n33474_, new_n1844_, new_n26620_ );
or   ( new_n33475_, new_n1846_, new_n26372_ );
and  ( new_n33476_, new_n33475_, new_n33474_ );
xor  ( new_n33477_, new_n33476_, new_n1586_ );
or   ( new_n33478_, new_n33477_, new_n33473_ );
and  ( new_n33479_, new_n33478_, new_n33472_ );
nor  ( new_n33480_, new_n33479_, new_n33463_ );
and  ( new_n33481_, new_n33479_, new_n33463_ );
or   ( new_n33482_, new_n897_, new_n28531_ );
or   ( new_n33483_, new_n899_, new_n28314_ );
and  ( new_n33484_, new_n33483_, new_n33482_ );
xor  ( new_n33485_, new_n33484_, new_n748_ );
or   ( new_n33486_, new_n755_, new_n29261_ );
or   ( new_n33487_, new_n757_, new_n29263_ );
and  ( new_n33488_, new_n33487_, new_n33486_ );
xor  ( new_n33489_, new_n33488_, new_n523_ );
nor  ( new_n33490_, new_n33489_, new_n33485_ );
and  ( new_n33491_, new_n33489_, new_n33485_ );
or   ( new_n33492_, new_n524_, new_n29619_ );
or   ( new_n33493_, new_n526_, new_n29474_ );
and  ( new_n33494_, new_n33493_, new_n33492_ );
xor  ( new_n33495_, new_n33494_, new_n403_ );
nor  ( new_n33496_, new_n33495_, new_n33491_ );
nor  ( new_n33497_, new_n33496_, new_n33490_ );
nor  ( new_n33498_, new_n33497_, new_n33481_ );
nor  ( new_n33499_, new_n33498_, new_n33480_ );
and  ( new_n33500_, new_n33446_, new_n33396_ );
or   ( new_n33501_, new_n33500_, new_n33499_ );
and  ( new_n33502_, new_n33501_, new_n33447_ );
nor  ( new_n33503_, new_n33502_, new_n33344_ );
and  ( new_n33504_, new_n33502_, new_n33344_ );
xnor ( new_n33505_, new_n33083_, new_n33079_ );
xor  ( new_n33506_, new_n33505_, new_n33089_ );
xnor ( new_n33507_, new_n33190_, new_n33186_ );
xor  ( new_n33508_, new_n33507_, new_n33196_ );
nor  ( new_n33509_, new_n33508_, new_n33506_ );
nand ( new_n33510_, new_n33508_, new_n33506_ );
xor  ( new_n33511_, new_n33208_, new_n33204_ );
xor  ( new_n33512_, new_n33511_, new_n33214_ );
and  ( new_n33513_, new_n33512_, new_n33510_ );
or   ( new_n33514_, new_n33513_, new_n33509_ );
xor  ( new_n33515_, new_n33233_, new_n33229_ );
xor  ( new_n33516_, new_n33515_, new_n33239_ );
or   ( new_n33517_, new_n409_, new_n30227_ );
or   ( new_n33518_, new_n411_, new_n30120_ );
and  ( new_n33519_, new_n33518_, new_n33517_ );
xor  ( new_n33520_, new_n33519_, new_n328_ );
or   ( new_n33521_, new_n337_, new_n30798_ );
or   ( new_n33522_, new_n340_, new_n30800_ );
and  ( new_n33523_, new_n33522_, new_n33521_ );
xor  ( new_n33524_, new_n33523_, new_n332_ );
or   ( new_n33525_, new_n33524_, new_n33520_ );
and  ( new_n33526_, new_n33524_, new_n33520_ );
or   ( new_n33527_, new_n317_, new_n31654_ );
or   ( new_n33528_, new_n320_, new_n31333_ );
and  ( new_n33529_, new_n33528_, new_n33527_ );
xor  ( new_n33530_, new_n33529_, new_n312_ );
or   ( new_n33531_, new_n33530_, new_n33526_ );
and  ( new_n33532_, new_n33531_, new_n33525_ );
or   ( new_n33533_, new_n33532_, new_n33516_ );
nand ( new_n33534_, new_n33532_, new_n33516_ );
xor  ( new_n33535_, new_n33174_, new_n33170_ );
xnor ( new_n33536_, new_n33535_, new_n33180_ );
nand ( new_n33537_, new_n33536_, new_n33534_ );
and  ( new_n33538_, new_n33537_, new_n33533_ );
and  ( new_n33539_, new_n33538_, new_n33514_ );
nor  ( new_n33540_, new_n33538_, new_n33514_ );
xnor ( new_n33541_, new_n33137_, new_n33133_ );
xor  ( new_n33542_, new_n33541_, new_n33143_ );
xnor ( new_n33543_, new_n33067_, new_n33063_ );
xor  ( new_n33544_, new_n33543_, new_n33073_ );
nor  ( new_n33545_, new_n33544_, new_n33542_ );
and  ( new_n33546_, new_n33544_, new_n33542_ );
xor  ( new_n33547_, new_n33101_, new_n33097_ );
xnor ( new_n33548_, new_n33547_, new_n33107_ );
nor  ( new_n33549_, new_n33548_, new_n33546_ );
nor  ( new_n33550_, new_n33549_, new_n33545_ );
nor  ( new_n33551_, new_n33550_, new_n33540_ );
nor  ( new_n33552_, new_n33551_, new_n33539_ );
not  ( new_n33553_, new_n33552_ );
nor  ( new_n33554_, new_n33553_, new_n33504_ );
nor  ( new_n33555_, new_n33554_, new_n33503_ );
nor  ( new_n33556_, new_n33555_, new_n33334_ );
nor  ( new_n33557_, new_n33556_, new_n33333_ );
not  ( new_n33558_, new_n33557_ );
or   ( new_n33559_, new_n33558_, new_n33304_ );
and  ( new_n33560_, new_n33559_, new_n33303_ );
xor  ( new_n33561_, new_n33001_, new_n32991_ );
xor  ( new_n33562_, new_n33561_, new_n33275_ );
or   ( new_n33563_, new_n33562_, new_n33560_ );
and  ( new_n33564_, new_n33562_, new_n33560_ );
xor  ( new_n33565_, new_n32981_, new_n32979_ );
xor  ( new_n33566_, new_n33565_, new_n32985_ );
not  ( new_n33567_, new_n33566_ );
or   ( new_n33568_, new_n33567_, new_n33564_ );
and  ( new_n33569_, new_n33568_, new_n33563_ );
or   ( new_n33570_, new_n33569_, new_n33290_ );
nand ( new_n33571_, new_n33569_, new_n33290_ );
xor  ( new_n33572_, new_n32974_, new_n32972_ );
nand ( new_n33573_, new_n33572_, new_n33571_ );
and  ( new_n33574_, new_n33573_, new_n33570_ );
nor  ( new_n33575_, new_n33574_, new_n33288_ );
xor  ( new_n33576_, new_n33562_, new_n33560_ );
xor  ( new_n33577_, new_n33576_, new_n33567_ );
xor  ( new_n33578_, new_n33039_, new_n33029_ );
xor  ( new_n33579_, new_n33578_, new_n33273_ );
xnor ( new_n33580_, new_n33023_, new_n33013_ );
xor  ( new_n33581_, new_n33580_, new_n33027_ );
xor  ( new_n33582_, new_n33538_, new_n33514_ );
xor  ( new_n33583_, new_n33582_, new_n33550_ );
xnor ( new_n33584_, new_n33446_, new_n33396_ );
xor  ( new_n33585_, new_n33584_, new_n33499_ );
nor  ( new_n33586_, new_n33585_, new_n33583_ );
nand ( new_n33587_, new_n33585_, new_n33583_ );
xor  ( new_n33588_, new_n33338_, new_n33336_ );
xor  ( new_n33589_, new_n33588_, new_n33342_ );
and  ( new_n33590_, new_n33589_, new_n33587_ );
or   ( new_n33591_, new_n33590_, new_n33586_ );
xor  ( new_n33592_, new_n33524_, new_n33520_ );
xor  ( new_n33593_, new_n33592_, new_n33530_ );
and  ( new_n33594_, new_n280_, RIbb33378_192 );
or   ( new_n33595_, new_n33594_, new_n277_ );
nand ( new_n33596_, new_n33594_, RIbb2f430_5 );
and  ( new_n33597_, new_n33596_, new_n33595_ );
nor  ( new_n33598_, new_n33597_, new_n33593_ );
nand ( new_n33599_, new_n33597_, new_n33593_ );
xor  ( new_n33600_, new_n33489_, new_n33485_ );
xnor ( new_n33601_, new_n33600_, new_n33495_ );
and  ( new_n33602_, new_n33601_, new_n33599_ );
or   ( new_n33603_, new_n33602_, new_n33598_ );
xnor ( new_n33604_, new_n33404_, new_n33400_ );
xor  ( new_n33605_, new_n33604_, new_n33410_ );
xnor ( new_n33606_, new_n33352_, new_n33348_ );
xor  ( new_n33607_, new_n33606_, new_n33358_ );
or   ( new_n33608_, new_n33607_, new_n33605_ );
and  ( new_n33609_, new_n33607_, new_n33605_ );
xor  ( new_n33610_, new_n33386_, new_n33382_ );
xnor ( new_n33611_, new_n33610_, new_n33392_ );
or   ( new_n33612_, new_n33611_, new_n33609_ );
and  ( new_n33613_, new_n33612_, new_n33608_ );
nor  ( new_n33614_, new_n33613_, new_n33603_ );
nand ( new_n33615_, new_n33613_, new_n33603_ );
xnor ( new_n33616_, new_n33368_, new_n33364_ );
xor  ( new_n33617_, new_n33616_, new_n33374_ );
xnor ( new_n33618_, new_n33471_, new_n33467_ );
xor  ( new_n33619_, new_n33618_, new_n33477_ );
nor  ( new_n33620_, new_n33619_, new_n33617_ );
nand ( new_n33621_, new_n33619_, new_n33617_ );
xor  ( new_n33622_, new_n33455_, new_n33451_ );
xor  ( new_n33623_, new_n33622_, new_n33461_ );
and  ( new_n33624_, new_n33623_, new_n33621_ );
or   ( new_n33625_, new_n33624_, new_n33620_ );
and  ( new_n33626_, new_n33625_, new_n33615_ );
or   ( new_n33627_, new_n33626_, new_n33614_ );
or   ( new_n33628_, new_n3117_, new_n25048_ );
or   ( new_n33629_, new_n3119_, new_n24925_ );
and  ( new_n33630_, new_n33629_, new_n33628_ );
xor  ( new_n33631_, new_n33630_, new_n2800_ );
or   ( new_n33632_, new_n2807_, new_n25486_ );
or   ( new_n33633_, new_n2809_, new_n25288_ );
and  ( new_n33634_, new_n33633_, new_n33632_ );
xor  ( new_n33635_, new_n33634_, new_n2424_ );
or   ( new_n33636_, new_n33635_, new_n33631_ );
and  ( new_n33637_, new_n33635_, new_n33631_ );
or   ( new_n33638_, new_n2425_, new_n26196_ );
or   ( new_n33639_, new_n2427_, new_n25813_ );
and  ( new_n33640_, new_n33639_, new_n33638_ );
xor  ( new_n33641_, new_n33640_, new_n2121_ );
or   ( new_n33642_, new_n33641_, new_n33637_ );
and  ( new_n33643_, new_n33642_, new_n33636_ );
or   ( new_n33644_, new_n4302_, new_n24006_ );
or   ( new_n33645_, new_n4304_, new_n23895_ );
and  ( new_n33646_, new_n33645_, new_n33644_ );
xor  ( new_n33647_, new_n33646_, new_n3895_ );
or   ( new_n33648_, new_n3896_, new_n24418_ );
or   ( new_n33649_, new_n3898_, new_n24227_ );
and  ( new_n33650_, new_n33649_, new_n33648_ );
xor  ( new_n33651_, new_n33650_, new_n3460_ );
or   ( new_n33652_, new_n33651_, new_n33647_ );
and  ( new_n33653_, new_n33651_, new_n33647_ );
or   ( new_n33654_, new_n3461_, new_n24927_ );
or   ( new_n33655_, new_n3463_, new_n24543_ );
and  ( new_n33656_, new_n33655_, new_n33654_ );
xor  ( new_n33657_, new_n33656_, new_n3116_ );
or   ( new_n33658_, new_n33657_, new_n33653_ );
and  ( new_n33659_, new_n33658_, new_n33652_ );
or   ( new_n33660_, new_n33659_, new_n33643_ );
and  ( new_n33661_, new_n33659_, new_n33643_ );
or   ( new_n33662_, new_n5604_, new_n23166_ );
or   ( new_n33663_, new_n5606_, new_n22973_ );
and  ( new_n33664_, new_n33663_, new_n33662_ );
xor  ( new_n33665_, new_n33664_, new_n5206_ );
or   ( new_n33666_, new_n5207_, new_n23370_ );
or   ( new_n33667_, new_n5209_, new_n23252_ );
and  ( new_n33668_, new_n33667_, new_n33666_ );
xor  ( new_n33669_, new_n33668_, new_n4708_ );
nor  ( new_n33670_, new_n33669_, new_n33665_ );
and  ( new_n33671_, new_n33669_, new_n33665_ );
or   ( new_n33672_, new_n4709_, new_n23733_ );
or   ( new_n33673_, new_n4711_, new_n23554_ );
and  ( new_n33674_, new_n33673_, new_n33672_ );
xor  ( new_n33675_, new_n33674_, new_n4295_ );
nor  ( new_n33676_, new_n33675_, new_n33671_ );
nor  ( new_n33677_, new_n33676_, new_n33670_ );
or   ( new_n33678_, new_n33677_, new_n33661_ );
and  ( new_n33679_, new_n33678_, new_n33660_ );
or   ( new_n33680_, new_n755_, new_n29474_ );
or   ( new_n33681_, new_n757_, new_n29261_ );
and  ( new_n33682_, new_n33681_, new_n33680_ );
xor  ( new_n33683_, new_n33682_, new_n523_ );
or   ( new_n33684_, new_n524_, new_n30120_ );
or   ( new_n33685_, new_n526_, new_n29619_ );
and  ( new_n33686_, new_n33685_, new_n33684_ );
xor  ( new_n33687_, new_n33686_, new_n403_ );
or   ( new_n33688_, new_n33687_, new_n33683_ );
and  ( new_n33689_, new_n33687_, new_n33683_ );
or   ( new_n33690_, new_n409_, new_n30800_ );
or   ( new_n33691_, new_n411_, new_n30227_ );
and  ( new_n33692_, new_n33691_, new_n33690_ );
xor  ( new_n33693_, new_n33692_, new_n328_ );
or   ( new_n33694_, new_n33693_, new_n33689_ );
and  ( new_n33695_, new_n33694_, new_n33688_ );
or   ( new_n33696_, new_n1364_, new_n27763_ );
or   ( new_n33697_, new_n1366_, new_n27602_ );
and  ( new_n33698_, new_n33697_, new_n33696_ );
xor  ( new_n33699_, new_n33698_, new_n1129_ );
or   ( new_n33700_, new_n1135_, new_n28314_ );
or   ( new_n33701_, new_n1137_, new_n28108_ );
and  ( new_n33702_, new_n33701_, new_n33700_ );
xor  ( new_n33703_, new_n33702_, new_n896_ );
or   ( new_n33704_, new_n33703_, new_n33699_ );
and  ( new_n33705_, new_n33703_, new_n33699_ );
or   ( new_n33706_, new_n897_, new_n29263_ );
or   ( new_n33707_, new_n899_, new_n28531_ );
and  ( new_n33708_, new_n33707_, new_n33706_ );
xor  ( new_n33709_, new_n33708_, new_n748_ );
or   ( new_n33710_, new_n33709_, new_n33705_ );
and  ( new_n33711_, new_n33710_, new_n33704_ );
or   ( new_n33712_, new_n33711_, new_n33695_ );
and  ( new_n33713_, new_n33711_, new_n33695_ );
or   ( new_n33714_, new_n2122_, new_n26372_ );
or   ( new_n33715_, new_n2124_, new_n26063_ );
and  ( new_n33716_, new_n33715_, new_n33714_ );
xor  ( new_n33717_, new_n33716_, new_n1843_ );
or   ( new_n33718_, new_n1844_, new_n26762_ );
or   ( new_n33719_, new_n1846_, new_n26620_ );
and  ( new_n33720_, new_n33719_, new_n33718_ );
xor  ( new_n33721_, new_n33720_, new_n1586_ );
nor  ( new_n33722_, new_n33721_, new_n33717_ );
and  ( new_n33723_, new_n33721_, new_n33717_ );
or   ( new_n33724_, new_n1593_, new_n27396_ );
or   ( new_n33725_, new_n1595_, new_n27085_ );
and  ( new_n33726_, new_n33725_, new_n33724_ );
xor  ( new_n33727_, new_n33726_, new_n1358_ );
nor  ( new_n33728_, new_n33727_, new_n33723_ );
nor  ( new_n33729_, new_n33728_, new_n33722_ );
or   ( new_n33730_, new_n33729_, new_n33713_ );
and  ( new_n33731_, new_n33730_, new_n33712_ );
or   ( new_n33732_, new_n33731_, new_n33679_ );
or   ( new_n33733_, new_n8874_, new_n21840_ );
or   ( new_n33734_, new_n8876_, new_n21842_ );
and  ( new_n33735_, new_n33734_, new_n33733_ );
xor  ( new_n33736_, new_n33735_, new_n8257_ );
or   ( new_n33737_, new_n8264_, new_n22098_ );
or   ( new_n33738_, new_n8266_, new_n21847_ );
and  ( new_n33739_, new_n33738_, new_n33737_ );
xor  ( new_n33740_, new_n33739_, new_n7725_ );
or   ( new_n33741_, new_n33740_, new_n33736_ );
and  ( new_n33742_, new_n33740_, new_n33736_ );
or   ( new_n33743_, new_n7732_, new_n22207_ );
or   ( new_n33744_, new_n7734_, new_n22129_ );
and  ( new_n33745_, new_n33744_, new_n33743_ );
xor  ( new_n33746_, new_n33745_, new_n7177_ );
or   ( new_n33747_, new_n33746_, new_n33742_ );
and  ( new_n33748_, new_n33747_, new_n33741_ );
or   ( new_n33749_, new_n10059_, new_n21685_ );
or   ( new_n33750_, new_n10061_, new_n21687_ );
and  ( new_n33751_, new_n33750_, new_n33749_ );
xor  ( new_n33752_, new_n33751_, new_n9421_ );
and  ( new_n33753_, RIbb318c0_135, RIbb2d888_64 );
or   ( new_n33754_, new_n21678_, RIbb2d888_64 );
and  ( new_n33755_, new_n33754_, RIbb2d900_63 );
or   ( new_n33756_, new_n33755_, new_n33753_ );
or   ( new_n33757_, new_n10770_, new_n21680_ );
and  ( new_n33758_, new_n33757_, new_n33756_ );
or   ( new_n33759_, new_n33758_, new_n33752_ );
and  ( new_n33760_, new_n33758_, new_n33752_ );
or   ( new_n33761_, new_n9422_, new_n21792_ );
or   ( new_n33762_, new_n9424_, new_n21751_ );
and  ( new_n33763_, new_n33762_, new_n33761_ );
xor  ( new_n33764_, new_n33763_, new_n8873_ );
or   ( new_n33765_, new_n33764_, new_n33760_ );
and  ( new_n33766_, new_n33765_, new_n33759_ );
or   ( new_n33767_, new_n33766_, new_n33748_ );
and  ( new_n33768_, new_n33766_, new_n33748_ );
or   ( new_n33769_, new_n7184_, new_n22423_ );
or   ( new_n33770_, new_n7186_, new_n22304_ );
and  ( new_n33771_, new_n33770_, new_n33769_ );
xor  ( new_n33772_, new_n33771_, new_n6638_ );
or   ( new_n33773_, new_n6645_, new_n22641_ );
or   ( new_n33774_, new_n6647_, new_n22590_ );
and  ( new_n33775_, new_n33774_, new_n33773_ );
xor  ( new_n33776_, new_n33775_, new_n6166_ );
nor  ( new_n33777_, new_n33776_, new_n33772_ );
and  ( new_n33778_, new_n33776_, new_n33772_ );
or   ( new_n33779_, new_n6173_, new_n22975_ );
or   ( new_n33780_, new_n6175_, new_n22829_ );
and  ( new_n33781_, new_n33780_, new_n33779_ );
xor  ( new_n33782_, new_n33781_, new_n5597_ );
nor  ( new_n33783_, new_n33782_, new_n33778_ );
nor  ( new_n33784_, new_n33783_, new_n33777_ );
or   ( new_n33785_, new_n33784_, new_n33768_ );
and  ( new_n33786_, new_n33785_, new_n33767_ );
and  ( new_n33787_, new_n33731_, new_n33679_ );
or   ( new_n33788_, new_n33787_, new_n33786_ );
and  ( new_n33789_, new_n33788_, new_n33732_ );
or   ( new_n33790_, new_n33789_, new_n33627_ );
and  ( new_n33791_, new_n33789_, new_n33627_ );
xnor ( new_n33792_, new_n33121_, new_n33115_ );
xor  ( new_n33793_, new_n33792_, new_n33127_ );
xnor ( new_n33794_, new_n33155_, new_n33151_ );
xor  ( new_n33795_, new_n33794_, new_n33161_ );
nor  ( new_n33796_, new_n33795_, new_n33793_ );
nand ( new_n33797_, new_n33795_, new_n33793_ );
xor  ( new_n33798_, new_n33544_, new_n33542_ );
xnor ( new_n33799_, new_n33798_, new_n33548_ );
and  ( new_n33800_, new_n33799_, new_n33797_ );
or   ( new_n33801_, new_n33800_, new_n33796_ );
or   ( new_n33802_, new_n33801_, new_n33791_ );
and  ( new_n33803_, new_n33802_, new_n33790_ );
or   ( new_n33804_, new_n33803_, new_n33591_ );
nand ( new_n33805_, new_n33803_, new_n33591_ );
xnor ( new_n33806_, new_n33145_, new_n33129_ );
xor  ( new_n33807_, new_n33806_, new_n33163_ );
xor  ( new_n33808_, new_n33479_, new_n33463_ );
xor  ( new_n33809_, new_n33808_, new_n33497_ );
xor  ( new_n33810_, new_n33508_, new_n33506_ );
xor  ( new_n33811_, new_n33810_, new_n33512_ );
nand ( new_n33812_, new_n33811_, new_n33809_ );
nor  ( new_n33813_, new_n33811_, new_n33809_ );
xor  ( new_n33814_, new_n33532_, new_n33516_ );
xor  ( new_n33815_, new_n33814_, new_n33536_ );
or   ( new_n33816_, new_n33815_, new_n33813_ );
and  ( new_n33817_, new_n33816_, new_n33812_ );
nor  ( new_n33818_, new_n33817_, new_n33807_ );
and  ( new_n33819_, new_n33817_, new_n33807_ );
xor  ( new_n33820_, new_n33314_, new_n33312_ );
xnor ( new_n33821_, new_n33820_, new_n33318_ );
not  ( new_n33822_, new_n33821_ );
nor  ( new_n33823_, new_n33822_, new_n33819_ );
nor  ( new_n33824_, new_n33823_, new_n33818_ );
nand ( new_n33825_, new_n33824_, new_n33805_ );
and  ( new_n33826_, new_n33825_, new_n33804_ );
nor  ( new_n33827_, new_n33826_, new_n33581_ );
xor  ( new_n33828_, new_n33502_, new_n33344_ );
xor  ( new_n33829_, new_n33828_, new_n33553_ );
xnor ( new_n33830_, new_n33308_, new_n33306_ );
xor  ( new_n33831_, new_n33830_, new_n33320_ );
nor  ( new_n33832_, new_n33831_, new_n33829_ );
nand ( new_n33833_, new_n33831_, new_n33829_ );
xor  ( new_n33834_, new_n33326_, new_n33324_ );
xor  ( new_n33835_, new_n33834_, new_n33330_ );
and  ( new_n33836_, new_n33835_, new_n33833_ );
or   ( new_n33837_, new_n33836_, new_n33832_ );
nand ( new_n33838_, new_n33826_, new_n33581_ );
and  ( new_n33839_, new_n33838_, new_n33837_ );
or   ( new_n33840_, new_n33839_, new_n33827_ );
or   ( new_n33841_, new_n33840_, new_n33579_ );
and  ( new_n33842_, new_n33840_, new_n33579_ );
xor  ( new_n33843_, new_n33221_, new_n33059_ );
xor  ( new_n33844_, new_n33843_, new_n33271_ );
xnor ( new_n33845_, new_n33332_, new_n33322_ );
xor  ( new_n33846_, new_n33845_, new_n33555_ );
or   ( new_n33847_, new_n33846_, new_n33844_ );
and  ( new_n33848_, new_n33846_, new_n33844_ );
xor  ( new_n33849_, new_n33296_, new_n33294_ );
xor  ( new_n33850_, new_n33849_, new_n33300_ );
or   ( new_n33851_, new_n33850_, new_n33848_ );
and  ( new_n33852_, new_n33851_, new_n33847_ );
or   ( new_n33853_, new_n33852_, new_n33842_ );
and  ( new_n33854_, new_n33853_, new_n33841_ );
nor  ( new_n33855_, new_n33854_, new_n33577_ );
xor  ( new_n33856_, new_n33569_, new_n33290_ );
xor  ( new_n33857_, new_n33856_, new_n33572_ );
and  ( new_n33858_, new_n33857_, new_n33855_ );
xnor ( new_n33859_, new_n33854_, new_n33577_ );
xor  ( new_n33860_, new_n33852_, new_n33579_ );
xor  ( new_n33861_, new_n33860_, new_n33840_ );
xor  ( new_n33862_, new_n33831_, new_n33829_ );
xor  ( new_n33863_, new_n33862_, new_n33835_ );
xor  ( new_n33864_, new_n33789_, new_n33627_ );
xor  ( new_n33865_, new_n33864_, new_n33801_ );
xor  ( new_n33866_, new_n33585_, new_n33583_ );
xor  ( new_n33867_, new_n33866_, new_n33589_ );
nand ( new_n33868_, new_n33867_, new_n33865_ );
nor  ( new_n33869_, new_n33867_, new_n33865_ );
xor  ( new_n33870_, new_n33817_, new_n33807_ );
xor  ( new_n33871_, new_n33870_, new_n33822_ );
or   ( new_n33872_, new_n33871_, new_n33869_ );
and  ( new_n33873_, new_n33872_, new_n33868_ );
or   ( new_n33874_, new_n33873_, new_n33863_ );
and  ( new_n33875_, new_n33873_, new_n33863_ );
xnor ( new_n33876_, new_n33376_, new_n33360_ );
xor  ( new_n33877_, new_n33876_, new_n33394_ );
xnor ( new_n33878_, new_n33607_, new_n33605_ );
xor  ( new_n33879_, new_n33878_, new_n33611_ );
xor  ( new_n33880_, new_n33619_, new_n33617_ );
xor  ( new_n33881_, new_n33880_, new_n33623_ );
nand ( new_n33882_, new_n33881_, new_n33879_ );
nor  ( new_n33883_, new_n33881_, new_n33879_ );
xor  ( new_n33884_, new_n33597_, new_n33593_ );
xor  ( new_n33885_, new_n33884_, new_n33601_ );
or   ( new_n33886_, new_n33885_, new_n33883_ );
and  ( new_n33887_, new_n33886_, new_n33882_ );
or   ( new_n33888_, new_n33887_, new_n33877_ );
and  ( new_n33889_, new_n33887_, new_n33877_ );
xnor ( new_n33890_, new_n33659_, new_n33643_ );
xor  ( new_n33891_, new_n33890_, new_n33677_ );
xnor ( new_n33892_, new_n33711_, new_n33695_ );
xor  ( new_n33893_, new_n33892_, new_n33729_ );
or   ( new_n33894_, new_n33893_, new_n33891_ );
and  ( new_n33895_, new_n33893_, new_n33891_ );
xor  ( new_n33896_, new_n33766_, new_n33748_ );
xnor ( new_n33897_, new_n33896_, new_n33784_ );
or   ( new_n33898_, new_n33897_, new_n33895_ );
and  ( new_n33899_, new_n33898_, new_n33894_ );
or   ( new_n33900_, new_n33899_, new_n33889_ );
and  ( new_n33901_, new_n33900_, new_n33888_ );
xnor ( new_n33902_, new_n33442_, new_n33426_ );
xor  ( new_n33903_, new_n33902_, new_n33412_ );
xnor ( new_n33904_, new_n33795_, new_n33793_ );
xor  ( new_n33905_, new_n33904_, new_n33799_ );
or   ( new_n33906_, new_n33905_, new_n33903_ );
and  ( new_n33907_, new_n33905_, new_n33903_ );
xor  ( new_n33908_, new_n33811_, new_n33809_ );
xor  ( new_n33909_, new_n33908_, new_n33815_ );
or   ( new_n33910_, new_n33909_, new_n33907_ );
and  ( new_n33911_, new_n33910_, new_n33906_ );
nor  ( new_n33912_, new_n33911_, new_n33901_ );
and  ( new_n33913_, new_n33911_, new_n33901_ );
xor  ( new_n33914_, new_n33422_, new_n33416_ );
xor  ( new_n33915_, new_n33914_, new_n278_ );
xnor ( new_n33916_, new_n33758_, new_n33752_ );
xor  ( new_n33917_, new_n33916_, new_n33764_ );
xnor ( new_n33918_, new_n33740_, new_n33736_ );
xor  ( new_n33919_, new_n33918_, new_n33746_ );
or   ( new_n33920_, new_n33919_, new_n33917_ );
and  ( new_n33921_, new_n33919_, new_n33917_ );
xor  ( new_n33922_, new_n33776_, new_n33772_ );
xnor ( new_n33923_, new_n33922_, new_n33782_ );
or   ( new_n33924_, new_n33923_, new_n33921_ );
and  ( new_n33925_, new_n33924_, new_n33920_ );
nor  ( new_n33926_, new_n33925_, new_n33915_ );
and  ( new_n33927_, new_n33925_, new_n33915_ );
xor  ( new_n33928_, new_n33434_, new_n33430_ );
xnor ( new_n33929_, new_n33928_, new_n33440_ );
nor  ( new_n33930_, new_n33929_, new_n33927_ );
or   ( new_n33931_, new_n33930_, new_n33926_ );
or   ( new_n33932_, new_n6173_, new_n22973_ );
or   ( new_n33933_, new_n6175_, new_n22975_ );
and  ( new_n33934_, new_n33933_, new_n33932_ );
xor  ( new_n33935_, new_n33934_, new_n5597_ );
or   ( new_n33936_, new_n5604_, new_n23252_ );
or   ( new_n33937_, new_n5606_, new_n23166_ );
and  ( new_n33938_, new_n33937_, new_n33936_ );
xor  ( new_n33939_, new_n33938_, new_n5206_ );
or   ( new_n33940_, new_n33939_, new_n33935_ );
and  ( new_n33941_, new_n33939_, new_n33935_ );
or   ( new_n33942_, new_n5207_, new_n23554_ );
or   ( new_n33943_, new_n5209_, new_n23370_ );
and  ( new_n33944_, new_n33943_, new_n33942_ );
xor  ( new_n33945_, new_n33944_, new_n4708_ );
or   ( new_n33946_, new_n33945_, new_n33941_ );
and  ( new_n33947_, new_n33946_, new_n33940_ );
or   ( new_n33948_, new_n3461_, new_n24925_ );
or   ( new_n33949_, new_n3463_, new_n24927_ );
and  ( new_n33950_, new_n33949_, new_n33948_ );
xor  ( new_n33951_, new_n33950_, new_n3116_ );
or   ( new_n33952_, new_n3117_, new_n25288_ );
or   ( new_n33953_, new_n3119_, new_n25048_ );
and  ( new_n33954_, new_n33953_, new_n33952_ );
xor  ( new_n33955_, new_n33954_, new_n2800_ );
or   ( new_n33956_, new_n33955_, new_n33951_ );
and  ( new_n33957_, new_n33955_, new_n33951_ );
or   ( new_n33958_, new_n2807_, new_n25813_ );
or   ( new_n33959_, new_n2809_, new_n25486_ );
and  ( new_n33960_, new_n33959_, new_n33958_ );
xor  ( new_n33961_, new_n33960_, new_n2424_ );
or   ( new_n33962_, new_n33961_, new_n33957_ );
and  ( new_n33963_, new_n33962_, new_n33956_ );
or   ( new_n33964_, new_n33963_, new_n33947_ );
and  ( new_n33965_, new_n33963_, new_n33947_ );
or   ( new_n33966_, new_n4709_, new_n23895_ );
or   ( new_n33967_, new_n4711_, new_n23733_ );
and  ( new_n33968_, new_n33967_, new_n33966_ );
xor  ( new_n33969_, new_n33968_, new_n4295_ );
or   ( new_n33970_, new_n4302_, new_n24227_ );
or   ( new_n33971_, new_n4304_, new_n24006_ );
and  ( new_n33972_, new_n33971_, new_n33970_ );
xor  ( new_n33973_, new_n33972_, new_n3895_ );
nor  ( new_n33974_, new_n33973_, new_n33969_ );
and  ( new_n33975_, new_n33973_, new_n33969_ );
or   ( new_n33976_, new_n3896_, new_n24543_ );
or   ( new_n33977_, new_n3898_, new_n24418_ );
and  ( new_n33978_, new_n33977_, new_n33976_ );
xor  ( new_n33979_, new_n33978_, new_n3460_ );
nor  ( new_n33980_, new_n33979_, new_n33975_ );
nor  ( new_n33981_, new_n33980_, new_n33974_ );
or   ( new_n33982_, new_n33981_, new_n33965_ );
and  ( new_n33983_, new_n33982_, new_n33964_ );
or   ( new_n33984_, new_n9422_, new_n21842_ );
or   ( new_n33985_, new_n9424_, new_n21792_ );
and  ( new_n33986_, new_n33985_, new_n33984_ );
xor  ( new_n33987_, new_n33986_, new_n8873_ );
or   ( new_n33988_, new_n8874_, new_n21847_ );
or   ( new_n33989_, new_n8876_, new_n21840_ );
and  ( new_n33990_, new_n33989_, new_n33988_ );
xor  ( new_n33991_, new_n33990_, new_n8257_ );
or   ( new_n33992_, new_n33991_, new_n33987_ );
and  ( new_n33993_, new_n33991_, new_n33987_ );
or   ( new_n33994_, new_n8264_, new_n22129_ );
or   ( new_n33995_, new_n8266_, new_n22098_ );
and  ( new_n33996_, new_n33995_, new_n33994_ );
xor  ( new_n33997_, new_n33996_, new_n7725_ );
or   ( new_n33998_, new_n33997_, new_n33993_ );
and  ( new_n33999_, new_n33998_, new_n33992_ );
or   ( new_n34000_, new_n10059_, new_n21751_ );
or   ( new_n34001_, new_n10061_, new_n21685_ );
and  ( new_n34002_, new_n34001_, new_n34000_ );
xor  ( new_n34003_, new_n34002_, new_n9421_ );
and  ( new_n34004_, RIbb31938_136, RIbb2d888_64 );
or   ( new_n34005_, new_n21687_, RIbb2d888_64 );
and  ( new_n34006_, new_n34005_, RIbb2d900_63 );
or   ( new_n34007_, new_n34006_, new_n34004_ );
or   ( new_n34008_, new_n10770_, new_n21678_ );
and  ( new_n34009_, new_n34008_, new_n34007_ );
nor  ( new_n34010_, new_n34009_, new_n34003_ );
and  ( new_n34011_, new_n34009_, new_n34003_ );
nor  ( new_n34012_, new_n34011_, new_n311_ );
nor  ( new_n34013_, new_n34012_, new_n34010_ );
or   ( new_n34014_, new_n7732_, new_n22304_ );
or   ( new_n34015_, new_n7734_, new_n22207_ );
and  ( new_n34016_, new_n34015_, new_n34014_ );
xor  ( new_n34017_, new_n34016_, new_n7177_ );
or   ( new_n34018_, new_n7184_, new_n22590_ );
or   ( new_n34019_, new_n7186_, new_n22423_ );
and  ( new_n34020_, new_n34019_, new_n34018_ );
xor  ( new_n34021_, new_n34020_, new_n6638_ );
or   ( new_n34022_, new_n34021_, new_n34017_ );
and  ( new_n34023_, new_n34021_, new_n34017_ );
or   ( new_n34024_, new_n6645_, new_n22829_ );
or   ( new_n34025_, new_n6647_, new_n22641_ );
and  ( new_n34026_, new_n34025_, new_n34024_ );
xor  ( new_n34027_, new_n34026_, new_n6166_ );
or   ( new_n34028_, new_n34027_, new_n34023_ );
and  ( new_n34029_, new_n34028_, new_n34022_ );
and  ( new_n34030_, new_n34029_, new_n34013_ );
or   ( new_n34031_, new_n34030_, new_n33999_ );
or   ( new_n34032_, new_n34029_, new_n34013_ );
and  ( new_n34033_, new_n34032_, new_n34031_ );
or   ( new_n34034_, new_n34033_, new_n33983_ );
or   ( new_n34035_, new_n897_, new_n29261_ );
or   ( new_n34036_, new_n899_, new_n29263_ );
and  ( new_n34037_, new_n34036_, new_n34035_ );
xor  ( new_n34038_, new_n34037_, new_n748_ );
or   ( new_n34039_, new_n755_, new_n29619_ );
or   ( new_n34040_, new_n757_, new_n29474_ );
and  ( new_n34041_, new_n34040_, new_n34039_ );
xor  ( new_n34042_, new_n34041_, new_n523_ );
or   ( new_n34043_, new_n34042_, new_n34038_ );
and  ( new_n34044_, new_n34042_, new_n34038_ );
or   ( new_n34045_, new_n524_, new_n30227_ );
or   ( new_n34046_, new_n526_, new_n30120_ );
and  ( new_n34047_, new_n34046_, new_n34045_ );
xor  ( new_n34048_, new_n34047_, new_n403_ );
or   ( new_n34049_, new_n34048_, new_n34044_ );
and  ( new_n34050_, new_n34049_, new_n34043_ );
or   ( new_n34051_, new_n1593_, new_n27602_ );
or   ( new_n34052_, new_n1595_, new_n27396_ );
and  ( new_n34053_, new_n34052_, new_n34051_ );
xor  ( new_n34054_, new_n34053_, new_n1358_ );
or   ( new_n34055_, new_n1364_, new_n28108_ );
or   ( new_n34056_, new_n1366_, new_n27763_ );
and  ( new_n34057_, new_n34056_, new_n34055_ );
xor  ( new_n34058_, new_n34057_, new_n1129_ );
or   ( new_n34059_, new_n34058_, new_n34054_ );
and  ( new_n34060_, new_n34058_, new_n34054_ );
or   ( new_n34061_, new_n1135_, new_n28531_ );
or   ( new_n34062_, new_n1137_, new_n28314_ );
and  ( new_n34063_, new_n34062_, new_n34061_ );
xor  ( new_n34064_, new_n34063_, new_n896_ );
or   ( new_n34065_, new_n34064_, new_n34060_ );
and  ( new_n34066_, new_n34065_, new_n34059_ );
nor  ( new_n34067_, new_n34066_, new_n34050_ );
and  ( new_n34068_, new_n34066_, new_n34050_ );
or   ( new_n34069_, new_n2425_, new_n26063_ );
or   ( new_n34070_, new_n2427_, new_n26196_ );
and  ( new_n34071_, new_n34070_, new_n34069_ );
xor  ( new_n34072_, new_n34071_, new_n2121_ );
or   ( new_n34073_, new_n2122_, new_n26620_ );
or   ( new_n34074_, new_n2124_, new_n26372_ );
and  ( new_n34075_, new_n34074_, new_n34073_ );
xor  ( new_n34076_, new_n34075_, new_n1843_ );
nor  ( new_n34077_, new_n34076_, new_n34072_ );
and  ( new_n34078_, new_n34076_, new_n34072_ );
or   ( new_n34079_, new_n1844_, new_n27085_ );
or   ( new_n34080_, new_n1846_, new_n26762_ );
and  ( new_n34081_, new_n34080_, new_n34079_ );
xor  ( new_n34082_, new_n34081_, new_n1586_ );
nor  ( new_n34083_, new_n34082_, new_n34078_ );
nor  ( new_n34084_, new_n34083_, new_n34077_ );
nor  ( new_n34085_, new_n34084_, new_n34068_ );
nor  ( new_n34086_, new_n34085_, new_n34067_ );
and  ( new_n34087_, new_n34033_, new_n33983_ );
or   ( new_n34088_, new_n34087_, new_n34086_ );
and  ( new_n34089_, new_n34088_, new_n34034_ );
and  ( new_n34090_, new_n34089_, new_n33931_ );
nor  ( new_n34091_, new_n34089_, new_n33931_ );
xnor ( new_n34092_, new_n33703_, new_n33699_ );
xor  ( new_n34093_, new_n34092_, new_n33709_ );
xnor ( new_n34094_, new_n33687_, new_n33683_ );
xor  ( new_n34095_, new_n34094_, new_n33693_ );
or   ( new_n34096_, new_n34095_, new_n34093_ );
and  ( new_n34097_, new_n34095_, new_n34093_ );
xor  ( new_n34098_, new_n33721_, new_n33717_ );
xnor ( new_n34099_, new_n34098_, new_n33727_ );
or   ( new_n34100_, new_n34099_, new_n34097_ );
and  ( new_n34101_, new_n34100_, new_n34096_ );
xnor ( new_n34102_, new_n33651_, new_n33647_ );
xor  ( new_n34103_, new_n34102_, new_n33657_ );
xnor ( new_n34104_, new_n33635_, new_n33631_ );
xor  ( new_n34105_, new_n34104_, new_n33641_ );
or   ( new_n34106_, new_n34105_, new_n34103_ );
and  ( new_n34107_, new_n34105_, new_n34103_ );
xor  ( new_n34108_, new_n33669_, new_n33665_ );
xnor ( new_n34109_, new_n34108_, new_n33675_ );
or   ( new_n34110_, new_n34109_, new_n34107_ );
and  ( new_n34111_, new_n34110_, new_n34106_ );
nor  ( new_n34112_, new_n34111_, new_n34101_ );
and  ( new_n34113_, new_n34111_, new_n34101_ );
or   ( new_n34114_, new_n337_, new_n31333_ );
or   ( new_n34115_, new_n340_, new_n30798_ );
and  ( new_n34116_, new_n34115_, new_n34114_ );
xor  ( new_n34117_, new_n34116_, new_n332_ );
or   ( new_n34118_, new_n409_, new_n30798_ );
or   ( new_n34119_, new_n411_, new_n30800_ );
and  ( new_n34120_, new_n34119_, new_n34118_ );
xor  ( new_n34121_, new_n34120_, new_n328_ );
or   ( new_n34122_, new_n337_, new_n31654_ );
or   ( new_n34123_, new_n340_, new_n31333_ );
and  ( new_n34124_, new_n34123_, new_n34122_ );
xor  ( new_n34125_, new_n34124_, new_n332_ );
or   ( new_n34126_, new_n34125_, new_n34121_ );
and  ( new_n34127_, new_n34125_, new_n34121_ );
and  ( new_n34128_, new_n314_, RIbb33378_192 );
nor  ( new_n34129_, new_n34128_, new_n311_ );
and  ( new_n34130_, new_n34128_, RIbb2f340_7 );
nor  ( new_n34131_, new_n34130_, new_n34129_ );
or   ( new_n34132_, new_n34131_, new_n34127_ );
and  ( new_n34133_, new_n34132_, new_n34126_ );
and  ( new_n34134_, new_n34133_, new_n34117_ );
nor  ( new_n34135_, new_n34133_, new_n34117_ );
or   ( new_n34136_, new_n317_, new_n31952_ );
or   ( new_n34137_, new_n320_, new_n31654_ );
and  ( new_n34138_, new_n34137_, new_n34136_ );
xor  ( new_n34139_, new_n34138_, new_n312_ );
not  ( new_n34140_, new_n34139_ );
nor  ( new_n34141_, new_n34140_, new_n34135_ );
nor  ( new_n34142_, new_n34141_, new_n34134_ );
nor  ( new_n34143_, new_n34142_, new_n34113_ );
nor  ( new_n34144_, new_n34143_, new_n34112_ );
nor  ( new_n34145_, new_n34144_, new_n34091_ );
nor  ( new_n34146_, new_n34145_, new_n34090_ );
nor  ( new_n34147_, new_n34146_, new_n33913_ );
nor  ( new_n34148_, new_n34147_, new_n33912_ );
or   ( new_n34149_, new_n34148_, new_n33875_ );
and  ( new_n34150_, new_n34149_, new_n33874_ );
xor  ( new_n34151_, new_n33826_, new_n33581_ );
xor  ( new_n34152_, new_n34151_, new_n33837_ );
or   ( new_n34153_, new_n34152_, new_n34150_ );
and  ( new_n34154_, new_n34152_, new_n34150_ );
xor  ( new_n34155_, new_n33846_, new_n33844_ );
xor  ( new_n34156_, new_n34155_, new_n33850_ );
or   ( new_n34157_, new_n34156_, new_n34154_ );
and  ( new_n34158_, new_n34157_, new_n34153_ );
or   ( new_n34159_, new_n34158_, new_n33861_ );
and  ( new_n34160_, new_n34158_, new_n33861_ );
xor  ( new_n34161_, new_n33302_, new_n33292_ );
xor  ( new_n34162_, new_n34161_, new_n33558_ );
or   ( new_n34163_, new_n34162_, new_n34160_ );
and  ( new_n34164_, new_n34163_, new_n34159_ );
nor  ( new_n34165_, new_n34164_, new_n33859_ );
xor  ( new_n34166_, new_n34152_, new_n34150_ );
xor  ( new_n34167_, new_n34166_, new_n34156_ );
xor  ( new_n34168_, new_n33867_, new_n33865_ );
xor  ( new_n34169_, new_n34168_, new_n33871_ );
xor  ( new_n34170_, new_n33731_, new_n33679_ );
xor  ( new_n34171_, new_n34170_, new_n33786_ );
xor  ( new_n34172_, new_n33613_, new_n33603_ );
xor  ( new_n34173_, new_n34172_, new_n33625_ );
nand ( new_n34174_, new_n34173_, new_n34171_ );
nor  ( new_n34175_, new_n34173_, new_n34171_ );
xor  ( new_n34176_, new_n33905_, new_n33903_ );
xor  ( new_n34177_, new_n34176_, new_n33909_ );
or   ( new_n34178_, new_n34177_, new_n34175_ );
and  ( new_n34179_, new_n34178_, new_n34174_ );
or   ( new_n34180_, new_n34179_, new_n34169_ );
and  ( new_n34181_, new_n34179_, new_n34169_ );
xnor ( new_n34182_, new_n33881_, new_n33879_ );
xor  ( new_n34183_, new_n34182_, new_n33885_ );
xnor ( new_n34184_, new_n33893_, new_n33891_ );
xor  ( new_n34185_, new_n34184_, new_n33897_ );
nand ( new_n34186_, new_n34185_, new_n34183_ );
nor  ( new_n34187_, new_n34185_, new_n34183_ );
xor  ( new_n34188_, new_n34133_, new_n34117_ );
xor  ( new_n34189_, new_n34188_, new_n34140_ );
xnor ( new_n34190_, new_n33963_, new_n33947_ );
xor  ( new_n34191_, new_n34190_, new_n33981_ );
or   ( new_n34192_, new_n34191_, new_n34189_ );
and  ( new_n34193_, new_n34191_, new_n34189_ );
xnor ( new_n34194_, new_n34066_, new_n34050_ );
xor  ( new_n34195_, new_n34194_, new_n34084_ );
or   ( new_n34196_, new_n34195_, new_n34193_ );
and  ( new_n34197_, new_n34196_, new_n34192_ );
or   ( new_n34198_, new_n34197_, new_n34187_ );
and  ( new_n34199_, new_n34198_, new_n34186_ );
xor  ( new_n34200_, new_n34111_, new_n34101_ );
xor  ( new_n34201_, new_n34200_, new_n34142_ );
xnor ( new_n34202_, new_n34033_, new_n33983_ );
xor  ( new_n34203_, new_n34202_, new_n34086_ );
or   ( new_n34204_, new_n34203_, new_n34201_ );
and  ( new_n34205_, new_n34203_, new_n34201_ );
xor  ( new_n34206_, new_n33925_, new_n33915_ );
xor  ( new_n34207_, new_n34206_, new_n33929_ );
or   ( new_n34208_, new_n34207_, new_n34205_ );
and  ( new_n34209_, new_n34208_, new_n34204_ );
and  ( new_n34210_, new_n34209_, new_n34199_ );
nor  ( new_n34211_, new_n34209_, new_n34199_ );
xnor ( new_n34212_, new_n34095_, new_n34093_ );
xor  ( new_n34213_, new_n34212_, new_n34099_ );
xnor ( new_n34214_, new_n33919_, new_n33917_ );
xor  ( new_n34215_, new_n34214_, new_n33923_ );
or   ( new_n34216_, new_n34215_, new_n34213_ );
and  ( new_n34217_, new_n34215_, new_n34213_ );
xor  ( new_n34218_, new_n34105_, new_n34103_ );
xnor ( new_n34219_, new_n34218_, new_n34109_ );
or   ( new_n34220_, new_n34219_, new_n34217_ );
and  ( new_n34221_, new_n34220_, new_n34216_ );
or   ( new_n34222_, new_n3117_, new_n25486_ );
or   ( new_n34223_, new_n3119_, new_n25288_ );
and  ( new_n34224_, new_n34223_, new_n34222_ );
xor  ( new_n34225_, new_n34224_, new_n2800_ );
or   ( new_n34226_, new_n2807_, new_n26196_ );
or   ( new_n34227_, new_n2809_, new_n25813_ );
and  ( new_n34228_, new_n34227_, new_n34226_ );
xor  ( new_n34229_, new_n34228_, new_n2424_ );
or   ( new_n34230_, new_n34229_, new_n34225_ );
and  ( new_n34231_, new_n34229_, new_n34225_ );
or   ( new_n34232_, new_n2425_, new_n26372_ );
or   ( new_n34233_, new_n2427_, new_n26063_ );
and  ( new_n34234_, new_n34233_, new_n34232_ );
xor  ( new_n34235_, new_n34234_, new_n2121_ );
or   ( new_n34236_, new_n34235_, new_n34231_ );
and  ( new_n34237_, new_n34236_, new_n34230_ );
or   ( new_n34238_, new_n5604_, new_n23370_ );
or   ( new_n34239_, new_n5606_, new_n23252_ );
and  ( new_n34240_, new_n34239_, new_n34238_ );
xor  ( new_n34241_, new_n34240_, new_n5206_ );
or   ( new_n34242_, new_n5207_, new_n23733_ );
or   ( new_n34243_, new_n5209_, new_n23554_ );
and  ( new_n34244_, new_n34243_, new_n34242_ );
xor  ( new_n34245_, new_n34244_, new_n4708_ );
or   ( new_n34246_, new_n34245_, new_n34241_ );
and  ( new_n34247_, new_n34245_, new_n34241_ );
or   ( new_n34248_, new_n4709_, new_n24006_ );
or   ( new_n34249_, new_n4711_, new_n23895_ );
and  ( new_n34250_, new_n34249_, new_n34248_ );
xor  ( new_n34251_, new_n34250_, new_n4295_ );
or   ( new_n34252_, new_n34251_, new_n34247_ );
and  ( new_n34253_, new_n34252_, new_n34246_ );
or   ( new_n34254_, new_n34253_, new_n34237_ );
and  ( new_n34255_, new_n34253_, new_n34237_ );
or   ( new_n34256_, new_n4302_, new_n24418_ );
or   ( new_n34257_, new_n4304_, new_n24227_ );
and  ( new_n34258_, new_n34257_, new_n34256_ );
xor  ( new_n34259_, new_n34258_, new_n3895_ );
or   ( new_n34260_, new_n3896_, new_n24927_ );
or   ( new_n34261_, new_n3898_, new_n24543_ );
and  ( new_n34262_, new_n34261_, new_n34260_ );
xor  ( new_n34263_, new_n34262_, new_n3460_ );
nor  ( new_n34264_, new_n34263_, new_n34259_ );
and  ( new_n34265_, new_n34263_, new_n34259_ );
or   ( new_n34266_, new_n3461_, new_n25048_ );
or   ( new_n34267_, new_n3463_, new_n24925_ );
and  ( new_n34268_, new_n34267_, new_n34266_ );
xor  ( new_n34269_, new_n34268_, new_n3116_ );
nor  ( new_n34270_, new_n34269_, new_n34265_ );
nor  ( new_n34271_, new_n34270_, new_n34264_ );
or   ( new_n34272_, new_n34271_, new_n34255_ );
and  ( new_n34273_, new_n34272_, new_n34254_ );
or   ( new_n34274_, new_n1364_, new_n28314_ );
or   ( new_n34275_, new_n1366_, new_n28108_ );
and  ( new_n34276_, new_n34275_, new_n34274_ );
xor  ( new_n34277_, new_n34276_, new_n1129_ );
or   ( new_n34278_, new_n1135_, new_n29263_ );
or   ( new_n34279_, new_n1137_, new_n28531_ );
and  ( new_n34280_, new_n34279_, new_n34278_ );
xor  ( new_n34281_, new_n34280_, new_n896_ );
or   ( new_n34282_, new_n34281_, new_n34277_ );
and  ( new_n34283_, new_n34281_, new_n34277_ );
or   ( new_n34284_, new_n897_, new_n29474_ );
or   ( new_n34285_, new_n899_, new_n29261_ );
and  ( new_n34286_, new_n34285_, new_n34284_ );
xor  ( new_n34287_, new_n34286_, new_n748_ );
or   ( new_n34288_, new_n34287_, new_n34283_ );
and  ( new_n34289_, new_n34288_, new_n34282_ );
or   ( new_n34290_, new_n755_, new_n30120_ );
or   ( new_n34291_, new_n757_, new_n29619_ );
and  ( new_n34292_, new_n34291_, new_n34290_ );
xor  ( new_n34293_, new_n34292_, new_n523_ );
or   ( new_n34294_, new_n524_, new_n30800_ );
or   ( new_n34295_, new_n526_, new_n30227_ );
and  ( new_n34296_, new_n34295_, new_n34294_ );
xor  ( new_n34297_, new_n34296_, new_n403_ );
or   ( new_n34298_, new_n34297_, new_n34293_ );
and  ( new_n34299_, new_n34297_, new_n34293_ );
or   ( new_n34300_, new_n409_, new_n31333_ );
or   ( new_n34301_, new_n411_, new_n30798_ );
and  ( new_n34302_, new_n34301_, new_n34300_ );
xor  ( new_n34303_, new_n34302_, new_n328_ );
or   ( new_n34304_, new_n34303_, new_n34299_ );
and  ( new_n34305_, new_n34304_, new_n34298_ );
or   ( new_n34306_, new_n34305_, new_n34289_ );
and  ( new_n34307_, new_n34305_, new_n34289_ );
or   ( new_n34308_, new_n2122_, new_n26762_ );
or   ( new_n34309_, new_n2124_, new_n26620_ );
and  ( new_n34310_, new_n34309_, new_n34308_ );
xor  ( new_n34311_, new_n34310_, new_n1843_ );
or   ( new_n34312_, new_n1844_, new_n27396_ );
or   ( new_n34313_, new_n1846_, new_n27085_ );
and  ( new_n34314_, new_n34313_, new_n34312_ );
xor  ( new_n34315_, new_n34314_, new_n1586_ );
nor  ( new_n34316_, new_n34315_, new_n34311_ );
and  ( new_n34317_, new_n34315_, new_n34311_ );
or   ( new_n34318_, new_n1593_, new_n27763_ );
or   ( new_n34319_, new_n1595_, new_n27602_ );
and  ( new_n34320_, new_n34319_, new_n34318_ );
xor  ( new_n34321_, new_n34320_, new_n1358_ );
nor  ( new_n34322_, new_n34321_, new_n34317_ );
nor  ( new_n34323_, new_n34322_, new_n34316_ );
or   ( new_n34324_, new_n34323_, new_n34307_ );
and  ( new_n34325_, new_n34324_, new_n34306_ );
or   ( new_n34326_, new_n34325_, new_n34273_ );
or   ( new_n34327_, new_n10059_, new_n21792_ );
or   ( new_n34328_, new_n10061_, new_n21751_ );
and  ( new_n34329_, new_n34328_, new_n34327_ );
xor  ( new_n34330_, new_n34329_, new_n9421_ );
and  ( new_n34331_, RIbb319b0_137, RIbb2d888_64 );
or   ( new_n34332_, new_n21685_, RIbb2d888_64 );
and  ( new_n34333_, new_n34332_, RIbb2d900_63 );
or   ( new_n34334_, new_n34333_, new_n34331_ );
or   ( new_n34335_, new_n10770_, new_n21687_ );
and  ( new_n34336_, new_n34335_, new_n34334_ );
or   ( new_n34337_, new_n34336_, new_n34330_ );
and  ( new_n34338_, new_n34336_, new_n34330_ );
or   ( new_n34339_, new_n9422_, new_n21840_ );
or   ( new_n34340_, new_n9424_, new_n21842_ );
and  ( new_n34341_, new_n34340_, new_n34339_ );
xor  ( new_n34342_, new_n34341_, new_n8873_ );
or   ( new_n34343_, new_n34342_, new_n34338_ );
and  ( new_n34344_, new_n34343_, new_n34337_ );
or   ( new_n34345_, new_n7184_, new_n22641_ );
or   ( new_n34346_, new_n7186_, new_n22590_ );
and  ( new_n34347_, new_n34346_, new_n34345_ );
xor  ( new_n34348_, new_n34347_, new_n6638_ );
or   ( new_n34349_, new_n6645_, new_n22975_ );
or   ( new_n34350_, new_n6647_, new_n22829_ );
and  ( new_n34351_, new_n34350_, new_n34349_ );
xor  ( new_n34352_, new_n34351_, new_n6166_ );
or   ( new_n34353_, new_n34352_, new_n34348_ );
and  ( new_n34354_, new_n34352_, new_n34348_ );
or   ( new_n34355_, new_n6173_, new_n23166_ );
or   ( new_n34356_, new_n6175_, new_n22973_ );
and  ( new_n34357_, new_n34356_, new_n34355_ );
xor  ( new_n34358_, new_n34357_, new_n5597_ );
or   ( new_n34359_, new_n34358_, new_n34354_ );
and  ( new_n34360_, new_n34359_, new_n34353_ );
nor  ( new_n34361_, new_n34360_, new_n34344_ );
and  ( new_n34362_, new_n34360_, new_n34344_ );
or   ( new_n34363_, new_n8874_, new_n22098_ );
or   ( new_n34364_, new_n8876_, new_n21847_ );
and  ( new_n34365_, new_n34364_, new_n34363_ );
xor  ( new_n34366_, new_n34365_, new_n8257_ );
or   ( new_n34367_, new_n8264_, new_n22207_ );
or   ( new_n34368_, new_n8266_, new_n22129_ );
and  ( new_n34369_, new_n34368_, new_n34367_ );
xor  ( new_n34370_, new_n34369_, new_n7725_ );
nor  ( new_n34371_, new_n34370_, new_n34366_ );
and  ( new_n34372_, new_n34370_, new_n34366_ );
or   ( new_n34373_, new_n7732_, new_n22423_ );
or   ( new_n34374_, new_n7734_, new_n22304_ );
and  ( new_n34375_, new_n34374_, new_n34373_ );
xor  ( new_n34376_, new_n34375_, new_n7177_ );
nor  ( new_n34377_, new_n34376_, new_n34372_ );
nor  ( new_n34378_, new_n34377_, new_n34371_ );
nor  ( new_n34379_, new_n34378_, new_n34362_ );
nor  ( new_n34380_, new_n34379_, new_n34361_ );
and  ( new_n34381_, new_n34325_, new_n34273_ );
or   ( new_n34382_, new_n34381_, new_n34380_ );
and  ( new_n34383_, new_n34382_, new_n34326_ );
nor  ( new_n34384_, new_n34383_, new_n34221_ );
and  ( new_n34385_, new_n34383_, new_n34221_ );
not  ( new_n34386_, new_n34385_ );
xnor ( new_n34387_, new_n33955_, new_n33951_ );
xor  ( new_n34388_, new_n34387_, new_n33961_ );
xnor ( new_n34389_, new_n33973_, new_n33969_ );
xor  ( new_n34390_, new_n34389_, new_n33979_ );
or   ( new_n34391_, new_n34390_, new_n34388_ );
and  ( new_n34392_, new_n34390_, new_n34388_ );
xor  ( new_n34393_, new_n34076_, new_n34072_ );
xnor ( new_n34394_, new_n34393_, new_n34082_ );
or   ( new_n34395_, new_n34394_, new_n34392_ );
and  ( new_n34396_, new_n34395_, new_n34391_ );
xnor ( new_n34397_, new_n34058_, new_n34054_ );
xor  ( new_n34398_, new_n34397_, new_n34064_ );
xnor ( new_n34399_, new_n34125_, new_n34121_ );
xor  ( new_n34400_, new_n34399_, new_n34131_ );
or   ( new_n34401_, new_n34400_, new_n34398_ );
and  ( new_n34402_, new_n34400_, new_n34398_ );
xor  ( new_n34403_, new_n34042_, new_n34038_ );
xnor ( new_n34404_, new_n34403_, new_n34048_ );
or   ( new_n34405_, new_n34404_, new_n34402_ );
and  ( new_n34406_, new_n34405_, new_n34401_ );
nor  ( new_n34407_, new_n34406_, new_n34396_ );
and  ( new_n34408_, new_n34406_, new_n34396_ );
xnor ( new_n34409_, new_n33991_, new_n33987_ );
xor  ( new_n34410_, new_n34409_, new_n33997_ );
xnor ( new_n34411_, new_n34021_, new_n34017_ );
xor  ( new_n34412_, new_n34411_, new_n34027_ );
nor  ( new_n34413_, new_n34412_, new_n34410_ );
and  ( new_n34414_, new_n34412_, new_n34410_ );
xor  ( new_n34415_, new_n33939_, new_n33935_ );
xnor ( new_n34416_, new_n34415_, new_n33945_ );
nor  ( new_n34417_, new_n34416_, new_n34414_ );
nor  ( new_n34418_, new_n34417_, new_n34413_ );
nor  ( new_n34419_, new_n34418_, new_n34408_ );
nor  ( new_n34420_, new_n34419_, new_n34407_ );
and  ( new_n34421_, new_n34420_, new_n34386_ );
nor  ( new_n34422_, new_n34421_, new_n34384_ );
nor  ( new_n34423_, new_n34422_, new_n34211_ );
nor  ( new_n34424_, new_n34423_, new_n34210_ );
not  ( new_n34425_, new_n34424_ );
or   ( new_n34426_, new_n34425_, new_n34181_ );
and  ( new_n34427_, new_n34426_, new_n34180_ );
xor  ( new_n34428_, new_n33803_, new_n33591_ );
xor  ( new_n34429_, new_n34428_, new_n33824_ );
or   ( new_n34430_, new_n34429_, new_n34427_ );
and  ( new_n34431_, new_n34429_, new_n34427_ );
xor  ( new_n34432_, new_n33873_, new_n33863_ );
xor  ( new_n34433_, new_n34432_, new_n34148_ );
or   ( new_n34434_, new_n34433_, new_n34431_ );
and  ( new_n34435_, new_n34434_, new_n34430_ );
nor  ( new_n34436_, new_n34435_, new_n34167_ );
xnor ( new_n34437_, new_n34158_, new_n33861_ );
xor  ( new_n34438_, new_n34437_, new_n34162_ );
and  ( new_n34439_, new_n34438_, new_n34436_ );
xor  ( new_n34440_, new_n33911_, new_n33901_ );
xor  ( new_n34441_, new_n34440_, new_n34146_ );
xor  ( new_n34442_, new_n34089_, new_n33931_ );
xor  ( new_n34443_, new_n34442_, new_n34144_ );
xnor ( new_n34444_, new_n34209_, new_n34199_ );
xor  ( new_n34445_, new_n34444_, new_n34422_ );
or   ( new_n34446_, new_n34445_, new_n34443_ );
and  ( new_n34447_, new_n34445_, new_n34443_ );
xor  ( new_n34448_, new_n34173_, new_n34171_ );
xor  ( new_n34449_, new_n34448_, new_n34177_ );
or   ( new_n34450_, new_n34449_, new_n34447_ );
and  ( new_n34451_, new_n34450_, new_n34446_ );
nor  ( new_n34452_, new_n34451_, new_n34441_ );
and  ( new_n34453_, new_n34451_, new_n34441_ );
xor  ( new_n34454_, new_n33887_, new_n33877_ );
xor  ( new_n34455_, new_n34454_, new_n33899_ );
xor  ( new_n34456_, new_n34383_, new_n34221_ );
xor  ( new_n34457_, new_n34456_, new_n34420_ );
xor  ( new_n34458_, new_n34203_, new_n34201_ );
xor  ( new_n34459_, new_n34458_, new_n34207_ );
or   ( new_n34460_, new_n34459_, new_n34457_ );
and  ( new_n34461_, new_n34459_, new_n34457_ );
xor  ( new_n34462_, new_n34185_, new_n34183_ );
xor  ( new_n34463_, new_n34462_, new_n34197_ );
or   ( new_n34464_, new_n34463_, new_n34461_ );
and  ( new_n34465_, new_n34464_, new_n34460_ );
nor  ( new_n34466_, new_n34465_, new_n34455_ );
and  ( new_n34467_, new_n34465_, new_n34455_ );
xnor ( new_n34468_, new_n34029_, new_n34013_ );
xor  ( new_n34469_, new_n34468_, new_n33999_ );
xnor ( new_n34470_, new_n34253_, new_n34237_ );
xor  ( new_n34471_, new_n34470_, new_n34271_ );
xnor ( new_n34472_, new_n34305_, new_n34289_ );
xor  ( new_n34473_, new_n34472_, new_n34323_ );
or   ( new_n34474_, new_n34473_, new_n34471_ );
and  ( new_n34475_, new_n34473_, new_n34471_ );
xor  ( new_n34476_, new_n34400_, new_n34398_ );
xnor ( new_n34477_, new_n34476_, new_n34404_ );
not  ( new_n34478_, new_n34477_ );
or   ( new_n34479_, new_n34478_, new_n34475_ );
and  ( new_n34480_, new_n34479_, new_n34474_ );
or   ( new_n34481_, new_n34480_, new_n34469_ );
and  ( new_n34482_, new_n34480_, new_n34469_ );
xor  ( new_n34483_, new_n34191_, new_n34189_ );
xor  ( new_n34484_, new_n34483_, new_n34195_ );
or   ( new_n34485_, new_n34484_, new_n34482_ );
and  ( new_n34486_, new_n34485_, new_n34481_ );
xor  ( new_n34487_, new_n34406_, new_n34396_ );
xor  ( new_n34488_, new_n34487_, new_n34418_ );
xnor ( new_n34489_, new_n34325_, new_n34273_ );
xor  ( new_n34490_, new_n34489_, new_n34380_ );
or   ( new_n34491_, new_n34490_, new_n34488_ );
and  ( new_n34492_, new_n34490_, new_n34488_ );
xnor ( new_n34493_, new_n34215_, new_n34213_ );
xor  ( new_n34494_, new_n34493_, new_n34219_ );
or   ( new_n34495_, new_n34494_, new_n34492_ );
and  ( new_n34496_, new_n34495_, new_n34491_ );
nor  ( new_n34497_, new_n34496_, new_n34486_ );
and  ( new_n34498_, new_n34496_, new_n34486_ );
xor  ( new_n34499_, new_n34009_, new_n34003_ );
xor  ( new_n34500_, new_n34499_, new_n311_ );
xnor ( new_n34501_, new_n34412_, new_n34410_ );
xor  ( new_n34502_, new_n34501_, new_n34416_ );
and  ( new_n34503_, new_n34502_, new_n34500_ );
or   ( new_n34504_, new_n34502_, new_n34500_ );
xor  ( new_n34505_, new_n34390_, new_n34388_ );
xnor ( new_n34506_, new_n34505_, new_n34394_ );
and  ( new_n34507_, new_n34506_, new_n34504_ );
or   ( new_n34508_, new_n34507_, new_n34503_ );
or   ( new_n34509_, new_n2425_, new_n26620_ );
or   ( new_n34510_, new_n2427_, new_n26372_ );
and  ( new_n34511_, new_n34510_, new_n34509_ );
xor  ( new_n34512_, new_n34511_, new_n2121_ );
or   ( new_n34513_, new_n2122_, new_n27085_ );
or   ( new_n34514_, new_n2124_, new_n26762_ );
and  ( new_n34515_, new_n34514_, new_n34513_ );
xor  ( new_n34516_, new_n34515_, new_n1843_ );
or   ( new_n34517_, new_n34516_, new_n34512_ );
and  ( new_n34518_, new_n34516_, new_n34512_ );
or   ( new_n34519_, new_n1844_, new_n27602_ );
or   ( new_n34520_, new_n1846_, new_n27396_ );
and  ( new_n34521_, new_n34520_, new_n34519_ );
xor  ( new_n34522_, new_n34521_, new_n1586_ );
or   ( new_n34523_, new_n34522_, new_n34518_ );
and  ( new_n34524_, new_n34523_, new_n34517_ );
or   ( new_n34525_, new_n897_, new_n29619_ );
or   ( new_n34526_, new_n899_, new_n29474_ );
and  ( new_n34527_, new_n34526_, new_n34525_ );
xor  ( new_n34528_, new_n34527_, new_n748_ );
or   ( new_n34529_, new_n755_, new_n30227_ );
or   ( new_n34530_, new_n757_, new_n30120_ );
and  ( new_n34531_, new_n34530_, new_n34529_ );
xor  ( new_n34532_, new_n34531_, new_n523_ );
or   ( new_n34533_, new_n34532_, new_n34528_ );
and  ( new_n34534_, new_n34532_, new_n34528_ );
or   ( new_n34535_, new_n524_, new_n30798_ );
or   ( new_n34536_, new_n526_, new_n30800_ );
and  ( new_n34537_, new_n34536_, new_n34535_ );
xor  ( new_n34538_, new_n34537_, new_n403_ );
or   ( new_n34539_, new_n34538_, new_n34534_ );
and  ( new_n34540_, new_n34539_, new_n34533_ );
or   ( new_n34541_, new_n34540_, new_n34524_ );
and  ( new_n34542_, new_n34540_, new_n34524_ );
or   ( new_n34543_, new_n1593_, new_n28108_ );
or   ( new_n34544_, new_n1595_, new_n27763_ );
and  ( new_n34545_, new_n34544_, new_n34543_ );
xor  ( new_n34546_, new_n34545_, new_n1358_ );
or   ( new_n34547_, new_n1364_, new_n28531_ );
or   ( new_n34548_, new_n1366_, new_n28314_ );
and  ( new_n34549_, new_n34548_, new_n34547_ );
xor  ( new_n34550_, new_n34549_, new_n1129_ );
nor  ( new_n34551_, new_n34550_, new_n34546_ );
and  ( new_n34552_, new_n34550_, new_n34546_ );
or   ( new_n34553_, new_n1135_, new_n29261_ );
or   ( new_n34554_, new_n1137_, new_n29263_ );
and  ( new_n34555_, new_n34554_, new_n34553_ );
xor  ( new_n34556_, new_n34555_, new_n896_ );
nor  ( new_n34557_, new_n34556_, new_n34552_ );
nor  ( new_n34558_, new_n34557_, new_n34551_ );
or   ( new_n34559_, new_n34558_, new_n34542_ );
and  ( new_n34560_, new_n34559_, new_n34541_ );
or   ( new_n34561_, new_n7732_, new_n22590_ );
or   ( new_n34562_, new_n7734_, new_n22423_ );
and  ( new_n34563_, new_n34562_, new_n34561_ );
xor  ( new_n34564_, new_n34563_, new_n7177_ );
or   ( new_n34565_, new_n7184_, new_n22829_ );
or   ( new_n34566_, new_n7186_, new_n22641_ );
and  ( new_n34567_, new_n34566_, new_n34565_ );
xor  ( new_n34568_, new_n34567_, new_n6638_ );
or   ( new_n34569_, new_n34568_, new_n34564_ );
and  ( new_n34570_, new_n34568_, new_n34564_ );
or   ( new_n34571_, new_n6645_, new_n22973_ );
or   ( new_n34572_, new_n6647_, new_n22975_ );
and  ( new_n34573_, new_n34572_, new_n34571_ );
xor  ( new_n34574_, new_n34573_, new_n6166_ );
or   ( new_n34575_, new_n34574_, new_n34570_ );
and  ( new_n34576_, new_n34575_, new_n34569_ );
or   ( new_n34577_, new_n10059_, new_n21842_ );
or   ( new_n34578_, new_n10061_, new_n21792_ );
and  ( new_n34579_, new_n34578_, new_n34577_ );
xor  ( new_n34580_, new_n34579_, new_n9421_ );
and  ( new_n34581_, RIbb31a28_138, RIbb2d888_64 );
or   ( new_n34582_, new_n21751_, RIbb2d888_64 );
and  ( new_n34583_, new_n34582_, RIbb2d900_63 );
or   ( new_n34584_, new_n34583_, new_n34581_ );
or   ( new_n34585_, new_n10770_, new_n21685_ );
and  ( new_n34586_, new_n34585_, new_n34584_ );
nor  ( new_n34587_, new_n34586_, new_n34580_ );
and  ( new_n34588_, new_n34586_, new_n34580_ );
nor  ( new_n34589_, new_n34588_, new_n331_ );
nor  ( new_n34590_, new_n34589_, new_n34587_ );
or   ( new_n34591_, new_n9422_, new_n21847_ );
or   ( new_n34592_, new_n9424_, new_n21840_ );
and  ( new_n34593_, new_n34592_, new_n34591_ );
xor  ( new_n34594_, new_n34593_, new_n8873_ );
or   ( new_n34595_, new_n8874_, new_n22129_ );
or   ( new_n34596_, new_n8876_, new_n22098_ );
and  ( new_n34597_, new_n34596_, new_n34595_ );
xor  ( new_n34598_, new_n34597_, new_n8257_ );
or   ( new_n34599_, new_n34598_, new_n34594_ );
and  ( new_n34600_, new_n34598_, new_n34594_ );
or   ( new_n34601_, new_n8264_, new_n22304_ );
or   ( new_n34602_, new_n8266_, new_n22207_ );
and  ( new_n34603_, new_n34602_, new_n34601_ );
xor  ( new_n34604_, new_n34603_, new_n7725_ );
or   ( new_n34605_, new_n34604_, new_n34600_ );
and  ( new_n34606_, new_n34605_, new_n34599_ );
and  ( new_n34607_, new_n34606_, new_n34590_ );
or   ( new_n34608_, new_n34607_, new_n34576_ );
or   ( new_n34609_, new_n34606_, new_n34590_ );
and  ( new_n34610_, new_n34609_, new_n34608_ );
or   ( new_n34611_, new_n34610_, new_n34560_ );
or   ( new_n34612_, new_n4709_, new_n24227_ );
or   ( new_n34613_, new_n4711_, new_n24006_ );
and  ( new_n34614_, new_n34613_, new_n34612_ );
xor  ( new_n34615_, new_n34614_, new_n4295_ );
or   ( new_n34616_, new_n4302_, new_n24543_ );
or   ( new_n34617_, new_n4304_, new_n24418_ );
and  ( new_n34618_, new_n34617_, new_n34616_ );
xor  ( new_n34619_, new_n34618_, new_n3895_ );
or   ( new_n34620_, new_n34619_, new_n34615_ );
and  ( new_n34621_, new_n34619_, new_n34615_ );
or   ( new_n34622_, new_n3896_, new_n24925_ );
or   ( new_n34623_, new_n3898_, new_n24927_ );
and  ( new_n34624_, new_n34623_, new_n34622_ );
xor  ( new_n34625_, new_n34624_, new_n3460_ );
or   ( new_n34626_, new_n34625_, new_n34621_ );
and  ( new_n34627_, new_n34626_, new_n34620_ );
or   ( new_n34628_, new_n3461_, new_n25288_ );
or   ( new_n34629_, new_n3463_, new_n25048_ );
and  ( new_n34630_, new_n34629_, new_n34628_ );
xor  ( new_n34631_, new_n34630_, new_n3116_ );
or   ( new_n34632_, new_n3117_, new_n25813_ );
or   ( new_n34633_, new_n3119_, new_n25486_ );
and  ( new_n34634_, new_n34633_, new_n34632_ );
xor  ( new_n34635_, new_n34634_, new_n2800_ );
or   ( new_n34636_, new_n34635_, new_n34631_ );
and  ( new_n34637_, new_n34635_, new_n34631_ );
or   ( new_n34638_, new_n2807_, new_n26063_ );
or   ( new_n34639_, new_n2809_, new_n26196_ );
and  ( new_n34640_, new_n34639_, new_n34638_ );
xor  ( new_n34641_, new_n34640_, new_n2424_ );
or   ( new_n34642_, new_n34641_, new_n34637_ );
and  ( new_n34643_, new_n34642_, new_n34636_ );
or   ( new_n34644_, new_n34643_, new_n34627_ );
and  ( new_n34645_, new_n34643_, new_n34627_ );
or   ( new_n34646_, new_n6173_, new_n23252_ );
or   ( new_n34647_, new_n6175_, new_n23166_ );
and  ( new_n34648_, new_n34647_, new_n34646_ );
xor  ( new_n34649_, new_n34648_, new_n5597_ );
or   ( new_n34650_, new_n5604_, new_n23554_ );
or   ( new_n34651_, new_n5606_, new_n23370_ );
and  ( new_n34652_, new_n34651_, new_n34650_ );
xor  ( new_n34653_, new_n34652_, new_n5206_ );
nor  ( new_n34654_, new_n34653_, new_n34649_ );
and  ( new_n34655_, new_n34653_, new_n34649_ );
or   ( new_n34656_, new_n5207_, new_n23895_ );
or   ( new_n34657_, new_n5209_, new_n23733_ );
and  ( new_n34658_, new_n34657_, new_n34656_ );
xor  ( new_n34659_, new_n34658_, new_n4708_ );
nor  ( new_n34660_, new_n34659_, new_n34655_ );
nor  ( new_n34661_, new_n34660_, new_n34654_ );
or   ( new_n34662_, new_n34661_, new_n34645_ );
and  ( new_n34663_, new_n34662_, new_n34644_ );
and  ( new_n34664_, new_n34610_, new_n34560_ );
or   ( new_n34665_, new_n34664_, new_n34663_ );
and  ( new_n34666_, new_n34665_, new_n34611_ );
and  ( new_n34667_, new_n34666_, new_n34508_ );
nor  ( new_n34668_, new_n34666_, new_n34508_ );
or   ( new_n34669_, new_n337_, new_n31952_ );
or   ( new_n34670_, new_n340_, new_n31654_ );
and  ( new_n34671_, new_n34670_, new_n34669_ );
xor  ( new_n34672_, new_n34671_, new_n331_ );
xnor ( new_n34673_, new_n34297_, new_n34293_ );
xor  ( new_n34674_, new_n34673_, new_n34303_ );
and  ( new_n34675_, new_n34674_, new_n34672_ );
or   ( new_n34676_, new_n34674_, new_n34672_ );
xor  ( new_n34677_, new_n34281_, new_n34277_ );
xnor ( new_n34678_, new_n34677_, new_n34287_ );
and  ( new_n34679_, new_n34678_, new_n34676_ );
or   ( new_n34680_, new_n34679_, new_n34675_ );
xnor ( new_n34681_, new_n34229_, new_n34225_ );
xor  ( new_n34682_, new_n34681_, new_n34235_ );
xnor ( new_n34683_, new_n34263_, new_n34259_ );
xor  ( new_n34684_, new_n34683_, new_n34269_ );
or   ( new_n34685_, new_n34684_, new_n34682_ );
and  ( new_n34686_, new_n34684_, new_n34682_ );
xor  ( new_n34687_, new_n34315_, new_n34311_ );
xnor ( new_n34688_, new_n34687_, new_n34321_ );
or   ( new_n34689_, new_n34688_, new_n34686_ );
and  ( new_n34690_, new_n34689_, new_n34685_ );
nor  ( new_n34691_, new_n34690_, new_n34680_ );
and  ( new_n34692_, new_n34690_, new_n34680_ );
xnor ( new_n34693_, new_n34245_, new_n34241_ );
xor  ( new_n34694_, new_n34693_, new_n34251_ );
xnor ( new_n34695_, new_n34352_, new_n34348_ );
xor  ( new_n34696_, new_n34695_, new_n34358_ );
nor  ( new_n34697_, new_n34696_, new_n34694_ );
and  ( new_n34698_, new_n34696_, new_n34694_ );
xor  ( new_n34699_, new_n34370_, new_n34366_ );
xnor ( new_n34700_, new_n34699_, new_n34376_ );
nor  ( new_n34701_, new_n34700_, new_n34698_ );
nor  ( new_n34702_, new_n34701_, new_n34697_ );
nor  ( new_n34703_, new_n34702_, new_n34692_ );
nor  ( new_n34704_, new_n34703_, new_n34691_ );
nor  ( new_n34705_, new_n34704_, new_n34668_ );
nor  ( new_n34706_, new_n34705_, new_n34667_ );
nor  ( new_n34707_, new_n34706_, new_n34498_ );
nor  ( new_n34708_, new_n34707_, new_n34497_ );
nor  ( new_n34709_, new_n34708_, new_n34467_ );
nor  ( new_n34710_, new_n34709_, new_n34466_ );
nor  ( new_n34711_, new_n34710_, new_n34453_ );
nor  ( new_n34712_, new_n34711_, new_n34452_ );
xnor ( new_n34713_, new_n34429_, new_n34427_ );
xnor ( new_n34714_, new_n34713_, new_n34433_ );
nor  ( new_n34715_, new_n34714_, new_n34712_ );
xor  ( new_n34716_, new_n34435_, new_n34167_ );
and  ( new_n34717_, new_n34716_, new_n34715_ );
xnor ( new_n34718_, new_n34714_, new_n34712_ );
xor  ( new_n34719_, new_n34451_, new_n34441_ );
xor  ( new_n34720_, new_n34719_, new_n34710_ );
xor  ( new_n34721_, new_n34459_, new_n34457_ );
xor  ( new_n34722_, new_n34721_, new_n34463_ );
xor  ( new_n34723_, new_n34666_, new_n34508_ );
xor  ( new_n34724_, new_n34723_, new_n34704_ );
xor  ( new_n34725_, new_n34480_, new_n34469_ );
xor  ( new_n34726_, new_n34725_, new_n34484_ );
or   ( new_n34727_, new_n34726_, new_n34724_ );
and  ( new_n34728_, new_n34726_, new_n34724_ );
xor  ( new_n34729_, new_n34490_, new_n34488_ );
xor  ( new_n34730_, new_n34729_, new_n34494_ );
or   ( new_n34731_, new_n34730_, new_n34728_ );
and  ( new_n34732_, new_n34731_, new_n34727_ );
or   ( new_n34733_, new_n34732_, new_n34722_ );
and  ( new_n34734_, new_n34732_, new_n34722_ );
xnor ( new_n34735_, new_n34360_, new_n34344_ );
xor  ( new_n34736_, new_n34735_, new_n34378_ );
xnor ( new_n34737_, new_n34540_, new_n34524_ );
xor  ( new_n34738_, new_n34737_, new_n34558_ );
xnor ( new_n34739_, new_n34643_, new_n34627_ );
xor  ( new_n34740_, new_n34739_, new_n34661_ );
or   ( new_n34741_, new_n34740_, new_n34738_ );
and  ( new_n34742_, new_n34740_, new_n34738_ );
xor  ( new_n34743_, new_n34674_, new_n34672_ );
xor  ( new_n34744_, new_n34743_, new_n34678_ );
or   ( new_n34745_, new_n34744_, new_n34742_ );
and  ( new_n34746_, new_n34745_, new_n34741_ );
or   ( new_n34747_, new_n34746_, new_n34736_ );
and  ( new_n34748_, new_n34746_, new_n34736_ );
xor  ( new_n34749_, new_n34473_, new_n34471_ );
xor  ( new_n34750_, new_n34749_, new_n34478_ );
or   ( new_n34751_, new_n34750_, new_n34748_ );
and  ( new_n34752_, new_n34751_, new_n34747_ );
xor  ( new_n34753_, new_n34610_, new_n34560_ );
xor  ( new_n34754_, new_n34753_, new_n34663_ );
xnor ( new_n34755_, new_n34690_, new_n34680_ );
xor  ( new_n34756_, new_n34755_, new_n34702_ );
nand ( new_n34757_, new_n34756_, new_n34754_ );
nor  ( new_n34758_, new_n34756_, new_n34754_ );
xnor ( new_n34759_, new_n34502_, new_n34500_ );
xor  ( new_n34760_, new_n34759_, new_n34506_ );
or   ( new_n34761_, new_n34760_, new_n34758_ );
and  ( new_n34762_, new_n34761_, new_n34757_ );
or   ( new_n34763_, new_n34762_, new_n34752_ );
and  ( new_n34764_, new_n34762_, new_n34752_ );
xor  ( new_n34765_, new_n34336_, new_n34330_ );
xor  ( new_n34766_, new_n34765_, new_n34342_ );
xnor ( new_n34767_, new_n34684_, new_n34682_ );
xor  ( new_n34768_, new_n34767_, new_n34688_ );
and  ( new_n34769_, new_n34768_, new_n34766_ );
or   ( new_n34770_, new_n34768_, new_n34766_ );
xor  ( new_n34771_, new_n34696_, new_n34694_ );
xnor ( new_n34772_, new_n34771_, new_n34700_ );
and  ( new_n34773_, new_n34772_, new_n34770_ );
or   ( new_n34774_, new_n34773_, new_n34769_ );
or   ( new_n34775_, new_n2122_, new_n27396_ );
or   ( new_n34776_, new_n2124_, new_n27085_ );
and  ( new_n34777_, new_n34776_, new_n34775_ );
xor  ( new_n34778_, new_n34777_, new_n1843_ );
or   ( new_n34779_, new_n1844_, new_n27763_ );
or   ( new_n34780_, new_n1846_, new_n27602_ );
and  ( new_n34781_, new_n34780_, new_n34779_ );
xor  ( new_n34782_, new_n34781_, new_n1586_ );
or   ( new_n34783_, new_n34782_, new_n34778_ );
and  ( new_n34784_, new_n34782_, new_n34778_ );
or   ( new_n34785_, new_n1593_, new_n28314_ );
or   ( new_n34786_, new_n1595_, new_n28108_ );
and  ( new_n34787_, new_n34786_, new_n34785_ );
xor  ( new_n34788_, new_n34787_, new_n1358_ );
or   ( new_n34789_, new_n34788_, new_n34784_ );
and  ( new_n34790_, new_n34789_, new_n34783_ );
or   ( new_n34791_, new_n755_, new_n30800_ );
or   ( new_n34792_, new_n757_, new_n30227_ );
and  ( new_n34793_, new_n34792_, new_n34791_ );
xor  ( new_n34794_, new_n34793_, new_n523_ );
or   ( new_n34795_, new_n524_, new_n31333_ );
or   ( new_n34796_, new_n526_, new_n30798_ );
and  ( new_n34797_, new_n34796_, new_n34795_ );
xor  ( new_n34798_, new_n34797_, new_n403_ );
or   ( new_n34799_, new_n34798_, new_n34794_ );
and  ( new_n34800_, new_n34798_, new_n34794_ );
or   ( new_n34801_, new_n409_, new_n31952_ );
or   ( new_n34802_, new_n411_, new_n31654_ );
and  ( new_n34803_, new_n34802_, new_n34801_ );
xor  ( new_n34804_, new_n34803_, new_n328_ );
or   ( new_n34805_, new_n34804_, new_n34800_ );
and  ( new_n34806_, new_n34805_, new_n34799_ );
or   ( new_n34807_, new_n34806_, new_n34790_ );
and  ( new_n34808_, new_n34806_, new_n34790_ );
or   ( new_n34809_, new_n1364_, new_n29263_ );
or   ( new_n34810_, new_n1366_, new_n28531_ );
and  ( new_n34811_, new_n34810_, new_n34809_ );
xor  ( new_n34812_, new_n34811_, new_n1129_ );
or   ( new_n34813_, new_n1135_, new_n29474_ );
or   ( new_n34814_, new_n1137_, new_n29261_ );
and  ( new_n34815_, new_n34814_, new_n34813_ );
xor  ( new_n34816_, new_n34815_, new_n896_ );
or   ( new_n34817_, new_n34816_, new_n34812_ );
and  ( new_n34818_, new_n34816_, new_n34812_ );
or   ( new_n34819_, new_n897_, new_n30120_ );
or   ( new_n34820_, new_n899_, new_n29619_ );
and  ( new_n34821_, new_n34820_, new_n34819_ );
xor  ( new_n34822_, new_n34821_, new_n748_ );
or   ( new_n34823_, new_n34822_, new_n34818_ );
and  ( new_n34824_, new_n34823_, new_n34817_ );
or   ( new_n34825_, new_n34824_, new_n34808_ );
and  ( new_n34826_, new_n34825_, new_n34807_ );
or   ( new_n34827_, new_n7184_, new_n22975_ );
or   ( new_n34828_, new_n7186_, new_n22829_ );
and  ( new_n34829_, new_n34828_, new_n34827_ );
xor  ( new_n34830_, new_n34829_, new_n6638_ );
or   ( new_n34831_, new_n6645_, new_n23166_ );
or   ( new_n34832_, new_n6647_, new_n22973_ );
and  ( new_n34833_, new_n34832_, new_n34831_ );
xor  ( new_n34834_, new_n34833_, new_n6166_ );
or   ( new_n34835_, new_n34834_, new_n34830_ );
and  ( new_n34836_, new_n34834_, new_n34830_ );
or   ( new_n34837_, new_n6173_, new_n23370_ );
or   ( new_n34838_, new_n6175_, new_n23252_ );
and  ( new_n34839_, new_n34838_, new_n34837_ );
xor  ( new_n34840_, new_n34839_, new_n5597_ );
or   ( new_n34841_, new_n34840_, new_n34836_ );
and  ( new_n34842_, new_n34841_, new_n34835_ );
or   ( new_n34843_, new_n8874_, new_n22207_ );
or   ( new_n34844_, new_n8876_, new_n22129_ );
and  ( new_n34845_, new_n34844_, new_n34843_ );
xor  ( new_n34846_, new_n34845_, new_n8257_ );
or   ( new_n34847_, new_n8264_, new_n22423_ );
or   ( new_n34848_, new_n8266_, new_n22304_ );
and  ( new_n34849_, new_n34848_, new_n34847_ );
xor  ( new_n34850_, new_n34849_, new_n7725_ );
or   ( new_n34851_, new_n34850_, new_n34846_ );
and  ( new_n34852_, new_n34850_, new_n34846_ );
or   ( new_n34853_, new_n7732_, new_n22641_ );
or   ( new_n34854_, new_n7734_, new_n22590_ );
and  ( new_n34855_, new_n34854_, new_n34853_ );
xor  ( new_n34856_, new_n34855_, new_n7177_ );
or   ( new_n34857_, new_n34856_, new_n34852_ );
and  ( new_n34858_, new_n34857_, new_n34851_ );
or   ( new_n34859_, new_n34858_, new_n34842_ );
and  ( new_n34860_, new_n34858_, new_n34842_ );
or   ( new_n34861_, new_n10059_, new_n21840_ );
or   ( new_n34862_, new_n10061_, new_n21842_ );
and  ( new_n34863_, new_n34862_, new_n34861_ );
xor  ( new_n34864_, new_n34863_, new_n9421_ );
and  ( new_n34865_, RIbb31aa0_139, RIbb2d888_64 );
or   ( new_n34866_, new_n21792_, RIbb2d888_64 );
and  ( new_n34867_, new_n34866_, RIbb2d900_63 );
or   ( new_n34868_, new_n34867_, new_n34865_ );
or   ( new_n34869_, new_n10770_, new_n21751_ );
and  ( new_n34870_, new_n34869_, new_n34868_ );
nor  ( new_n34871_, new_n34870_, new_n34864_ );
and  ( new_n34872_, new_n34870_, new_n34864_ );
or   ( new_n34873_, new_n9422_, new_n22098_ );
or   ( new_n34874_, new_n9424_, new_n21847_ );
and  ( new_n34875_, new_n34874_, new_n34873_ );
xor  ( new_n34876_, new_n34875_, new_n8873_ );
nor  ( new_n34877_, new_n34876_, new_n34872_ );
nor  ( new_n34878_, new_n34877_, new_n34871_ );
or   ( new_n34879_, new_n34878_, new_n34860_ );
and  ( new_n34880_, new_n34879_, new_n34859_ );
or   ( new_n34881_, new_n34880_, new_n34826_ );
or   ( new_n34882_, new_n4302_, new_n24927_ );
or   ( new_n34883_, new_n4304_, new_n24543_ );
and  ( new_n34884_, new_n34883_, new_n34882_ );
xor  ( new_n34885_, new_n34884_, new_n3895_ );
or   ( new_n34886_, new_n3896_, new_n25048_ );
or   ( new_n34887_, new_n3898_, new_n24925_ );
and  ( new_n34888_, new_n34887_, new_n34886_ );
xor  ( new_n34889_, new_n34888_, new_n3460_ );
or   ( new_n34890_, new_n34889_, new_n34885_ );
and  ( new_n34891_, new_n34889_, new_n34885_ );
or   ( new_n34892_, new_n3461_, new_n25486_ );
or   ( new_n34893_, new_n3463_, new_n25288_ );
and  ( new_n34894_, new_n34893_, new_n34892_ );
xor  ( new_n34895_, new_n34894_, new_n3116_ );
or   ( new_n34896_, new_n34895_, new_n34891_ );
and  ( new_n34897_, new_n34896_, new_n34890_ );
or   ( new_n34898_, new_n3117_, new_n26196_ );
or   ( new_n34899_, new_n3119_, new_n25813_ );
and  ( new_n34900_, new_n34899_, new_n34898_ );
xor  ( new_n34901_, new_n34900_, new_n2800_ );
or   ( new_n34902_, new_n2807_, new_n26372_ );
or   ( new_n34903_, new_n2809_, new_n26063_ );
and  ( new_n34904_, new_n34903_, new_n34902_ );
xor  ( new_n34905_, new_n34904_, new_n2424_ );
or   ( new_n34906_, new_n34905_, new_n34901_ );
and  ( new_n34907_, new_n34905_, new_n34901_ );
or   ( new_n34908_, new_n2425_, new_n26762_ );
or   ( new_n34909_, new_n2427_, new_n26620_ );
and  ( new_n34910_, new_n34909_, new_n34908_ );
xor  ( new_n34911_, new_n34910_, new_n2121_ );
or   ( new_n34912_, new_n34911_, new_n34907_ );
and  ( new_n34913_, new_n34912_, new_n34906_ );
nor  ( new_n34914_, new_n34913_, new_n34897_ );
and  ( new_n34915_, new_n34913_, new_n34897_ );
or   ( new_n34916_, new_n5604_, new_n23733_ );
or   ( new_n34917_, new_n5606_, new_n23554_ );
and  ( new_n34918_, new_n34917_, new_n34916_ );
xor  ( new_n34919_, new_n34918_, new_n5206_ );
or   ( new_n34920_, new_n5207_, new_n24006_ );
or   ( new_n34921_, new_n5209_, new_n23895_ );
and  ( new_n34922_, new_n34921_, new_n34920_ );
xor  ( new_n34923_, new_n34922_, new_n4708_ );
nor  ( new_n34924_, new_n34923_, new_n34919_ );
and  ( new_n34925_, new_n34923_, new_n34919_ );
or   ( new_n34926_, new_n4709_, new_n24418_ );
or   ( new_n34927_, new_n4711_, new_n24227_ );
and  ( new_n34928_, new_n34927_, new_n34926_ );
xor  ( new_n34929_, new_n34928_, new_n4295_ );
nor  ( new_n34930_, new_n34929_, new_n34925_ );
nor  ( new_n34931_, new_n34930_, new_n34924_ );
nor  ( new_n34932_, new_n34931_, new_n34915_ );
nor  ( new_n34933_, new_n34932_, new_n34914_ );
and  ( new_n34934_, new_n34880_, new_n34826_ );
or   ( new_n34935_, new_n34934_, new_n34933_ );
and  ( new_n34936_, new_n34935_, new_n34881_ );
and  ( new_n34937_, new_n34936_, new_n34774_ );
nor  ( new_n34938_, new_n34936_, new_n34774_ );
xnor ( new_n34939_, new_n34635_, new_n34631_ );
xor  ( new_n34940_, new_n34939_, new_n34641_ );
xnor ( new_n34941_, new_n34516_, new_n34512_ );
xor  ( new_n34942_, new_n34941_, new_n34522_ );
nor  ( new_n34943_, new_n34942_, new_n34940_ );
nand ( new_n34944_, new_n34942_, new_n34940_ );
xor  ( new_n34945_, new_n34550_, new_n34546_ );
xor  ( new_n34946_, new_n34945_, new_n34556_ );
and  ( new_n34947_, new_n34946_, new_n34944_ );
or   ( new_n34948_, new_n34947_, new_n34943_ );
or   ( new_n34949_, new_n409_, new_n31654_ );
or   ( new_n34950_, new_n411_, new_n31333_ );
and  ( new_n34951_, new_n34950_, new_n34949_ );
xor  ( new_n34952_, new_n34951_, new_n328_ );
and  ( new_n34953_, new_n334_, RIbb33378_192 );
or   ( new_n34954_, new_n34953_, new_n331_ );
or   ( new_n34955_, new_n13845_, new_n31952_ );
and  ( new_n34956_, new_n34955_, new_n34954_ );
or   ( new_n34957_, new_n34956_, new_n34952_ );
nand ( new_n34958_, new_n34956_, new_n34952_ );
xor  ( new_n34959_, new_n34532_, new_n34528_ );
xnor ( new_n34960_, new_n34959_, new_n34538_ );
nand ( new_n34961_, new_n34960_, new_n34958_ );
and  ( new_n34962_, new_n34961_, new_n34957_ );
and  ( new_n34963_, new_n34962_, new_n34948_ );
nor  ( new_n34964_, new_n34962_, new_n34948_ );
xnor ( new_n34965_, new_n34568_, new_n34564_ );
xor  ( new_n34966_, new_n34965_, new_n34574_ );
xnor ( new_n34967_, new_n34619_, new_n34615_ );
xor  ( new_n34968_, new_n34967_, new_n34625_ );
nor  ( new_n34969_, new_n34968_, new_n34966_ );
and  ( new_n34970_, new_n34968_, new_n34966_ );
xor  ( new_n34971_, new_n34653_, new_n34649_ );
xnor ( new_n34972_, new_n34971_, new_n34659_ );
nor  ( new_n34973_, new_n34972_, new_n34970_ );
nor  ( new_n34974_, new_n34973_, new_n34969_ );
nor  ( new_n34975_, new_n34974_, new_n34964_ );
nor  ( new_n34976_, new_n34975_, new_n34963_ );
nor  ( new_n34977_, new_n34976_, new_n34938_ );
nor  ( new_n34978_, new_n34977_, new_n34937_ );
or   ( new_n34979_, new_n34978_, new_n34764_ );
and  ( new_n34980_, new_n34979_, new_n34763_ );
or   ( new_n34981_, new_n34980_, new_n34734_ );
and  ( new_n34982_, new_n34981_, new_n34733_ );
xor  ( new_n34983_, new_n34465_, new_n34455_ );
xor  ( new_n34984_, new_n34983_, new_n34708_ );
or   ( new_n34985_, new_n34984_, new_n34982_ );
and  ( new_n34986_, new_n34984_, new_n34982_ );
xor  ( new_n34987_, new_n34445_, new_n34443_ );
xor  ( new_n34988_, new_n34987_, new_n34449_ );
or   ( new_n34989_, new_n34988_, new_n34986_ );
and  ( new_n34990_, new_n34989_, new_n34985_ );
or   ( new_n34991_, new_n34990_, new_n34720_ );
and  ( new_n34992_, new_n34990_, new_n34720_ );
xor  ( new_n34993_, new_n34179_, new_n34169_ );
xor  ( new_n34994_, new_n34993_, new_n34425_ );
or   ( new_n34995_, new_n34994_, new_n34992_ );
and  ( new_n34996_, new_n34995_, new_n34991_ );
nor  ( new_n34997_, new_n34996_, new_n34718_ );
xor  ( new_n34998_, new_n34984_, new_n34982_ );
xor  ( new_n34999_, new_n34998_, new_n34988_ );
xnor ( new_n35000_, new_n34936_, new_n34774_ );
xor  ( new_n35001_, new_n35000_, new_n34976_ );
xnor ( new_n35002_, new_n34746_, new_n34736_ );
xor  ( new_n35003_, new_n35002_, new_n34750_ );
nor  ( new_n35004_, new_n35003_, new_n35001_ );
nand ( new_n35005_, new_n35003_, new_n35001_ );
xor  ( new_n35006_, new_n34756_, new_n34754_ );
xor  ( new_n35007_, new_n35006_, new_n34760_ );
and  ( new_n35008_, new_n35007_, new_n35005_ );
or   ( new_n35009_, new_n35008_, new_n35004_ );
xor  ( new_n35010_, new_n34726_, new_n34724_ );
xor  ( new_n35011_, new_n35010_, new_n34730_ );
nor  ( new_n35012_, new_n35011_, new_n35009_ );
and  ( new_n35013_, new_n35011_, new_n35009_ );
xnor ( new_n35014_, new_n34858_, new_n34842_ );
xor  ( new_n35015_, new_n35014_, new_n34878_ );
xnor ( new_n35016_, new_n34913_, new_n34897_ );
xor  ( new_n35017_, new_n35016_, new_n34931_ );
or   ( new_n35018_, new_n35017_, new_n35015_ );
xor  ( new_n35019_, new_n34806_, new_n34790_ );
xor  ( new_n35020_, new_n35019_, new_n34824_ );
xor  ( new_n35021_, new_n34942_, new_n34940_ );
xor  ( new_n35022_, new_n35021_, new_n34946_ );
nand ( new_n35023_, new_n35022_, new_n35020_ );
nor  ( new_n35024_, new_n35022_, new_n35020_ );
xor  ( new_n35025_, new_n34956_, new_n34952_ );
xor  ( new_n35026_, new_n35025_, new_n34960_ );
or   ( new_n35027_, new_n35026_, new_n35024_ );
and  ( new_n35028_, new_n35027_, new_n35023_ );
or   ( new_n35029_, new_n35028_, new_n35018_ );
and  ( new_n35030_, new_n35028_, new_n35018_ );
xnor ( new_n35031_, new_n34606_, new_n34590_ );
xor  ( new_n35032_, new_n35031_, new_n34576_ );
or   ( new_n35033_, new_n35032_, new_n35030_ );
and  ( new_n35034_, new_n35033_, new_n35029_ );
xnor ( new_n35035_, new_n34962_, new_n34948_ );
xor  ( new_n35036_, new_n35035_, new_n34974_ );
xnor ( new_n35037_, new_n34740_, new_n34738_ );
xor  ( new_n35038_, new_n35037_, new_n34744_ );
nand ( new_n35039_, new_n35038_, new_n35036_ );
nor  ( new_n35040_, new_n35038_, new_n35036_ );
xor  ( new_n35041_, new_n34768_, new_n34766_ );
xnor ( new_n35042_, new_n35041_, new_n34772_ );
or   ( new_n35043_, new_n35042_, new_n35040_ );
and  ( new_n35044_, new_n35043_, new_n35039_ );
nor  ( new_n35045_, new_n35044_, new_n35034_ );
and  ( new_n35046_, new_n35044_, new_n35034_ );
xnor ( new_n35047_, new_n34598_, new_n34594_ );
xor  ( new_n35048_, new_n35047_, new_n34604_ );
xor  ( new_n35049_, new_n34586_, new_n34580_ );
xor  ( new_n35050_, new_n35049_, new_n332_ );
nor  ( new_n35051_, new_n35050_, new_n35048_ );
nand ( new_n35052_, new_n35050_, new_n35048_ );
xor  ( new_n35053_, new_n34968_, new_n34966_ );
xnor ( new_n35054_, new_n35053_, new_n34972_ );
and  ( new_n35055_, new_n35054_, new_n35052_ );
or   ( new_n35056_, new_n35055_, new_n35051_ );
or   ( new_n35057_, new_n6173_, new_n23554_ );
or   ( new_n35058_, new_n6175_, new_n23370_ );
and  ( new_n35059_, new_n35058_, new_n35057_ );
xor  ( new_n35060_, new_n35059_, new_n5597_ );
or   ( new_n35061_, new_n5604_, new_n23895_ );
or   ( new_n35062_, new_n5606_, new_n23733_ );
and  ( new_n35063_, new_n35062_, new_n35061_ );
xor  ( new_n35064_, new_n35063_, new_n5206_ );
or   ( new_n35065_, new_n35064_, new_n35060_ );
and  ( new_n35066_, new_n35064_, new_n35060_ );
or   ( new_n35067_, new_n5207_, new_n24227_ );
or   ( new_n35068_, new_n5209_, new_n24006_ );
and  ( new_n35069_, new_n35068_, new_n35067_ );
xor  ( new_n35070_, new_n35069_, new_n4708_ );
or   ( new_n35071_, new_n35070_, new_n35066_ );
and  ( new_n35072_, new_n35071_, new_n35065_ );
or   ( new_n35073_, new_n3461_, new_n25813_ );
or   ( new_n35074_, new_n3463_, new_n25486_ );
and  ( new_n35075_, new_n35074_, new_n35073_ );
xor  ( new_n35076_, new_n35075_, new_n3116_ );
or   ( new_n35077_, new_n3117_, new_n26063_ );
or   ( new_n35078_, new_n3119_, new_n26196_ );
and  ( new_n35079_, new_n35078_, new_n35077_ );
xor  ( new_n35080_, new_n35079_, new_n2800_ );
or   ( new_n35081_, new_n35080_, new_n35076_ );
and  ( new_n35082_, new_n35080_, new_n35076_ );
or   ( new_n35083_, new_n2807_, new_n26620_ );
or   ( new_n35084_, new_n2809_, new_n26372_ );
and  ( new_n35085_, new_n35084_, new_n35083_ );
xor  ( new_n35086_, new_n35085_, new_n2424_ );
or   ( new_n35087_, new_n35086_, new_n35082_ );
and  ( new_n35088_, new_n35087_, new_n35081_ );
or   ( new_n35089_, new_n35088_, new_n35072_ );
and  ( new_n35090_, new_n35088_, new_n35072_ );
or   ( new_n35091_, new_n4709_, new_n24543_ );
or   ( new_n35092_, new_n4711_, new_n24418_ );
and  ( new_n35093_, new_n35092_, new_n35091_ );
xor  ( new_n35094_, new_n35093_, new_n4295_ );
or   ( new_n35095_, new_n4302_, new_n24925_ );
or   ( new_n35096_, new_n4304_, new_n24927_ );
and  ( new_n35097_, new_n35096_, new_n35095_ );
xor  ( new_n35098_, new_n35097_, new_n3895_ );
or   ( new_n35099_, new_n35098_, new_n35094_ );
and  ( new_n35100_, new_n35098_, new_n35094_ );
or   ( new_n35101_, new_n3896_, new_n25288_ );
or   ( new_n35102_, new_n3898_, new_n25048_ );
and  ( new_n35103_, new_n35102_, new_n35101_ );
xor  ( new_n35104_, new_n35103_, new_n3460_ );
or   ( new_n35105_, new_n35104_, new_n35100_ );
and  ( new_n35106_, new_n35105_, new_n35099_ );
or   ( new_n35107_, new_n35106_, new_n35090_ );
and  ( new_n35108_, new_n35107_, new_n35089_ );
or   ( new_n35109_, new_n9422_, new_n22129_ );
or   ( new_n35110_, new_n9424_, new_n22098_ );
and  ( new_n35111_, new_n35110_, new_n35109_ );
xor  ( new_n35112_, new_n35111_, new_n8873_ );
or   ( new_n35113_, new_n8874_, new_n22304_ );
or   ( new_n35114_, new_n8876_, new_n22207_ );
and  ( new_n35115_, new_n35114_, new_n35113_ );
xor  ( new_n35116_, new_n35115_, new_n8257_ );
nor  ( new_n35117_, new_n35116_, new_n35112_ );
and  ( new_n35118_, new_n35116_, new_n35112_ );
or   ( new_n35119_, new_n8264_, new_n22590_ );
or   ( new_n35120_, new_n8266_, new_n22423_ );
and  ( new_n35121_, new_n35120_, new_n35119_ );
xor  ( new_n35122_, new_n35121_, new_n7725_ );
nor  ( new_n35123_, new_n35122_, new_n35118_ );
nor  ( new_n35124_, new_n35123_, new_n35117_ );
or   ( new_n35125_, new_n10059_, new_n21847_ );
or   ( new_n35126_, new_n10061_, new_n21840_ );
and  ( new_n35127_, new_n35126_, new_n35125_ );
xor  ( new_n35128_, new_n35127_, new_n9421_ );
and  ( new_n35129_, RIbb31b18_140, RIbb2d888_64 );
or   ( new_n35130_, new_n21842_, RIbb2d888_64 );
and  ( new_n35131_, new_n35130_, RIbb2d900_63 );
or   ( new_n35132_, new_n35131_, new_n35129_ );
or   ( new_n35133_, new_n10770_, new_n21792_ );
and  ( new_n35134_, new_n35133_, new_n35132_ );
nor  ( new_n35135_, new_n35134_, new_n35128_ );
and  ( new_n35136_, new_n35134_, new_n35128_ );
nor  ( new_n35137_, new_n35136_, new_n327_ );
nor  ( new_n35138_, new_n35137_, new_n35135_ );
or   ( new_n35139_, new_n7732_, new_n22829_ );
or   ( new_n35140_, new_n7734_, new_n22641_ );
and  ( new_n35141_, new_n35140_, new_n35139_ );
xor  ( new_n35142_, new_n35141_, new_n7177_ );
or   ( new_n35143_, new_n7184_, new_n22973_ );
or   ( new_n35144_, new_n7186_, new_n22975_ );
and  ( new_n35145_, new_n35144_, new_n35143_ );
xor  ( new_n35146_, new_n35145_, new_n6638_ );
or   ( new_n35147_, new_n35146_, new_n35142_ );
and  ( new_n35148_, new_n35146_, new_n35142_ );
or   ( new_n35149_, new_n6645_, new_n23252_ );
or   ( new_n35150_, new_n6647_, new_n23166_ );
and  ( new_n35151_, new_n35150_, new_n35149_ );
xor  ( new_n35152_, new_n35151_, new_n6166_ );
or   ( new_n35153_, new_n35152_, new_n35148_ );
and  ( new_n35154_, new_n35153_, new_n35147_ );
and  ( new_n35155_, new_n35154_, new_n35138_ );
or   ( new_n35156_, new_n35155_, new_n35124_ );
or   ( new_n35157_, new_n35154_, new_n35138_ );
and  ( new_n35158_, new_n35157_, new_n35156_ );
or   ( new_n35159_, new_n35158_, new_n35108_ );
or   ( new_n35160_, new_n2425_, new_n27085_ );
or   ( new_n35161_, new_n2427_, new_n26762_ );
and  ( new_n35162_, new_n35161_, new_n35160_ );
xor  ( new_n35163_, new_n35162_, new_n2121_ );
or   ( new_n35164_, new_n2122_, new_n27602_ );
or   ( new_n35165_, new_n2124_, new_n27396_ );
and  ( new_n35166_, new_n35165_, new_n35164_ );
xor  ( new_n35167_, new_n35166_, new_n1843_ );
or   ( new_n35168_, new_n35167_, new_n35163_ );
and  ( new_n35169_, new_n35167_, new_n35163_ );
or   ( new_n35170_, new_n1844_, new_n28108_ );
or   ( new_n35171_, new_n1846_, new_n27763_ );
and  ( new_n35172_, new_n35171_, new_n35170_ );
xor  ( new_n35173_, new_n35172_, new_n1586_ );
or   ( new_n35174_, new_n35173_, new_n35169_ );
and  ( new_n35175_, new_n35174_, new_n35168_ );
or   ( new_n35176_, new_n897_, new_n30227_ );
or   ( new_n35177_, new_n899_, new_n30120_ );
and  ( new_n35178_, new_n35177_, new_n35176_ );
xor  ( new_n35179_, new_n35178_, new_n748_ );
or   ( new_n35180_, new_n755_, new_n30798_ );
or   ( new_n35181_, new_n757_, new_n30800_ );
and  ( new_n35182_, new_n35181_, new_n35180_ );
xor  ( new_n35183_, new_n35182_, new_n523_ );
or   ( new_n35184_, new_n35183_, new_n35179_ );
and  ( new_n35185_, new_n35183_, new_n35179_ );
or   ( new_n35186_, new_n524_, new_n31654_ );
or   ( new_n35187_, new_n526_, new_n31333_ );
and  ( new_n35188_, new_n35187_, new_n35186_ );
xor  ( new_n35189_, new_n35188_, new_n403_ );
or   ( new_n35190_, new_n35189_, new_n35185_ );
and  ( new_n35191_, new_n35190_, new_n35184_ );
nor  ( new_n35192_, new_n35191_, new_n35175_ );
and  ( new_n35193_, new_n35191_, new_n35175_ );
or   ( new_n35194_, new_n1593_, new_n28531_ );
or   ( new_n35195_, new_n1595_, new_n28314_ );
and  ( new_n35196_, new_n35195_, new_n35194_ );
xor  ( new_n35197_, new_n35196_, new_n1358_ );
or   ( new_n35198_, new_n1364_, new_n29261_ );
or   ( new_n35199_, new_n1366_, new_n29263_ );
and  ( new_n35200_, new_n35199_, new_n35198_ );
xor  ( new_n35201_, new_n35200_, new_n1129_ );
nor  ( new_n35202_, new_n35201_, new_n35197_ );
and  ( new_n35203_, new_n35201_, new_n35197_ );
or   ( new_n35204_, new_n1135_, new_n29619_ );
or   ( new_n35205_, new_n1137_, new_n29474_ );
and  ( new_n35206_, new_n35205_, new_n35204_ );
xor  ( new_n35207_, new_n35206_, new_n896_ );
nor  ( new_n35208_, new_n35207_, new_n35203_ );
nor  ( new_n35209_, new_n35208_, new_n35202_ );
nor  ( new_n35210_, new_n35209_, new_n35193_ );
nor  ( new_n35211_, new_n35210_, new_n35192_ );
and  ( new_n35212_, new_n35158_, new_n35108_ );
or   ( new_n35213_, new_n35212_, new_n35211_ );
and  ( new_n35214_, new_n35213_, new_n35159_ );
and  ( new_n35215_, new_n35214_, new_n35056_ );
nor  ( new_n35216_, new_n35214_, new_n35056_ );
xnor ( new_n35217_, new_n34798_, new_n34794_ );
xor  ( new_n35218_, new_n35217_, new_n34804_ );
xnor ( new_n35219_, new_n34782_, new_n34778_ );
xor  ( new_n35220_, new_n35219_, new_n34788_ );
or   ( new_n35221_, new_n35220_, new_n35218_ );
and  ( new_n35222_, new_n35220_, new_n35218_ );
xor  ( new_n35223_, new_n34816_, new_n34812_ );
xnor ( new_n35224_, new_n35223_, new_n34822_ );
or   ( new_n35225_, new_n35224_, new_n35222_ );
and  ( new_n35226_, new_n35225_, new_n35221_ );
xnor ( new_n35227_, new_n34850_, new_n34846_ );
xor  ( new_n35228_, new_n35227_, new_n34856_ );
xnor ( new_n35229_, new_n34834_, new_n34830_ );
xor  ( new_n35230_, new_n35229_, new_n34840_ );
or   ( new_n35231_, new_n35230_, new_n35228_ );
and  ( new_n35232_, new_n35230_, new_n35228_ );
xor  ( new_n35233_, new_n34870_, new_n34864_ );
xnor ( new_n35234_, new_n35233_, new_n34876_ );
or   ( new_n35235_, new_n35234_, new_n35232_ );
and  ( new_n35236_, new_n35235_, new_n35231_ );
nor  ( new_n35237_, new_n35236_, new_n35226_ );
and  ( new_n35238_, new_n35236_, new_n35226_ );
xnor ( new_n35239_, new_n34905_, new_n34901_ );
xor  ( new_n35240_, new_n35239_, new_n34911_ );
xnor ( new_n35241_, new_n34889_, new_n34885_ );
xor  ( new_n35242_, new_n35241_, new_n34895_ );
nor  ( new_n35243_, new_n35242_, new_n35240_ );
and  ( new_n35244_, new_n35242_, new_n35240_ );
xor  ( new_n35245_, new_n34923_, new_n34919_ );
xnor ( new_n35246_, new_n35245_, new_n34929_ );
nor  ( new_n35247_, new_n35246_, new_n35244_ );
nor  ( new_n35248_, new_n35247_, new_n35243_ );
nor  ( new_n35249_, new_n35248_, new_n35238_ );
nor  ( new_n35250_, new_n35249_, new_n35237_ );
nor  ( new_n35251_, new_n35250_, new_n35216_ );
nor  ( new_n35252_, new_n35251_, new_n35215_ );
nor  ( new_n35253_, new_n35252_, new_n35046_ );
nor  ( new_n35254_, new_n35253_, new_n35045_ );
nor  ( new_n35255_, new_n35254_, new_n35013_ );
or   ( new_n35256_, new_n35255_, new_n35012_ );
xnor ( new_n35257_, new_n34496_, new_n34486_ );
xor  ( new_n35258_, new_n35257_, new_n34706_ );
nand ( new_n35259_, new_n35258_, new_n35256_ );
nor  ( new_n35260_, new_n35258_, new_n35256_ );
xor  ( new_n35261_, new_n34732_, new_n34722_ );
xor  ( new_n35262_, new_n35261_, new_n34980_ );
or   ( new_n35263_, new_n35262_, new_n35260_ );
and  ( new_n35264_, new_n35263_, new_n35259_ );
nor  ( new_n35265_, new_n35264_, new_n34999_ );
xnor ( new_n35266_, new_n34990_, new_n34720_ );
xor  ( new_n35267_, new_n35266_, new_n34994_ );
and  ( new_n35268_, new_n35267_, new_n35265_ );
xor  ( new_n35269_, new_n35258_, new_n35256_ );
xor  ( new_n35270_, new_n35269_, new_n35262_ );
xor  ( new_n35271_, new_n35017_, new_n35015_ );
xnor ( new_n35272_, new_n35022_, new_n35020_ );
xor  ( new_n35273_, new_n35272_, new_n35026_ );
and  ( new_n35274_, new_n35273_, new_n35271_ );
nor  ( new_n35275_, new_n35273_, new_n35271_ );
xor  ( new_n35276_, new_n35088_, new_n35072_ );
xor  ( new_n35277_, new_n35276_, new_n35106_ );
xor  ( new_n35278_, new_n35154_, new_n35138_ );
xor  ( new_n35279_, new_n35278_, new_n35124_ );
and  ( new_n35280_, new_n35279_, new_n35277_ );
nor  ( new_n35281_, new_n35279_, new_n35277_ );
xor  ( new_n35282_, new_n35191_, new_n35175_ );
xnor ( new_n35283_, new_n35282_, new_n35209_ );
nor  ( new_n35284_, new_n35283_, new_n35281_ );
nor  ( new_n35285_, new_n35284_, new_n35280_ );
nor  ( new_n35286_, new_n35285_, new_n35275_ );
nor  ( new_n35287_, new_n35286_, new_n35274_ );
xnor ( new_n35288_, new_n35242_, new_n35240_ );
xor  ( new_n35289_, new_n35288_, new_n35246_ );
xnor ( new_n35290_, new_n35220_, new_n35218_ );
xor  ( new_n35291_, new_n35290_, new_n35224_ );
nor  ( new_n35292_, new_n35291_, new_n35289_ );
and  ( new_n35293_, new_n35291_, new_n35289_ );
xor  ( new_n35294_, new_n35230_, new_n35228_ );
xnor ( new_n35295_, new_n35294_, new_n35234_ );
nor  ( new_n35296_, new_n35295_, new_n35293_ );
nor  ( new_n35297_, new_n35296_, new_n35292_ );
or   ( new_n35298_, new_n5604_, new_n24006_ );
or   ( new_n35299_, new_n5606_, new_n23895_ );
and  ( new_n35300_, new_n35299_, new_n35298_ );
xor  ( new_n35301_, new_n35300_, new_n5206_ );
or   ( new_n35302_, new_n5207_, new_n24418_ );
or   ( new_n35303_, new_n5209_, new_n24227_ );
and  ( new_n35304_, new_n35303_, new_n35302_ );
xor  ( new_n35305_, new_n35304_, new_n4708_ );
or   ( new_n35306_, new_n35305_, new_n35301_ );
and  ( new_n35307_, new_n35305_, new_n35301_ );
or   ( new_n35308_, new_n4709_, new_n24927_ );
or   ( new_n35309_, new_n4711_, new_n24543_ );
and  ( new_n35310_, new_n35309_, new_n35308_ );
xor  ( new_n35311_, new_n35310_, new_n4295_ );
or   ( new_n35312_, new_n35311_, new_n35307_ );
and  ( new_n35313_, new_n35312_, new_n35306_ );
or   ( new_n35314_, new_n4302_, new_n25048_ );
or   ( new_n35315_, new_n4304_, new_n24925_ );
and  ( new_n35316_, new_n35315_, new_n35314_ );
xor  ( new_n35317_, new_n35316_, new_n3895_ );
or   ( new_n35318_, new_n3896_, new_n25486_ );
or   ( new_n35319_, new_n3898_, new_n25288_ );
and  ( new_n35320_, new_n35319_, new_n35318_ );
xor  ( new_n35321_, new_n35320_, new_n3460_ );
or   ( new_n35322_, new_n35321_, new_n35317_ );
and  ( new_n35323_, new_n35321_, new_n35317_ );
or   ( new_n35324_, new_n3461_, new_n26196_ );
or   ( new_n35325_, new_n3463_, new_n25813_ );
and  ( new_n35326_, new_n35325_, new_n35324_ );
xor  ( new_n35327_, new_n35326_, new_n3116_ );
or   ( new_n35328_, new_n35327_, new_n35323_ );
and  ( new_n35329_, new_n35328_, new_n35322_ );
or   ( new_n35330_, new_n35329_, new_n35313_ );
and  ( new_n35331_, new_n35329_, new_n35313_ );
or   ( new_n35332_, new_n3117_, new_n26372_ );
or   ( new_n35333_, new_n3119_, new_n26063_ );
and  ( new_n35334_, new_n35333_, new_n35332_ );
xor  ( new_n35335_, new_n35334_, new_n2800_ );
or   ( new_n35336_, new_n2807_, new_n26762_ );
or   ( new_n35337_, new_n2809_, new_n26620_ );
and  ( new_n35338_, new_n35337_, new_n35336_ );
xor  ( new_n35339_, new_n35338_, new_n2424_ );
or   ( new_n35340_, new_n35339_, new_n35335_ );
and  ( new_n35341_, new_n35339_, new_n35335_ );
or   ( new_n35342_, new_n2425_, new_n27396_ );
or   ( new_n35343_, new_n2427_, new_n27085_ );
and  ( new_n35344_, new_n35343_, new_n35342_ );
xor  ( new_n35345_, new_n35344_, new_n2121_ );
or   ( new_n35346_, new_n35345_, new_n35341_ );
and  ( new_n35347_, new_n35346_, new_n35340_ );
or   ( new_n35348_, new_n35347_, new_n35331_ );
and  ( new_n35349_, new_n35348_, new_n35330_ );
or   ( new_n35350_, new_n1364_, new_n29474_ );
or   ( new_n35351_, new_n1366_, new_n29261_ );
and  ( new_n35352_, new_n35351_, new_n35350_ );
xor  ( new_n35353_, new_n35352_, new_n1129_ );
or   ( new_n35354_, new_n1135_, new_n30120_ );
or   ( new_n35355_, new_n1137_, new_n29619_ );
and  ( new_n35356_, new_n35355_, new_n35354_ );
xor  ( new_n35357_, new_n35356_, new_n896_ );
nor  ( new_n35358_, new_n35357_, new_n35353_ );
and  ( new_n35359_, new_n35357_, new_n35353_ );
or   ( new_n35360_, new_n897_, new_n30800_ );
or   ( new_n35361_, new_n899_, new_n30227_ );
and  ( new_n35362_, new_n35361_, new_n35360_ );
xor  ( new_n35363_, new_n35362_, new_n748_ );
nor  ( new_n35364_, new_n35363_, new_n35359_ );
nor  ( new_n35365_, new_n35364_, new_n35358_ );
or   ( new_n35366_, new_n755_, new_n31333_ );
or   ( new_n35367_, new_n757_, new_n30798_ );
and  ( new_n35368_, new_n35367_, new_n35366_ );
xor  ( new_n35369_, new_n35368_, new_n523_ );
or   ( new_n35370_, new_n524_, new_n31952_ );
or   ( new_n35371_, new_n526_, new_n31654_ );
and  ( new_n35372_, new_n35371_, new_n35370_ );
xor  ( new_n35373_, new_n35372_, new_n403_ );
and  ( new_n35374_, new_n35373_, new_n35369_ );
or   ( new_n35375_, new_n2122_, new_n27763_ );
or   ( new_n35376_, new_n2124_, new_n27602_ );
and  ( new_n35377_, new_n35376_, new_n35375_ );
xor  ( new_n35378_, new_n35377_, new_n1843_ );
or   ( new_n35379_, new_n1844_, new_n28314_ );
or   ( new_n35380_, new_n1846_, new_n28108_ );
and  ( new_n35381_, new_n35380_, new_n35379_ );
xor  ( new_n35382_, new_n35381_, new_n1586_ );
or   ( new_n35383_, new_n35382_, new_n35378_ );
and  ( new_n35384_, new_n35382_, new_n35378_ );
or   ( new_n35385_, new_n1593_, new_n29263_ );
or   ( new_n35386_, new_n1595_, new_n28531_ );
and  ( new_n35387_, new_n35386_, new_n35385_ );
xor  ( new_n35388_, new_n35387_, new_n1358_ );
or   ( new_n35389_, new_n35388_, new_n35384_ );
and  ( new_n35390_, new_n35389_, new_n35383_ );
and  ( new_n35391_, new_n35390_, new_n35374_ );
or   ( new_n35392_, new_n35391_, new_n35365_ );
or   ( new_n35393_, new_n35390_, new_n35374_ );
and  ( new_n35394_, new_n35393_, new_n35392_ );
nor  ( new_n35395_, new_n35394_, new_n35349_ );
or   ( new_n35396_, new_n10059_, new_n22098_ );
or   ( new_n35397_, new_n10061_, new_n21847_ );
and  ( new_n35398_, new_n35397_, new_n35396_ );
xor  ( new_n35399_, new_n35398_, new_n9421_ );
and  ( new_n35400_, RIbb31b90_141, RIbb2d888_64 );
or   ( new_n35401_, new_n21840_, RIbb2d888_64 );
and  ( new_n35402_, new_n35401_, RIbb2d900_63 );
or   ( new_n35403_, new_n35402_, new_n35400_ );
or   ( new_n35404_, new_n10770_, new_n21842_ );
and  ( new_n35405_, new_n35404_, new_n35403_ );
or   ( new_n35406_, new_n35405_, new_n35399_ );
and  ( new_n35407_, new_n35405_, new_n35399_ );
or   ( new_n35408_, new_n9422_, new_n22207_ );
or   ( new_n35409_, new_n9424_, new_n22129_ );
and  ( new_n35410_, new_n35409_, new_n35408_ );
xor  ( new_n35411_, new_n35410_, new_n8873_ );
or   ( new_n35412_, new_n35411_, new_n35407_ );
and  ( new_n35413_, new_n35412_, new_n35406_ );
or   ( new_n35414_, new_n7184_, new_n23166_ );
or   ( new_n35415_, new_n7186_, new_n22973_ );
and  ( new_n35416_, new_n35415_, new_n35414_ );
xor  ( new_n35417_, new_n35416_, new_n6638_ );
or   ( new_n35418_, new_n6645_, new_n23370_ );
or   ( new_n35419_, new_n6647_, new_n23252_ );
and  ( new_n35420_, new_n35419_, new_n35418_ );
xor  ( new_n35421_, new_n35420_, new_n6166_ );
or   ( new_n35422_, new_n35421_, new_n35417_ );
and  ( new_n35423_, new_n35421_, new_n35417_ );
or   ( new_n35424_, new_n6173_, new_n23733_ );
or   ( new_n35425_, new_n6175_, new_n23554_ );
and  ( new_n35426_, new_n35425_, new_n35424_ );
xor  ( new_n35427_, new_n35426_, new_n5597_ );
or   ( new_n35428_, new_n35427_, new_n35423_ );
and  ( new_n35429_, new_n35428_, new_n35422_ );
nor  ( new_n35430_, new_n35429_, new_n35413_ );
and  ( new_n35431_, new_n35429_, new_n35413_ );
or   ( new_n35432_, new_n8874_, new_n22423_ );
or   ( new_n35433_, new_n8876_, new_n22304_ );
and  ( new_n35434_, new_n35433_, new_n35432_ );
xor  ( new_n35435_, new_n35434_, new_n8257_ );
or   ( new_n35436_, new_n8264_, new_n22641_ );
or   ( new_n35437_, new_n8266_, new_n22590_ );
and  ( new_n35438_, new_n35437_, new_n35436_ );
xor  ( new_n35439_, new_n35438_, new_n7725_ );
nor  ( new_n35440_, new_n35439_, new_n35435_ );
and  ( new_n35441_, new_n35439_, new_n35435_ );
or   ( new_n35442_, new_n7732_, new_n22975_ );
or   ( new_n35443_, new_n7734_, new_n22829_ );
and  ( new_n35444_, new_n35443_, new_n35442_ );
xor  ( new_n35445_, new_n35444_, new_n7177_ );
nor  ( new_n35446_, new_n35445_, new_n35441_ );
nor  ( new_n35447_, new_n35446_, new_n35440_ );
nor  ( new_n35448_, new_n35447_, new_n35431_ );
nor  ( new_n35449_, new_n35448_, new_n35430_ );
and  ( new_n35450_, new_n35394_, new_n35349_ );
nor  ( new_n35451_, new_n35450_, new_n35449_ );
nor  ( new_n35452_, new_n35451_, new_n35395_ );
and  ( new_n35453_, new_n35452_, new_n35297_ );
nor  ( new_n35454_, new_n35452_, new_n35297_ );
and  ( new_n35455_, new_n371_, RIbb33378_192 );
or   ( new_n35456_, new_n35455_, new_n328_ );
nand ( new_n35457_, new_n35455_, new_n325_ );
and  ( new_n35458_, new_n35457_, new_n35456_ );
xnor ( new_n35459_, new_n35201_, new_n35197_ );
xor  ( new_n35460_, new_n35459_, new_n35207_ );
or   ( new_n35461_, new_n35460_, new_n35458_ );
and  ( new_n35462_, new_n35460_, new_n35458_ );
xor  ( new_n35463_, new_n35183_, new_n35179_ );
xnor ( new_n35464_, new_n35463_, new_n35189_ );
or   ( new_n35465_, new_n35464_, new_n35462_ );
and  ( new_n35466_, new_n35465_, new_n35461_ );
xnor ( new_n35467_, new_n35116_, new_n35112_ );
xor  ( new_n35468_, new_n35467_, new_n35122_ );
xnor ( new_n35469_, new_n35146_, new_n35142_ );
xor  ( new_n35470_, new_n35469_, new_n35152_ );
or   ( new_n35471_, new_n35470_, new_n35468_ );
and  ( new_n35472_, new_n35470_, new_n35468_ );
xor  ( new_n35473_, new_n35064_, new_n35060_ );
xnor ( new_n35474_, new_n35473_, new_n35070_ );
or   ( new_n35475_, new_n35474_, new_n35472_ );
and  ( new_n35476_, new_n35475_, new_n35471_ );
nor  ( new_n35477_, new_n35476_, new_n35466_ );
and  ( new_n35478_, new_n35476_, new_n35466_ );
xnor ( new_n35479_, new_n35167_, new_n35163_ );
xor  ( new_n35480_, new_n35479_, new_n35173_ );
xnor ( new_n35481_, new_n35080_, new_n35076_ );
xor  ( new_n35482_, new_n35481_, new_n35086_ );
nor  ( new_n35483_, new_n35482_, new_n35480_ );
and  ( new_n35484_, new_n35482_, new_n35480_ );
xor  ( new_n35485_, new_n35098_, new_n35094_ );
xnor ( new_n35486_, new_n35485_, new_n35104_ );
nor  ( new_n35487_, new_n35486_, new_n35484_ );
nor  ( new_n35488_, new_n35487_, new_n35483_ );
nor  ( new_n35489_, new_n35488_, new_n35478_ );
nor  ( new_n35490_, new_n35489_, new_n35477_ );
nor  ( new_n35491_, new_n35490_, new_n35454_ );
nor  ( new_n35492_, new_n35491_, new_n35453_ );
and  ( new_n35493_, new_n35492_, new_n35287_ );
not  ( new_n35494_, new_n35493_ );
xor  ( new_n35495_, new_n35236_, new_n35226_ );
xor  ( new_n35496_, new_n35495_, new_n35248_ );
xnor ( new_n35497_, new_n35158_, new_n35108_ );
xor  ( new_n35498_, new_n35497_, new_n35211_ );
nor  ( new_n35499_, new_n35498_, new_n35496_ );
and  ( new_n35500_, new_n35498_, new_n35496_ );
xor  ( new_n35501_, new_n35050_, new_n35048_ );
xnor ( new_n35502_, new_n35501_, new_n35054_ );
nor  ( new_n35503_, new_n35502_, new_n35500_ );
nor  ( new_n35504_, new_n35503_, new_n35499_ );
not  ( new_n35505_, new_n35504_ );
and  ( new_n35506_, new_n35505_, new_n35494_ );
nor  ( new_n35507_, new_n35492_, new_n35287_ );
nor  ( new_n35508_, new_n35507_, new_n35506_ );
xor  ( new_n35509_, new_n35003_, new_n35001_ );
xor  ( new_n35510_, new_n35509_, new_n35007_ );
and  ( new_n35511_, new_n35510_, new_n35508_ );
xnor ( new_n35512_, new_n34880_, new_n34826_ );
xor  ( new_n35513_, new_n35512_, new_n34933_ );
xor  ( new_n35514_, new_n35028_, new_n35018_ );
xor  ( new_n35515_, new_n35514_, new_n35032_ );
nor  ( new_n35516_, new_n35515_, new_n35513_ );
and  ( new_n35517_, new_n35515_, new_n35513_ );
xor  ( new_n35518_, new_n35038_, new_n35036_ );
xnor ( new_n35519_, new_n35518_, new_n35042_ );
not  ( new_n35520_, new_n35519_ );
nor  ( new_n35521_, new_n35520_, new_n35517_ );
nor  ( new_n35522_, new_n35521_, new_n35516_ );
nor  ( new_n35523_, new_n35522_, new_n35511_ );
nor  ( new_n35524_, new_n35510_, new_n35508_ );
or   ( new_n35525_, new_n35524_, new_n35523_ );
xnor ( new_n35526_, new_n34762_, new_n34752_ );
xor  ( new_n35527_, new_n35526_, new_n34978_ );
nand ( new_n35528_, new_n35527_, new_n35525_ );
nor  ( new_n35529_, new_n35527_, new_n35525_ );
xor  ( new_n35530_, new_n35011_, new_n35009_ );
xor  ( new_n35531_, new_n35530_, new_n35254_ );
or   ( new_n35532_, new_n35531_, new_n35529_ );
and  ( new_n35533_, new_n35532_, new_n35528_ );
nor  ( new_n35534_, new_n35533_, new_n35270_ );
xor  ( new_n35535_, new_n35264_, new_n34999_ );
and  ( new_n35536_, new_n35535_, new_n35534_ );
xor  ( new_n35537_, new_n35492_, new_n35287_ );
nor  ( new_n35538_, new_n35537_, new_n35505_ );
not  ( new_n35539_, new_n35507_ );
and  ( new_n35540_, new_n35539_, new_n35506_ );
nor  ( new_n35541_, new_n35540_, new_n35538_ );
xor  ( new_n35542_, new_n35515_, new_n35513_ );
xor  ( new_n35543_, new_n35542_, new_n35519_ );
nand ( new_n35544_, new_n35543_, new_n35541_ );
xnor ( new_n35545_, new_n35452_, new_n35297_ );
xor  ( new_n35546_, new_n35545_, new_n35490_ );
xnor ( new_n35547_, new_n35498_, new_n35496_ );
xor  ( new_n35548_, new_n35547_, new_n35502_ );
nor  ( new_n35549_, new_n35548_, new_n35546_ );
nand ( new_n35550_, new_n35548_, new_n35546_ );
xor  ( new_n35551_, new_n35273_, new_n35271_ );
xor  ( new_n35552_, new_n35551_, new_n35285_ );
and  ( new_n35553_, new_n35552_, new_n35550_ );
or   ( new_n35554_, new_n35553_, new_n35549_ );
xor  ( new_n35555_, new_n35214_, new_n35056_ );
xor  ( new_n35556_, new_n35555_, new_n35250_ );
or   ( new_n35557_, new_n35556_, new_n35554_ );
and  ( new_n35558_, new_n35556_, new_n35554_ );
xor  ( new_n35559_, new_n35394_, new_n35349_ );
xnor ( new_n35560_, new_n35559_, new_n35449_ );
not  ( new_n35561_, new_n35560_ );
xnor ( new_n35562_, new_n35476_, new_n35466_ );
xor  ( new_n35563_, new_n35562_, new_n35488_ );
and  ( new_n35564_, new_n35563_, new_n35561_ );
xnor ( new_n35565_, new_n35321_, new_n35317_ );
xor  ( new_n35566_, new_n35565_, new_n35327_ );
xnor ( new_n35567_, new_n35305_, new_n35301_ );
xor  ( new_n35568_, new_n35567_, new_n35311_ );
or   ( new_n35569_, new_n35568_, new_n35566_ );
and  ( new_n35570_, new_n35568_, new_n35566_ );
xor  ( new_n35571_, new_n35339_, new_n35335_ );
xnor ( new_n35572_, new_n35571_, new_n35345_ );
or   ( new_n35573_, new_n35572_, new_n35570_ );
and  ( new_n35574_, new_n35573_, new_n35569_ );
xnor ( new_n35575_, new_n35357_, new_n35353_ );
xor  ( new_n35576_, new_n35575_, new_n35363_ );
xnor ( new_n35577_, new_n35382_, new_n35378_ );
xor  ( new_n35578_, new_n35577_, new_n35388_ );
or   ( new_n35579_, new_n35578_, new_n35576_ );
nand ( new_n35580_, new_n35578_, new_n35576_ );
xor  ( new_n35581_, new_n35373_, new_n35369_ );
nand ( new_n35582_, new_n35581_, new_n35580_ );
and  ( new_n35583_, new_n35582_, new_n35579_ );
nor  ( new_n35584_, new_n35583_, new_n35574_ );
nand ( new_n35585_, new_n35583_, new_n35574_ );
xnor ( new_n35586_, new_n35421_, new_n35417_ );
xor  ( new_n35587_, new_n35586_, new_n35427_ );
xnor ( new_n35588_, new_n35405_, new_n35399_ );
xor  ( new_n35589_, new_n35588_, new_n35411_ );
nor  ( new_n35590_, new_n35589_, new_n35587_ );
nand ( new_n35591_, new_n35589_, new_n35587_ );
xor  ( new_n35592_, new_n35439_, new_n35435_ );
xor  ( new_n35593_, new_n35592_, new_n35445_ );
and  ( new_n35594_, new_n35593_, new_n35591_ );
or   ( new_n35595_, new_n35594_, new_n35590_ );
and  ( new_n35596_, new_n35595_, new_n35585_ );
or   ( new_n35597_, new_n35596_, new_n35584_ );
or   ( new_n35598_, new_n6173_, new_n23895_ );
or   ( new_n35599_, new_n6175_, new_n23733_ );
and  ( new_n35600_, new_n35599_, new_n35598_ );
xor  ( new_n35601_, new_n35600_, new_n5597_ );
or   ( new_n35602_, new_n5604_, new_n24227_ );
or   ( new_n35603_, new_n5606_, new_n24006_ );
and  ( new_n35604_, new_n35603_, new_n35602_ );
xor  ( new_n35605_, new_n35604_, new_n5206_ );
or   ( new_n35606_, new_n35605_, new_n35601_ );
and  ( new_n35607_, new_n35605_, new_n35601_ );
or   ( new_n35608_, new_n5207_, new_n24543_ );
or   ( new_n35609_, new_n5209_, new_n24418_ );
and  ( new_n35610_, new_n35609_, new_n35608_ );
xor  ( new_n35611_, new_n35610_, new_n4708_ );
or   ( new_n35612_, new_n35611_, new_n35607_ );
and  ( new_n35613_, new_n35612_, new_n35606_ );
or   ( new_n35614_, new_n4709_, new_n24925_ );
or   ( new_n35615_, new_n4711_, new_n24927_ );
and  ( new_n35616_, new_n35615_, new_n35614_ );
xor  ( new_n35617_, new_n35616_, new_n4295_ );
or   ( new_n35618_, new_n4302_, new_n25288_ );
or   ( new_n35619_, new_n4304_, new_n25048_ );
and  ( new_n35620_, new_n35619_, new_n35618_ );
xor  ( new_n35621_, new_n35620_, new_n3895_ );
or   ( new_n35622_, new_n35621_, new_n35617_ );
and  ( new_n35623_, new_n35621_, new_n35617_ );
or   ( new_n35624_, new_n3896_, new_n25813_ );
or   ( new_n35625_, new_n3898_, new_n25486_ );
and  ( new_n35626_, new_n35625_, new_n35624_ );
xor  ( new_n35627_, new_n35626_, new_n3460_ );
or   ( new_n35628_, new_n35627_, new_n35623_ );
and  ( new_n35629_, new_n35628_, new_n35622_ );
or   ( new_n35630_, new_n35629_, new_n35613_ );
and  ( new_n35631_, new_n35629_, new_n35613_ );
or   ( new_n35632_, new_n3461_, new_n26063_ );
or   ( new_n35633_, new_n3463_, new_n26196_ );
and  ( new_n35634_, new_n35633_, new_n35632_ );
xor  ( new_n35635_, new_n35634_, new_n3116_ );
or   ( new_n35636_, new_n3117_, new_n26620_ );
or   ( new_n35637_, new_n3119_, new_n26372_ );
and  ( new_n35638_, new_n35637_, new_n35636_ );
xor  ( new_n35639_, new_n35638_, new_n2800_ );
or   ( new_n35640_, new_n35639_, new_n35635_ );
and  ( new_n35641_, new_n35639_, new_n35635_ );
or   ( new_n35642_, new_n2807_, new_n27085_ );
or   ( new_n35643_, new_n2809_, new_n26762_ );
and  ( new_n35644_, new_n35643_, new_n35642_ );
xor  ( new_n35645_, new_n35644_, new_n2424_ );
or   ( new_n35646_, new_n35645_, new_n35641_ );
and  ( new_n35647_, new_n35646_, new_n35640_ );
or   ( new_n35648_, new_n35647_, new_n35631_ );
and  ( new_n35649_, new_n35648_, new_n35630_ );
or   ( new_n35650_, new_n7732_, new_n22973_ );
or   ( new_n35651_, new_n7734_, new_n22975_ );
and  ( new_n35652_, new_n35651_, new_n35650_ );
xor  ( new_n35653_, new_n35652_, new_n7177_ );
or   ( new_n35654_, new_n7184_, new_n23252_ );
or   ( new_n35655_, new_n7186_, new_n23166_ );
and  ( new_n35656_, new_n35655_, new_n35654_ );
xor  ( new_n35657_, new_n35656_, new_n6638_ );
nor  ( new_n35658_, new_n35657_, new_n35653_ );
and  ( new_n35659_, new_n35657_, new_n35653_ );
or   ( new_n35660_, new_n6645_, new_n23554_ );
or   ( new_n35661_, new_n6647_, new_n23370_ );
and  ( new_n35662_, new_n35661_, new_n35660_ );
xor  ( new_n35663_, new_n35662_, new_n6166_ );
nor  ( new_n35664_, new_n35663_, new_n35659_ );
nor  ( new_n35665_, new_n35664_, new_n35658_ );
or   ( new_n35666_, new_n10059_, new_n22129_ );
or   ( new_n35667_, new_n10061_, new_n22098_ );
and  ( new_n35668_, new_n35667_, new_n35666_ );
xor  ( new_n35669_, new_n35668_, new_n9421_ );
and  ( new_n35670_, RIbb31c08_142, RIbb2d888_64 );
or   ( new_n35671_, new_n21847_, RIbb2d888_64 );
and  ( new_n35672_, new_n35671_, RIbb2d900_63 );
or   ( new_n35673_, new_n35672_, new_n35670_ );
or   ( new_n35674_, new_n10770_, new_n21840_ );
and  ( new_n35675_, new_n35674_, new_n35673_ );
nor  ( new_n35676_, new_n35675_, new_n35669_ );
and  ( new_n35677_, new_n35675_, new_n35669_ );
nor  ( new_n35678_, new_n35677_, new_n402_ );
nor  ( new_n35679_, new_n35678_, new_n35676_ );
or   ( new_n35680_, new_n9422_, new_n22304_ );
or   ( new_n35681_, new_n9424_, new_n22207_ );
and  ( new_n35682_, new_n35681_, new_n35680_ );
xor  ( new_n35683_, new_n35682_, new_n8873_ );
or   ( new_n35684_, new_n8874_, new_n22590_ );
or   ( new_n35685_, new_n8876_, new_n22423_ );
and  ( new_n35686_, new_n35685_, new_n35684_ );
xor  ( new_n35687_, new_n35686_, new_n8257_ );
or   ( new_n35688_, new_n35687_, new_n35683_ );
and  ( new_n35689_, new_n35687_, new_n35683_ );
or   ( new_n35690_, new_n8264_, new_n22829_ );
or   ( new_n35691_, new_n8266_, new_n22641_ );
and  ( new_n35692_, new_n35691_, new_n35690_ );
xor  ( new_n35693_, new_n35692_, new_n7725_ );
or   ( new_n35694_, new_n35693_, new_n35689_ );
and  ( new_n35695_, new_n35694_, new_n35688_ );
and  ( new_n35696_, new_n35695_, new_n35679_ );
or   ( new_n35697_, new_n35696_, new_n35665_ );
or   ( new_n35698_, new_n35695_, new_n35679_ );
and  ( new_n35699_, new_n35698_, new_n35697_ );
or   ( new_n35700_, new_n35699_, new_n35649_ );
and  ( new_n35701_, new_n35699_, new_n35649_ );
or   ( new_n35702_, new_n1593_, new_n29261_ );
or   ( new_n35703_, new_n1595_, new_n29263_ );
and  ( new_n35704_, new_n35703_, new_n35702_ );
xor  ( new_n35705_, new_n35704_, new_n1358_ );
or   ( new_n35706_, new_n1364_, new_n29619_ );
or   ( new_n35707_, new_n1366_, new_n29474_ );
and  ( new_n35708_, new_n35707_, new_n35706_ );
xor  ( new_n35709_, new_n35708_, new_n1129_ );
nor  ( new_n35710_, new_n35709_, new_n35705_ );
and  ( new_n35711_, new_n35709_, new_n35705_ );
or   ( new_n35712_, new_n1135_, new_n30227_ );
or   ( new_n35713_, new_n1137_, new_n30120_ );
and  ( new_n35714_, new_n35713_, new_n35712_ );
xor  ( new_n35715_, new_n35714_, new_n896_ );
nor  ( new_n35716_, new_n35715_, new_n35711_ );
nor  ( new_n35717_, new_n35716_, new_n35710_ );
or   ( new_n35718_, new_n2425_, new_n27602_ );
or   ( new_n35719_, new_n2427_, new_n27396_ );
and  ( new_n35720_, new_n35719_, new_n35718_ );
xor  ( new_n35721_, new_n35720_, new_n2121_ );
or   ( new_n35722_, new_n2122_, new_n28108_ );
or   ( new_n35723_, new_n2124_, new_n27763_ );
and  ( new_n35724_, new_n35723_, new_n35722_ );
xor  ( new_n35725_, new_n35724_, new_n1843_ );
or   ( new_n35726_, new_n35725_, new_n35721_ );
and  ( new_n35727_, new_n35725_, new_n35721_ );
or   ( new_n35728_, new_n1844_, new_n28531_ );
or   ( new_n35729_, new_n1846_, new_n28314_ );
and  ( new_n35730_, new_n35729_, new_n35728_ );
xor  ( new_n35731_, new_n35730_, new_n1586_ );
or   ( new_n35732_, new_n35731_, new_n35727_ );
and  ( new_n35733_, new_n35732_, new_n35726_ );
and  ( new_n35734_, new_n35733_, new_n35717_ );
or   ( new_n35735_, new_n35733_, new_n35717_ );
or   ( new_n35736_, new_n897_, new_n30798_ );
or   ( new_n35737_, new_n899_, new_n30800_ );
and  ( new_n35738_, new_n35737_, new_n35736_ );
xor  ( new_n35739_, new_n35738_, new_n748_ );
or   ( new_n35740_, new_n755_, new_n31654_ );
or   ( new_n35741_, new_n757_, new_n31333_ );
and  ( new_n35742_, new_n35741_, new_n35740_ );
xor  ( new_n35743_, new_n35742_, new_n523_ );
and  ( new_n35744_, new_n35743_, new_n35739_ );
or   ( new_n35745_, new_n35743_, new_n35739_ );
and  ( new_n35746_, new_n454_, RIbb33378_192 );
nor  ( new_n35747_, new_n35746_, new_n403_ );
and  ( new_n35748_, new_n35746_, new_n400_ );
or   ( new_n35749_, new_n35748_, new_n35747_ );
and  ( new_n35750_, new_n35749_, new_n35745_ );
or   ( new_n35751_, new_n35750_, new_n35744_ );
and  ( new_n35752_, new_n35751_, new_n35735_ );
or   ( new_n35753_, new_n35752_, new_n35734_ );
or   ( new_n35754_, new_n35753_, new_n35701_ );
and  ( new_n35755_, new_n35754_, new_n35700_ );
or   ( new_n35756_, new_n35755_, new_n35597_ );
and  ( new_n35757_, new_n35755_, new_n35597_ );
xor  ( new_n35758_, new_n35134_, new_n35128_ );
xor  ( new_n35759_, new_n35758_, new_n327_ );
xnor ( new_n35760_, new_n35470_, new_n35468_ );
xor  ( new_n35761_, new_n35760_, new_n35474_ );
and  ( new_n35762_, new_n35761_, new_n35759_ );
or   ( new_n35763_, new_n35761_, new_n35759_ );
xor  ( new_n35764_, new_n35482_, new_n35480_ );
xnor ( new_n35765_, new_n35764_, new_n35486_ );
and  ( new_n35766_, new_n35765_, new_n35763_ );
or   ( new_n35767_, new_n35766_, new_n35762_ );
or   ( new_n35768_, new_n35767_, new_n35757_ );
and  ( new_n35769_, new_n35768_, new_n35756_ );
and  ( new_n35770_, new_n35769_, new_n35564_ );
nor  ( new_n35771_, new_n35769_, new_n35564_ );
xor  ( new_n35772_, new_n35291_, new_n35289_ );
xor  ( new_n35773_, new_n35772_, new_n35295_ );
xnor ( new_n35774_, new_n35279_, new_n35277_ );
xor  ( new_n35775_, new_n35774_, new_n35283_ );
and  ( new_n35776_, new_n35775_, new_n35773_ );
nor  ( new_n35777_, new_n35775_, new_n35773_ );
xor  ( new_n35778_, new_n35329_, new_n35313_ );
xor  ( new_n35779_, new_n35778_, new_n35347_ );
xor  ( new_n35780_, new_n35390_, new_n35374_ );
xor  ( new_n35781_, new_n35780_, new_n35365_ );
and  ( new_n35782_, new_n35781_, new_n35779_ );
nor  ( new_n35783_, new_n35781_, new_n35779_ );
xor  ( new_n35784_, new_n35460_, new_n35458_ );
xnor ( new_n35785_, new_n35784_, new_n35464_ );
not  ( new_n35786_, new_n35785_ );
nor  ( new_n35787_, new_n35786_, new_n35783_ );
nor  ( new_n35788_, new_n35787_, new_n35782_ );
nor  ( new_n35789_, new_n35788_, new_n35777_ );
nor  ( new_n35790_, new_n35789_, new_n35776_ );
nor  ( new_n35791_, new_n35790_, new_n35771_ );
nor  ( new_n35792_, new_n35791_, new_n35770_ );
or   ( new_n35793_, new_n35792_, new_n35558_ );
and  ( new_n35794_, new_n35793_, new_n35557_ );
nor  ( new_n35795_, new_n35794_, new_n35544_ );
nand ( new_n35796_, new_n35794_, new_n35544_ );
xor  ( new_n35797_, new_n35044_, new_n35034_ );
xnor ( new_n35798_, new_n35797_, new_n35252_ );
and  ( new_n35799_, new_n35798_, new_n35796_ );
or   ( new_n35800_, new_n35799_, new_n35795_ );
xnor ( new_n35801_, new_n35527_, new_n35525_ );
xor  ( new_n35802_, new_n35801_, new_n35531_ );
and  ( new_n35803_, new_n35802_, new_n35800_ );
xor  ( new_n35804_, new_n35533_, new_n35270_ );
and  ( new_n35805_, new_n35804_, new_n35803_ );
xor  ( new_n35806_, new_n35794_, new_n35544_ );
xnor ( new_n35807_, new_n35806_, new_n35798_ );
xor  ( new_n35808_, new_n35510_, new_n35508_ );
xor  ( new_n35809_, new_n35808_, new_n35522_ );
nor  ( new_n35810_, new_n35809_, new_n35807_ );
xor  ( new_n35811_, new_n35802_, new_n35800_ );
and  ( new_n35812_, new_n35811_, new_n35810_ );
xnor ( new_n35813_, new_n35809_, new_n35807_ );
xor  ( new_n35814_, new_n35629_, new_n35613_ );
xor  ( new_n35815_, new_n35814_, new_n35647_ );
xor  ( new_n35816_, new_n35695_, new_n35679_ );
xor  ( new_n35817_, new_n35816_, new_n35665_ );
nor  ( new_n35818_, new_n35817_, new_n35815_ );
nand ( new_n35819_, new_n35817_, new_n35815_ );
xnor ( new_n35820_, new_n35733_, new_n35717_ );
xor  ( new_n35821_, new_n35820_, new_n35751_ );
and  ( new_n35822_, new_n35821_, new_n35819_ );
or   ( new_n35823_, new_n35822_, new_n35818_ );
xnor ( new_n35824_, new_n35429_, new_n35413_ );
xor  ( new_n35825_, new_n35824_, new_n35447_ );
nor  ( new_n35826_, new_n35825_, new_n35823_ );
and  ( new_n35827_, new_n35825_, new_n35823_ );
xor  ( new_n35828_, new_n35781_, new_n35779_ );
xor  ( new_n35829_, new_n35828_, new_n35785_ );
not  ( new_n35830_, new_n35829_ );
nor  ( new_n35831_, new_n35830_, new_n35827_ );
nor  ( new_n35832_, new_n35831_, new_n35826_ );
xor  ( new_n35833_, new_n35589_, new_n35587_ );
xor  ( new_n35834_, new_n35833_, new_n35593_ );
xnor ( new_n35835_, new_n35568_, new_n35566_ );
xor  ( new_n35836_, new_n35835_, new_n35572_ );
or   ( new_n35837_, new_n35836_, new_n35834_ );
and  ( new_n35838_, new_n35836_, new_n35834_ );
xor  ( new_n35839_, new_n35578_, new_n35576_ );
xor  ( new_n35840_, new_n35839_, new_n35581_ );
or   ( new_n35841_, new_n35840_, new_n35838_ );
and  ( new_n35842_, new_n35841_, new_n35837_ );
or   ( new_n35843_, new_n10059_, new_n22207_ );
or   ( new_n35844_, new_n10061_, new_n22129_ );
and  ( new_n35845_, new_n35844_, new_n35843_ );
xor  ( new_n35846_, new_n35845_, new_n9421_ );
and  ( new_n35847_, RIbb31c80_143, RIbb2d888_64 );
or   ( new_n35848_, new_n22098_, RIbb2d888_64 );
and  ( new_n35849_, new_n35848_, RIbb2d900_63 );
or   ( new_n35850_, new_n35849_, new_n35847_ );
or   ( new_n35851_, new_n10770_, new_n21847_ );
and  ( new_n35852_, new_n35851_, new_n35850_ );
or   ( new_n35853_, new_n35852_, new_n35846_ );
and  ( new_n35854_, new_n35852_, new_n35846_ );
or   ( new_n35855_, new_n9422_, new_n22423_ );
or   ( new_n35856_, new_n9424_, new_n22304_ );
and  ( new_n35857_, new_n35856_, new_n35855_ );
xor  ( new_n35858_, new_n35857_, new_n8873_ );
or   ( new_n35859_, new_n35858_, new_n35854_ );
and  ( new_n35860_, new_n35859_, new_n35853_ );
or   ( new_n35861_, new_n7184_, new_n23370_ );
or   ( new_n35862_, new_n7186_, new_n23252_ );
and  ( new_n35863_, new_n35862_, new_n35861_ );
xor  ( new_n35864_, new_n35863_, new_n6638_ );
or   ( new_n35865_, new_n6645_, new_n23733_ );
or   ( new_n35866_, new_n6647_, new_n23554_ );
and  ( new_n35867_, new_n35866_, new_n35865_ );
xor  ( new_n35868_, new_n35867_, new_n6166_ );
or   ( new_n35869_, new_n35868_, new_n35864_ );
and  ( new_n35870_, new_n35868_, new_n35864_ );
or   ( new_n35871_, new_n6173_, new_n24006_ );
or   ( new_n35872_, new_n6175_, new_n23895_ );
and  ( new_n35873_, new_n35872_, new_n35871_ );
xor  ( new_n35874_, new_n35873_, new_n5597_ );
or   ( new_n35875_, new_n35874_, new_n35870_ );
and  ( new_n35876_, new_n35875_, new_n35869_ );
or   ( new_n35877_, new_n35876_, new_n35860_ );
and  ( new_n35878_, new_n35876_, new_n35860_ );
or   ( new_n35879_, new_n8874_, new_n22641_ );
or   ( new_n35880_, new_n8876_, new_n22590_ );
and  ( new_n35881_, new_n35880_, new_n35879_ );
xor  ( new_n35882_, new_n35881_, new_n8257_ );
or   ( new_n35883_, new_n8264_, new_n22975_ );
or   ( new_n35884_, new_n8266_, new_n22829_ );
and  ( new_n35885_, new_n35884_, new_n35883_ );
xor  ( new_n35886_, new_n35885_, new_n7725_ );
nor  ( new_n35887_, new_n35886_, new_n35882_ );
and  ( new_n35888_, new_n35886_, new_n35882_ );
or   ( new_n35889_, new_n7732_, new_n23166_ );
or   ( new_n35890_, new_n7734_, new_n22973_ );
and  ( new_n35891_, new_n35890_, new_n35889_ );
xor  ( new_n35892_, new_n35891_, new_n7177_ );
nor  ( new_n35893_, new_n35892_, new_n35888_ );
nor  ( new_n35894_, new_n35893_, new_n35887_ );
or   ( new_n35895_, new_n35894_, new_n35878_ );
and  ( new_n35896_, new_n35895_, new_n35877_ );
xor  ( new_n35897_, new_n35743_, new_n35739_ );
xor  ( new_n35898_, new_n35897_, new_n35749_ );
or   ( new_n35899_, new_n1364_, new_n30120_ );
or   ( new_n35900_, new_n1366_, new_n29619_ );
and  ( new_n35901_, new_n35900_, new_n35899_ );
xor  ( new_n35902_, new_n35901_, new_n1129_ );
or   ( new_n35903_, new_n1135_, new_n30800_ );
or   ( new_n35904_, new_n1137_, new_n30227_ );
and  ( new_n35905_, new_n35904_, new_n35903_ );
xor  ( new_n35906_, new_n35905_, new_n896_ );
or   ( new_n35907_, new_n35906_, new_n35902_ );
and  ( new_n35908_, new_n35906_, new_n35902_ );
or   ( new_n35909_, new_n897_, new_n31333_ );
or   ( new_n35910_, new_n899_, new_n30798_ );
and  ( new_n35911_, new_n35910_, new_n35909_ );
xor  ( new_n35912_, new_n35911_, new_n748_ );
or   ( new_n35913_, new_n35912_, new_n35908_ );
and  ( new_n35914_, new_n35913_, new_n35907_ );
or   ( new_n35915_, new_n35914_, new_n35898_ );
and  ( new_n35916_, new_n35914_, new_n35898_ );
or   ( new_n35917_, new_n2122_, new_n28314_ );
or   ( new_n35918_, new_n2124_, new_n28108_ );
and  ( new_n35919_, new_n35918_, new_n35917_ );
xor  ( new_n35920_, new_n35919_, new_n1843_ );
or   ( new_n35921_, new_n1844_, new_n29263_ );
or   ( new_n35922_, new_n1846_, new_n28531_ );
and  ( new_n35923_, new_n35922_, new_n35921_ );
xor  ( new_n35924_, new_n35923_, new_n1586_ );
nor  ( new_n35925_, new_n35924_, new_n35920_ );
and  ( new_n35926_, new_n35924_, new_n35920_ );
or   ( new_n35927_, new_n1593_, new_n29474_ );
or   ( new_n35928_, new_n1595_, new_n29261_ );
and  ( new_n35929_, new_n35928_, new_n35927_ );
xor  ( new_n35930_, new_n35929_, new_n1358_ );
nor  ( new_n35931_, new_n35930_, new_n35926_ );
nor  ( new_n35932_, new_n35931_, new_n35925_ );
or   ( new_n35933_, new_n35932_, new_n35916_ );
and  ( new_n35934_, new_n35933_, new_n35915_ );
or   ( new_n35935_, new_n35934_, new_n35896_ );
and  ( new_n35936_, new_n35934_, new_n35896_ );
or   ( new_n35937_, new_n5604_, new_n24418_ );
or   ( new_n35938_, new_n5606_, new_n24227_ );
and  ( new_n35939_, new_n35938_, new_n35937_ );
xor  ( new_n35940_, new_n35939_, new_n5206_ );
or   ( new_n35941_, new_n5207_, new_n24927_ );
or   ( new_n35942_, new_n5209_, new_n24543_ );
and  ( new_n35943_, new_n35942_, new_n35941_ );
xor  ( new_n35944_, new_n35943_, new_n4708_ );
or   ( new_n35945_, new_n35944_, new_n35940_ );
and  ( new_n35946_, new_n35944_, new_n35940_ );
or   ( new_n35947_, new_n4709_, new_n25048_ );
or   ( new_n35948_, new_n4711_, new_n24925_ );
and  ( new_n35949_, new_n35948_, new_n35947_ );
xor  ( new_n35950_, new_n35949_, new_n4295_ );
or   ( new_n35951_, new_n35950_, new_n35946_ );
and  ( new_n35952_, new_n35951_, new_n35945_ );
or   ( new_n35953_, new_n4302_, new_n25486_ );
or   ( new_n35954_, new_n4304_, new_n25288_ );
and  ( new_n35955_, new_n35954_, new_n35953_ );
xor  ( new_n35956_, new_n35955_, new_n3895_ );
or   ( new_n35957_, new_n3896_, new_n26196_ );
or   ( new_n35958_, new_n3898_, new_n25813_ );
and  ( new_n35959_, new_n35958_, new_n35957_ );
xor  ( new_n35960_, new_n35959_, new_n3460_ );
or   ( new_n35961_, new_n35960_, new_n35956_ );
and  ( new_n35962_, new_n35960_, new_n35956_ );
or   ( new_n35963_, new_n3461_, new_n26372_ );
or   ( new_n35964_, new_n3463_, new_n26063_ );
and  ( new_n35965_, new_n35964_, new_n35963_ );
xor  ( new_n35966_, new_n35965_, new_n3116_ );
or   ( new_n35967_, new_n35966_, new_n35962_ );
and  ( new_n35968_, new_n35967_, new_n35961_ );
nor  ( new_n35969_, new_n35968_, new_n35952_ );
and  ( new_n35970_, new_n35968_, new_n35952_ );
or   ( new_n35971_, new_n3117_, new_n26762_ );
or   ( new_n35972_, new_n3119_, new_n26620_ );
and  ( new_n35973_, new_n35972_, new_n35971_ );
xor  ( new_n35974_, new_n35973_, new_n2800_ );
or   ( new_n35975_, new_n2807_, new_n27396_ );
or   ( new_n35976_, new_n2809_, new_n27085_ );
and  ( new_n35977_, new_n35976_, new_n35975_ );
xor  ( new_n35978_, new_n35977_, new_n2424_ );
nor  ( new_n35979_, new_n35978_, new_n35974_ );
and  ( new_n35980_, new_n35978_, new_n35974_ );
or   ( new_n35981_, new_n2425_, new_n27763_ );
or   ( new_n35982_, new_n2427_, new_n27602_ );
and  ( new_n35983_, new_n35982_, new_n35981_ );
xor  ( new_n35984_, new_n35983_, new_n2121_ );
nor  ( new_n35985_, new_n35984_, new_n35980_ );
nor  ( new_n35986_, new_n35985_, new_n35979_ );
nor  ( new_n35987_, new_n35986_, new_n35970_ );
nor  ( new_n35988_, new_n35987_, new_n35969_ );
or   ( new_n35989_, new_n35988_, new_n35936_ );
and  ( new_n35990_, new_n35989_, new_n35935_ );
and  ( new_n35991_, new_n35990_, new_n35842_ );
nor  ( new_n35992_, new_n35990_, new_n35842_ );
xor  ( new_n35993_, new_n35687_, new_n35683_ );
xnor ( new_n35994_, new_n35993_, new_n35693_ );
xor  ( new_n35995_, new_n35675_, new_n35669_ );
xor  ( new_n35996_, new_n35995_, new_n403_ );
or   ( new_n35997_, new_n35996_, new_n35994_ );
xnor ( new_n35998_, new_n35725_, new_n35721_ );
xor  ( new_n35999_, new_n35998_, new_n35731_ );
xnor ( new_n36000_, new_n35639_, new_n35635_ );
xor  ( new_n36001_, new_n36000_, new_n35645_ );
or   ( new_n36002_, new_n36001_, new_n35999_ );
and  ( new_n36003_, new_n36001_, new_n35999_ );
xor  ( new_n36004_, new_n35709_, new_n35705_ );
xnor ( new_n36005_, new_n36004_, new_n35715_ );
or   ( new_n36006_, new_n36005_, new_n36003_ );
and  ( new_n36007_, new_n36006_, new_n36002_ );
nor  ( new_n36008_, new_n36007_, new_n35997_ );
and  ( new_n36009_, new_n36007_, new_n35997_ );
xnor ( new_n36010_, new_n35621_, new_n35617_ );
xor  ( new_n36011_, new_n36010_, new_n35627_ );
xnor ( new_n36012_, new_n35605_, new_n35601_ );
xor  ( new_n36013_, new_n36012_, new_n35611_ );
nor  ( new_n36014_, new_n36013_, new_n36011_ );
and  ( new_n36015_, new_n36013_, new_n36011_ );
xor  ( new_n36016_, new_n35657_, new_n35653_ );
xnor ( new_n36017_, new_n36016_, new_n35663_ );
nor  ( new_n36018_, new_n36017_, new_n36015_ );
nor  ( new_n36019_, new_n36018_, new_n36014_ );
nor  ( new_n36020_, new_n36019_, new_n36009_ );
nor  ( new_n36021_, new_n36020_, new_n36008_ );
nor  ( new_n36022_, new_n36021_, new_n35992_ );
nor  ( new_n36023_, new_n36022_, new_n35991_ );
and  ( new_n36024_, new_n36023_, new_n35832_ );
xor  ( new_n36025_, new_n35699_, new_n35649_ );
xor  ( new_n36026_, new_n36025_, new_n35753_ );
xor  ( new_n36027_, new_n35583_, new_n35574_ );
xor  ( new_n36028_, new_n36027_, new_n35595_ );
and  ( new_n36029_, new_n36028_, new_n36026_ );
nor  ( new_n36030_, new_n36028_, new_n36026_ );
xor  ( new_n36031_, new_n35761_, new_n35759_ );
xnor ( new_n36032_, new_n36031_, new_n35765_ );
nor  ( new_n36033_, new_n36032_, new_n36030_ );
nor  ( new_n36034_, new_n36033_, new_n36029_ );
nor  ( new_n36035_, new_n36034_, new_n36024_ );
nor  ( new_n36036_, new_n36023_, new_n35832_ );
nor  ( new_n36037_, new_n36036_, new_n36035_ );
xor  ( new_n36038_, new_n35548_, new_n35546_ );
xor  ( new_n36039_, new_n36038_, new_n35552_ );
and  ( new_n36040_, new_n36039_, new_n36037_ );
xor  ( new_n36041_, new_n35755_, new_n35597_ );
xor  ( new_n36042_, new_n36041_, new_n35767_ );
xnor ( new_n36043_, new_n35775_, new_n35773_ );
xor  ( new_n36044_, new_n36043_, new_n35788_ );
and  ( new_n36045_, new_n36044_, new_n36042_ );
nor  ( new_n36046_, new_n36044_, new_n36042_ );
xor  ( new_n36047_, new_n35563_, new_n35561_ );
not  ( new_n36048_, new_n36047_ );
nor  ( new_n36049_, new_n36048_, new_n36046_ );
nor  ( new_n36050_, new_n36049_, new_n36045_ );
nor  ( new_n36051_, new_n36050_, new_n36040_ );
nor  ( new_n36052_, new_n36039_, new_n36037_ );
or   ( new_n36053_, new_n36052_, new_n36051_ );
xnor ( new_n36054_, new_n35556_, new_n35554_ );
xor  ( new_n36055_, new_n36054_, new_n35792_ );
nand ( new_n36056_, new_n36055_, new_n36053_ );
nor  ( new_n36057_, new_n36055_, new_n36053_ );
xnor ( new_n36058_, new_n35543_, new_n35541_ );
or   ( new_n36059_, new_n36058_, new_n36057_ );
and  ( new_n36060_, new_n36059_, new_n36056_ );
nor  ( new_n36061_, new_n36060_, new_n35813_ );
xor  ( new_n36062_, new_n36055_, new_n36053_ );
xor  ( new_n36063_, new_n36062_, new_n36058_ );
xnor ( new_n36064_, new_n36023_, new_n35832_ );
nand ( new_n36065_, new_n36064_, new_n36034_ );
or   ( new_n36066_, new_n36034_, new_n36024_ );
or   ( new_n36067_, new_n36036_, new_n36066_ );
and  ( new_n36068_, new_n36067_, new_n36065_ );
xor  ( new_n36069_, new_n36028_, new_n36026_ );
xor  ( new_n36070_, new_n36069_, new_n36032_ );
xnor ( new_n36071_, new_n36001_, new_n35999_ );
xor  ( new_n36072_, new_n36071_, new_n36005_ );
xnor ( new_n36073_, new_n36013_, new_n36011_ );
xor  ( new_n36074_, new_n36073_, new_n36017_ );
or   ( new_n36075_, new_n36074_, new_n36072_ );
and  ( new_n36076_, new_n36074_, new_n36072_ );
xor  ( new_n36077_, new_n35996_, new_n35994_ );
or   ( new_n36078_, new_n36077_, new_n36076_ );
and  ( new_n36079_, new_n36078_, new_n36075_ );
or   ( new_n36080_, new_n6173_, new_n24227_ );
or   ( new_n36081_, new_n6175_, new_n24006_ );
and  ( new_n36082_, new_n36081_, new_n36080_ );
xor  ( new_n36083_, new_n36082_, new_n5597_ );
or   ( new_n36084_, new_n5604_, new_n24543_ );
or   ( new_n36085_, new_n5606_, new_n24418_ );
and  ( new_n36086_, new_n36085_, new_n36084_ );
xor  ( new_n36087_, new_n36086_, new_n5206_ );
or   ( new_n36088_, new_n36087_, new_n36083_ );
and  ( new_n36089_, new_n36087_, new_n36083_ );
or   ( new_n36090_, new_n5207_, new_n24925_ );
or   ( new_n36091_, new_n5209_, new_n24927_ );
and  ( new_n36092_, new_n36091_, new_n36090_ );
xor  ( new_n36093_, new_n36092_, new_n4708_ );
or   ( new_n36094_, new_n36093_, new_n36089_ );
and  ( new_n36095_, new_n36094_, new_n36088_ );
or   ( new_n36096_, new_n4709_, new_n25288_ );
or   ( new_n36097_, new_n4711_, new_n25048_ );
and  ( new_n36098_, new_n36097_, new_n36096_ );
xor  ( new_n36099_, new_n36098_, new_n4295_ );
or   ( new_n36100_, new_n4302_, new_n25813_ );
or   ( new_n36101_, new_n4304_, new_n25486_ );
and  ( new_n36102_, new_n36101_, new_n36100_ );
xor  ( new_n36103_, new_n36102_, new_n3895_ );
or   ( new_n36104_, new_n36103_, new_n36099_ );
and  ( new_n36105_, new_n36103_, new_n36099_ );
or   ( new_n36106_, new_n3896_, new_n26063_ );
or   ( new_n36107_, new_n3898_, new_n26196_ );
and  ( new_n36108_, new_n36107_, new_n36106_ );
xor  ( new_n36109_, new_n36108_, new_n3460_ );
or   ( new_n36110_, new_n36109_, new_n36105_ );
and  ( new_n36111_, new_n36110_, new_n36104_ );
or   ( new_n36112_, new_n36111_, new_n36095_ );
and  ( new_n36113_, new_n36111_, new_n36095_ );
or   ( new_n36114_, new_n3461_, new_n26620_ );
or   ( new_n36115_, new_n3463_, new_n26372_ );
and  ( new_n36116_, new_n36115_, new_n36114_ );
xor  ( new_n36117_, new_n36116_, new_n3116_ );
or   ( new_n36118_, new_n3117_, new_n27085_ );
or   ( new_n36119_, new_n3119_, new_n26762_ );
and  ( new_n36120_, new_n36119_, new_n36118_ );
xor  ( new_n36121_, new_n36120_, new_n2800_ );
nor  ( new_n36122_, new_n36121_, new_n36117_ );
and  ( new_n36123_, new_n36121_, new_n36117_ );
or   ( new_n36124_, new_n2807_, new_n27602_ );
or   ( new_n36125_, new_n2809_, new_n27396_ );
and  ( new_n36126_, new_n36125_, new_n36124_ );
xor  ( new_n36127_, new_n36126_, new_n2424_ );
nor  ( new_n36128_, new_n36127_, new_n36123_ );
nor  ( new_n36129_, new_n36128_, new_n36122_ );
or   ( new_n36130_, new_n36129_, new_n36113_ );
and  ( new_n36131_, new_n36130_, new_n36112_ );
or   ( new_n36132_, new_n755_, new_n31952_ );
or   ( new_n36133_, new_n757_, new_n31654_ );
and  ( new_n36134_, new_n36133_, new_n36132_ );
xor  ( new_n36135_, new_n36134_, new_n523_ );
or   ( new_n36136_, new_n2425_, new_n28108_ );
or   ( new_n36137_, new_n2427_, new_n27763_ );
and  ( new_n36138_, new_n36137_, new_n36136_ );
xor  ( new_n36139_, new_n36138_, new_n2121_ );
or   ( new_n36140_, new_n2122_, new_n28531_ );
or   ( new_n36141_, new_n2124_, new_n28314_ );
and  ( new_n36142_, new_n36141_, new_n36140_ );
xor  ( new_n36143_, new_n36142_, new_n1843_ );
or   ( new_n36144_, new_n36143_, new_n36139_ );
and  ( new_n36145_, new_n36143_, new_n36139_ );
or   ( new_n36146_, new_n1844_, new_n29261_ );
or   ( new_n36147_, new_n1846_, new_n29263_ );
and  ( new_n36148_, new_n36147_, new_n36146_ );
xor  ( new_n36149_, new_n36148_, new_n1586_ );
or   ( new_n36150_, new_n36149_, new_n36145_ );
and  ( new_n36151_, new_n36150_, new_n36144_ );
or   ( new_n36152_, new_n36151_, new_n36135_ );
and  ( new_n36153_, new_n36151_, new_n36135_ );
or   ( new_n36154_, new_n1593_, new_n29619_ );
or   ( new_n36155_, new_n1595_, new_n29474_ );
and  ( new_n36156_, new_n36155_, new_n36154_ );
xor  ( new_n36157_, new_n36156_, new_n1358_ );
or   ( new_n36158_, new_n1364_, new_n30227_ );
or   ( new_n36159_, new_n1366_, new_n30120_ );
and  ( new_n36160_, new_n36159_, new_n36158_ );
xor  ( new_n36161_, new_n36160_, new_n1129_ );
nor  ( new_n36162_, new_n36161_, new_n36157_ );
and  ( new_n36163_, new_n36161_, new_n36157_ );
or   ( new_n36164_, new_n1135_, new_n30798_ );
or   ( new_n36165_, new_n1137_, new_n30800_ );
and  ( new_n36166_, new_n36165_, new_n36164_ );
xor  ( new_n36167_, new_n36166_, new_n896_ );
nor  ( new_n36168_, new_n36167_, new_n36163_ );
nor  ( new_n36169_, new_n36168_, new_n36162_ );
or   ( new_n36170_, new_n36169_, new_n36153_ );
and  ( new_n36171_, new_n36170_, new_n36152_ );
or   ( new_n36172_, new_n36171_, new_n36131_ );
and  ( new_n36173_, new_n36171_, new_n36131_ );
or   ( new_n36174_, new_n7732_, new_n23252_ );
or   ( new_n36175_, new_n7734_, new_n23166_ );
and  ( new_n36176_, new_n36175_, new_n36174_ );
xor  ( new_n36177_, new_n36176_, new_n7177_ );
or   ( new_n36178_, new_n7184_, new_n23554_ );
or   ( new_n36179_, new_n7186_, new_n23370_ );
and  ( new_n36180_, new_n36179_, new_n36178_ );
xor  ( new_n36181_, new_n36180_, new_n6638_ );
nor  ( new_n36182_, new_n36181_, new_n36177_ );
and  ( new_n36183_, new_n36181_, new_n36177_ );
or   ( new_n36184_, new_n6645_, new_n23895_ );
or   ( new_n36185_, new_n6647_, new_n23733_ );
and  ( new_n36186_, new_n36185_, new_n36184_ );
xor  ( new_n36187_, new_n36186_, new_n6166_ );
nor  ( new_n36188_, new_n36187_, new_n36183_ );
nor  ( new_n36189_, new_n36188_, new_n36182_ );
or   ( new_n36190_, new_n10059_, new_n22304_ );
or   ( new_n36191_, new_n10061_, new_n22207_ );
and  ( new_n36192_, new_n36191_, new_n36190_ );
xor  ( new_n36193_, new_n36192_, new_n9421_ );
and  ( new_n36194_, RIbb31cf8_144, RIbb2d888_64 );
or   ( new_n36195_, new_n22129_, RIbb2d888_64 );
and  ( new_n36196_, new_n36195_, RIbb2d900_63 );
or   ( new_n36197_, new_n36196_, new_n36194_ );
or   ( new_n36198_, new_n10770_, new_n22098_ );
and  ( new_n36199_, new_n36198_, new_n36197_ );
nor  ( new_n36200_, new_n36199_, new_n36193_ );
and  ( new_n36201_, new_n36199_, new_n36193_ );
nor  ( new_n36202_, new_n36201_, new_n522_ );
nor  ( new_n36203_, new_n36202_, new_n36200_ );
or   ( new_n36204_, new_n9422_, new_n22590_ );
or   ( new_n36205_, new_n9424_, new_n22423_ );
and  ( new_n36206_, new_n36205_, new_n36204_ );
xor  ( new_n36207_, new_n36206_, new_n8873_ );
or   ( new_n36208_, new_n8874_, new_n22829_ );
or   ( new_n36209_, new_n8876_, new_n22641_ );
and  ( new_n36210_, new_n36209_, new_n36208_ );
xor  ( new_n36211_, new_n36210_, new_n8257_ );
nor  ( new_n36212_, new_n36211_, new_n36207_ );
and  ( new_n36213_, new_n36211_, new_n36207_ );
or   ( new_n36214_, new_n8264_, new_n22973_ );
or   ( new_n36215_, new_n8266_, new_n22975_ );
and  ( new_n36216_, new_n36215_, new_n36214_ );
xor  ( new_n36217_, new_n36216_, new_n7725_ );
nor  ( new_n36218_, new_n36217_, new_n36213_ );
nor  ( new_n36219_, new_n36218_, new_n36212_ );
and  ( new_n36220_, new_n36219_, new_n36203_ );
nor  ( new_n36221_, new_n36220_, new_n36189_ );
nor  ( new_n36222_, new_n36219_, new_n36203_ );
nor  ( new_n36223_, new_n36222_, new_n36221_ );
or   ( new_n36224_, new_n36223_, new_n36173_ );
and  ( new_n36225_, new_n36224_, new_n36172_ );
nand ( new_n36226_, new_n36225_, new_n36079_ );
nor  ( new_n36227_, new_n36225_, new_n36079_ );
xor  ( new_n36228_, new_n35852_, new_n35846_ );
xnor ( new_n36229_, new_n36228_, new_n35858_ );
xnor ( new_n36230_, new_n35886_, new_n35882_ );
xor  ( new_n36231_, new_n36230_, new_n35892_ );
or   ( new_n36232_, new_n36231_, new_n36229_ );
xnor ( new_n36233_, new_n35906_, new_n35902_ );
xor  ( new_n36234_, new_n36233_, new_n35912_ );
xnor ( new_n36235_, new_n35978_, new_n35974_ );
xor  ( new_n36236_, new_n36235_, new_n35984_ );
or   ( new_n36237_, new_n36236_, new_n36234_ );
and  ( new_n36238_, new_n36236_, new_n36234_ );
xor  ( new_n36239_, new_n35924_, new_n35920_ );
xnor ( new_n36240_, new_n36239_, new_n35930_ );
or   ( new_n36241_, new_n36240_, new_n36238_ );
and  ( new_n36242_, new_n36241_, new_n36237_ );
or   ( new_n36243_, new_n36242_, new_n36232_ );
and  ( new_n36244_, new_n36242_, new_n36232_ );
xnor ( new_n36245_, new_n35960_, new_n35956_ );
xor  ( new_n36246_, new_n36245_, new_n35966_ );
xnor ( new_n36247_, new_n35944_, new_n35940_ );
xor  ( new_n36248_, new_n36247_, new_n35950_ );
nor  ( new_n36249_, new_n36248_, new_n36246_ );
and  ( new_n36250_, new_n36248_, new_n36246_ );
xor  ( new_n36251_, new_n35868_, new_n35864_ );
xnor ( new_n36252_, new_n36251_, new_n35874_ );
nor  ( new_n36253_, new_n36252_, new_n36250_ );
nor  ( new_n36254_, new_n36253_, new_n36249_ );
or   ( new_n36255_, new_n36254_, new_n36244_ );
and  ( new_n36256_, new_n36255_, new_n36243_ );
or   ( new_n36257_, new_n36256_, new_n36227_ );
and  ( new_n36258_, new_n36257_, new_n36226_ );
nand ( new_n36259_, new_n36258_, new_n36070_ );
or   ( new_n36260_, new_n36258_, new_n36070_ );
xnor ( new_n36261_, new_n35836_, new_n35834_ );
xor  ( new_n36262_, new_n36261_, new_n35840_ );
xor  ( new_n36263_, new_n35817_, new_n35815_ );
xor  ( new_n36264_, new_n36263_, new_n35821_ );
nor  ( new_n36265_, new_n36264_, new_n36262_ );
and  ( new_n36266_, new_n36264_, new_n36262_ );
xnor ( new_n36267_, new_n35876_, new_n35860_ );
xor  ( new_n36268_, new_n36267_, new_n35894_ );
xnor ( new_n36269_, new_n35968_, new_n35952_ );
xor  ( new_n36270_, new_n36269_, new_n35986_ );
nor  ( new_n36271_, new_n36270_, new_n36268_ );
and  ( new_n36272_, new_n36270_, new_n36268_ );
xor  ( new_n36273_, new_n35914_, new_n35898_ );
xnor ( new_n36274_, new_n36273_, new_n35932_ );
nor  ( new_n36275_, new_n36274_, new_n36272_ );
nor  ( new_n36276_, new_n36275_, new_n36271_ );
nor  ( new_n36277_, new_n36276_, new_n36266_ );
nor  ( new_n36278_, new_n36277_, new_n36265_ );
nand ( new_n36279_, new_n36278_, new_n36260_ );
and  ( new_n36280_, new_n36279_, new_n36259_ );
and  ( new_n36281_, new_n36280_, new_n36068_ );
or   ( new_n36282_, new_n36280_, new_n36068_ );
xor  ( new_n36283_, new_n36044_, new_n36042_ );
xor  ( new_n36284_, new_n36283_, new_n36047_ );
and  ( new_n36285_, new_n36284_, new_n36282_ );
or   ( new_n36286_, new_n36285_, new_n36281_ );
xnor ( new_n36287_, new_n35769_, new_n35564_ );
xor  ( new_n36288_, new_n36287_, new_n35790_ );
nand ( new_n36289_, new_n36288_, new_n36286_ );
nor  ( new_n36290_, new_n36288_, new_n36286_ );
xor  ( new_n36291_, new_n36039_, new_n36037_ );
xor  ( new_n36292_, new_n36291_, new_n36050_ );
or   ( new_n36293_, new_n36292_, new_n36290_ );
and  ( new_n36294_, new_n36293_, new_n36289_ );
nor  ( new_n36295_, new_n36294_, new_n36063_ );
xor  ( new_n36296_, new_n36288_, new_n36286_ );
xor  ( new_n36297_, new_n36296_, new_n36292_ );
xor  ( new_n36298_, new_n35990_, new_n35842_ );
xnor ( new_n36299_, new_n36298_, new_n36021_ );
xor  ( new_n36300_, new_n36258_, new_n36070_ );
xnor ( new_n36301_, new_n36300_, new_n36278_ );
nand ( new_n36302_, new_n36301_, new_n36299_ );
xor  ( new_n36303_, new_n35825_, new_n35823_ );
xor  ( new_n36304_, new_n36303_, new_n35830_ );
xor  ( new_n36305_, new_n36225_, new_n36079_ );
xor  ( new_n36306_, new_n36305_, new_n36256_ );
xnor ( new_n36307_, new_n35934_, new_n35896_ );
xor  ( new_n36308_, new_n36307_, new_n35988_ );
or   ( new_n36309_, new_n36308_, new_n36306_ );
and  ( new_n36310_, new_n36308_, new_n36306_ );
xor  ( new_n36311_, new_n36264_, new_n36262_ );
xor  ( new_n36312_, new_n36311_, new_n36276_ );
or   ( new_n36313_, new_n36312_, new_n36310_ );
and  ( new_n36314_, new_n36313_, new_n36309_ );
or   ( new_n36315_, new_n36314_, new_n36304_ );
and  ( new_n36316_, new_n36314_, new_n36304_ );
xnor ( new_n36317_, new_n36111_, new_n36095_ );
xor  ( new_n36318_, new_n36317_, new_n36129_ );
xnor ( new_n36319_, new_n36151_, new_n36135_ );
xor  ( new_n36320_, new_n36319_, new_n36169_ );
nor  ( new_n36321_, new_n36320_, new_n36318_ );
nand ( new_n36322_, new_n36320_, new_n36318_ );
xnor ( new_n36323_, new_n36219_, new_n36203_ );
xnor ( new_n36324_, new_n36323_, new_n36189_ );
and  ( new_n36325_, new_n36324_, new_n36322_ );
or   ( new_n36326_, new_n36325_, new_n36321_ );
xnor ( new_n36327_, new_n36270_, new_n36268_ );
xor  ( new_n36328_, new_n36327_, new_n36274_ );
and  ( new_n36329_, new_n36328_, new_n36326_ );
nor  ( new_n36330_, new_n36328_, new_n36326_ );
xor  ( new_n36331_, new_n36074_, new_n36072_ );
xnor ( new_n36332_, new_n36331_, new_n36077_ );
nor  ( new_n36333_, new_n36332_, new_n36330_ );
or   ( new_n36334_, new_n36333_, new_n36329_ );
xnor ( new_n36335_, new_n36007_, new_n35997_ );
xor  ( new_n36336_, new_n36335_, new_n36019_ );
and  ( new_n36337_, new_n36336_, new_n36334_ );
nor  ( new_n36338_, new_n36336_, new_n36334_ );
not  ( new_n36339_, new_n36338_ );
and  ( new_n36340_, new_n660_, RIbb33378_192 );
or   ( new_n36341_, new_n36340_, new_n523_ );
nand ( new_n36342_, new_n36340_, new_n520_ );
and  ( new_n36343_, new_n36342_, new_n36341_ );
xnor ( new_n36344_, new_n36161_, new_n36157_ );
xor  ( new_n36345_, new_n36344_, new_n36167_ );
or   ( new_n36346_, new_n36345_, new_n36343_ );
and  ( new_n36347_, new_n36345_, new_n36343_ );
xor  ( new_n36348_, new_n36143_, new_n36139_ );
xnor ( new_n36349_, new_n36348_, new_n36149_ );
or   ( new_n36350_, new_n36349_, new_n36347_ );
and  ( new_n36351_, new_n36350_, new_n36346_ );
xnor ( new_n36352_, new_n36181_, new_n36177_ );
xor  ( new_n36353_, new_n36352_, new_n36187_ );
xnor ( new_n36354_, new_n36211_, new_n36207_ );
xor  ( new_n36355_, new_n36354_, new_n36217_ );
or   ( new_n36356_, new_n36355_, new_n36353_ );
and  ( new_n36357_, new_n36355_, new_n36353_ );
xor  ( new_n36358_, new_n36199_, new_n36193_ );
xor  ( new_n36359_, new_n36358_, new_n523_ );
or   ( new_n36360_, new_n36359_, new_n36357_ );
and  ( new_n36361_, new_n36360_, new_n36356_ );
nor  ( new_n36362_, new_n36361_, new_n36351_ );
and  ( new_n36363_, new_n36361_, new_n36351_ );
xnor ( new_n36364_, new_n36103_, new_n36099_ );
xor  ( new_n36365_, new_n36364_, new_n36109_ );
xnor ( new_n36366_, new_n36087_, new_n36083_ );
xor  ( new_n36367_, new_n36366_, new_n36093_ );
nor  ( new_n36368_, new_n36367_, new_n36365_ );
and  ( new_n36369_, new_n36367_, new_n36365_ );
xor  ( new_n36370_, new_n36121_, new_n36117_ );
xnor ( new_n36371_, new_n36370_, new_n36127_ );
nor  ( new_n36372_, new_n36371_, new_n36369_ );
nor  ( new_n36373_, new_n36372_, new_n36368_ );
nor  ( new_n36374_, new_n36373_, new_n36363_ );
or   ( new_n36375_, new_n36374_, new_n36362_ );
or   ( new_n36376_, new_n3117_, new_n27396_ );
or   ( new_n36377_, new_n3119_, new_n27085_ );
and  ( new_n36378_, new_n36377_, new_n36376_ );
xor  ( new_n36379_, new_n36378_, new_n2800_ );
or   ( new_n36380_, new_n2807_, new_n27763_ );
or   ( new_n36381_, new_n2809_, new_n27602_ );
and  ( new_n36382_, new_n36381_, new_n36380_ );
xor  ( new_n36383_, new_n36382_, new_n2424_ );
or   ( new_n36384_, new_n36383_, new_n36379_ );
and  ( new_n36385_, new_n36383_, new_n36379_ );
or   ( new_n36386_, new_n2425_, new_n28314_ );
or   ( new_n36387_, new_n2427_, new_n28108_ );
and  ( new_n36388_, new_n36387_, new_n36386_ );
xor  ( new_n36389_, new_n36388_, new_n2121_ );
or   ( new_n36390_, new_n36389_, new_n36385_ );
and  ( new_n36391_, new_n36390_, new_n36384_ );
or   ( new_n36392_, new_n4302_, new_n26196_ );
or   ( new_n36393_, new_n4304_, new_n25813_ );
and  ( new_n36394_, new_n36393_, new_n36392_ );
xor  ( new_n36395_, new_n36394_, new_n3895_ );
or   ( new_n36396_, new_n3896_, new_n26372_ );
or   ( new_n36397_, new_n3898_, new_n26063_ );
and  ( new_n36398_, new_n36397_, new_n36396_ );
xor  ( new_n36399_, new_n36398_, new_n3460_ );
or   ( new_n36400_, new_n36399_, new_n36395_ );
and  ( new_n36401_, new_n36399_, new_n36395_ );
or   ( new_n36402_, new_n3461_, new_n26762_ );
or   ( new_n36403_, new_n3463_, new_n26620_ );
and  ( new_n36404_, new_n36403_, new_n36402_ );
xor  ( new_n36405_, new_n36404_, new_n3116_ );
or   ( new_n36406_, new_n36405_, new_n36401_ );
and  ( new_n36407_, new_n36406_, new_n36400_ );
or   ( new_n36408_, new_n36407_, new_n36391_ );
and  ( new_n36409_, new_n36407_, new_n36391_ );
or   ( new_n36410_, new_n5604_, new_n24927_ );
or   ( new_n36411_, new_n5606_, new_n24543_ );
and  ( new_n36412_, new_n36411_, new_n36410_ );
xor  ( new_n36413_, new_n36412_, new_n5206_ );
or   ( new_n36414_, new_n5207_, new_n25048_ );
or   ( new_n36415_, new_n5209_, new_n24925_ );
and  ( new_n36416_, new_n36415_, new_n36414_ );
xor  ( new_n36417_, new_n36416_, new_n4708_ );
nor  ( new_n36418_, new_n36417_, new_n36413_ );
and  ( new_n36419_, new_n36417_, new_n36413_ );
or   ( new_n36420_, new_n4709_, new_n25486_ );
or   ( new_n36421_, new_n4711_, new_n25288_ );
and  ( new_n36422_, new_n36421_, new_n36420_ );
xor  ( new_n36423_, new_n36422_, new_n4295_ );
nor  ( new_n36424_, new_n36423_, new_n36419_ );
nor  ( new_n36425_, new_n36424_, new_n36418_ );
or   ( new_n36426_, new_n36425_, new_n36409_ );
and  ( new_n36427_, new_n36426_, new_n36408_ );
or   ( new_n36428_, new_n897_, new_n31654_ );
or   ( new_n36429_, new_n899_, new_n31333_ );
and  ( new_n36430_, new_n36429_, new_n36428_ );
xor  ( new_n36431_, new_n36430_, new_n748_ );
or   ( new_n36432_, new_n2122_, new_n29263_ );
or   ( new_n36433_, new_n2124_, new_n28531_ );
and  ( new_n36434_, new_n36433_, new_n36432_ );
xor  ( new_n36435_, new_n36434_, new_n1843_ );
or   ( new_n36436_, new_n1844_, new_n29474_ );
or   ( new_n36437_, new_n1846_, new_n29261_ );
and  ( new_n36438_, new_n36437_, new_n36436_ );
xor  ( new_n36439_, new_n36438_, new_n1586_ );
or   ( new_n36440_, new_n36439_, new_n36435_ );
and  ( new_n36441_, new_n36439_, new_n36435_ );
or   ( new_n36442_, new_n1593_, new_n30120_ );
or   ( new_n36443_, new_n1595_, new_n29619_ );
and  ( new_n36444_, new_n36443_, new_n36442_ );
xor  ( new_n36445_, new_n36444_, new_n1358_ );
or   ( new_n36446_, new_n36445_, new_n36441_ );
and  ( new_n36447_, new_n36446_, new_n36440_ );
or   ( new_n36448_, new_n36447_, new_n36431_ );
and  ( new_n36449_, new_n36447_, new_n36431_ );
or   ( new_n36450_, new_n1364_, new_n30800_ );
or   ( new_n36451_, new_n1366_, new_n30227_ );
and  ( new_n36452_, new_n36451_, new_n36450_ );
xor  ( new_n36453_, new_n36452_, new_n1129_ );
or   ( new_n36454_, new_n1135_, new_n31333_ );
or   ( new_n36455_, new_n1137_, new_n30798_ );
and  ( new_n36456_, new_n36455_, new_n36454_ );
xor  ( new_n36457_, new_n36456_, new_n896_ );
nor  ( new_n36458_, new_n36457_, new_n36453_ );
and  ( new_n36459_, new_n36457_, new_n36453_ );
or   ( new_n36460_, new_n897_, new_n31952_ );
or   ( new_n36461_, new_n899_, new_n31654_ );
and  ( new_n36462_, new_n36461_, new_n36460_ );
xor  ( new_n36463_, new_n36462_, new_n748_ );
nor  ( new_n36464_, new_n36463_, new_n36459_ );
nor  ( new_n36465_, new_n36464_, new_n36458_ );
or   ( new_n36466_, new_n36465_, new_n36449_ );
and  ( new_n36467_, new_n36466_, new_n36448_ );
or   ( new_n36468_, new_n36467_, new_n36427_ );
and  ( new_n36469_, new_n36467_, new_n36427_ );
or   ( new_n36470_, new_n8874_, new_n22975_ );
or   ( new_n36471_, new_n8876_, new_n22829_ );
and  ( new_n36472_, new_n36471_, new_n36470_ );
xor  ( new_n36473_, new_n36472_, new_n8257_ );
or   ( new_n36474_, new_n8264_, new_n23166_ );
or   ( new_n36475_, new_n8266_, new_n22973_ );
and  ( new_n36476_, new_n36475_, new_n36474_ );
xor  ( new_n36477_, new_n36476_, new_n7725_ );
or   ( new_n36478_, new_n36477_, new_n36473_ );
and  ( new_n36479_, new_n36477_, new_n36473_ );
or   ( new_n36480_, new_n7732_, new_n23370_ );
or   ( new_n36481_, new_n7734_, new_n23252_ );
and  ( new_n36482_, new_n36481_, new_n36480_ );
xor  ( new_n36483_, new_n36482_, new_n7177_ );
or   ( new_n36484_, new_n36483_, new_n36479_ );
and  ( new_n36485_, new_n36484_, new_n36478_ );
or   ( new_n36486_, new_n10059_, new_n22423_ );
or   ( new_n36487_, new_n10061_, new_n22304_ );
and  ( new_n36488_, new_n36487_, new_n36486_ );
xor  ( new_n36489_, new_n36488_, new_n9421_ );
and  ( new_n36490_, RIbb31d70_145, RIbb2d888_64 );
or   ( new_n36491_, new_n22207_, RIbb2d888_64 );
and  ( new_n36492_, new_n36491_, RIbb2d900_63 );
or   ( new_n36493_, new_n36492_, new_n36490_ );
or   ( new_n36494_, new_n10770_, new_n22129_ );
and  ( new_n36495_, new_n36494_, new_n36493_ );
or   ( new_n36496_, new_n36495_, new_n36489_ );
and  ( new_n36497_, new_n36495_, new_n36489_ );
or   ( new_n36498_, new_n9422_, new_n22641_ );
or   ( new_n36499_, new_n9424_, new_n22590_ );
and  ( new_n36500_, new_n36499_, new_n36498_ );
xor  ( new_n36501_, new_n36500_, new_n8873_ );
or   ( new_n36502_, new_n36501_, new_n36497_ );
and  ( new_n36503_, new_n36502_, new_n36496_ );
nor  ( new_n36504_, new_n36503_, new_n36485_ );
and  ( new_n36505_, new_n36503_, new_n36485_ );
or   ( new_n36506_, new_n7184_, new_n23733_ );
or   ( new_n36507_, new_n7186_, new_n23554_ );
and  ( new_n36508_, new_n36507_, new_n36506_ );
xor  ( new_n36509_, new_n36508_, new_n6638_ );
or   ( new_n36510_, new_n6645_, new_n24006_ );
or   ( new_n36511_, new_n6647_, new_n23895_ );
and  ( new_n36512_, new_n36511_, new_n36510_ );
xor  ( new_n36513_, new_n36512_, new_n6166_ );
nor  ( new_n36514_, new_n36513_, new_n36509_ );
and  ( new_n36515_, new_n36513_, new_n36509_ );
or   ( new_n36516_, new_n6173_, new_n24418_ );
or   ( new_n36517_, new_n6175_, new_n24227_ );
and  ( new_n36518_, new_n36517_, new_n36516_ );
xor  ( new_n36519_, new_n36518_, new_n5597_ );
nor  ( new_n36520_, new_n36519_, new_n36515_ );
nor  ( new_n36521_, new_n36520_, new_n36514_ );
nor  ( new_n36522_, new_n36521_, new_n36505_ );
nor  ( new_n36523_, new_n36522_, new_n36504_ );
or   ( new_n36524_, new_n36523_, new_n36469_ );
and  ( new_n36525_, new_n36524_, new_n36468_ );
nor  ( new_n36526_, new_n36525_, new_n36375_ );
and  ( new_n36527_, new_n36525_, new_n36375_ );
xnor ( new_n36528_, new_n36236_, new_n36234_ );
xor  ( new_n36529_, new_n36528_, new_n36240_ );
xnor ( new_n36530_, new_n36248_, new_n36246_ );
xor  ( new_n36531_, new_n36530_, new_n36252_ );
nor  ( new_n36532_, new_n36531_, new_n36529_ );
and  ( new_n36533_, new_n36531_, new_n36529_ );
xor  ( new_n36534_, new_n36231_, new_n36229_ );
nor  ( new_n36535_, new_n36534_, new_n36533_ );
nor  ( new_n36536_, new_n36535_, new_n36532_ );
nor  ( new_n36537_, new_n36536_, new_n36527_ );
nor  ( new_n36538_, new_n36537_, new_n36526_ );
and  ( new_n36539_, new_n36538_, new_n36339_ );
nor  ( new_n36540_, new_n36539_, new_n36337_ );
or   ( new_n36541_, new_n36540_, new_n36316_ );
and  ( new_n36542_, new_n36541_, new_n36315_ );
or   ( new_n36543_, new_n36542_, new_n36302_ );
and  ( new_n36544_, new_n36542_, new_n36302_ );
xnor ( new_n36545_, new_n36280_, new_n36068_ );
xor  ( new_n36546_, new_n36545_, new_n36284_ );
or   ( new_n36547_, new_n36546_, new_n36544_ );
and  ( new_n36548_, new_n36547_, new_n36543_ );
nor  ( new_n36549_, new_n36548_, new_n36297_ );
xor  ( new_n36550_, new_n36542_, new_n36302_ );
xor  ( new_n36551_, new_n36550_, new_n36546_ );
xor  ( new_n36552_, new_n36308_, new_n36306_ );
xor  ( new_n36553_, new_n36552_, new_n36312_ );
xnor ( new_n36554_, new_n36525_, new_n36375_ );
xor  ( new_n36555_, new_n36554_, new_n36536_ );
xnor ( new_n36556_, new_n36171_, new_n36131_ );
xor  ( new_n36557_, new_n36556_, new_n36223_ );
or   ( new_n36558_, new_n36557_, new_n36555_ );
and  ( new_n36559_, new_n36557_, new_n36555_ );
xor  ( new_n36560_, new_n36328_, new_n36326_ );
xor  ( new_n36561_, new_n36560_, new_n36332_ );
or   ( new_n36562_, new_n36561_, new_n36559_ );
and  ( new_n36563_, new_n36562_, new_n36558_ );
nor  ( new_n36564_, new_n36563_, new_n36553_ );
and  ( new_n36565_, new_n36563_, new_n36553_ );
xor  ( new_n36566_, new_n36361_, new_n36351_ );
xor  ( new_n36567_, new_n36566_, new_n36373_ );
xnor ( new_n36568_, new_n36320_, new_n36318_ );
xor  ( new_n36569_, new_n36568_, new_n36324_ );
nor  ( new_n36570_, new_n36569_, new_n36567_ );
and  ( new_n36571_, new_n36569_, new_n36567_ );
xor  ( new_n36572_, new_n36531_, new_n36529_ );
xnor ( new_n36573_, new_n36572_, new_n36534_ );
nor  ( new_n36574_, new_n36573_, new_n36571_ );
or   ( new_n36575_, new_n36574_, new_n36570_ );
xnor ( new_n36576_, new_n36242_, new_n36232_ );
xor  ( new_n36577_, new_n36576_, new_n36254_ );
and  ( new_n36578_, new_n36577_, new_n36575_ );
nor  ( new_n36579_, new_n36577_, new_n36575_ );
xor  ( new_n36580_, new_n36367_, new_n36365_ );
xor  ( new_n36581_, new_n36580_, new_n36371_ );
xnor ( new_n36582_, new_n36447_, new_n36431_ );
xor  ( new_n36583_, new_n36582_, new_n36465_ );
or   ( new_n36584_, new_n36583_, new_n36581_ );
nand ( new_n36585_, new_n36583_, new_n36581_ );
xor  ( new_n36586_, new_n36345_, new_n36343_ );
xnor ( new_n36587_, new_n36586_, new_n36349_ );
nand ( new_n36588_, new_n36587_, new_n36585_ );
and  ( new_n36589_, new_n36588_, new_n36584_ );
xor  ( new_n36590_, new_n36355_, new_n36353_ );
xor  ( new_n36591_, new_n36590_, new_n36359_ );
xnor ( new_n36592_, new_n36477_, new_n36473_ );
xor  ( new_n36593_, new_n36592_, new_n36483_ );
xnor ( new_n36594_, new_n36417_, new_n36413_ );
xor  ( new_n36595_, new_n36594_, new_n36423_ );
or   ( new_n36596_, new_n36595_, new_n36593_ );
and  ( new_n36597_, new_n36595_, new_n36593_ );
xor  ( new_n36598_, new_n36513_, new_n36509_ );
xnor ( new_n36599_, new_n36598_, new_n36519_ );
or   ( new_n36600_, new_n36599_, new_n36597_ );
and  ( new_n36601_, new_n36600_, new_n36596_ );
or   ( new_n36602_, new_n36601_, new_n36591_ );
and  ( new_n36603_, new_n36601_, new_n36591_ );
xnor ( new_n36604_, new_n36439_, new_n36435_ );
xor  ( new_n36605_, new_n36604_, new_n36445_ );
xnor ( new_n36606_, new_n36399_, new_n36395_ );
xor  ( new_n36607_, new_n36606_, new_n36405_ );
nor  ( new_n36608_, new_n36607_, new_n36605_ );
and  ( new_n36609_, new_n36607_, new_n36605_ );
xor  ( new_n36610_, new_n36383_, new_n36379_ );
xnor ( new_n36611_, new_n36610_, new_n36389_ );
nor  ( new_n36612_, new_n36611_, new_n36609_ );
nor  ( new_n36613_, new_n36612_, new_n36608_ );
or   ( new_n36614_, new_n36613_, new_n36603_ );
and  ( new_n36615_, new_n36614_, new_n36602_ );
nor  ( new_n36616_, new_n36615_, new_n36589_ );
and  ( new_n36617_, new_n36615_, new_n36589_ );
or   ( new_n36618_, new_n4709_, new_n25813_ );
or   ( new_n36619_, new_n4711_, new_n25486_ );
and  ( new_n36620_, new_n36619_, new_n36618_ );
xor  ( new_n36621_, new_n36620_, new_n4295_ );
or   ( new_n36622_, new_n4302_, new_n26063_ );
or   ( new_n36623_, new_n4304_, new_n26196_ );
and  ( new_n36624_, new_n36623_, new_n36622_ );
xor  ( new_n36625_, new_n36624_, new_n3895_ );
or   ( new_n36626_, new_n36625_, new_n36621_ );
and  ( new_n36627_, new_n36625_, new_n36621_ );
or   ( new_n36628_, new_n3896_, new_n26620_ );
or   ( new_n36629_, new_n3898_, new_n26372_ );
and  ( new_n36630_, new_n36629_, new_n36628_ );
xor  ( new_n36631_, new_n36630_, new_n3460_ );
or   ( new_n36632_, new_n36631_, new_n36627_ );
and  ( new_n36633_, new_n36632_, new_n36626_ );
or   ( new_n36634_, new_n3461_, new_n27085_ );
or   ( new_n36635_, new_n3463_, new_n26762_ );
and  ( new_n36636_, new_n36635_, new_n36634_ );
xor  ( new_n36637_, new_n36636_, new_n3116_ );
or   ( new_n36638_, new_n3117_, new_n27602_ );
or   ( new_n36639_, new_n3119_, new_n27396_ );
and  ( new_n36640_, new_n36639_, new_n36638_ );
xor  ( new_n36641_, new_n36640_, new_n2800_ );
or   ( new_n36642_, new_n36641_, new_n36637_ );
and  ( new_n36643_, new_n36641_, new_n36637_ );
or   ( new_n36644_, new_n2807_, new_n28108_ );
or   ( new_n36645_, new_n2809_, new_n27763_ );
and  ( new_n36646_, new_n36645_, new_n36644_ );
xor  ( new_n36647_, new_n36646_, new_n2424_ );
or   ( new_n36648_, new_n36647_, new_n36643_ );
and  ( new_n36649_, new_n36648_, new_n36642_ );
or   ( new_n36650_, new_n36649_, new_n36633_ );
and  ( new_n36651_, new_n36649_, new_n36633_ );
or   ( new_n36652_, new_n6173_, new_n24543_ );
or   ( new_n36653_, new_n6175_, new_n24418_ );
and  ( new_n36654_, new_n36653_, new_n36652_ );
xor  ( new_n36655_, new_n36654_, new_n5597_ );
or   ( new_n36656_, new_n5604_, new_n24925_ );
or   ( new_n36657_, new_n5606_, new_n24927_ );
and  ( new_n36658_, new_n36657_, new_n36656_ );
xor  ( new_n36659_, new_n36658_, new_n5206_ );
or   ( new_n36660_, new_n36659_, new_n36655_ );
and  ( new_n36661_, new_n36659_, new_n36655_ );
or   ( new_n36662_, new_n5207_, new_n25288_ );
or   ( new_n36663_, new_n5209_, new_n25048_ );
and  ( new_n36664_, new_n36663_, new_n36662_ );
xor  ( new_n36665_, new_n36664_, new_n4708_ );
or   ( new_n36666_, new_n36665_, new_n36661_ );
and  ( new_n36667_, new_n36666_, new_n36660_ );
or   ( new_n36668_, new_n36667_, new_n36651_ );
and  ( new_n36669_, new_n36668_, new_n36650_ );
xor  ( new_n36670_, new_n36457_, new_n36453_ );
xor  ( new_n36671_, new_n36670_, new_n36463_ );
or   ( new_n36672_, new_n2425_, new_n28531_ );
or   ( new_n36673_, new_n2427_, new_n28314_ );
and  ( new_n36674_, new_n36673_, new_n36672_ );
xor  ( new_n36675_, new_n36674_, new_n2121_ );
or   ( new_n36676_, new_n2122_, new_n29261_ );
or   ( new_n36677_, new_n2124_, new_n29263_ );
and  ( new_n36678_, new_n36677_, new_n36676_ );
xor  ( new_n36679_, new_n36678_, new_n1843_ );
or   ( new_n36680_, new_n36679_, new_n36675_ );
and  ( new_n36681_, new_n36679_, new_n36675_ );
or   ( new_n36682_, new_n1844_, new_n29619_ );
or   ( new_n36683_, new_n1846_, new_n29474_ );
and  ( new_n36684_, new_n36683_, new_n36682_ );
xor  ( new_n36685_, new_n36684_, new_n1586_ );
or   ( new_n36686_, new_n36685_, new_n36681_ );
and  ( new_n36687_, new_n36686_, new_n36680_ );
or   ( new_n36688_, new_n36687_, new_n36671_ );
and  ( new_n36689_, new_n36687_, new_n36671_ );
or   ( new_n36690_, new_n1593_, new_n30227_ );
or   ( new_n36691_, new_n1595_, new_n30120_ );
and  ( new_n36692_, new_n36691_, new_n36690_ );
xor  ( new_n36693_, new_n36692_, new_n1358_ );
or   ( new_n36694_, new_n1364_, new_n30798_ );
or   ( new_n36695_, new_n1366_, new_n30800_ );
and  ( new_n36696_, new_n36695_, new_n36694_ );
xor  ( new_n36697_, new_n36696_, new_n1129_ );
nor  ( new_n36698_, new_n36697_, new_n36693_ );
and  ( new_n36699_, new_n36697_, new_n36693_ );
or   ( new_n36700_, new_n1135_, new_n31654_ );
or   ( new_n36701_, new_n1137_, new_n31333_ );
and  ( new_n36702_, new_n36701_, new_n36700_ );
xor  ( new_n36703_, new_n36702_, new_n896_ );
nor  ( new_n36704_, new_n36703_, new_n36699_ );
nor  ( new_n36705_, new_n36704_, new_n36698_ );
or   ( new_n36706_, new_n36705_, new_n36689_ );
and  ( new_n36707_, new_n36706_, new_n36688_ );
nor  ( new_n36708_, new_n36707_, new_n36669_ );
and  ( new_n36709_, new_n36707_, new_n36669_ );
or   ( new_n36710_, new_n9422_, new_n22829_ );
or   ( new_n36711_, new_n9424_, new_n22641_ );
and  ( new_n36712_, new_n36711_, new_n36710_ );
xor  ( new_n36713_, new_n36712_, new_n8873_ );
or   ( new_n36714_, new_n8874_, new_n22973_ );
or   ( new_n36715_, new_n8876_, new_n22975_ );
and  ( new_n36716_, new_n36715_, new_n36714_ );
xor  ( new_n36717_, new_n36716_, new_n8257_ );
nor  ( new_n36718_, new_n36717_, new_n36713_ );
and  ( new_n36719_, new_n36717_, new_n36713_ );
or   ( new_n36720_, new_n8264_, new_n23252_ );
or   ( new_n36721_, new_n8266_, new_n23166_ );
and  ( new_n36722_, new_n36721_, new_n36720_ );
xor  ( new_n36723_, new_n36722_, new_n7725_ );
nor  ( new_n36724_, new_n36723_, new_n36719_ );
nor  ( new_n36725_, new_n36724_, new_n36718_ );
or   ( new_n36726_, new_n10059_, new_n22590_ );
or   ( new_n36727_, new_n10061_, new_n22423_ );
and  ( new_n36728_, new_n36727_, new_n36726_ );
xor  ( new_n36729_, new_n36728_, new_n9421_ );
and  ( new_n36730_, RIbb31de8_146, RIbb2d888_64 );
or   ( new_n36731_, new_n22304_, RIbb2d888_64 );
and  ( new_n36732_, new_n36731_, RIbb2d900_63 );
or   ( new_n36733_, new_n36732_, new_n36730_ );
or   ( new_n36734_, new_n10770_, new_n22207_ );
and  ( new_n36735_, new_n36734_, new_n36733_ );
nor  ( new_n36736_, new_n36735_, new_n36729_ );
and  ( new_n36737_, new_n36735_, new_n36729_ );
nor  ( new_n36738_, new_n36737_, new_n747_ );
nor  ( new_n36739_, new_n36738_, new_n36736_ );
or   ( new_n36740_, new_n7732_, new_n23554_ );
or   ( new_n36741_, new_n7734_, new_n23370_ );
and  ( new_n36742_, new_n36741_, new_n36740_ );
xor  ( new_n36743_, new_n36742_, new_n7177_ );
or   ( new_n36744_, new_n7184_, new_n23895_ );
or   ( new_n36745_, new_n7186_, new_n23733_ );
and  ( new_n36746_, new_n36745_, new_n36744_ );
xor  ( new_n36747_, new_n36746_, new_n6638_ );
nor  ( new_n36748_, new_n36747_, new_n36743_ );
and  ( new_n36749_, new_n36747_, new_n36743_ );
or   ( new_n36750_, new_n6645_, new_n24227_ );
or   ( new_n36751_, new_n6647_, new_n24006_ );
and  ( new_n36752_, new_n36751_, new_n36750_ );
xor  ( new_n36753_, new_n36752_, new_n6166_ );
nor  ( new_n36754_, new_n36753_, new_n36749_ );
nor  ( new_n36755_, new_n36754_, new_n36748_ );
and  ( new_n36756_, new_n36755_, new_n36739_ );
nor  ( new_n36757_, new_n36756_, new_n36725_ );
nor  ( new_n36758_, new_n36755_, new_n36739_ );
nor  ( new_n36759_, new_n36758_, new_n36757_ );
nor  ( new_n36760_, new_n36759_, new_n36709_ );
nor  ( new_n36761_, new_n36760_, new_n36708_ );
not  ( new_n36762_, new_n36761_ );
nor  ( new_n36763_, new_n36762_, new_n36617_ );
nor  ( new_n36764_, new_n36763_, new_n36616_ );
nor  ( new_n36765_, new_n36764_, new_n36579_ );
nor  ( new_n36766_, new_n36765_, new_n36578_ );
nor  ( new_n36767_, new_n36766_, new_n36565_ );
or   ( new_n36768_, new_n36767_, new_n36564_ );
xnor ( new_n36769_, new_n36314_, new_n36304_ );
xor  ( new_n36770_, new_n36769_, new_n36540_ );
nand ( new_n36771_, new_n36770_, new_n36768_ );
nor  ( new_n36772_, new_n36770_, new_n36768_ );
xnor ( new_n36773_, new_n36301_, new_n36299_ );
or   ( new_n36774_, new_n36773_, new_n36772_ );
and  ( new_n36775_, new_n36774_, new_n36771_ );
nor  ( new_n36776_, new_n36775_, new_n36551_ );
xor  ( new_n36777_, new_n36770_, new_n36768_ );
xor  ( new_n36778_, new_n36777_, new_n36773_ );
xor  ( new_n36779_, new_n36557_, new_n36555_ );
xor  ( new_n36780_, new_n36779_, new_n36561_ );
xnor ( new_n36781_, new_n36467_, new_n36427_ );
xor  ( new_n36782_, new_n36781_, new_n36523_ );
xor  ( new_n36783_, new_n36615_, new_n36589_ );
xor  ( new_n36784_, new_n36783_, new_n36762_ );
or   ( new_n36785_, new_n36784_, new_n36782_ );
and  ( new_n36786_, new_n36784_, new_n36782_ );
xor  ( new_n36787_, new_n36569_, new_n36567_ );
xor  ( new_n36788_, new_n36787_, new_n36573_ );
or   ( new_n36789_, new_n36788_, new_n36786_ );
and  ( new_n36790_, new_n36789_, new_n36785_ );
nor  ( new_n36791_, new_n36790_, new_n36780_ );
nand ( new_n36792_, new_n36790_, new_n36780_ );
xor  ( new_n36793_, new_n36601_, new_n36591_ );
xnor ( new_n36794_, new_n36793_, new_n36613_ );
not  ( new_n36795_, new_n36794_ );
xnor ( new_n36796_, new_n36707_, new_n36669_ );
xor  ( new_n36797_, new_n36796_, new_n36759_ );
or   ( new_n36798_, new_n36797_, new_n36795_ );
xnor ( new_n36799_, new_n36495_, new_n36489_ );
xor  ( new_n36800_, new_n36799_, new_n36501_ );
xnor ( new_n36801_, new_n36717_, new_n36713_ );
xor  ( new_n36802_, new_n36801_, new_n36723_ );
xnor ( new_n36803_, new_n36659_, new_n36655_ );
xor  ( new_n36804_, new_n36803_, new_n36665_ );
or   ( new_n36805_, new_n36804_, new_n36802_ );
and  ( new_n36806_, new_n36804_, new_n36802_ );
xor  ( new_n36807_, new_n36747_, new_n36743_ );
xnor ( new_n36808_, new_n36807_, new_n36753_ );
or   ( new_n36809_, new_n36808_, new_n36806_ );
and  ( new_n36810_, new_n36809_, new_n36805_ );
nor  ( new_n36811_, new_n36810_, new_n36800_ );
and  ( new_n36812_, new_n36810_, new_n36800_ );
xnor ( new_n36813_, new_n36641_, new_n36637_ );
xor  ( new_n36814_, new_n36813_, new_n36647_ );
xnor ( new_n36815_, new_n36679_, new_n36675_ );
xor  ( new_n36816_, new_n36815_, new_n36685_ );
nor  ( new_n36817_, new_n36816_, new_n36814_ );
and  ( new_n36818_, new_n36816_, new_n36814_ );
xor  ( new_n36819_, new_n36625_, new_n36621_ );
xnor ( new_n36820_, new_n36819_, new_n36631_ );
nor  ( new_n36821_, new_n36820_, new_n36818_ );
nor  ( new_n36822_, new_n36821_, new_n36817_ );
nor  ( new_n36823_, new_n36822_, new_n36812_ );
nor  ( new_n36824_, new_n36823_, new_n36811_ );
or   ( new_n36825_, new_n7184_, new_n24006_ );
or   ( new_n36826_, new_n7186_, new_n23895_ );
and  ( new_n36827_, new_n36826_, new_n36825_ );
xor  ( new_n36828_, new_n36827_, new_n6638_ );
or   ( new_n36829_, new_n6645_, new_n24418_ );
or   ( new_n36830_, new_n6647_, new_n24227_ );
and  ( new_n36831_, new_n36830_, new_n36829_ );
xor  ( new_n36832_, new_n36831_, new_n6166_ );
or   ( new_n36833_, new_n36832_, new_n36828_ );
and  ( new_n36834_, new_n36832_, new_n36828_ );
or   ( new_n36835_, new_n6173_, new_n24927_ );
or   ( new_n36836_, new_n6175_, new_n24543_ );
and  ( new_n36837_, new_n36836_, new_n36835_ );
xor  ( new_n36838_, new_n36837_, new_n5597_ );
or   ( new_n36839_, new_n36838_, new_n36834_ );
and  ( new_n36840_, new_n36839_, new_n36833_ );
or   ( new_n36841_, new_n8874_, new_n23166_ );
or   ( new_n36842_, new_n8876_, new_n22973_ );
and  ( new_n36843_, new_n36842_, new_n36841_ );
xor  ( new_n36844_, new_n36843_, new_n8257_ );
or   ( new_n36845_, new_n8264_, new_n23370_ );
or   ( new_n36846_, new_n8266_, new_n23252_ );
and  ( new_n36847_, new_n36846_, new_n36845_ );
xor  ( new_n36848_, new_n36847_, new_n7725_ );
or   ( new_n36849_, new_n36848_, new_n36844_ );
and  ( new_n36850_, new_n36848_, new_n36844_ );
or   ( new_n36851_, new_n7732_, new_n23733_ );
or   ( new_n36852_, new_n7734_, new_n23554_ );
and  ( new_n36853_, new_n36852_, new_n36851_ );
xor  ( new_n36854_, new_n36853_, new_n7177_ );
or   ( new_n36855_, new_n36854_, new_n36850_ );
and  ( new_n36856_, new_n36855_, new_n36849_ );
nor  ( new_n36857_, new_n36856_, new_n36840_ );
and  ( new_n36858_, new_n36856_, new_n36840_ );
or   ( new_n36859_, new_n10059_, new_n22641_ );
or   ( new_n36860_, new_n10061_, new_n22590_ );
and  ( new_n36861_, new_n36860_, new_n36859_ );
xor  ( new_n36862_, new_n36861_, new_n9421_ );
and  ( new_n36863_, RIbb31e60_147, RIbb2d888_64 );
or   ( new_n36864_, new_n22423_, RIbb2d888_64 );
and  ( new_n36865_, new_n36864_, RIbb2d900_63 );
or   ( new_n36866_, new_n36865_, new_n36863_ );
or   ( new_n36867_, new_n10770_, new_n22304_ );
and  ( new_n36868_, new_n36867_, new_n36866_ );
nor  ( new_n36869_, new_n36868_, new_n36862_ );
and  ( new_n36870_, new_n36868_, new_n36862_ );
or   ( new_n36871_, new_n9422_, new_n22975_ );
or   ( new_n36872_, new_n9424_, new_n22829_ );
and  ( new_n36873_, new_n36872_, new_n36871_ );
xor  ( new_n36874_, new_n36873_, new_n8873_ );
nor  ( new_n36875_, new_n36874_, new_n36870_ );
nor  ( new_n36876_, new_n36875_, new_n36869_ );
nor  ( new_n36877_, new_n36876_, new_n36858_ );
nor  ( new_n36878_, new_n36877_, new_n36857_ );
or   ( new_n36879_, new_n4302_, new_n26372_ );
or   ( new_n36880_, new_n4304_, new_n26063_ );
and  ( new_n36881_, new_n36880_, new_n36879_ );
xor  ( new_n36882_, new_n36881_, new_n3895_ );
or   ( new_n36883_, new_n3896_, new_n26762_ );
or   ( new_n36884_, new_n3898_, new_n26620_ );
and  ( new_n36885_, new_n36884_, new_n36883_ );
xor  ( new_n36886_, new_n36885_, new_n3460_ );
or   ( new_n36887_, new_n36886_, new_n36882_ );
and  ( new_n36888_, new_n36886_, new_n36882_ );
or   ( new_n36889_, new_n3461_, new_n27396_ );
or   ( new_n36890_, new_n3463_, new_n27085_ );
and  ( new_n36891_, new_n36890_, new_n36889_ );
xor  ( new_n36892_, new_n36891_, new_n3116_ );
or   ( new_n36893_, new_n36892_, new_n36888_ );
and  ( new_n36894_, new_n36893_, new_n36887_ );
or   ( new_n36895_, new_n5604_, new_n25048_ );
or   ( new_n36896_, new_n5606_, new_n24925_ );
and  ( new_n36897_, new_n36896_, new_n36895_ );
xor  ( new_n36898_, new_n36897_, new_n5206_ );
or   ( new_n36899_, new_n5207_, new_n25486_ );
or   ( new_n36900_, new_n5209_, new_n25288_ );
and  ( new_n36901_, new_n36900_, new_n36899_ );
xor  ( new_n36902_, new_n36901_, new_n4708_ );
or   ( new_n36903_, new_n36902_, new_n36898_ );
and  ( new_n36904_, new_n36902_, new_n36898_ );
or   ( new_n36905_, new_n4709_, new_n26196_ );
or   ( new_n36906_, new_n4711_, new_n25813_ );
and  ( new_n36907_, new_n36906_, new_n36905_ );
xor  ( new_n36908_, new_n36907_, new_n4295_ );
or   ( new_n36909_, new_n36908_, new_n36904_ );
and  ( new_n36910_, new_n36909_, new_n36903_ );
nor  ( new_n36911_, new_n36910_, new_n36894_ );
and  ( new_n36912_, new_n36910_, new_n36894_ );
or   ( new_n36913_, new_n3117_, new_n27763_ );
or   ( new_n36914_, new_n3119_, new_n27602_ );
and  ( new_n36915_, new_n36914_, new_n36913_ );
xor  ( new_n36916_, new_n36915_, new_n2800_ );
or   ( new_n36917_, new_n2807_, new_n28314_ );
or   ( new_n36918_, new_n2809_, new_n28108_ );
and  ( new_n36919_, new_n36918_, new_n36917_ );
xor  ( new_n36920_, new_n36919_, new_n2424_ );
nor  ( new_n36921_, new_n36920_, new_n36916_ );
and  ( new_n36922_, new_n36920_, new_n36916_ );
or   ( new_n36923_, new_n2425_, new_n29263_ );
or   ( new_n36924_, new_n2427_, new_n28531_ );
and  ( new_n36925_, new_n36924_, new_n36923_ );
xor  ( new_n36926_, new_n36925_, new_n2121_ );
nor  ( new_n36927_, new_n36926_, new_n36922_ );
nor  ( new_n36928_, new_n36927_, new_n36921_ );
nor  ( new_n36929_, new_n36928_, new_n36912_ );
nor  ( new_n36930_, new_n36929_, new_n36911_ );
and  ( new_n36931_, new_n36930_, new_n36878_ );
nor  ( new_n36932_, new_n36930_, new_n36878_ );
and  ( new_n36933_, new_n820_, RIbb33378_192 );
or   ( new_n36934_, new_n36933_, new_n748_ );
nand ( new_n36935_, new_n36933_, new_n745_ );
and  ( new_n36936_, new_n36935_, new_n36934_ );
xnor ( new_n36937_, new_n36697_, new_n36693_ );
xor  ( new_n36938_, new_n36937_, new_n36703_ );
nor  ( new_n36939_, new_n36938_, new_n36936_ );
and  ( new_n36940_, new_n36938_, new_n36936_ );
not  ( new_n36941_, new_n36940_ );
or   ( new_n36942_, new_n2122_, new_n29474_ );
or   ( new_n36943_, new_n2124_, new_n29261_ );
and  ( new_n36944_, new_n36943_, new_n36942_ );
xor  ( new_n36945_, new_n36944_, new_n1843_ );
or   ( new_n36946_, new_n1844_, new_n30120_ );
or   ( new_n36947_, new_n1846_, new_n29619_ );
and  ( new_n36948_, new_n36947_, new_n36946_ );
xor  ( new_n36949_, new_n36948_, new_n1586_ );
nor  ( new_n36950_, new_n36949_, new_n36945_ );
and  ( new_n36951_, new_n36949_, new_n36945_ );
or   ( new_n36952_, new_n1593_, new_n30800_ );
or   ( new_n36953_, new_n1595_, new_n30227_ );
and  ( new_n36954_, new_n36953_, new_n36952_ );
xor  ( new_n36955_, new_n36954_, new_n1358_ );
nor  ( new_n36956_, new_n36955_, new_n36951_ );
nor  ( new_n36957_, new_n36956_, new_n36950_ );
and  ( new_n36958_, new_n36957_, new_n36941_ );
nor  ( new_n36959_, new_n36958_, new_n36939_ );
nor  ( new_n36960_, new_n36959_, new_n36932_ );
nor  ( new_n36961_, new_n36960_, new_n36931_ );
and  ( new_n36962_, new_n36961_, new_n36824_ );
xnor ( new_n36963_, new_n36607_, new_n36605_ );
xor  ( new_n36964_, new_n36963_, new_n36611_ );
xnor ( new_n36965_, new_n36595_, new_n36593_ );
xor  ( new_n36966_, new_n36965_, new_n36599_ );
and  ( new_n36967_, new_n36966_, new_n36964_ );
nor  ( new_n36968_, new_n36966_, new_n36964_ );
xor  ( new_n36969_, new_n36687_, new_n36671_ );
xnor ( new_n36970_, new_n36969_, new_n36705_ );
nor  ( new_n36971_, new_n36970_, new_n36968_ );
nor  ( new_n36972_, new_n36971_, new_n36967_ );
nor  ( new_n36973_, new_n36972_, new_n36962_ );
nor  ( new_n36974_, new_n36961_, new_n36824_ );
nor  ( new_n36975_, new_n36974_, new_n36973_ );
nor  ( new_n36976_, new_n36975_, new_n36798_ );
and  ( new_n36977_, new_n36975_, new_n36798_ );
xnor ( new_n36978_, new_n36503_, new_n36485_ );
xor  ( new_n36979_, new_n36978_, new_n36521_ );
xnor ( new_n36980_, new_n36407_, new_n36391_ );
xor  ( new_n36981_, new_n36980_, new_n36425_ );
nor  ( new_n36982_, new_n36981_, new_n36979_ );
and  ( new_n36983_, new_n36981_, new_n36979_ );
xor  ( new_n36984_, new_n36583_, new_n36581_ );
xor  ( new_n36985_, new_n36984_, new_n36587_ );
not  ( new_n36986_, new_n36985_ );
nor  ( new_n36987_, new_n36986_, new_n36983_ );
nor  ( new_n36988_, new_n36987_, new_n36982_ );
nor  ( new_n36989_, new_n36988_, new_n36977_ );
nor  ( new_n36990_, new_n36989_, new_n36976_ );
not  ( new_n36991_, new_n36990_ );
and  ( new_n36992_, new_n36991_, new_n36792_ );
or   ( new_n36993_, new_n36992_, new_n36791_ );
xor  ( new_n36994_, new_n36336_, new_n36334_ );
xor  ( new_n36995_, new_n36994_, new_n36538_ );
nand ( new_n36996_, new_n36995_, new_n36993_ );
nor  ( new_n36997_, new_n36995_, new_n36993_ );
xor  ( new_n36998_, new_n36563_, new_n36553_ );
xor  ( new_n36999_, new_n36998_, new_n36766_ );
or   ( new_n37000_, new_n36999_, new_n36997_ );
and  ( new_n37001_, new_n37000_, new_n36996_ );
nor  ( new_n37002_, new_n37001_, new_n36778_ );
xor  ( new_n37003_, new_n36995_, new_n36993_ );
xor  ( new_n37004_, new_n37003_, new_n36999_ );
xor  ( new_n37005_, new_n36784_, new_n36782_ );
xor  ( new_n37006_, new_n37005_, new_n36788_ );
xnor ( new_n37007_, new_n36961_, new_n36824_ );
and  ( new_n37008_, new_n37007_, new_n36972_ );
not  ( new_n37009_, new_n36974_ );
and  ( new_n37010_, new_n37009_, new_n36973_ );
or   ( new_n37011_, new_n37010_, new_n37008_ );
xor  ( new_n37012_, new_n36981_, new_n36979_ );
xor  ( new_n37013_, new_n37012_, new_n36986_ );
or   ( new_n37014_, new_n37013_, new_n37011_ );
nand ( new_n37015_, new_n37013_, new_n37011_ );
xor  ( new_n37016_, new_n36797_, new_n36795_ );
nand ( new_n37017_, new_n37016_, new_n37015_ );
and  ( new_n37018_, new_n37017_, new_n37014_ );
nor  ( new_n37019_, new_n37018_, new_n37006_ );
nand ( new_n37020_, new_n37018_, new_n37006_ );
xnor ( new_n37021_, new_n36930_, new_n36878_ );
xor  ( new_n37022_, new_n37021_, new_n36959_ );
xnor ( new_n37023_, new_n36810_, new_n36800_ );
xor  ( new_n37024_, new_n37023_, new_n36822_ );
nand ( new_n37025_, new_n37024_, new_n37022_ );
or   ( new_n37026_, new_n10059_, new_n22829_ );
or   ( new_n37027_, new_n10061_, new_n22641_ );
and  ( new_n37028_, new_n37027_, new_n37026_ );
xor  ( new_n37029_, new_n37028_, new_n9421_ );
and  ( new_n37030_, RIbb31ed8_148, RIbb2d888_64 );
or   ( new_n37031_, new_n22590_, RIbb2d888_64 );
and  ( new_n37032_, new_n37031_, RIbb2d900_63 );
or   ( new_n37033_, new_n37032_, new_n37030_ );
or   ( new_n37034_, new_n10770_, new_n22423_ );
and  ( new_n37035_, new_n37034_, new_n37033_ );
or   ( new_n37036_, new_n37035_, new_n37029_ );
and  ( new_n37037_, new_n37035_, new_n37029_ );
or   ( new_n37038_, new_n37037_, new_n895_ );
and  ( new_n37039_, new_n37038_, new_n37036_ );
or   ( new_n37040_, new_n7732_, new_n23895_ );
or   ( new_n37041_, new_n7734_, new_n23733_ );
and  ( new_n37042_, new_n37041_, new_n37040_ );
xor  ( new_n37043_, new_n37042_, new_n7177_ );
or   ( new_n37044_, new_n7184_, new_n24227_ );
or   ( new_n37045_, new_n7186_, new_n24006_ );
and  ( new_n37046_, new_n37045_, new_n37044_ );
xor  ( new_n37047_, new_n37046_, new_n6638_ );
or   ( new_n37048_, new_n37047_, new_n37043_ );
and  ( new_n37049_, new_n37047_, new_n37043_ );
or   ( new_n37050_, new_n6645_, new_n24543_ );
or   ( new_n37051_, new_n6647_, new_n24418_ );
and  ( new_n37052_, new_n37051_, new_n37050_ );
xor  ( new_n37053_, new_n37052_, new_n6166_ );
or   ( new_n37054_, new_n37053_, new_n37049_ );
and  ( new_n37055_, new_n37054_, new_n37048_ );
or   ( new_n37056_, new_n37055_, new_n37039_ );
and  ( new_n37057_, new_n37055_, new_n37039_ );
or   ( new_n37058_, new_n9422_, new_n22973_ );
or   ( new_n37059_, new_n9424_, new_n22975_ );
and  ( new_n37060_, new_n37059_, new_n37058_ );
xor  ( new_n37061_, new_n37060_, new_n8873_ );
or   ( new_n37062_, new_n8874_, new_n23252_ );
or   ( new_n37063_, new_n8876_, new_n23166_ );
and  ( new_n37064_, new_n37063_, new_n37062_ );
xor  ( new_n37065_, new_n37064_, new_n8257_ );
nor  ( new_n37066_, new_n37065_, new_n37061_ );
and  ( new_n37067_, new_n37065_, new_n37061_ );
or   ( new_n37068_, new_n8264_, new_n23554_ );
or   ( new_n37069_, new_n8266_, new_n23370_ );
and  ( new_n37070_, new_n37069_, new_n37068_ );
xor  ( new_n37071_, new_n37070_, new_n7725_ );
nor  ( new_n37072_, new_n37071_, new_n37067_ );
nor  ( new_n37073_, new_n37072_, new_n37066_ );
or   ( new_n37074_, new_n37073_, new_n37057_ );
and  ( new_n37075_, new_n37074_, new_n37056_ );
or   ( new_n37076_, new_n1364_, new_n31333_ );
or   ( new_n37077_, new_n1366_, new_n30798_ );
and  ( new_n37078_, new_n37077_, new_n37076_ );
xor  ( new_n37079_, new_n37078_, new_n1128_ );
or   ( new_n37080_, new_n1593_, new_n30798_ );
or   ( new_n37081_, new_n1595_, new_n30800_ );
and  ( new_n37082_, new_n37081_, new_n37080_ );
xor  ( new_n37083_, new_n37082_, new_n1358_ );
or   ( new_n37084_, new_n1364_, new_n31654_ );
or   ( new_n37085_, new_n1366_, new_n31333_ );
and  ( new_n37086_, new_n37085_, new_n37084_ );
xor  ( new_n37087_, new_n37086_, new_n1129_ );
nand ( new_n37088_, new_n37087_, new_n37083_ );
nor  ( new_n37089_, new_n37087_, new_n37083_ );
and  ( new_n37090_, new_n1040_, RIbb33378_192 );
nor  ( new_n37091_, new_n37090_, new_n896_ );
and  ( new_n37092_, new_n37090_, new_n893_ );
nor  ( new_n37093_, new_n37092_, new_n37091_ );
or   ( new_n37094_, new_n37093_, new_n37089_ );
and  ( new_n37095_, new_n37094_, new_n37088_ );
nand ( new_n37096_, new_n37095_, new_n37079_ );
nor  ( new_n37097_, new_n37095_, new_n37079_ );
or   ( new_n37098_, new_n2425_, new_n29261_ );
or   ( new_n37099_, new_n2427_, new_n29263_ );
and  ( new_n37100_, new_n37099_, new_n37098_ );
xor  ( new_n37101_, new_n37100_, new_n2121_ );
or   ( new_n37102_, new_n2122_, new_n29619_ );
or   ( new_n37103_, new_n2124_, new_n29474_ );
and  ( new_n37104_, new_n37103_, new_n37102_ );
xor  ( new_n37105_, new_n37104_, new_n1843_ );
nor  ( new_n37106_, new_n37105_, new_n37101_ );
and  ( new_n37107_, new_n37105_, new_n37101_ );
or   ( new_n37108_, new_n1844_, new_n30227_ );
or   ( new_n37109_, new_n1846_, new_n30120_ );
and  ( new_n37110_, new_n37109_, new_n37108_ );
xor  ( new_n37111_, new_n37110_, new_n1586_ );
nor  ( new_n37112_, new_n37111_, new_n37107_ );
nor  ( new_n37113_, new_n37112_, new_n37106_ );
or   ( new_n37114_, new_n37113_, new_n37097_ );
and  ( new_n37115_, new_n37114_, new_n37096_ );
nor  ( new_n37116_, new_n37115_, new_n37075_ );
nand ( new_n37117_, new_n37115_, new_n37075_ );
or   ( new_n37118_, new_n4709_, new_n26063_ );
or   ( new_n37119_, new_n4711_, new_n26196_ );
and  ( new_n37120_, new_n37119_, new_n37118_ );
xor  ( new_n37121_, new_n37120_, new_n4295_ );
or   ( new_n37122_, new_n4302_, new_n26620_ );
or   ( new_n37123_, new_n4304_, new_n26372_ );
and  ( new_n37124_, new_n37123_, new_n37122_ );
xor  ( new_n37125_, new_n37124_, new_n3895_ );
or   ( new_n37126_, new_n37125_, new_n37121_ );
and  ( new_n37127_, new_n37125_, new_n37121_ );
or   ( new_n37128_, new_n3896_, new_n27085_ );
or   ( new_n37129_, new_n3898_, new_n26762_ );
and  ( new_n37130_, new_n37129_, new_n37128_ );
xor  ( new_n37131_, new_n37130_, new_n3460_ );
or   ( new_n37132_, new_n37131_, new_n37127_ );
and  ( new_n37133_, new_n37132_, new_n37126_ );
or   ( new_n37134_, new_n6173_, new_n24925_ );
or   ( new_n37135_, new_n6175_, new_n24927_ );
and  ( new_n37136_, new_n37135_, new_n37134_ );
xor  ( new_n37137_, new_n37136_, new_n5597_ );
or   ( new_n37138_, new_n5604_, new_n25288_ );
or   ( new_n37139_, new_n5606_, new_n25048_ );
and  ( new_n37140_, new_n37139_, new_n37138_ );
xor  ( new_n37141_, new_n37140_, new_n5206_ );
or   ( new_n37142_, new_n37141_, new_n37137_ );
and  ( new_n37143_, new_n37141_, new_n37137_ );
or   ( new_n37144_, new_n5207_, new_n25813_ );
or   ( new_n37145_, new_n5209_, new_n25486_ );
and  ( new_n37146_, new_n37145_, new_n37144_ );
xor  ( new_n37147_, new_n37146_, new_n4708_ );
or   ( new_n37148_, new_n37147_, new_n37143_ );
and  ( new_n37149_, new_n37148_, new_n37142_ );
nor  ( new_n37150_, new_n37149_, new_n37133_ );
nand ( new_n37151_, new_n37149_, new_n37133_ );
or   ( new_n37152_, new_n3461_, new_n27602_ );
or   ( new_n37153_, new_n3463_, new_n27396_ );
and  ( new_n37154_, new_n37153_, new_n37152_ );
xor  ( new_n37155_, new_n37154_, new_n3116_ );
or   ( new_n37156_, new_n3117_, new_n28108_ );
or   ( new_n37157_, new_n3119_, new_n27763_ );
and  ( new_n37158_, new_n37157_, new_n37156_ );
xor  ( new_n37159_, new_n37158_, new_n2800_ );
nor  ( new_n37160_, new_n37159_, new_n37155_ );
and  ( new_n37161_, new_n37159_, new_n37155_ );
or   ( new_n37162_, new_n2807_, new_n28531_ );
or   ( new_n37163_, new_n2809_, new_n28314_ );
and  ( new_n37164_, new_n37163_, new_n37162_ );
xor  ( new_n37165_, new_n37164_, new_n2424_ );
nor  ( new_n37166_, new_n37165_, new_n37161_ );
or   ( new_n37167_, new_n37166_, new_n37160_ );
and  ( new_n37168_, new_n37167_, new_n37151_ );
or   ( new_n37169_, new_n37168_, new_n37150_ );
and  ( new_n37170_, new_n37169_, new_n37117_ );
or   ( new_n37171_, new_n37170_, new_n37116_ );
or   ( new_n37172_, new_n1135_, new_n31952_ );
or   ( new_n37173_, new_n1137_, new_n31654_ );
and  ( new_n37174_, new_n37173_, new_n37172_ );
xor  ( new_n37175_, new_n37174_, new_n895_ );
xnor ( new_n37176_, new_n36920_, new_n36916_ );
xor  ( new_n37177_, new_n37176_, new_n36926_ );
and  ( new_n37178_, new_n37177_, new_n37175_ );
or   ( new_n37179_, new_n37177_, new_n37175_ );
xnor ( new_n37180_, new_n36949_, new_n36945_ );
xor  ( new_n37181_, new_n37180_, new_n36955_ );
and  ( new_n37182_, new_n37181_, new_n37179_ );
or   ( new_n37183_, new_n37182_, new_n37178_ );
xnor ( new_n37184_, new_n36902_, new_n36898_ );
xor  ( new_n37185_, new_n37184_, new_n36908_ );
xnor ( new_n37186_, new_n36886_, new_n36882_ );
xor  ( new_n37187_, new_n37186_, new_n36892_ );
or   ( new_n37188_, new_n37187_, new_n37185_ );
and  ( new_n37189_, new_n37187_, new_n37185_ );
xor  ( new_n37190_, new_n36832_, new_n36828_ );
xnor ( new_n37191_, new_n37190_, new_n36838_ );
or   ( new_n37192_, new_n37191_, new_n37189_ );
and  ( new_n37193_, new_n37192_, new_n37188_ );
or   ( new_n37194_, new_n37193_, new_n37183_ );
and  ( new_n37195_, new_n37193_, new_n37183_ );
xor  ( new_n37196_, new_n36735_, new_n36729_ );
xor  ( new_n37197_, new_n37196_, new_n748_ );
or   ( new_n37198_, new_n37197_, new_n37195_ );
and  ( new_n37199_, new_n37198_, new_n37194_ );
or   ( new_n37200_, new_n37199_, new_n37171_ );
and  ( new_n37201_, new_n37199_, new_n37171_ );
xor  ( new_n37202_, new_n36938_, new_n36936_ );
xor  ( new_n37203_, new_n37202_, new_n36957_ );
xnor ( new_n37204_, new_n36804_, new_n36802_ );
xor  ( new_n37205_, new_n37204_, new_n36808_ );
nor  ( new_n37206_, new_n37205_, new_n37203_ );
nand ( new_n37207_, new_n37205_, new_n37203_ );
xor  ( new_n37208_, new_n36816_, new_n36814_ );
xnor ( new_n37209_, new_n37208_, new_n36820_ );
not  ( new_n37210_, new_n37209_ );
and  ( new_n37211_, new_n37210_, new_n37207_ );
or   ( new_n37212_, new_n37211_, new_n37206_ );
or   ( new_n37213_, new_n37212_, new_n37201_ );
and  ( new_n37214_, new_n37213_, new_n37200_ );
nor  ( new_n37215_, new_n37214_, new_n37025_ );
and  ( new_n37216_, new_n37214_, new_n37025_ );
xor  ( new_n37217_, new_n36649_, new_n36633_ );
xor  ( new_n37218_, new_n37217_, new_n36667_ );
xor  ( new_n37219_, new_n36755_, new_n36739_ );
xor  ( new_n37220_, new_n37219_, new_n36725_ );
and  ( new_n37221_, new_n37220_, new_n37218_ );
nor  ( new_n37222_, new_n37220_, new_n37218_ );
xor  ( new_n37223_, new_n36966_, new_n36964_ );
xnor ( new_n37224_, new_n37223_, new_n36970_ );
not  ( new_n37225_, new_n37224_ );
nor  ( new_n37226_, new_n37225_, new_n37222_ );
nor  ( new_n37227_, new_n37226_, new_n37221_ );
nor  ( new_n37228_, new_n37227_, new_n37216_ );
nor  ( new_n37229_, new_n37228_, new_n37215_ );
not  ( new_n37230_, new_n37229_ );
and  ( new_n37231_, new_n37230_, new_n37020_ );
or   ( new_n37232_, new_n37231_, new_n37019_ );
xnor ( new_n37233_, new_n36577_, new_n36575_ );
xor  ( new_n37234_, new_n37233_, new_n36764_ );
nand ( new_n37235_, new_n37234_, new_n37232_ );
or   ( new_n37236_, new_n37234_, new_n37232_ );
xor  ( new_n37237_, new_n36790_, new_n36780_ );
xor  ( new_n37238_, new_n37237_, new_n36991_ );
nand ( new_n37239_, new_n37238_, new_n37236_ );
and  ( new_n37240_, new_n37239_, new_n37235_ );
nor  ( new_n37241_, new_n37240_, new_n37004_ );
xor  ( new_n37242_, new_n37013_, new_n37011_ );
xor  ( new_n37243_, new_n37242_, new_n37016_ );
xnor ( new_n37244_, new_n36910_, new_n36894_ );
xor  ( new_n37245_, new_n37244_, new_n36928_ );
xnor ( new_n37246_, new_n37055_, new_n37039_ );
xor  ( new_n37247_, new_n37246_, new_n37073_ );
xor  ( new_n37248_, new_n37149_, new_n37133_ );
xor  ( new_n37249_, new_n37248_, new_n37167_ );
or   ( new_n37250_, new_n37249_, new_n37247_ );
and  ( new_n37251_, new_n37249_, new_n37247_ );
xor  ( new_n37252_, new_n37095_, new_n37079_ );
xnor ( new_n37253_, new_n37252_, new_n37113_ );
or   ( new_n37254_, new_n37253_, new_n37251_ );
and  ( new_n37255_, new_n37254_, new_n37250_ );
nor  ( new_n37256_, new_n37255_, new_n37245_ );
and  ( new_n37257_, new_n37255_, new_n37245_ );
xor  ( new_n37258_, new_n36856_, new_n36840_ );
xnor ( new_n37259_, new_n37258_, new_n36876_ );
nor  ( new_n37260_, new_n37259_, new_n37257_ );
or   ( new_n37261_, new_n37260_, new_n37256_ );
xnor ( new_n37262_, new_n36848_, new_n36844_ );
xor  ( new_n37263_, new_n37262_, new_n36854_ );
xor  ( new_n37264_, new_n37035_, new_n37029_ );
xor  ( new_n37265_, new_n37264_, new_n896_ );
xnor ( new_n37266_, new_n37047_, new_n37043_ );
xor  ( new_n37267_, new_n37266_, new_n37053_ );
or   ( new_n37268_, new_n37267_, new_n37265_ );
and  ( new_n37269_, new_n37267_, new_n37265_ );
xnor ( new_n37270_, new_n37065_, new_n37061_ );
xor  ( new_n37271_, new_n37270_, new_n37071_ );
or   ( new_n37272_, new_n37271_, new_n37269_ );
and  ( new_n37273_, new_n37272_, new_n37268_ );
nor  ( new_n37274_, new_n37273_, new_n37263_ );
nand ( new_n37275_, new_n37273_, new_n37263_ );
xnor ( new_n37276_, new_n37141_, new_n37137_ );
xor  ( new_n37277_, new_n37276_, new_n37147_ );
xnor ( new_n37278_, new_n37125_, new_n37121_ );
xor  ( new_n37279_, new_n37278_, new_n37131_ );
nor  ( new_n37280_, new_n37279_, new_n37277_ );
nand ( new_n37281_, new_n37279_, new_n37277_ );
xor  ( new_n37282_, new_n37159_, new_n37155_ );
xor  ( new_n37283_, new_n37282_, new_n37165_ );
and  ( new_n37284_, new_n37283_, new_n37281_ );
or   ( new_n37285_, new_n37284_, new_n37280_ );
and  ( new_n37286_, new_n37285_, new_n37275_ );
or   ( new_n37287_, new_n37286_, new_n37274_ );
or   ( new_n37288_, new_n8874_, new_n23370_ );
or   ( new_n37289_, new_n8876_, new_n23252_ );
and  ( new_n37290_, new_n37289_, new_n37288_ );
xor  ( new_n37291_, new_n37290_, new_n8257_ );
or   ( new_n37292_, new_n8264_, new_n23733_ );
or   ( new_n37293_, new_n8266_, new_n23554_ );
and  ( new_n37294_, new_n37293_, new_n37292_ );
xor  ( new_n37295_, new_n37294_, new_n7725_ );
or   ( new_n37296_, new_n37295_, new_n37291_ );
and  ( new_n37297_, new_n37295_, new_n37291_ );
or   ( new_n37298_, new_n7732_, new_n24006_ );
or   ( new_n37299_, new_n7734_, new_n23895_ );
and  ( new_n37300_, new_n37299_, new_n37298_ );
xor  ( new_n37301_, new_n37300_, new_n7177_ );
or   ( new_n37302_, new_n37301_, new_n37297_ );
and  ( new_n37303_, new_n37302_, new_n37296_ );
or   ( new_n37304_, new_n10059_, new_n22975_ );
or   ( new_n37305_, new_n10061_, new_n22829_ );
and  ( new_n37306_, new_n37305_, new_n37304_ );
xor  ( new_n37307_, new_n37306_, new_n9421_ );
and  ( new_n37308_, RIbb31f50_149, RIbb2d888_64 );
or   ( new_n37309_, new_n22641_, RIbb2d888_64 );
and  ( new_n37310_, new_n37309_, RIbb2d900_63 );
or   ( new_n37311_, new_n37310_, new_n37308_ );
or   ( new_n37312_, new_n10770_, new_n22590_ );
and  ( new_n37313_, new_n37312_, new_n37311_ );
or   ( new_n37314_, new_n37313_, new_n37307_ );
and  ( new_n37315_, new_n37313_, new_n37307_ );
or   ( new_n37316_, new_n9422_, new_n23166_ );
or   ( new_n37317_, new_n9424_, new_n22973_ );
and  ( new_n37318_, new_n37317_, new_n37316_ );
xor  ( new_n37319_, new_n37318_, new_n8873_ );
or   ( new_n37320_, new_n37319_, new_n37315_ );
and  ( new_n37321_, new_n37320_, new_n37314_ );
or   ( new_n37322_, new_n37321_, new_n37303_ );
and  ( new_n37323_, new_n37321_, new_n37303_ );
or   ( new_n37324_, new_n7184_, new_n24418_ );
or   ( new_n37325_, new_n7186_, new_n24227_ );
and  ( new_n37326_, new_n37325_, new_n37324_ );
xor  ( new_n37327_, new_n37326_, new_n6638_ );
or   ( new_n37328_, new_n6645_, new_n24927_ );
or   ( new_n37329_, new_n6647_, new_n24543_ );
and  ( new_n37330_, new_n37329_, new_n37328_ );
xor  ( new_n37331_, new_n37330_, new_n6166_ );
or   ( new_n37332_, new_n37331_, new_n37327_ );
and  ( new_n37333_, new_n37331_, new_n37327_ );
or   ( new_n37334_, new_n6173_, new_n25048_ );
or   ( new_n37335_, new_n6175_, new_n24925_ );
and  ( new_n37336_, new_n37335_, new_n37334_ );
xor  ( new_n37337_, new_n37336_, new_n5597_ );
or   ( new_n37338_, new_n37337_, new_n37333_ );
and  ( new_n37339_, new_n37338_, new_n37332_ );
or   ( new_n37340_, new_n37339_, new_n37323_ );
and  ( new_n37341_, new_n37340_, new_n37322_ );
xor  ( new_n37342_, new_n37105_, new_n37101_ );
xor  ( new_n37343_, new_n37342_, new_n37111_ );
or   ( new_n37344_, new_n2122_, new_n30120_ );
or   ( new_n37345_, new_n2124_, new_n29619_ );
and  ( new_n37346_, new_n37345_, new_n37344_ );
xor  ( new_n37347_, new_n37346_, new_n1843_ );
or   ( new_n37348_, new_n1844_, new_n30800_ );
or   ( new_n37349_, new_n1846_, new_n30227_ );
and  ( new_n37350_, new_n37349_, new_n37348_ );
xor  ( new_n37351_, new_n37350_, new_n1586_ );
or   ( new_n37352_, new_n37351_, new_n37347_ );
and  ( new_n37353_, new_n37351_, new_n37347_ );
or   ( new_n37354_, new_n1593_, new_n31333_ );
or   ( new_n37355_, new_n1595_, new_n30798_ );
and  ( new_n37356_, new_n37355_, new_n37354_ );
xor  ( new_n37357_, new_n37356_, new_n1358_ );
or   ( new_n37358_, new_n37357_, new_n37353_ );
and  ( new_n37359_, new_n37358_, new_n37352_ );
or   ( new_n37360_, new_n37359_, new_n37343_ );
and  ( new_n37361_, new_n37359_, new_n37343_ );
xor  ( new_n37362_, new_n37087_, new_n37083_ );
xnor ( new_n37363_, new_n37362_, new_n37093_ );
or   ( new_n37364_, new_n37363_, new_n37361_ );
and  ( new_n37365_, new_n37364_, new_n37360_ );
or   ( new_n37366_, new_n37365_, new_n37341_ );
and  ( new_n37367_, new_n37365_, new_n37341_ );
or   ( new_n37368_, new_n3117_, new_n28314_ );
or   ( new_n37369_, new_n3119_, new_n28108_ );
and  ( new_n37370_, new_n37369_, new_n37368_ );
xor  ( new_n37371_, new_n37370_, new_n2800_ );
or   ( new_n37372_, new_n2807_, new_n29263_ );
or   ( new_n37373_, new_n2809_, new_n28531_ );
and  ( new_n37374_, new_n37373_, new_n37372_ );
xor  ( new_n37375_, new_n37374_, new_n2424_ );
or   ( new_n37376_, new_n37375_, new_n37371_ );
and  ( new_n37377_, new_n37375_, new_n37371_ );
or   ( new_n37378_, new_n2425_, new_n29474_ );
or   ( new_n37379_, new_n2427_, new_n29261_ );
and  ( new_n37380_, new_n37379_, new_n37378_ );
xor  ( new_n37381_, new_n37380_, new_n2121_ );
or   ( new_n37382_, new_n37381_, new_n37377_ );
and  ( new_n37383_, new_n37382_, new_n37376_ );
or   ( new_n37384_, new_n4302_, new_n26762_ );
or   ( new_n37385_, new_n4304_, new_n26620_ );
and  ( new_n37386_, new_n37385_, new_n37384_ );
xor  ( new_n37387_, new_n37386_, new_n3895_ );
or   ( new_n37388_, new_n3896_, new_n27396_ );
or   ( new_n37389_, new_n3898_, new_n27085_ );
and  ( new_n37390_, new_n37389_, new_n37388_ );
xor  ( new_n37391_, new_n37390_, new_n3460_ );
or   ( new_n37392_, new_n37391_, new_n37387_ );
and  ( new_n37393_, new_n37391_, new_n37387_ );
or   ( new_n37394_, new_n3461_, new_n27763_ );
or   ( new_n37395_, new_n3463_, new_n27602_ );
and  ( new_n37396_, new_n37395_, new_n37394_ );
xor  ( new_n37397_, new_n37396_, new_n3116_ );
or   ( new_n37398_, new_n37397_, new_n37393_ );
and  ( new_n37399_, new_n37398_, new_n37392_ );
nor  ( new_n37400_, new_n37399_, new_n37383_ );
and  ( new_n37401_, new_n37399_, new_n37383_ );
or   ( new_n37402_, new_n5604_, new_n25486_ );
or   ( new_n37403_, new_n5606_, new_n25288_ );
and  ( new_n37404_, new_n37403_, new_n37402_ );
xor  ( new_n37405_, new_n37404_, new_n5206_ );
or   ( new_n37406_, new_n5207_, new_n26196_ );
or   ( new_n37407_, new_n5209_, new_n25813_ );
and  ( new_n37408_, new_n37407_, new_n37406_ );
xor  ( new_n37409_, new_n37408_, new_n4708_ );
nor  ( new_n37410_, new_n37409_, new_n37405_ );
and  ( new_n37411_, new_n37409_, new_n37405_ );
or   ( new_n37412_, new_n4709_, new_n26372_ );
or   ( new_n37413_, new_n4711_, new_n26063_ );
and  ( new_n37414_, new_n37413_, new_n37412_ );
xor  ( new_n37415_, new_n37414_, new_n4295_ );
nor  ( new_n37416_, new_n37415_, new_n37411_ );
nor  ( new_n37417_, new_n37416_, new_n37410_ );
nor  ( new_n37418_, new_n37417_, new_n37401_ );
nor  ( new_n37419_, new_n37418_, new_n37400_ );
or   ( new_n37420_, new_n37419_, new_n37367_ );
and  ( new_n37421_, new_n37420_, new_n37366_ );
or   ( new_n37422_, new_n37421_, new_n37287_ );
nand ( new_n37423_, new_n37421_, new_n37287_ );
xnor ( new_n37424_, new_n36868_, new_n36862_ );
xor  ( new_n37425_, new_n37424_, new_n36874_ );
xor  ( new_n37426_, new_n37177_, new_n37175_ );
xor  ( new_n37427_, new_n37426_, new_n37181_ );
nor  ( new_n37428_, new_n37427_, new_n37425_ );
and  ( new_n37429_, new_n37427_, new_n37425_ );
xor  ( new_n37430_, new_n37187_, new_n37185_ );
xnor ( new_n37431_, new_n37430_, new_n37191_ );
not  ( new_n37432_, new_n37431_ );
nor  ( new_n37433_, new_n37432_, new_n37429_ );
nor  ( new_n37434_, new_n37433_, new_n37428_ );
nand ( new_n37435_, new_n37434_, new_n37423_ );
and  ( new_n37436_, new_n37435_, new_n37422_ );
or   ( new_n37437_, new_n37436_, new_n37261_ );
nand ( new_n37438_, new_n37436_, new_n37261_ );
xor  ( new_n37439_, new_n37193_, new_n37183_ );
xor  ( new_n37440_, new_n37439_, new_n37197_ );
xor  ( new_n37441_, new_n37115_, new_n37075_ );
xor  ( new_n37442_, new_n37441_, new_n37169_ );
nor  ( new_n37443_, new_n37442_, new_n37440_ );
and  ( new_n37444_, new_n37442_, new_n37440_ );
xor  ( new_n37445_, new_n37205_, new_n37203_ );
xor  ( new_n37446_, new_n37445_, new_n37210_ );
nor  ( new_n37447_, new_n37446_, new_n37444_ );
nor  ( new_n37448_, new_n37447_, new_n37443_ );
nand ( new_n37449_, new_n37448_, new_n37438_ );
and  ( new_n37450_, new_n37449_, new_n37437_ );
or   ( new_n37451_, new_n37450_, new_n37243_ );
nand ( new_n37452_, new_n37450_, new_n37243_ );
xor  ( new_n37453_, new_n37199_, new_n37171_ );
xor  ( new_n37454_, new_n37453_, new_n37212_ );
xor  ( new_n37455_, new_n37220_, new_n37218_ );
xor  ( new_n37456_, new_n37455_, new_n37225_ );
nor  ( new_n37457_, new_n37456_, new_n37454_ );
and  ( new_n37458_, new_n37456_, new_n37454_ );
xor  ( new_n37459_, new_n37024_, new_n37022_ );
not  ( new_n37460_, new_n37459_ );
nor  ( new_n37461_, new_n37460_, new_n37458_ );
nor  ( new_n37462_, new_n37461_, new_n37457_ );
nand ( new_n37463_, new_n37462_, new_n37452_ );
and  ( new_n37464_, new_n37463_, new_n37451_ );
xnor ( new_n37465_, new_n36975_, new_n36798_ );
xor  ( new_n37466_, new_n37465_, new_n36988_ );
or   ( new_n37467_, new_n37466_, new_n37464_ );
and  ( new_n37468_, new_n37466_, new_n37464_ );
xor  ( new_n37469_, new_n37018_, new_n37006_ );
xor  ( new_n37470_, new_n37469_, new_n37230_ );
or   ( new_n37471_, new_n37470_, new_n37468_ );
and  ( new_n37472_, new_n37471_, new_n37467_ );
xor  ( new_n37473_, new_n37234_, new_n37232_ );
xor  ( new_n37474_, new_n37473_, new_n37238_ );
and  ( new_n37475_, new_n37474_, new_n37472_ );
xnor ( new_n37476_, new_n37466_, new_n37464_ );
xor  ( new_n37477_, new_n37476_, new_n37470_ );
xnor ( new_n37478_, new_n37442_, new_n37440_ );
xor  ( new_n37479_, new_n37478_, new_n37446_ );
or   ( new_n37480_, new_n6173_, new_n25288_ );
or   ( new_n37481_, new_n6175_, new_n25048_ );
and  ( new_n37482_, new_n37481_, new_n37480_ );
xor  ( new_n37483_, new_n37482_, new_n5597_ );
or   ( new_n37484_, new_n5604_, new_n25813_ );
or   ( new_n37485_, new_n5606_, new_n25486_ );
and  ( new_n37486_, new_n37485_, new_n37484_ );
xor  ( new_n37487_, new_n37486_, new_n5206_ );
or   ( new_n37488_, new_n37487_, new_n37483_ );
and  ( new_n37489_, new_n37487_, new_n37483_ );
or   ( new_n37490_, new_n5207_, new_n26063_ );
or   ( new_n37491_, new_n5209_, new_n26196_ );
and  ( new_n37492_, new_n37491_, new_n37490_ );
xor  ( new_n37493_, new_n37492_, new_n4708_ );
or   ( new_n37494_, new_n37493_, new_n37489_ );
and  ( new_n37495_, new_n37494_, new_n37488_ );
or   ( new_n37496_, new_n3461_, new_n28108_ );
or   ( new_n37497_, new_n3463_, new_n27763_ );
and  ( new_n37498_, new_n37497_, new_n37496_ );
xor  ( new_n37499_, new_n37498_, new_n3116_ );
or   ( new_n37500_, new_n3117_, new_n28531_ );
or   ( new_n37501_, new_n3119_, new_n28314_ );
and  ( new_n37502_, new_n37501_, new_n37500_ );
xor  ( new_n37503_, new_n37502_, new_n2800_ );
or   ( new_n37504_, new_n37503_, new_n37499_ );
and  ( new_n37505_, new_n37503_, new_n37499_ );
or   ( new_n37506_, new_n2807_, new_n29261_ );
or   ( new_n37507_, new_n2809_, new_n29263_ );
and  ( new_n37508_, new_n37507_, new_n37506_ );
xor  ( new_n37509_, new_n37508_, new_n2424_ );
or   ( new_n37510_, new_n37509_, new_n37505_ );
and  ( new_n37511_, new_n37510_, new_n37504_ );
or   ( new_n37512_, new_n37511_, new_n37495_ );
and  ( new_n37513_, new_n37511_, new_n37495_ );
or   ( new_n37514_, new_n4709_, new_n26620_ );
or   ( new_n37515_, new_n4711_, new_n26372_ );
and  ( new_n37516_, new_n37515_, new_n37514_ );
xor  ( new_n37517_, new_n37516_, new_n4295_ );
or   ( new_n37518_, new_n4302_, new_n27085_ );
or   ( new_n37519_, new_n4304_, new_n26762_ );
and  ( new_n37520_, new_n37519_, new_n37518_ );
xor  ( new_n37521_, new_n37520_, new_n3895_ );
nor  ( new_n37522_, new_n37521_, new_n37517_ );
and  ( new_n37523_, new_n37521_, new_n37517_ );
or   ( new_n37524_, new_n3896_, new_n27602_ );
or   ( new_n37525_, new_n3898_, new_n27396_ );
and  ( new_n37526_, new_n37525_, new_n37524_ );
xor  ( new_n37527_, new_n37526_, new_n3460_ );
nor  ( new_n37528_, new_n37527_, new_n37523_ );
nor  ( new_n37529_, new_n37528_, new_n37522_ );
or   ( new_n37530_, new_n37529_, new_n37513_ );
and  ( new_n37531_, new_n37530_, new_n37512_ );
or   ( new_n37532_, new_n1593_, new_n31654_ );
or   ( new_n37533_, new_n1595_, new_n31333_ );
and  ( new_n37534_, new_n37533_, new_n37532_ );
xor  ( new_n37535_, new_n37534_, new_n1358_ );
not  ( new_n37536_, new_n37535_ );
and  ( new_n37537_, new_n1251_, RIbb33378_192 );
or   ( new_n37538_, new_n37537_, new_n1129_ );
nand ( new_n37539_, new_n37537_, new_n1126_ );
and  ( new_n37540_, new_n37539_, new_n37538_ );
nor  ( new_n37541_, new_n37540_, new_n37536_ );
or   ( new_n37542_, new_n1364_, new_n31952_ );
or   ( new_n37543_, new_n1366_, new_n31654_ );
and  ( new_n37544_, new_n37543_, new_n37542_ );
xor  ( new_n37545_, new_n37544_, new_n1129_ );
or   ( new_n37546_, new_n37545_, new_n37541_ );
and  ( new_n37547_, new_n37545_, new_n37541_ );
or   ( new_n37548_, new_n2425_, new_n29619_ );
or   ( new_n37549_, new_n2427_, new_n29474_ );
and  ( new_n37550_, new_n37549_, new_n37548_ );
xor  ( new_n37551_, new_n37550_, new_n2121_ );
or   ( new_n37552_, new_n2122_, new_n30227_ );
or   ( new_n37553_, new_n2124_, new_n30120_ );
and  ( new_n37554_, new_n37553_, new_n37552_ );
xor  ( new_n37555_, new_n37554_, new_n1843_ );
nor  ( new_n37556_, new_n37555_, new_n37551_ );
and  ( new_n37557_, new_n37555_, new_n37551_ );
or   ( new_n37558_, new_n1844_, new_n30798_ );
or   ( new_n37559_, new_n1846_, new_n30800_ );
and  ( new_n37560_, new_n37559_, new_n37558_ );
xor  ( new_n37561_, new_n37560_, new_n1586_ );
nor  ( new_n37562_, new_n37561_, new_n37557_ );
nor  ( new_n37563_, new_n37562_, new_n37556_ );
or   ( new_n37564_, new_n37563_, new_n37547_ );
and  ( new_n37565_, new_n37564_, new_n37546_ );
nor  ( new_n37566_, new_n37565_, new_n37531_ );
nand ( new_n37567_, new_n37565_, new_n37531_ );
or   ( new_n37568_, new_n10059_, new_n22973_ );
or   ( new_n37569_, new_n10061_, new_n22975_ );
and  ( new_n37570_, new_n37569_, new_n37568_ );
xor  ( new_n37571_, new_n37570_, new_n9421_ );
and  ( new_n37572_, RIbb31fc8_150, RIbb2d888_64 );
or   ( new_n37573_, new_n22829_, RIbb2d888_64 );
and  ( new_n37574_, new_n37573_, RIbb2d900_63 );
or   ( new_n37575_, new_n37574_, new_n37572_ );
or   ( new_n37576_, new_n10770_, new_n22641_ );
and  ( new_n37577_, new_n37576_, new_n37575_ );
or   ( new_n37578_, new_n37577_, new_n37571_ );
and  ( new_n37579_, new_n37577_, new_n37571_ );
or   ( new_n37580_, new_n37579_, new_n1128_ );
and  ( new_n37581_, new_n37580_, new_n37578_ );
or   ( new_n37582_, new_n7732_, new_n24227_ );
or   ( new_n37583_, new_n7734_, new_n24006_ );
and  ( new_n37584_, new_n37583_, new_n37582_ );
xor  ( new_n37585_, new_n37584_, new_n7177_ );
or   ( new_n37586_, new_n7184_, new_n24543_ );
or   ( new_n37587_, new_n7186_, new_n24418_ );
and  ( new_n37588_, new_n37587_, new_n37586_ );
xor  ( new_n37589_, new_n37588_, new_n6638_ );
or   ( new_n37590_, new_n37589_, new_n37585_ );
and  ( new_n37591_, new_n37589_, new_n37585_ );
or   ( new_n37592_, new_n6645_, new_n24925_ );
or   ( new_n37593_, new_n6647_, new_n24927_ );
and  ( new_n37594_, new_n37593_, new_n37592_ );
xor  ( new_n37595_, new_n37594_, new_n6166_ );
or   ( new_n37596_, new_n37595_, new_n37591_ );
and  ( new_n37597_, new_n37596_, new_n37590_ );
nor  ( new_n37598_, new_n37597_, new_n37581_ );
and  ( new_n37599_, new_n37597_, new_n37581_ );
or   ( new_n37600_, new_n9422_, new_n23252_ );
or   ( new_n37601_, new_n9424_, new_n23166_ );
and  ( new_n37602_, new_n37601_, new_n37600_ );
xor  ( new_n37603_, new_n37602_, new_n8873_ );
or   ( new_n37604_, new_n8874_, new_n23554_ );
or   ( new_n37605_, new_n8876_, new_n23370_ );
and  ( new_n37606_, new_n37605_, new_n37604_ );
xor  ( new_n37607_, new_n37606_, new_n8257_ );
nor  ( new_n37608_, new_n37607_, new_n37603_ );
and  ( new_n37609_, new_n37607_, new_n37603_ );
or   ( new_n37610_, new_n8264_, new_n23895_ );
or   ( new_n37611_, new_n8266_, new_n23733_ );
and  ( new_n37612_, new_n37611_, new_n37610_ );
xor  ( new_n37613_, new_n37612_, new_n7725_ );
nor  ( new_n37614_, new_n37613_, new_n37609_ );
nor  ( new_n37615_, new_n37614_, new_n37608_ );
nor  ( new_n37616_, new_n37615_, new_n37599_ );
nor  ( new_n37617_, new_n37616_, new_n37598_ );
not  ( new_n37618_, new_n37617_ );
and  ( new_n37619_, new_n37618_, new_n37567_ );
or   ( new_n37620_, new_n37619_, new_n37566_ );
xor  ( new_n37621_, new_n37267_, new_n37265_ );
xor  ( new_n37622_, new_n37621_, new_n37271_ );
xnor ( new_n37623_, new_n37391_, new_n37387_ );
xor  ( new_n37624_, new_n37623_, new_n37397_ );
xnor ( new_n37625_, new_n37351_, new_n37347_ );
xor  ( new_n37626_, new_n37625_, new_n37357_ );
or   ( new_n37627_, new_n37626_, new_n37624_ );
and  ( new_n37628_, new_n37626_, new_n37624_ );
xnor ( new_n37629_, new_n37375_, new_n37371_ );
xor  ( new_n37630_, new_n37629_, new_n37381_ );
or   ( new_n37631_, new_n37630_, new_n37628_ );
and  ( new_n37632_, new_n37631_, new_n37627_ );
or   ( new_n37633_, new_n37632_, new_n37622_ );
and  ( new_n37634_, new_n37632_, new_n37622_ );
xnor ( new_n37635_, new_n37295_, new_n37291_ );
xor  ( new_n37636_, new_n37635_, new_n37301_ );
xnor ( new_n37637_, new_n37409_, new_n37405_ );
xor  ( new_n37638_, new_n37637_, new_n37415_ );
nor  ( new_n37639_, new_n37638_, new_n37636_ );
and  ( new_n37640_, new_n37638_, new_n37636_ );
xor  ( new_n37641_, new_n37331_, new_n37327_ );
xnor ( new_n37642_, new_n37641_, new_n37337_ );
nor  ( new_n37643_, new_n37642_, new_n37640_ );
nor  ( new_n37644_, new_n37643_, new_n37639_ );
or   ( new_n37645_, new_n37644_, new_n37634_ );
and  ( new_n37646_, new_n37645_, new_n37633_ );
nand ( new_n37647_, new_n37646_, new_n37620_ );
or   ( new_n37648_, new_n37646_, new_n37620_ );
xor  ( new_n37649_, new_n37399_, new_n37383_ );
xor  ( new_n37650_, new_n37649_, new_n37417_ );
xor  ( new_n37651_, new_n37279_, new_n37277_ );
xor  ( new_n37652_, new_n37651_, new_n37283_ );
and  ( new_n37653_, new_n37652_, new_n37650_ );
nor  ( new_n37654_, new_n37652_, new_n37650_ );
xor  ( new_n37655_, new_n37359_, new_n37343_ );
xnor ( new_n37656_, new_n37655_, new_n37363_ );
nor  ( new_n37657_, new_n37656_, new_n37654_ );
nor  ( new_n37658_, new_n37657_, new_n37653_ );
nand ( new_n37659_, new_n37658_, new_n37648_ );
and  ( new_n37660_, new_n37659_, new_n37647_ );
nor  ( new_n37661_, new_n37660_, new_n37479_ );
nand ( new_n37662_, new_n37660_, new_n37479_ );
xnor ( new_n37663_, new_n37249_, new_n37247_ );
xor  ( new_n37664_, new_n37663_, new_n37253_ );
xor  ( new_n37665_, new_n37273_, new_n37263_ );
xor  ( new_n37666_, new_n37665_, new_n37285_ );
nand ( new_n37667_, new_n37666_, new_n37664_ );
nor  ( new_n37668_, new_n37666_, new_n37664_ );
xor  ( new_n37669_, new_n37427_, new_n37425_ );
xor  ( new_n37670_, new_n37669_, new_n37432_ );
or   ( new_n37671_, new_n37670_, new_n37668_ );
and  ( new_n37672_, new_n37671_, new_n37667_ );
and  ( new_n37673_, new_n37672_, new_n37662_ );
or   ( new_n37674_, new_n37673_, new_n37661_ );
xor  ( new_n37675_, new_n37436_, new_n37261_ );
xor  ( new_n37676_, new_n37675_, new_n37448_ );
nor  ( new_n37677_, new_n37676_, new_n37674_ );
and  ( new_n37678_, new_n37676_, new_n37674_ );
xor  ( new_n37679_, new_n37456_, new_n37454_ );
xor  ( new_n37680_, new_n37679_, new_n37460_ );
nor  ( new_n37681_, new_n37680_, new_n37678_ );
or   ( new_n37682_, new_n37681_, new_n37677_ );
xnor ( new_n37683_, new_n37214_, new_n37025_ );
xor  ( new_n37684_, new_n37683_, new_n37227_ );
nand ( new_n37685_, new_n37684_, new_n37682_ );
nor  ( new_n37686_, new_n37684_, new_n37682_ );
xor  ( new_n37687_, new_n37450_, new_n37243_ );
xor  ( new_n37688_, new_n37687_, new_n37462_ );
or   ( new_n37689_, new_n37688_, new_n37686_ );
and  ( new_n37690_, new_n37689_, new_n37685_ );
nor  ( new_n37691_, new_n37690_, new_n37477_ );
xor  ( new_n37692_, new_n37684_, new_n37682_ );
xor  ( new_n37693_, new_n37692_, new_n37688_ );
xor  ( new_n37694_, new_n37421_, new_n37287_ );
xor  ( new_n37695_, new_n37694_, new_n37434_ );
xor  ( new_n37696_, new_n37660_, new_n37479_ );
xor  ( new_n37697_, new_n37696_, new_n37672_ );
or   ( new_n37698_, new_n37697_, new_n37695_ );
xor  ( new_n37699_, new_n37646_, new_n37620_ );
xor  ( new_n37700_, new_n37699_, new_n37658_ );
xnor ( new_n37701_, new_n37666_, new_n37664_ );
xnor ( new_n37702_, new_n37701_, new_n37670_ );
or   ( new_n37703_, new_n37702_, new_n37700_ );
xor  ( new_n37704_, new_n37321_, new_n37303_ );
xor  ( new_n37705_, new_n37704_, new_n37339_ );
xnor ( new_n37706_, new_n37632_, new_n37622_ );
xor  ( new_n37707_, new_n37706_, new_n37644_ );
nand ( new_n37708_, new_n37707_, new_n37705_ );
nor  ( new_n37709_, new_n37707_, new_n37705_ );
xor  ( new_n37710_, new_n37652_, new_n37650_ );
xor  ( new_n37711_, new_n37710_, new_n37656_ );
or   ( new_n37712_, new_n37711_, new_n37709_ );
and  ( new_n37713_, new_n37712_, new_n37708_ );
xnor ( new_n37714_, new_n37365_, new_n37341_ );
xor  ( new_n37715_, new_n37714_, new_n37419_ );
or   ( new_n37716_, new_n37715_, new_n37713_ );
and  ( new_n37717_, new_n37715_, new_n37713_ );
xnor ( new_n37718_, new_n37313_, new_n37307_ );
xor  ( new_n37719_, new_n37718_, new_n37319_ );
xnor ( new_n37720_, new_n37503_, new_n37499_ );
xor  ( new_n37721_, new_n37720_, new_n37509_ );
xnor ( new_n37722_, new_n37487_, new_n37483_ );
xor  ( new_n37723_, new_n37722_, new_n37493_ );
or   ( new_n37724_, new_n37723_, new_n37721_ );
and  ( new_n37725_, new_n37723_, new_n37721_ );
xor  ( new_n37726_, new_n37521_, new_n37517_ );
xnor ( new_n37727_, new_n37726_, new_n37527_ );
or   ( new_n37728_, new_n37727_, new_n37725_ );
and  ( new_n37729_, new_n37728_, new_n37724_ );
nor  ( new_n37730_, new_n37729_, new_n37719_ );
and  ( new_n37731_, new_n37729_, new_n37719_ );
xor  ( new_n37732_, new_n37577_, new_n37571_ );
xor  ( new_n37733_, new_n37732_, new_n1129_ );
xnor ( new_n37734_, new_n37589_, new_n37585_ );
xor  ( new_n37735_, new_n37734_, new_n37595_ );
nor  ( new_n37736_, new_n37735_, new_n37733_ );
and  ( new_n37737_, new_n37735_, new_n37733_ );
xor  ( new_n37738_, new_n37607_, new_n37603_ );
xnor ( new_n37739_, new_n37738_, new_n37613_ );
nor  ( new_n37740_, new_n37739_, new_n37737_ );
nor  ( new_n37741_, new_n37740_, new_n37736_ );
nor  ( new_n37742_, new_n37741_, new_n37731_ );
or   ( new_n37743_, new_n37742_, new_n37730_ );
xor  ( new_n37744_, new_n37626_, new_n37624_ );
xor  ( new_n37745_, new_n37744_, new_n37630_ );
xnor ( new_n37746_, new_n37545_, new_n37541_ );
xor  ( new_n37747_, new_n37746_, new_n37563_ );
nand ( new_n37748_, new_n37747_, new_n37745_ );
nor  ( new_n37749_, new_n37747_, new_n37745_ );
xor  ( new_n37750_, new_n37638_, new_n37636_ );
xnor ( new_n37751_, new_n37750_, new_n37642_ );
or   ( new_n37752_, new_n37751_, new_n37749_ );
and  ( new_n37753_, new_n37752_, new_n37748_ );
nor  ( new_n37754_, new_n37753_, new_n37743_ );
nand ( new_n37755_, new_n37753_, new_n37743_ );
or   ( new_n37756_, new_n3117_, new_n29263_ );
or   ( new_n37757_, new_n3119_, new_n28531_ );
and  ( new_n37758_, new_n37757_, new_n37756_ );
xor  ( new_n37759_, new_n37758_, new_n2800_ );
or   ( new_n37760_, new_n2807_, new_n29474_ );
or   ( new_n37761_, new_n2809_, new_n29261_ );
and  ( new_n37762_, new_n37761_, new_n37760_ );
xor  ( new_n37763_, new_n37762_, new_n2424_ );
or   ( new_n37764_, new_n37763_, new_n37759_ );
and  ( new_n37765_, new_n37763_, new_n37759_ );
or   ( new_n37766_, new_n2425_, new_n30120_ );
or   ( new_n37767_, new_n2427_, new_n29619_ );
and  ( new_n37768_, new_n37767_, new_n37766_ );
xor  ( new_n37769_, new_n37768_, new_n2121_ );
or   ( new_n37770_, new_n37769_, new_n37765_ );
and  ( new_n37771_, new_n37770_, new_n37764_ );
or   ( new_n37772_, new_n4302_, new_n27396_ );
or   ( new_n37773_, new_n4304_, new_n27085_ );
and  ( new_n37774_, new_n37773_, new_n37772_ );
xor  ( new_n37775_, new_n37774_, new_n3895_ );
or   ( new_n37776_, new_n3896_, new_n27763_ );
or   ( new_n37777_, new_n3898_, new_n27602_ );
and  ( new_n37778_, new_n37777_, new_n37776_ );
xor  ( new_n37779_, new_n37778_, new_n3460_ );
or   ( new_n37780_, new_n37779_, new_n37775_ );
and  ( new_n37781_, new_n37779_, new_n37775_ );
or   ( new_n37782_, new_n3461_, new_n28314_ );
or   ( new_n37783_, new_n3463_, new_n28108_ );
and  ( new_n37784_, new_n37783_, new_n37782_ );
xor  ( new_n37785_, new_n37784_, new_n3116_ );
or   ( new_n37786_, new_n37785_, new_n37781_ );
and  ( new_n37787_, new_n37786_, new_n37780_ );
or   ( new_n37788_, new_n37787_, new_n37771_ );
and  ( new_n37789_, new_n37787_, new_n37771_ );
or   ( new_n37790_, new_n5604_, new_n26196_ );
or   ( new_n37791_, new_n5606_, new_n25813_ );
and  ( new_n37792_, new_n37791_, new_n37790_ );
xor  ( new_n37793_, new_n37792_, new_n5206_ );
or   ( new_n37794_, new_n5207_, new_n26372_ );
or   ( new_n37795_, new_n5209_, new_n26063_ );
and  ( new_n37796_, new_n37795_, new_n37794_ );
xor  ( new_n37797_, new_n37796_, new_n4708_ );
or   ( new_n37798_, new_n37797_, new_n37793_ );
and  ( new_n37799_, new_n37797_, new_n37793_ );
or   ( new_n37800_, new_n4709_, new_n26762_ );
or   ( new_n37801_, new_n4711_, new_n26620_ );
and  ( new_n37802_, new_n37801_, new_n37800_ );
xor  ( new_n37803_, new_n37802_, new_n4295_ );
or   ( new_n37804_, new_n37803_, new_n37799_ );
and  ( new_n37805_, new_n37804_, new_n37798_ );
or   ( new_n37806_, new_n37805_, new_n37789_ );
and  ( new_n37807_, new_n37806_, new_n37788_ );
xor  ( new_n37808_, new_n37555_, new_n37551_ );
xor  ( new_n37809_, new_n37808_, new_n37561_ );
or   ( new_n37810_, new_n2122_, new_n30800_ );
or   ( new_n37811_, new_n2124_, new_n30227_ );
and  ( new_n37812_, new_n37811_, new_n37810_ );
xor  ( new_n37813_, new_n37812_, new_n1843_ );
or   ( new_n37814_, new_n1844_, new_n31333_ );
or   ( new_n37815_, new_n1846_, new_n30798_ );
and  ( new_n37816_, new_n37815_, new_n37814_ );
xor  ( new_n37817_, new_n37816_, new_n1586_ );
or   ( new_n37818_, new_n37817_, new_n37813_ );
and  ( new_n37819_, new_n37817_, new_n37813_ );
or   ( new_n37820_, new_n1593_, new_n31952_ );
or   ( new_n37821_, new_n1595_, new_n31654_ );
and  ( new_n37822_, new_n37821_, new_n37820_ );
xor  ( new_n37823_, new_n37822_, new_n1358_ );
or   ( new_n37824_, new_n37823_, new_n37819_ );
and  ( new_n37825_, new_n37824_, new_n37818_ );
or   ( new_n37826_, new_n37825_, new_n37809_ );
and  ( new_n37827_, new_n37825_, new_n37809_ );
xor  ( new_n37828_, new_n37540_, new_n37536_ );
or   ( new_n37829_, new_n37828_, new_n37827_ );
and  ( new_n37830_, new_n37829_, new_n37826_ );
nor  ( new_n37831_, new_n37830_, new_n37807_ );
nand ( new_n37832_, new_n37830_, new_n37807_ );
or   ( new_n37833_, new_n8874_, new_n23733_ );
or   ( new_n37834_, new_n8876_, new_n23554_ );
and  ( new_n37835_, new_n37834_, new_n37833_ );
xor  ( new_n37836_, new_n37835_, new_n8257_ );
or   ( new_n37837_, new_n8264_, new_n24006_ );
or   ( new_n37838_, new_n8266_, new_n23895_ );
and  ( new_n37839_, new_n37838_, new_n37837_ );
xor  ( new_n37840_, new_n37839_, new_n7725_ );
or   ( new_n37841_, new_n37840_, new_n37836_ );
and  ( new_n37842_, new_n37840_, new_n37836_ );
or   ( new_n37843_, new_n7732_, new_n24418_ );
or   ( new_n37844_, new_n7734_, new_n24227_ );
and  ( new_n37845_, new_n37844_, new_n37843_ );
xor  ( new_n37846_, new_n37845_, new_n7177_ );
or   ( new_n37847_, new_n37846_, new_n37842_ );
and  ( new_n37848_, new_n37847_, new_n37841_ );
or   ( new_n37849_, new_n7184_, new_n24927_ );
or   ( new_n37850_, new_n7186_, new_n24543_ );
and  ( new_n37851_, new_n37850_, new_n37849_ );
xor  ( new_n37852_, new_n37851_, new_n6638_ );
or   ( new_n37853_, new_n6645_, new_n25048_ );
or   ( new_n37854_, new_n6647_, new_n24925_ );
and  ( new_n37855_, new_n37854_, new_n37853_ );
xor  ( new_n37856_, new_n37855_, new_n6166_ );
or   ( new_n37857_, new_n37856_, new_n37852_ );
and  ( new_n37858_, new_n37856_, new_n37852_ );
or   ( new_n37859_, new_n6173_, new_n25486_ );
or   ( new_n37860_, new_n6175_, new_n25288_ );
and  ( new_n37861_, new_n37860_, new_n37859_ );
xor  ( new_n37862_, new_n37861_, new_n5597_ );
or   ( new_n37863_, new_n37862_, new_n37858_ );
and  ( new_n37864_, new_n37863_, new_n37857_ );
nor  ( new_n37865_, new_n37864_, new_n37848_ );
nand ( new_n37866_, new_n37864_, new_n37848_ );
or   ( new_n37867_, new_n10059_, new_n23166_ );
or   ( new_n37868_, new_n10061_, new_n22973_ );
and  ( new_n37869_, new_n37868_, new_n37867_ );
xor  ( new_n37870_, new_n37869_, new_n9421_ );
and  ( new_n37871_, RIbb32040_151, RIbb2d888_64 );
or   ( new_n37872_, new_n22975_, RIbb2d888_64 );
and  ( new_n37873_, new_n37872_, RIbb2d900_63 );
or   ( new_n37874_, new_n37873_, new_n37871_ );
or   ( new_n37875_, new_n10770_, new_n22829_ );
and  ( new_n37876_, new_n37875_, new_n37874_ );
nor  ( new_n37877_, new_n37876_, new_n37870_ );
nand ( new_n37878_, new_n37876_, new_n37870_ );
or   ( new_n37879_, new_n9422_, new_n23370_ );
or   ( new_n37880_, new_n9424_, new_n23252_ );
and  ( new_n37881_, new_n37880_, new_n37879_ );
xor  ( new_n37882_, new_n37881_, new_n8872_ );
and  ( new_n37883_, new_n37882_, new_n37878_ );
or   ( new_n37884_, new_n37883_, new_n37877_ );
and  ( new_n37885_, new_n37884_, new_n37866_ );
or   ( new_n37886_, new_n37885_, new_n37865_ );
and  ( new_n37887_, new_n37886_, new_n37832_ );
or   ( new_n37888_, new_n37887_, new_n37831_ );
and  ( new_n37889_, new_n37888_, new_n37755_ );
or   ( new_n37890_, new_n37889_, new_n37754_ );
or   ( new_n37891_, new_n37890_, new_n37717_ );
and  ( new_n37892_, new_n37891_, new_n37716_ );
or   ( new_n37893_, new_n37892_, new_n37703_ );
and  ( new_n37894_, new_n37892_, new_n37703_ );
xor  ( new_n37895_, new_n37255_, new_n37245_ );
xor  ( new_n37896_, new_n37895_, new_n37259_ );
or   ( new_n37897_, new_n37896_, new_n37894_ );
and  ( new_n37898_, new_n37897_, new_n37893_ );
or   ( new_n37899_, new_n37898_, new_n37698_ );
and  ( new_n37900_, new_n37898_, new_n37698_ );
xor  ( new_n37901_, new_n37676_, new_n37674_ );
xor  ( new_n37902_, new_n37901_, new_n37680_ );
or   ( new_n37903_, new_n37902_, new_n37900_ );
and  ( new_n37904_, new_n37903_, new_n37899_ );
nor  ( new_n37905_, new_n37904_, new_n37693_ );
xor  ( new_n37906_, new_n37898_, new_n37698_ );
xor  ( new_n37907_, new_n37906_, new_n37902_ );
xor  ( new_n37908_, new_n37892_, new_n37703_ );
xor  ( new_n37909_, new_n37908_, new_n37896_ );
xnor ( new_n37910_, new_n37511_, new_n37495_ );
xor  ( new_n37911_, new_n37910_, new_n37529_ );
xnor ( new_n37912_, new_n37597_, new_n37581_ );
xor  ( new_n37913_, new_n37912_, new_n37615_ );
nor  ( new_n37914_, new_n37913_, new_n37911_ );
and  ( new_n37915_, new_n37913_, new_n37911_ );
xor  ( new_n37916_, new_n37747_, new_n37745_ );
xnor ( new_n37917_, new_n37916_, new_n37751_ );
nor  ( new_n37918_, new_n37917_, new_n37915_ );
or   ( new_n37919_, new_n37918_, new_n37914_ );
xor  ( new_n37920_, new_n37817_, new_n37813_ );
xor  ( new_n37921_, new_n37920_, new_n37823_ );
or   ( new_n37922_, new_n2425_, new_n30227_ );
or   ( new_n37923_, new_n2427_, new_n30120_ );
and  ( new_n37924_, new_n37923_, new_n37922_ );
xor  ( new_n37925_, new_n37924_, new_n2121_ );
or   ( new_n37926_, new_n2122_, new_n30798_ );
or   ( new_n37927_, new_n2124_, new_n30800_ );
and  ( new_n37928_, new_n37927_, new_n37926_ );
xor  ( new_n37929_, new_n37928_, new_n1843_ );
or   ( new_n37930_, new_n37929_, new_n37925_ );
and  ( new_n37931_, new_n37929_, new_n37925_ );
or   ( new_n37932_, new_n1844_, new_n31654_ );
or   ( new_n37933_, new_n1846_, new_n31333_ );
and  ( new_n37934_, new_n37933_, new_n37932_ );
xor  ( new_n37935_, new_n37934_, new_n1586_ );
or   ( new_n37936_, new_n37935_, new_n37931_ );
and  ( new_n37937_, new_n37936_, new_n37930_ );
or   ( new_n37938_, new_n37937_, new_n37921_ );
nand ( new_n37939_, new_n37937_, new_n37921_ );
xor  ( new_n37940_, new_n37763_, new_n37759_ );
xnor ( new_n37941_, new_n37940_, new_n37769_ );
nand ( new_n37942_, new_n37941_, new_n37939_ );
and  ( new_n37943_, new_n37942_, new_n37938_ );
or   ( new_n37944_, new_n7732_, new_n24543_ );
or   ( new_n37945_, new_n7734_, new_n24418_ );
and  ( new_n37946_, new_n37945_, new_n37944_ );
xor  ( new_n37947_, new_n37946_, new_n7177_ );
or   ( new_n37948_, new_n7184_, new_n24925_ );
or   ( new_n37949_, new_n7186_, new_n24927_ );
and  ( new_n37950_, new_n37949_, new_n37948_ );
xor  ( new_n37951_, new_n37950_, new_n6638_ );
or   ( new_n37952_, new_n37951_, new_n37947_ );
and  ( new_n37953_, new_n37951_, new_n37947_ );
or   ( new_n37954_, new_n6645_, new_n25288_ );
or   ( new_n37955_, new_n6647_, new_n25048_ );
and  ( new_n37956_, new_n37955_, new_n37954_ );
xor  ( new_n37957_, new_n37956_, new_n6166_ );
or   ( new_n37958_, new_n37957_, new_n37953_ );
and  ( new_n37959_, new_n37958_, new_n37952_ );
or   ( new_n37960_, new_n10059_, new_n23252_ );
or   ( new_n37961_, new_n10061_, new_n23166_ );
and  ( new_n37962_, new_n37961_, new_n37960_ );
xor  ( new_n37963_, new_n37962_, new_n9421_ );
and  ( new_n37964_, RIbb320b8_152, RIbb2d888_64 );
or   ( new_n37965_, new_n22973_, RIbb2d888_64 );
and  ( new_n37966_, new_n37965_, RIbb2d900_63 );
or   ( new_n37967_, new_n37966_, new_n37964_ );
or   ( new_n37968_, new_n10770_, new_n22975_ );
and  ( new_n37969_, new_n37968_, new_n37967_ );
nor  ( new_n37970_, new_n37969_, new_n37963_ );
and  ( new_n37971_, new_n37969_, new_n37963_ );
nor  ( new_n37972_, new_n37971_, new_n1357_ );
nor  ( new_n37973_, new_n37972_, new_n37970_ );
or   ( new_n37974_, new_n9422_, new_n23554_ );
or   ( new_n37975_, new_n9424_, new_n23370_ );
and  ( new_n37976_, new_n37975_, new_n37974_ );
xor  ( new_n37977_, new_n37976_, new_n8873_ );
or   ( new_n37978_, new_n8874_, new_n23895_ );
or   ( new_n37979_, new_n8876_, new_n23733_ );
and  ( new_n37980_, new_n37979_, new_n37978_ );
xor  ( new_n37981_, new_n37980_, new_n8257_ );
or   ( new_n37982_, new_n37981_, new_n37977_ );
and  ( new_n37983_, new_n37981_, new_n37977_ );
or   ( new_n37984_, new_n8264_, new_n24227_ );
or   ( new_n37985_, new_n8266_, new_n24006_ );
and  ( new_n37986_, new_n37985_, new_n37984_ );
xor  ( new_n37987_, new_n37986_, new_n7725_ );
or   ( new_n37988_, new_n37987_, new_n37983_ );
and  ( new_n37989_, new_n37988_, new_n37982_ );
and  ( new_n37990_, new_n37989_, new_n37973_ );
or   ( new_n37991_, new_n37990_, new_n37959_ );
or   ( new_n37992_, new_n37989_, new_n37973_ );
and  ( new_n37993_, new_n37992_, new_n37991_ );
nor  ( new_n37994_, new_n37993_, new_n37943_ );
nand ( new_n37995_, new_n37993_, new_n37943_ );
or   ( new_n37996_, new_n6173_, new_n25813_ );
or   ( new_n37997_, new_n6175_, new_n25486_ );
and  ( new_n37998_, new_n37997_, new_n37996_ );
xor  ( new_n37999_, new_n37998_, new_n5597_ );
or   ( new_n38000_, new_n5604_, new_n26063_ );
or   ( new_n38001_, new_n5606_, new_n26196_ );
and  ( new_n38002_, new_n38001_, new_n38000_ );
xor  ( new_n38003_, new_n38002_, new_n5206_ );
or   ( new_n38004_, new_n38003_, new_n37999_ );
and  ( new_n38005_, new_n38003_, new_n37999_ );
or   ( new_n38006_, new_n5207_, new_n26620_ );
or   ( new_n38007_, new_n5209_, new_n26372_ );
and  ( new_n38008_, new_n38007_, new_n38006_ );
xor  ( new_n38009_, new_n38008_, new_n4708_ );
or   ( new_n38010_, new_n38009_, new_n38005_ );
and  ( new_n38011_, new_n38010_, new_n38004_ );
or   ( new_n38012_, new_n3461_, new_n28531_ );
or   ( new_n38013_, new_n3463_, new_n28314_ );
and  ( new_n38014_, new_n38013_, new_n38012_ );
xor  ( new_n38015_, new_n38014_, new_n3116_ );
or   ( new_n38016_, new_n3117_, new_n29261_ );
or   ( new_n38017_, new_n3119_, new_n29263_ );
and  ( new_n38018_, new_n38017_, new_n38016_ );
xor  ( new_n38019_, new_n38018_, new_n2800_ );
or   ( new_n38020_, new_n38019_, new_n38015_ );
and  ( new_n38021_, new_n38019_, new_n38015_ );
or   ( new_n38022_, new_n2807_, new_n29619_ );
or   ( new_n38023_, new_n2809_, new_n29474_ );
and  ( new_n38024_, new_n38023_, new_n38022_ );
xor  ( new_n38025_, new_n38024_, new_n2424_ );
or   ( new_n38026_, new_n38025_, new_n38021_ );
and  ( new_n38027_, new_n38026_, new_n38020_ );
nor  ( new_n38028_, new_n38027_, new_n38011_ );
and  ( new_n38029_, new_n38027_, new_n38011_ );
or   ( new_n38030_, new_n4709_, new_n27085_ );
or   ( new_n38031_, new_n4711_, new_n26762_ );
and  ( new_n38032_, new_n38031_, new_n38030_ );
xor  ( new_n38033_, new_n38032_, new_n4295_ );
or   ( new_n38034_, new_n4302_, new_n27602_ );
or   ( new_n38035_, new_n4304_, new_n27396_ );
and  ( new_n38036_, new_n38035_, new_n38034_ );
xor  ( new_n38037_, new_n38036_, new_n3895_ );
nor  ( new_n38038_, new_n38037_, new_n38033_ );
and  ( new_n38039_, new_n38037_, new_n38033_ );
or   ( new_n38040_, new_n3896_, new_n28108_ );
or   ( new_n38041_, new_n3898_, new_n27763_ );
and  ( new_n38042_, new_n38041_, new_n38040_ );
xor  ( new_n38043_, new_n38042_, new_n3460_ );
nor  ( new_n38044_, new_n38043_, new_n38039_ );
nor  ( new_n38045_, new_n38044_, new_n38038_ );
nor  ( new_n38046_, new_n38045_, new_n38029_ );
nor  ( new_n38047_, new_n38046_, new_n38028_ );
not  ( new_n38048_, new_n38047_ );
and  ( new_n38049_, new_n38048_, new_n37995_ );
or   ( new_n38050_, new_n38049_, new_n37994_ );
xor  ( new_n38051_, new_n37840_, new_n37836_ );
xnor ( new_n38052_, new_n38051_, new_n37846_ );
xor  ( new_n38053_, new_n37876_, new_n37870_ );
xor  ( new_n38054_, new_n38053_, new_n37882_ );
or   ( new_n38055_, new_n38054_, new_n38052_ );
xnor ( new_n38056_, new_n37779_, new_n37775_ );
xor  ( new_n38057_, new_n38056_, new_n37785_ );
xnor ( new_n38058_, new_n37856_, new_n37852_ );
xor  ( new_n38059_, new_n38058_, new_n37862_ );
or   ( new_n38060_, new_n38059_, new_n38057_ );
and  ( new_n38061_, new_n38059_, new_n38057_ );
xnor ( new_n38062_, new_n37797_, new_n37793_ );
xor  ( new_n38063_, new_n38062_, new_n37803_ );
or   ( new_n38064_, new_n38063_, new_n38061_ );
and  ( new_n38065_, new_n38064_, new_n38060_ );
or   ( new_n38066_, new_n38065_, new_n38055_ );
and  ( new_n38067_, new_n38065_, new_n38055_ );
xor  ( new_n38068_, new_n37735_, new_n37733_ );
xor  ( new_n38069_, new_n38068_, new_n37739_ );
or   ( new_n38070_, new_n38069_, new_n38067_ );
and  ( new_n38071_, new_n38070_, new_n38066_ );
nand ( new_n38072_, new_n38071_, new_n38050_ );
or   ( new_n38073_, new_n38071_, new_n38050_ );
xor  ( new_n38074_, new_n37787_, new_n37771_ );
xor  ( new_n38075_, new_n38074_, new_n37805_ );
xnor ( new_n38076_, new_n37723_, new_n37721_ );
xor  ( new_n38077_, new_n38076_, new_n37727_ );
and  ( new_n38078_, new_n38077_, new_n38075_ );
nor  ( new_n38079_, new_n38077_, new_n38075_ );
xor  ( new_n38080_, new_n37825_, new_n37809_ );
xnor ( new_n38081_, new_n38080_, new_n37828_ );
nor  ( new_n38082_, new_n38081_, new_n38079_ );
nor  ( new_n38083_, new_n38082_, new_n38078_ );
nand ( new_n38084_, new_n38083_, new_n38073_ );
and  ( new_n38085_, new_n38084_, new_n38072_ );
nor  ( new_n38086_, new_n38085_, new_n37919_ );
nand ( new_n38087_, new_n38085_, new_n37919_ );
xor  ( new_n38088_, new_n37565_, new_n37531_ );
xor  ( new_n38089_, new_n38088_, new_n37618_ );
and  ( new_n38090_, new_n38089_, new_n38087_ );
or   ( new_n38091_, new_n38090_, new_n38086_ );
xor  ( new_n38092_, new_n37715_, new_n37713_ );
xor  ( new_n38093_, new_n38092_, new_n37890_ );
or   ( new_n38094_, new_n38093_, new_n38091_ );
and  ( new_n38095_, new_n38093_, new_n38091_ );
xnor ( new_n38096_, new_n37702_, new_n37700_ );
or   ( new_n38097_, new_n38096_, new_n38095_ );
and  ( new_n38098_, new_n38097_, new_n38094_ );
or   ( new_n38099_, new_n38098_, new_n37909_ );
and  ( new_n38100_, new_n38098_, new_n37909_ );
xnor ( new_n38101_, new_n37697_, new_n37695_ );
or   ( new_n38102_, new_n38101_, new_n38100_ );
and  ( new_n38103_, new_n38102_, new_n38099_ );
nor  ( new_n38104_, new_n38103_, new_n37907_ );
xor  ( new_n38105_, new_n38098_, new_n37909_ );
xor  ( new_n38106_, new_n38105_, new_n38101_ );
xor  ( new_n38107_, new_n38085_, new_n37919_ );
xor  ( new_n38108_, new_n38107_, new_n38089_ );
xor  ( new_n38109_, new_n37753_, new_n37743_ );
xor  ( new_n38110_, new_n38109_, new_n37888_ );
or   ( new_n38111_, new_n38110_, new_n38108_ );
xor  ( new_n38112_, new_n37707_, new_n37705_ );
xor  ( new_n38113_, new_n38112_, new_n37711_ );
xor  ( new_n38114_, new_n37729_, new_n37719_ );
xor  ( new_n38115_, new_n38114_, new_n37741_ );
and  ( new_n38116_, new_n1474_, RIbb33378_192 );
or   ( new_n38117_, new_n38116_, new_n1358_ );
nand ( new_n38118_, new_n38116_, new_n1355_ );
and  ( new_n38119_, new_n38118_, new_n38117_ );
xnor ( new_n38120_, new_n37929_, new_n37925_ );
xor  ( new_n38121_, new_n38120_, new_n37935_ );
nor  ( new_n38122_, new_n38121_, new_n38119_ );
nand ( new_n38123_, new_n38121_, new_n38119_ );
xor  ( new_n38124_, new_n38019_, new_n38015_ );
xnor ( new_n38125_, new_n38124_, new_n38025_ );
not  ( new_n38126_, new_n38125_ );
and  ( new_n38127_, new_n38126_, new_n38123_ );
or   ( new_n38128_, new_n38127_, new_n38122_ );
or   ( new_n38129_, new_n8874_, new_n24006_ );
or   ( new_n38130_, new_n8876_, new_n23895_ );
and  ( new_n38131_, new_n38130_, new_n38129_ );
xor  ( new_n38132_, new_n38131_, new_n8257_ );
or   ( new_n38133_, new_n8264_, new_n24418_ );
or   ( new_n38134_, new_n8266_, new_n24227_ );
and  ( new_n38135_, new_n38134_, new_n38133_ );
xor  ( new_n38136_, new_n38135_, new_n7725_ );
or   ( new_n38137_, new_n38136_, new_n38132_ );
and  ( new_n38138_, new_n38136_, new_n38132_ );
or   ( new_n38139_, new_n7732_, new_n24927_ );
or   ( new_n38140_, new_n7734_, new_n24543_ );
and  ( new_n38141_, new_n38140_, new_n38139_ );
xor  ( new_n38142_, new_n38141_, new_n7177_ );
or   ( new_n38143_, new_n38142_, new_n38138_ );
and  ( new_n38144_, new_n38143_, new_n38137_ );
or   ( new_n38145_, new_n10059_, new_n23370_ );
or   ( new_n38146_, new_n10061_, new_n23252_ );
and  ( new_n38147_, new_n38146_, new_n38145_ );
xor  ( new_n38148_, new_n38147_, new_n9421_ );
and  ( new_n38149_, RIbb32130_153, RIbb2d888_64 );
or   ( new_n38150_, new_n23166_, RIbb2d888_64 );
and  ( new_n38151_, new_n38150_, RIbb2d900_63 );
or   ( new_n38152_, new_n38151_, new_n38149_ );
or   ( new_n38153_, new_n10770_, new_n22973_ );
and  ( new_n38154_, new_n38153_, new_n38152_ );
or   ( new_n38155_, new_n38154_, new_n38148_ );
and  ( new_n38156_, new_n38154_, new_n38148_ );
or   ( new_n38157_, new_n9422_, new_n23733_ );
or   ( new_n38158_, new_n9424_, new_n23554_ );
and  ( new_n38159_, new_n38158_, new_n38157_ );
xor  ( new_n38160_, new_n38159_, new_n8873_ );
or   ( new_n38161_, new_n38160_, new_n38156_ );
and  ( new_n38162_, new_n38161_, new_n38155_ );
or   ( new_n38163_, new_n38162_, new_n38144_ );
and  ( new_n38164_, new_n38162_, new_n38144_ );
or   ( new_n38165_, new_n7184_, new_n25048_ );
or   ( new_n38166_, new_n7186_, new_n24925_ );
and  ( new_n38167_, new_n38166_, new_n38165_ );
xor  ( new_n38168_, new_n38167_, new_n6638_ );
or   ( new_n38169_, new_n6645_, new_n25486_ );
or   ( new_n38170_, new_n6647_, new_n25288_ );
and  ( new_n38171_, new_n38170_, new_n38169_ );
xor  ( new_n38172_, new_n38171_, new_n6166_ );
nor  ( new_n38173_, new_n38172_, new_n38168_ );
and  ( new_n38174_, new_n38172_, new_n38168_ );
or   ( new_n38175_, new_n6173_, new_n26196_ );
or   ( new_n38176_, new_n6175_, new_n25813_ );
and  ( new_n38177_, new_n38176_, new_n38175_ );
xor  ( new_n38178_, new_n38177_, new_n5597_ );
nor  ( new_n38179_, new_n38178_, new_n38174_ );
nor  ( new_n38180_, new_n38179_, new_n38173_ );
or   ( new_n38181_, new_n38180_, new_n38164_ );
and  ( new_n38182_, new_n38181_, new_n38163_ );
nor  ( new_n38183_, new_n38182_, new_n38128_ );
nand ( new_n38184_, new_n38182_, new_n38128_ );
or   ( new_n38185_, new_n5604_, new_n26372_ );
or   ( new_n38186_, new_n5606_, new_n26063_ );
and  ( new_n38187_, new_n38186_, new_n38185_ );
xor  ( new_n38188_, new_n38187_, new_n5206_ );
or   ( new_n38189_, new_n5207_, new_n26762_ );
or   ( new_n38190_, new_n5209_, new_n26620_ );
and  ( new_n38191_, new_n38190_, new_n38189_ );
xor  ( new_n38192_, new_n38191_, new_n4708_ );
or   ( new_n38193_, new_n38192_, new_n38188_ );
and  ( new_n38194_, new_n38192_, new_n38188_ );
or   ( new_n38195_, new_n4709_, new_n27396_ );
or   ( new_n38196_, new_n4711_, new_n27085_ );
and  ( new_n38197_, new_n38196_, new_n38195_ );
xor  ( new_n38198_, new_n38197_, new_n4295_ );
or   ( new_n38199_, new_n38198_, new_n38194_ );
and  ( new_n38200_, new_n38199_, new_n38193_ );
or   ( new_n38201_, new_n4302_, new_n27763_ );
or   ( new_n38202_, new_n4304_, new_n27602_ );
and  ( new_n38203_, new_n38202_, new_n38201_ );
xor  ( new_n38204_, new_n38203_, new_n3895_ );
or   ( new_n38205_, new_n3896_, new_n28314_ );
or   ( new_n38206_, new_n3898_, new_n28108_ );
and  ( new_n38207_, new_n38206_, new_n38205_ );
xor  ( new_n38208_, new_n38207_, new_n3460_ );
or   ( new_n38209_, new_n38208_, new_n38204_ );
and  ( new_n38210_, new_n38208_, new_n38204_ );
or   ( new_n38211_, new_n3461_, new_n29263_ );
or   ( new_n38212_, new_n3463_, new_n28531_ );
and  ( new_n38213_, new_n38212_, new_n38211_ );
xor  ( new_n38214_, new_n38213_, new_n3116_ );
or   ( new_n38215_, new_n38214_, new_n38210_ );
and  ( new_n38216_, new_n38215_, new_n38209_ );
nor  ( new_n38217_, new_n38216_, new_n38200_ );
nand ( new_n38218_, new_n38216_, new_n38200_ );
or   ( new_n38219_, new_n3117_, new_n29474_ );
or   ( new_n38220_, new_n3119_, new_n29261_ );
and  ( new_n38221_, new_n38220_, new_n38219_ );
xor  ( new_n38222_, new_n38221_, new_n2800_ );
or   ( new_n38223_, new_n2807_, new_n30120_ );
or   ( new_n38224_, new_n2809_, new_n29619_ );
and  ( new_n38225_, new_n38224_, new_n38223_ );
xor  ( new_n38226_, new_n38225_, new_n2424_ );
nor  ( new_n38227_, new_n38226_, new_n38222_ );
nand ( new_n38228_, new_n38226_, new_n38222_ );
or   ( new_n38229_, new_n2425_, new_n30800_ );
or   ( new_n38230_, new_n2427_, new_n30227_ );
and  ( new_n38231_, new_n38230_, new_n38229_ );
xor  ( new_n38232_, new_n38231_, new_n2121_ );
not  ( new_n38233_, new_n38232_ );
and  ( new_n38234_, new_n38233_, new_n38228_ );
or   ( new_n38235_, new_n38234_, new_n38227_ );
and  ( new_n38236_, new_n38235_, new_n38218_ );
or   ( new_n38237_, new_n38236_, new_n38217_ );
and  ( new_n38238_, new_n38237_, new_n38184_ );
or   ( new_n38239_, new_n38238_, new_n38183_ );
xnor ( new_n38240_, new_n37989_, new_n37973_ );
xor  ( new_n38241_, new_n38240_, new_n37959_ );
xnor ( new_n38242_, new_n38027_, new_n38011_ );
xor  ( new_n38243_, new_n38242_, new_n38045_ );
or   ( new_n38244_, new_n38243_, new_n38241_ );
and  ( new_n38245_, new_n38243_, new_n38241_ );
xor  ( new_n38246_, new_n37937_, new_n37921_ );
xor  ( new_n38247_, new_n38246_, new_n37941_ );
or   ( new_n38248_, new_n38247_, new_n38245_ );
and  ( new_n38249_, new_n38248_, new_n38244_ );
and  ( new_n38250_, new_n38249_, new_n38239_ );
or   ( new_n38251_, new_n38249_, new_n38239_ );
xor  ( new_n38252_, new_n38059_, new_n38057_ );
xor  ( new_n38253_, new_n38252_, new_n38063_ );
xnor ( new_n38254_, new_n37951_, new_n37947_ );
xor  ( new_n38255_, new_n38254_, new_n37957_ );
xnor ( new_n38256_, new_n38003_, new_n37999_ );
xor  ( new_n38257_, new_n38256_, new_n38009_ );
or   ( new_n38258_, new_n38257_, new_n38255_ );
and  ( new_n38259_, new_n38257_, new_n38255_ );
xor  ( new_n38260_, new_n38037_, new_n38033_ );
xnor ( new_n38261_, new_n38260_, new_n38043_ );
or   ( new_n38262_, new_n38261_, new_n38259_ );
and  ( new_n38263_, new_n38262_, new_n38258_ );
nor  ( new_n38264_, new_n38263_, new_n38253_ );
and  ( new_n38265_, new_n38263_, new_n38253_ );
xor  ( new_n38266_, new_n38054_, new_n38052_ );
not  ( new_n38267_, new_n38266_ );
nor  ( new_n38268_, new_n38267_, new_n38265_ );
nor  ( new_n38269_, new_n38268_, new_n38264_ );
and  ( new_n38270_, new_n38269_, new_n38251_ );
or   ( new_n38271_, new_n38270_, new_n38250_ );
or   ( new_n38272_, new_n38271_, new_n38115_ );
and  ( new_n38273_, new_n38271_, new_n38115_ );
xor  ( new_n38274_, new_n37864_, new_n37848_ );
xor  ( new_n38275_, new_n38274_, new_n37884_ );
xor  ( new_n38276_, new_n38065_, new_n38055_ );
xor  ( new_n38277_, new_n38276_, new_n38069_ );
or   ( new_n38278_, new_n38277_, new_n38275_ );
and  ( new_n38279_, new_n38277_, new_n38275_ );
xor  ( new_n38280_, new_n38077_, new_n38075_ );
xor  ( new_n38281_, new_n38280_, new_n38081_ );
or   ( new_n38282_, new_n38281_, new_n38279_ );
and  ( new_n38283_, new_n38282_, new_n38278_ );
or   ( new_n38284_, new_n38283_, new_n38273_ );
and  ( new_n38285_, new_n38284_, new_n38272_ );
and  ( new_n38286_, new_n38285_, new_n38113_ );
xor  ( new_n38287_, new_n38071_, new_n38050_ );
xor  ( new_n38288_, new_n38287_, new_n38083_ );
xor  ( new_n38289_, new_n37830_, new_n37807_ );
xor  ( new_n38290_, new_n38289_, new_n37886_ );
or   ( new_n38291_, new_n38290_, new_n38288_ );
and  ( new_n38292_, new_n38290_, new_n38288_ );
xor  ( new_n38293_, new_n37913_, new_n37911_ );
xor  ( new_n38294_, new_n38293_, new_n37917_ );
or   ( new_n38295_, new_n38294_, new_n38292_ );
and  ( new_n38296_, new_n38295_, new_n38291_ );
or   ( new_n38297_, new_n38296_, new_n38286_ );
or   ( new_n38298_, new_n38285_, new_n38113_ );
and  ( new_n38299_, new_n38298_, new_n38297_ );
or   ( new_n38300_, new_n38299_, new_n38111_ );
and  ( new_n38301_, new_n38299_, new_n38111_ );
xor  ( new_n38302_, new_n38093_, new_n38091_ );
xor  ( new_n38303_, new_n38302_, new_n38096_ );
or   ( new_n38304_, new_n38303_, new_n38301_ );
and  ( new_n38305_, new_n38304_, new_n38300_ );
nor  ( new_n38306_, new_n38305_, new_n38106_ );
xor  ( new_n38307_, new_n38299_, new_n38111_ );
xor  ( new_n38308_, new_n38307_, new_n38303_ );
xor  ( new_n38309_, new_n38285_, new_n38113_ );
xor  ( new_n38310_, new_n38309_, new_n38296_ );
xor  ( new_n38311_, new_n38249_, new_n38239_ );
xor  ( new_n38312_, new_n38311_, new_n38269_ );
xor  ( new_n38313_, new_n38277_, new_n38275_ );
xor  ( new_n38314_, new_n38313_, new_n38281_ );
or   ( new_n38315_, new_n38314_, new_n38312_ );
xnor ( new_n38316_, new_n37981_, new_n37977_ );
xor  ( new_n38317_, new_n38316_, new_n37987_ );
xnor ( new_n38318_, new_n38208_, new_n38204_ );
xor  ( new_n38319_, new_n38318_, new_n38214_ );
xnor ( new_n38320_, new_n38192_, new_n38188_ );
xor  ( new_n38321_, new_n38320_, new_n38198_ );
or   ( new_n38322_, new_n38321_, new_n38319_ );
and  ( new_n38323_, new_n38321_, new_n38319_ );
xor  ( new_n38324_, new_n38226_, new_n38222_ );
xor  ( new_n38325_, new_n38324_, new_n38233_ );
or   ( new_n38326_, new_n38325_, new_n38323_ );
and  ( new_n38327_, new_n38326_, new_n38322_ );
nor  ( new_n38328_, new_n38327_, new_n38317_ );
and  ( new_n38329_, new_n38327_, new_n38317_ );
xnor ( new_n38330_, new_n38154_, new_n38148_ );
xor  ( new_n38331_, new_n38330_, new_n38160_ );
xnor ( new_n38332_, new_n38136_, new_n38132_ );
xor  ( new_n38333_, new_n38332_, new_n38142_ );
nor  ( new_n38334_, new_n38333_, new_n38331_ );
and  ( new_n38335_, new_n38333_, new_n38331_ );
xor  ( new_n38336_, new_n38172_, new_n38168_ );
xnor ( new_n38337_, new_n38336_, new_n38178_ );
nor  ( new_n38338_, new_n38337_, new_n38335_ );
nor  ( new_n38339_, new_n38338_, new_n38334_ );
nor  ( new_n38340_, new_n38339_, new_n38329_ );
nor  ( new_n38341_, new_n38340_, new_n38328_ );
or   ( new_n38342_, new_n3461_, new_n29261_ );
or   ( new_n38343_, new_n3463_, new_n29263_ );
and  ( new_n38344_, new_n38343_, new_n38342_ );
xor  ( new_n38345_, new_n38344_, new_n3116_ );
or   ( new_n38346_, new_n3117_, new_n29619_ );
or   ( new_n38347_, new_n3119_, new_n29474_ );
and  ( new_n38348_, new_n38347_, new_n38346_ );
xor  ( new_n38349_, new_n38348_, new_n2800_ );
or   ( new_n38350_, new_n38349_, new_n38345_ );
and  ( new_n38351_, new_n38349_, new_n38345_ );
or   ( new_n38352_, new_n2807_, new_n30227_ );
or   ( new_n38353_, new_n2809_, new_n30120_ );
and  ( new_n38354_, new_n38353_, new_n38352_ );
xor  ( new_n38355_, new_n38354_, new_n2424_ );
or   ( new_n38356_, new_n38355_, new_n38351_ );
and  ( new_n38357_, new_n38356_, new_n38350_ );
or   ( new_n38358_, new_n6173_, new_n26063_ );
or   ( new_n38359_, new_n6175_, new_n26196_ );
and  ( new_n38360_, new_n38359_, new_n38358_ );
xor  ( new_n38361_, new_n38360_, new_n5597_ );
or   ( new_n38362_, new_n5604_, new_n26620_ );
or   ( new_n38363_, new_n5606_, new_n26372_ );
and  ( new_n38364_, new_n38363_, new_n38362_ );
xor  ( new_n38365_, new_n38364_, new_n5206_ );
or   ( new_n38366_, new_n38365_, new_n38361_ );
and  ( new_n38367_, new_n38365_, new_n38361_ );
or   ( new_n38368_, new_n5207_, new_n27085_ );
or   ( new_n38369_, new_n5209_, new_n26762_ );
and  ( new_n38370_, new_n38369_, new_n38368_ );
xor  ( new_n38371_, new_n38370_, new_n4708_ );
or   ( new_n38372_, new_n38371_, new_n38367_ );
and  ( new_n38373_, new_n38372_, new_n38366_ );
nor  ( new_n38374_, new_n38373_, new_n38357_ );
and  ( new_n38375_, new_n38373_, new_n38357_ );
or   ( new_n38376_, new_n4709_, new_n27602_ );
or   ( new_n38377_, new_n4711_, new_n27396_ );
and  ( new_n38378_, new_n38377_, new_n38376_ );
xor  ( new_n38379_, new_n38378_, new_n4295_ );
or   ( new_n38380_, new_n4302_, new_n28108_ );
or   ( new_n38381_, new_n4304_, new_n27763_ );
and  ( new_n38382_, new_n38381_, new_n38380_ );
xor  ( new_n38383_, new_n38382_, new_n3895_ );
nor  ( new_n38384_, new_n38383_, new_n38379_ );
and  ( new_n38385_, new_n38383_, new_n38379_ );
or   ( new_n38386_, new_n3896_, new_n28531_ );
or   ( new_n38387_, new_n3898_, new_n28314_ );
and  ( new_n38388_, new_n38387_, new_n38386_ );
xor  ( new_n38389_, new_n38388_, new_n3460_ );
nor  ( new_n38390_, new_n38389_, new_n38385_ );
nor  ( new_n38391_, new_n38390_, new_n38384_ );
nor  ( new_n38392_, new_n38391_, new_n38375_ );
nor  ( new_n38393_, new_n38392_, new_n38374_ );
or   ( new_n38394_, new_n10059_, new_n23554_ );
or   ( new_n38395_, new_n10061_, new_n23370_ );
and  ( new_n38396_, new_n38395_, new_n38394_ );
xor  ( new_n38397_, new_n38396_, new_n9421_ );
and  ( new_n38398_, RIbb321a8_154, RIbb2d888_64 );
or   ( new_n38399_, new_n23252_, RIbb2d888_64 );
and  ( new_n38400_, new_n38399_, RIbb2d900_63 );
or   ( new_n38401_, new_n38400_, new_n38398_ );
or   ( new_n38402_, new_n10770_, new_n23166_ );
and  ( new_n38403_, new_n38402_, new_n38401_ );
or   ( new_n38404_, new_n38403_, new_n38397_ );
and  ( new_n38405_, new_n38403_, new_n38397_ );
or   ( new_n38406_, new_n38405_, new_n1585_ );
and  ( new_n38407_, new_n38406_, new_n38404_ );
or   ( new_n38408_, new_n7732_, new_n24925_ );
or   ( new_n38409_, new_n7734_, new_n24927_ );
and  ( new_n38410_, new_n38409_, new_n38408_ );
xor  ( new_n38411_, new_n38410_, new_n7177_ );
or   ( new_n38412_, new_n7184_, new_n25288_ );
or   ( new_n38413_, new_n7186_, new_n25048_ );
and  ( new_n38414_, new_n38413_, new_n38412_ );
xor  ( new_n38415_, new_n38414_, new_n6638_ );
or   ( new_n38416_, new_n38415_, new_n38411_ );
and  ( new_n38417_, new_n38415_, new_n38411_ );
or   ( new_n38418_, new_n6645_, new_n25813_ );
or   ( new_n38419_, new_n6647_, new_n25486_ );
and  ( new_n38420_, new_n38419_, new_n38418_ );
xor  ( new_n38421_, new_n38420_, new_n6166_ );
or   ( new_n38422_, new_n38421_, new_n38417_ );
and  ( new_n38423_, new_n38422_, new_n38416_ );
nor  ( new_n38424_, new_n38423_, new_n38407_ );
and  ( new_n38425_, new_n38423_, new_n38407_ );
or   ( new_n38426_, new_n9422_, new_n23895_ );
or   ( new_n38427_, new_n9424_, new_n23733_ );
and  ( new_n38428_, new_n38427_, new_n38426_ );
xor  ( new_n38429_, new_n38428_, new_n8873_ );
or   ( new_n38430_, new_n8874_, new_n24227_ );
or   ( new_n38431_, new_n8876_, new_n24006_ );
and  ( new_n38432_, new_n38431_, new_n38430_ );
xor  ( new_n38433_, new_n38432_, new_n8257_ );
nor  ( new_n38434_, new_n38433_, new_n38429_ );
and  ( new_n38435_, new_n38433_, new_n38429_ );
or   ( new_n38436_, new_n8264_, new_n24543_ );
or   ( new_n38437_, new_n8266_, new_n24418_ );
and  ( new_n38438_, new_n38437_, new_n38436_ );
xor  ( new_n38439_, new_n38438_, new_n7725_ );
nor  ( new_n38440_, new_n38439_, new_n38435_ );
nor  ( new_n38441_, new_n38440_, new_n38434_ );
nor  ( new_n38442_, new_n38441_, new_n38425_ );
nor  ( new_n38443_, new_n38442_, new_n38424_ );
and  ( new_n38444_, new_n38443_, new_n38393_ );
nor  ( new_n38445_, new_n38443_, new_n38393_ );
or   ( new_n38446_, new_n2122_, new_n31333_ );
or   ( new_n38447_, new_n2124_, new_n30798_ );
and  ( new_n38448_, new_n38447_, new_n38446_ );
xor  ( new_n38449_, new_n38448_, new_n1842_ );
or   ( new_n38450_, new_n2425_, new_n30798_ );
or   ( new_n38451_, new_n2427_, new_n30800_ );
and  ( new_n38452_, new_n38451_, new_n38450_ );
xor  ( new_n38453_, new_n38452_, new_n2121_ );
or   ( new_n38454_, new_n2122_, new_n31654_ );
or   ( new_n38455_, new_n2124_, new_n31333_ );
and  ( new_n38456_, new_n38455_, new_n38454_ );
xor  ( new_n38457_, new_n38456_, new_n1843_ );
nand ( new_n38458_, new_n38457_, new_n38453_ );
nor  ( new_n38459_, new_n38457_, new_n38453_ );
and  ( new_n38460_, new_n1739_, RIbb33378_192 );
or   ( new_n38461_, new_n38460_, new_n1586_ );
nand ( new_n38462_, new_n38460_, new_n1583_ );
and  ( new_n38463_, new_n38462_, new_n38461_ );
or   ( new_n38464_, new_n38463_, new_n38459_ );
and  ( new_n38465_, new_n38464_, new_n38458_ );
nor  ( new_n38466_, new_n38465_, new_n38449_ );
and  ( new_n38467_, new_n38465_, new_n38449_ );
not  ( new_n38468_, new_n38467_ );
or   ( new_n38469_, new_n1844_, new_n31952_ );
or   ( new_n38470_, new_n1846_, new_n31654_ );
and  ( new_n38471_, new_n38470_, new_n38469_ );
xor  ( new_n38472_, new_n38471_, new_n1586_ );
and  ( new_n38473_, new_n38472_, new_n38468_ );
nor  ( new_n38474_, new_n38473_, new_n38466_ );
nor  ( new_n38475_, new_n38474_, new_n38445_ );
nor  ( new_n38476_, new_n38475_, new_n38444_ );
and  ( new_n38477_, new_n38476_, new_n38341_ );
not  ( new_n38478_, new_n38477_ );
xor  ( new_n38479_, new_n37969_, new_n37963_ );
xor  ( new_n38480_, new_n38479_, new_n1357_ );
xnor ( new_n38481_, new_n38257_, new_n38255_ );
xor  ( new_n38482_, new_n38481_, new_n38261_ );
and  ( new_n38483_, new_n38482_, new_n38480_ );
nor  ( new_n38484_, new_n38482_, new_n38480_ );
xor  ( new_n38485_, new_n38121_, new_n38119_ );
xor  ( new_n38486_, new_n38485_, new_n38126_ );
not  ( new_n38487_, new_n38486_ );
nor  ( new_n38488_, new_n38487_, new_n38484_ );
nor  ( new_n38489_, new_n38488_, new_n38483_ );
not  ( new_n38490_, new_n38489_ );
and  ( new_n38491_, new_n38490_, new_n38478_ );
nor  ( new_n38492_, new_n38476_, new_n38341_ );
nor  ( new_n38493_, new_n38492_, new_n38491_ );
xor  ( new_n38494_, new_n38243_, new_n38241_ );
xor  ( new_n38495_, new_n38494_, new_n38247_ );
xor  ( new_n38496_, new_n38182_, new_n38128_ );
xor  ( new_n38497_, new_n38496_, new_n38237_ );
or   ( new_n38498_, new_n38497_, new_n38495_ );
nand ( new_n38499_, new_n38497_, new_n38495_ );
xor  ( new_n38500_, new_n38263_, new_n38253_ );
xor  ( new_n38501_, new_n38500_, new_n38266_ );
nand ( new_n38502_, new_n38501_, new_n38499_ );
and  ( new_n38503_, new_n38502_, new_n38498_ );
and  ( new_n38504_, new_n38503_, new_n38493_ );
xor  ( new_n38505_, new_n37993_, new_n37943_ );
xor  ( new_n38506_, new_n38505_, new_n38048_ );
or   ( new_n38507_, new_n38506_, new_n38504_ );
or   ( new_n38508_, new_n38503_, new_n38493_ );
and  ( new_n38509_, new_n38508_, new_n38507_ );
or   ( new_n38510_, new_n38509_, new_n38315_ );
and  ( new_n38511_, new_n38509_, new_n38315_ );
xor  ( new_n38512_, new_n38290_, new_n38288_ );
xor  ( new_n38513_, new_n38512_, new_n38294_ );
or   ( new_n38514_, new_n38513_, new_n38511_ );
and  ( new_n38515_, new_n38514_, new_n38510_ );
or   ( new_n38516_, new_n38515_, new_n38310_ );
and  ( new_n38517_, new_n38515_, new_n38310_ );
xnor ( new_n38518_, new_n38110_, new_n38108_ );
or   ( new_n38519_, new_n38518_, new_n38517_ );
and  ( new_n38520_, new_n38519_, new_n38516_ );
nor  ( new_n38521_, new_n38520_, new_n38308_ );
xor  ( new_n38522_, new_n38515_, new_n38310_ );
xor  ( new_n38523_, new_n38522_, new_n38518_ );
xor  ( new_n38524_, new_n38283_, new_n38115_ );
xor  ( new_n38525_, new_n38524_, new_n38271_ );
xor  ( new_n38526_, new_n38423_, new_n38407_ );
xor  ( new_n38527_, new_n38526_, new_n38441_ );
xor  ( new_n38528_, new_n38465_, new_n38449_ );
xor  ( new_n38529_, new_n38528_, new_n38472_ );
and  ( new_n38530_, new_n38529_, new_n38527_ );
nor  ( new_n38531_, new_n38529_, new_n38527_ );
xor  ( new_n38532_, new_n38373_, new_n38357_ );
xnor ( new_n38533_, new_n38532_, new_n38391_ );
nor  ( new_n38534_, new_n38533_, new_n38531_ );
nor  ( new_n38535_, new_n38534_, new_n38530_ );
or   ( new_n38536_, new_n8874_, new_n24418_ );
or   ( new_n38537_, new_n8876_, new_n24227_ );
and  ( new_n38538_, new_n38537_, new_n38536_ );
xor  ( new_n38539_, new_n38538_, new_n8257_ );
or   ( new_n38540_, new_n8264_, new_n24927_ );
or   ( new_n38541_, new_n8266_, new_n24543_ );
and  ( new_n38542_, new_n38541_, new_n38540_ );
xor  ( new_n38543_, new_n38542_, new_n7725_ );
or   ( new_n38544_, new_n38543_, new_n38539_ );
and  ( new_n38545_, new_n38543_, new_n38539_ );
or   ( new_n38546_, new_n7732_, new_n25048_ );
or   ( new_n38547_, new_n7734_, new_n24925_ );
and  ( new_n38548_, new_n38547_, new_n38546_ );
xor  ( new_n38549_, new_n38548_, new_n7177_ );
or   ( new_n38550_, new_n38549_, new_n38545_ );
and  ( new_n38551_, new_n38550_, new_n38544_ );
or   ( new_n38552_, new_n7184_, new_n25486_ );
or   ( new_n38553_, new_n7186_, new_n25288_ );
and  ( new_n38554_, new_n38553_, new_n38552_ );
xor  ( new_n38555_, new_n38554_, new_n6638_ );
or   ( new_n38556_, new_n6645_, new_n26196_ );
or   ( new_n38557_, new_n6647_, new_n25813_ );
and  ( new_n38558_, new_n38557_, new_n38556_ );
xor  ( new_n38559_, new_n38558_, new_n6166_ );
or   ( new_n38560_, new_n38559_, new_n38555_ );
and  ( new_n38561_, new_n38559_, new_n38555_ );
or   ( new_n38562_, new_n6173_, new_n26372_ );
or   ( new_n38563_, new_n6175_, new_n26063_ );
and  ( new_n38564_, new_n38563_, new_n38562_ );
xor  ( new_n38565_, new_n38564_, new_n5597_ );
or   ( new_n38566_, new_n38565_, new_n38561_ );
and  ( new_n38567_, new_n38566_, new_n38560_ );
nor  ( new_n38568_, new_n38567_, new_n38551_ );
and  ( new_n38569_, new_n38567_, new_n38551_ );
or   ( new_n38570_, new_n10059_, new_n23733_ );
or   ( new_n38571_, new_n10061_, new_n23554_ );
and  ( new_n38572_, new_n38571_, new_n38570_ );
xor  ( new_n38573_, new_n38572_, new_n9421_ );
and  ( new_n38574_, RIbb32220_155, RIbb2d888_64 );
or   ( new_n38575_, new_n23370_, RIbb2d888_64 );
and  ( new_n38576_, new_n38575_, RIbb2d900_63 );
or   ( new_n38577_, new_n38576_, new_n38574_ );
or   ( new_n38578_, new_n10770_, new_n23252_ );
and  ( new_n38579_, new_n38578_, new_n38577_ );
nor  ( new_n38580_, new_n38579_, new_n38573_ );
and  ( new_n38581_, new_n38579_, new_n38573_ );
or   ( new_n38582_, new_n9422_, new_n24006_ );
or   ( new_n38583_, new_n9424_, new_n23895_ );
and  ( new_n38584_, new_n38583_, new_n38582_ );
xor  ( new_n38585_, new_n38584_, new_n8873_ );
nor  ( new_n38586_, new_n38585_, new_n38581_ );
nor  ( new_n38587_, new_n38586_, new_n38580_ );
nor  ( new_n38588_, new_n38587_, new_n38569_ );
nor  ( new_n38589_, new_n38588_, new_n38568_ );
or   ( new_n38590_, new_n5604_, new_n26762_ );
or   ( new_n38591_, new_n5606_, new_n26620_ );
and  ( new_n38592_, new_n38591_, new_n38590_ );
xor  ( new_n38593_, new_n38592_, new_n5206_ );
or   ( new_n38594_, new_n5207_, new_n27396_ );
or   ( new_n38595_, new_n5209_, new_n27085_ );
and  ( new_n38596_, new_n38595_, new_n38594_ );
xor  ( new_n38597_, new_n38596_, new_n4708_ );
or   ( new_n38598_, new_n38597_, new_n38593_ );
and  ( new_n38599_, new_n38597_, new_n38593_ );
or   ( new_n38600_, new_n4709_, new_n27763_ );
or   ( new_n38601_, new_n4711_, new_n27602_ );
and  ( new_n38602_, new_n38601_, new_n38600_ );
xor  ( new_n38603_, new_n38602_, new_n4295_ );
or   ( new_n38604_, new_n38603_, new_n38599_ );
and  ( new_n38605_, new_n38604_, new_n38598_ );
or   ( new_n38606_, new_n3117_, new_n30120_ );
or   ( new_n38607_, new_n3119_, new_n29619_ );
and  ( new_n38608_, new_n38607_, new_n38606_ );
xor  ( new_n38609_, new_n38608_, new_n2800_ );
or   ( new_n38610_, new_n2807_, new_n30800_ );
or   ( new_n38611_, new_n2809_, new_n30227_ );
and  ( new_n38612_, new_n38611_, new_n38610_ );
xor  ( new_n38613_, new_n38612_, new_n2424_ );
or   ( new_n38614_, new_n38613_, new_n38609_ );
and  ( new_n38615_, new_n38613_, new_n38609_ );
or   ( new_n38616_, new_n2425_, new_n31333_ );
or   ( new_n38617_, new_n2427_, new_n30798_ );
and  ( new_n38618_, new_n38617_, new_n38616_ );
xor  ( new_n38619_, new_n38618_, new_n2121_ );
or   ( new_n38620_, new_n38619_, new_n38615_ );
and  ( new_n38621_, new_n38620_, new_n38614_ );
nor  ( new_n38622_, new_n38621_, new_n38605_ );
and  ( new_n38623_, new_n38621_, new_n38605_ );
or   ( new_n38624_, new_n4302_, new_n28314_ );
or   ( new_n38625_, new_n4304_, new_n28108_ );
and  ( new_n38626_, new_n38625_, new_n38624_ );
xor  ( new_n38627_, new_n38626_, new_n3895_ );
or   ( new_n38628_, new_n3896_, new_n29263_ );
or   ( new_n38629_, new_n3898_, new_n28531_ );
and  ( new_n38630_, new_n38629_, new_n38628_ );
xor  ( new_n38631_, new_n38630_, new_n3460_ );
nor  ( new_n38632_, new_n38631_, new_n38627_ );
and  ( new_n38633_, new_n38631_, new_n38627_ );
or   ( new_n38634_, new_n3461_, new_n29474_ );
or   ( new_n38635_, new_n3463_, new_n29261_ );
and  ( new_n38636_, new_n38635_, new_n38634_ );
xor  ( new_n38637_, new_n38636_, new_n3116_ );
nor  ( new_n38638_, new_n38637_, new_n38633_ );
nor  ( new_n38639_, new_n38638_, new_n38632_ );
nor  ( new_n38640_, new_n38639_, new_n38623_ );
nor  ( new_n38641_, new_n38640_, new_n38622_ );
and  ( new_n38642_, new_n38641_, new_n38589_ );
nor  ( new_n38643_, new_n38641_, new_n38589_ );
xor  ( new_n38644_, new_n38457_, new_n38453_ );
xor  ( new_n38645_, new_n38644_, new_n38463_ );
xnor ( new_n38646_, new_n38349_, new_n38345_ );
xor  ( new_n38647_, new_n38646_, new_n38355_ );
nor  ( new_n38648_, new_n38647_, new_n38645_ );
and  ( new_n38649_, new_n38647_, new_n38645_ );
xor  ( new_n38650_, new_n38383_, new_n38379_ );
xnor ( new_n38651_, new_n38650_, new_n38389_ );
nor  ( new_n38652_, new_n38651_, new_n38649_ );
nor  ( new_n38653_, new_n38652_, new_n38648_ );
nor  ( new_n38654_, new_n38653_, new_n38643_ );
nor  ( new_n38655_, new_n38654_, new_n38642_ );
and  ( new_n38656_, new_n38655_, new_n38535_ );
not  ( new_n38657_, new_n38656_ );
xor  ( new_n38658_, new_n38333_, new_n38331_ );
xor  ( new_n38659_, new_n38658_, new_n38337_ );
xnor ( new_n38660_, new_n38365_, new_n38361_ );
xor  ( new_n38661_, new_n38660_, new_n38371_ );
xnor ( new_n38662_, new_n38415_, new_n38411_ );
xor  ( new_n38663_, new_n38662_, new_n38421_ );
or   ( new_n38664_, new_n38663_, new_n38661_ );
and  ( new_n38665_, new_n38663_, new_n38661_ );
xnor ( new_n38666_, new_n38433_, new_n38429_ );
xor  ( new_n38667_, new_n38666_, new_n38439_ );
or   ( new_n38668_, new_n38667_, new_n38665_ );
and  ( new_n38669_, new_n38668_, new_n38664_ );
nor  ( new_n38670_, new_n38669_, new_n38659_ );
and  ( new_n38671_, new_n38669_, new_n38659_ );
xor  ( new_n38672_, new_n38321_, new_n38319_ );
xnor ( new_n38673_, new_n38672_, new_n38325_ );
not  ( new_n38674_, new_n38673_ );
nor  ( new_n38675_, new_n38674_, new_n38671_ );
nor  ( new_n38676_, new_n38675_, new_n38670_ );
not  ( new_n38677_, new_n38676_ );
and  ( new_n38678_, new_n38677_, new_n38657_ );
nor  ( new_n38679_, new_n38655_, new_n38535_ );
or   ( new_n38680_, new_n38679_, new_n38678_ );
xor  ( new_n38681_, new_n38497_, new_n38495_ );
xor  ( new_n38682_, new_n38681_, new_n38501_ );
or   ( new_n38683_, new_n38682_, new_n38680_ );
nand ( new_n38684_, new_n38682_, new_n38680_ );
xnor ( new_n38685_, new_n38162_, new_n38144_ );
xor  ( new_n38686_, new_n38685_, new_n38180_ );
xor  ( new_n38687_, new_n38216_, new_n38200_ );
xor  ( new_n38688_, new_n38687_, new_n38235_ );
nor  ( new_n38689_, new_n38688_, new_n38686_ );
and  ( new_n38690_, new_n38688_, new_n38686_ );
xor  ( new_n38691_, new_n38482_, new_n38480_ );
xor  ( new_n38692_, new_n38691_, new_n38486_ );
not  ( new_n38693_, new_n38692_ );
nor  ( new_n38694_, new_n38693_, new_n38690_ );
nor  ( new_n38695_, new_n38694_, new_n38689_ );
nand ( new_n38696_, new_n38695_, new_n38684_ );
and  ( new_n38697_, new_n38696_, new_n38683_ );
xnor ( new_n38698_, new_n38503_, new_n38493_ );
xor  ( new_n38699_, new_n38698_, new_n38506_ );
nand ( new_n38700_, new_n38699_, new_n38697_ );
nor  ( new_n38701_, new_n38699_, new_n38697_ );
xnor ( new_n38702_, new_n38314_, new_n38312_ );
or   ( new_n38703_, new_n38702_, new_n38701_ );
and  ( new_n38704_, new_n38703_, new_n38700_ );
or   ( new_n38705_, new_n38704_, new_n38525_ );
and  ( new_n38706_, new_n38704_, new_n38525_ );
xor  ( new_n38707_, new_n38509_, new_n38315_ );
xor  ( new_n38708_, new_n38707_, new_n38513_ );
or   ( new_n38709_, new_n38708_, new_n38706_ );
and  ( new_n38710_, new_n38709_, new_n38705_ );
nor  ( new_n38711_, new_n38710_, new_n38523_ );
xor  ( new_n38712_, new_n38655_, new_n38535_ );
or   ( new_n38713_, new_n38712_, new_n38677_ );
not  ( new_n38714_, new_n38678_ );
or   ( new_n38715_, new_n38679_, new_n38714_ );
and  ( new_n38716_, new_n38715_, new_n38713_ );
xnor ( new_n38717_, new_n38443_, new_n38393_ );
xor  ( new_n38718_, new_n38717_, new_n38474_ );
nand ( new_n38719_, new_n38718_, new_n38716_ );
nor  ( new_n38720_, new_n38718_, new_n38716_ );
xor  ( new_n38721_, new_n38688_, new_n38686_ );
xor  ( new_n38722_, new_n38721_, new_n38693_ );
or   ( new_n38723_, new_n38722_, new_n38720_ );
and  ( new_n38724_, new_n38723_, new_n38719_ );
or   ( new_n38725_, new_n2122_, new_n31952_ );
or   ( new_n38726_, new_n2124_, new_n31654_ );
and  ( new_n38727_, new_n38726_, new_n38725_ );
xor  ( new_n38728_, new_n38727_, new_n1842_ );
xnor ( new_n38729_, new_n38613_, new_n38609_ );
xor  ( new_n38730_, new_n38729_, new_n38619_ );
nand ( new_n38731_, new_n38730_, new_n38728_ );
or   ( new_n38732_, new_n38730_, new_n38728_ );
xor  ( new_n38733_, new_n38631_, new_n38627_ );
xnor ( new_n38734_, new_n38733_, new_n38637_ );
nand ( new_n38735_, new_n38734_, new_n38732_ );
and  ( new_n38736_, new_n38735_, new_n38731_ );
or   ( new_n38737_, new_n7732_, new_n25288_ );
or   ( new_n38738_, new_n7734_, new_n25048_ );
and  ( new_n38739_, new_n38738_, new_n38737_ );
xor  ( new_n38740_, new_n38739_, new_n7177_ );
or   ( new_n38741_, new_n7184_, new_n25813_ );
or   ( new_n38742_, new_n7186_, new_n25486_ );
and  ( new_n38743_, new_n38742_, new_n38741_ );
xor  ( new_n38744_, new_n38743_, new_n6638_ );
nor  ( new_n38745_, new_n38744_, new_n38740_ );
and  ( new_n38746_, new_n38744_, new_n38740_ );
or   ( new_n38747_, new_n6645_, new_n26063_ );
or   ( new_n38748_, new_n6647_, new_n26196_ );
and  ( new_n38749_, new_n38748_, new_n38747_ );
xor  ( new_n38750_, new_n38749_, new_n6166_ );
nor  ( new_n38751_, new_n38750_, new_n38746_ );
nor  ( new_n38752_, new_n38751_, new_n38745_ );
or   ( new_n38753_, new_n10059_, new_n23895_ );
or   ( new_n38754_, new_n10061_, new_n23733_ );
and  ( new_n38755_, new_n38754_, new_n38753_ );
xor  ( new_n38756_, new_n38755_, new_n9421_ );
and  ( new_n38757_, RIbb32298_156, RIbb2d888_64 );
or   ( new_n38758_, new_n23554_, RIbb2d888_64 );
and  ( new_n38759_, new_n38758_, RIbb2d900_63 );
or   ( new_n38760_, new_n38759_, new_n38757_ );
or   ( new_n38761_, new_n10770_, new_n23370_ );
and  ( new_n38762_, new_n38761_, new_n38760_ );
nor  ( new_n38763_, new_n38762_, new_n38756_ );
and  ( new_n38764_, new_n38762_, new_n38756_ );
nor  ( new_n38765_, new_n38764_, new_n1842_ );
nor  ( new_n38766_, new_n38765_, new_n38763_ );
or   ( new_n38767_, new_n9422_, new_n24227_ );
or   ( new_n38768_, new_n9424_, new_n24006_ );
and  ( new_n38769_, new_n38768_, new_n38767_ );
xor  ( new_n38770_, new_n38769_, new_n8873_ );
or   ( new_n38771_, new_n8874_, new_n24543_ );
or   ( new_n38772_, new_n8876_, new_n24418_ );
and  ( new_n38773_, new_n38772_, new_n38771_ );
xor  ( new_n38774_, new_n38773_, new_n8257_ );
or   ( new_n38775_, new_n38774_, new_n38770_ );
and  ( new_n38776_, new_n38774_, new_n38770_ );
or   ( new_n38777_, new_n8264_, new_n24925_ );
or   ( new_n38778_, new_n8266_, new_n24927_ );
and  ( new_n38779_, new_n38778_, new_n38777_ );
xor  ( new_n38780_, new_n38779_, new_n7725_ );
or   ( new_n38781_, new_n38780_, new_n38776_ );
and  ( new_n38782_, new_n38781_, new_n38775_ );
and  ( new_n38783_, new_n38782_, new_n38766_ );
or   ( new_n38784_, new_n38783_, new_n38752_ );
or   ( new_n38785_, new_n38782_, new_n38766_ );
and  ( new_n38786_, new_n38785_, new_n38784_ );
nor  ( new_n38787_, new_n38786_, new_n38736_ );
nand ( new_n38788_, new_n38786_, new_n38736_ );
or   ( new_n38789_, new_n6173_, new_n26620_ );
or   ( new_n38790_, new_n6175_, new_n26372_ );
and  ( new_n38791_, new_n38790_, new_n38789_ );
xor  ( new_n38792_, new_n38791_, new_n5597_ );
or   ( new_n38793_, new_n5604_, new_n27085_ );
or   ( new_n38794_, new_n5606_, new_n26762_ );
and  ( new_n38795_, new_n38794_, new_n38793_ );
xor  ( new_n38796_, new_n38795_, new_n5206_ );
or   ( new_n38797_, new_n38796_, new_n38792_ );
and  ( new_n38798_, new_n38796_, new_n38792_ );
or   ( new_n38799_, new_n5207_, new_n27602_ );
or   ( new_n38800_, new_n5209_, new_n27396_ );
and  ( new_n38801_, new_n38800_, new_n38799_ );
xor  ( new_n38802_, new_n38801_, new_n4708_ );
or   ( new_n38803_, new_n38802_, new_n38798_ );
and  ( new_n38804_, new_n38803_, new_n38797_ );
or   ( new_n38805_, new_n3461_, new_n29619_ );
or   ( new_n38806_, new_n3463_, new_n29474_ );
and  ( new_n38807_, new_n38806_, new_n38805_ );
xor  ( new_n38808_, new_n38807_, new_n3116_ );
or   ( new_n38809_, new_n3117_, new_n30227_ );
or   ( new_n38810_, new_n3119_, new_n30120_ );
and  ( new_n38811_, new_n38810_, new_n38809_ );
xor  ( new_n38812_, new_n38811_, new_n2800_ );
or   ( new_n38813_, new_n38812_, new_n38808_ );
and  ( new_n38814_, new_n38812_, new_n38808_ );
or   ( new_n38815_, new_n2807_, new_n30798_ );
or   ( new_n38816_, new_n2809_, new_n30800_ );
and  ( new_n38817_, new_n38816_, new_n38815_ );
xor  ( new_n38818_, new_n38817_, new_n2424_ );
or   ( new_n38819_, new_n38818_, new_n38814_ );
and  ( new_n38820_, new_n38819_, new_n38813_ );
nor  ( new_n38821_, new_n38820_, new_n38804_ );
and  ( new_n38822_, new_n38820_, new_n38804_ );
or   ( new_n38823_, new_n4709_, new_n28108_ );
or   ( new_n38824_, new_n4711_, new_n27763_ );
and  ( new_n38825_, new_n38824_, new_n38823_ );
xor  ( new_n38826_, new_n38825_, new_n4295_ );
or   ( new_n38827_, new_n4302_, new_n28531_ );
or   ( new_n38828_, new_n4304_, new_n28314_ );
and  ( new_n38829_, new_n38828_, new_n38827_ );
xor  ( new_n38830_, new_n38829_, new_n3895_ );
nor  ( new_n38831_, new_n38830_, new_n38826_ );
and  ( new_n38832_, new_n38830_, new_n38826_ );
or   ( new_n38833_, new_n3896_, new_n29261_ );
or   ( new_n38834_, new_n3898_, new_n29263_ );
and  ( new_n38835_, new_n38834_, new_n38833_ );
xor  ( new_n38836_, new_n38835_, new_n3460_ );
nor  ( new_n38837_, new_n38836_, new_n38832_ );
nor  ( new_n38838_, new_n38837_, new_n38831_ );
nor  ( new_n38839_, new_n38838_, new_n38822_ );
or   ( new_n38840_, new_n38839_, new_n38821_ );
and  ( new_n38841_, new_n38840_, new_n38788_ );
or   ( new_n38842_, new_n38841_, new_n38787_ );
xor  ( new_n38843_, new_n38403_, new_n38397_ );
xor  ( new_n38844_, new_n38843_, new_n1586_ );
xnor ( new_n38845_, new_n38559_, new_n38555_ );
xor  ( new_n38846_, new_n38845_, new_n38565_ );
xnor ( new_n38847_, new_n38597_, new_n38593_ );
xor  ( new_n38848_, new_n38847_, new_n38603_ );
or   ( new_n38849_, new_n38848_, new_n38846_ );
and  ( new_n38850_, new_n38848_, new_n38846_ );
xor  ( new_n38851_, new_n38543_, new_n38539_ );
xnor ( new_n38852_, new_n38851_, new_n38549_ );
or   ( new_n38853_, new_n38852_, new_n38850_ );
and  ( new_n38854_, new_n38853_, new_n38849_ );
or   ( new_n38855_, new_n38854_, new_n38844_ );
and  ( new_n38856_, new_n38854_, new_n38844_ );
xor  ( new_n38857_, new_n38663_, new_n38661_ );
xor  ( new_n38858_, new_n38857_, new_n38667_ );
or   ( new_n38859_, new_n38858_, new_n38856_ );
and  ( new_n38860_, new_n38859_, new_n38855_ );
and  ( new_n38861_, new_n38860_, new_n38842_ );
or   ( new_n38862_, new_n38860_, new_n38842_ );
xnor ( new_n38863_, new_n38621_, new_n38605_ );
xor  ( new_n38864_, new_n38863_, new_n38639_ );
xnor ( new_n38865_, new_n38567_, new_n38551_ );
xor  ( new_n38866_, new_n38865_, new_n38587_ );
or   ( new_n38867_, new_n38866_, new_n38864_ );
and  ( new_n38868_, new_n38866_, new_n38864_ );
xor  ( new_n38869_, new_n38647_, new_n38645_ );
xnor ( new_n38870_, new_n38869_, new_n38651_ );
not  ( new_n38871_, new_n38870_ );
or   ( new_n38872_, new_n38871_, new_n38868_ );
and  ( new_n38873_, new_n38872_, new_n38867_ );
and  ( new_n38874_, new_n38873_, new_n38862_ );
or   ( new_n38875_, new_n38874_, new_n38861_ );
xnor ( new_n38876_, new_n38641_, new_n38589_ );
xor  ( new_n38877_, new_n38876_, new_n38653_ );
xnor ( new_n38878_, new_n38529_, new_n38527_ );
xor  ( new_n38879_, new_n38878_, new_n38533_ );
nand ( new_n38880_, new_n38879_, new_n38877_ );
nor  ( new_n38881_, new_n38879_, new_n38877_ );
xor  ( new_n38882_, new_n38669_, new_n38659_ );
xor  ( new_n38883_, new_n38882_, new_n38674_ );
or   ( new_n38884_, new_n38883_, new_n38881_ );
and  ( new_n38885_, new_n38884_, new_n38880_ );
or   ( new_n38886_, new_n38885_, new_n38875_ );
and  ( new_n38887_, new_n38885_, new_n38875_ );
xor  ( new_n38888_, new_n38327_, new_n38317_ );
xor  ( new_n38889_, new_n38888_, new_n38339_ );
or   ( new_n38890_, new_n38889_, new_n38887_ );
and  ( new_n38891_, new_n38890_, new_n38886_ );
nor  ( new_n38892_, new_n38891_, new_n38724_ );
and  ( new_n38893_, new_n38891_, new_n38724_ );
xor  ( new_n38894_, new_n38476_, new_n38341_ );
nor  ( new_n38895_, new_n38894_, new_n38490_ );
not  ( new_n38896_, new_n38492_ );
and  ( new_n38897_, new_n38896_, new_n38491_ );
nor  ( new_n38898_, new_n38897_, new_n38895_ );
not  ( new_n38899_, new_n38898_ );
nor  ( new_n38900_, new_n38899_, new_n38893_ );
nor  ( new_n38901_, new_n38900_, new_n38892_ );
xor  ( new_n38902_, new_n38699_, new_n38697_ );
xor  ( new_n38903_, new_n38902_, new_n38702_ );
or   ( new_n38904_, new_n38903_, new_n38901_ );
xor  ( new_n38905_, new_n38704_, new_n38525_ );
xor  ( new_n38906_, new_n38905_, new_n38708_ );
nor  ( new_n38907_, new_n38906_, new_n38904_ );
xnor ( new_n38908_, new_n38903_, new_n38901_ );
xor  ( new_n38909_, new_n38891_, new_n38724_ );
xor  ( new_n38910_, new_n38909_, new_n38899_ );
xnor ( new_n38911_, new_n38879_, new_n38877_ );
xor  ( new_n38912_, new_n38911_, new_n38883_ );
or   ( new_n38913_, new_n8874_, new_n24927_ );
or   ( new_n38914_, new_n8876_, new_n24543_ );
and  ( new_n38915_, new_n38914_, new_n38913_ );
xor  ( new_n38916_, new_n38915_, new_n8257_ );
or   ( new_n38917_, new_n8264_, new_n25048_ );
or   ( new_n38918_, new_n8266_, new_n24925_ );
and  ( new_n38919_, new_n38918_, new_n38917_ );
xor  ( new_n38920_, new_n38919_, new_n7725_ );
or   ( new_n38921_, new_n38920_, new_n38916_ );
and  ( new_n38922_, new_n38920_, new_n38916_ );
or   ( new_n38923_, new_n7732_, new_n25486_ );
or   ( new_n38924_, new_n7734_, new_n25288_ );
and  ( new_n38925_, new_n38924_, new_n38923_ );
xor  ( new_n38926_, new_n38925_, new_n7177_ );
or   ( new_n38927_, new_n38926_, new_n38922_ );
and  ( new_n38928_, new_n38927_, new_n38921_ );
or   ( new_n38929_, new_n10059_, new_n24006_ );
or   ( new_n38930_, new_n10061_, new_n23895_ );
and  ( new_n38931_, new_n38930_, new_n38929_ );
xor  ( new_n38932_, new_n38931_, new_n9421_ );
and  ( new_n38933_, RIbb32310_157, RIbb2d888_64 );
or   ( new_n38934_, new_n23733_, RIbb2d888_64 );
and  ( new_n38935_, new_n38934_, RIbb2d900_63 );
or   ( new_n38936_, new_n38935_, new_n38933_ );
or   ( new_n38937_, new_n10770_, new_n23554_ );
and  ( new_n38938_, new_n38937_, new_n38936_ );
or   ( new_n38939_, new_n38938_, new_n38932_ );
and  ( new_n38940_, new_n38938_, new_n38932_ );
or   ( new_n38941_, new_n9422_, new_n24418_ );
or   ( new_n38942_, new_n9424_, new_n24227_ );
and  ( new_n38943_, new_n38942_, new_n38941_ );
xor  ( new_n38944_, new_n38943_, new_n8873_ );
or   ( new_n38945_, new_n38944_, new_n38940_ );
and  ( new_n38946_, new_n38945_, new_n38939_ );
or   ( new_n38947_, new_n38946_, new_n38928_ );
and  ( new_n38948_, new_n38946_, new_n38928_ );
or   ( new_n38949_, new_n7184_, new_n26196_ );
or   ( new_n38950_, new_n7186_, new_n25813_ );
and  ( new_n38951_, new_n38950_, new_n38949_ );
xor  ( new_n38952_, new_n38951_, new_n6638_ );
or   ( new_n38953_, new_n6645_, new_n26372_ );
or   ( new_n38954_, new_n6647_, new_n26063_ );
and  ( new_n38955_, new_n38954_, new_n38953_ );
xor  ( new_n38956_, new_n38955_, new_n6166_ );
nor  ( new_n38957_, new_n38956_, new_n38952_ );
and  ( new_n38958_, new_n38956_, new_n38952_ );
or   ( new_n38959_, new_n6173_, new_n26762_ );
or   ( new_n38960_, new_n6175_, new_n26620_ );
and  ( new_n38961_, new_n38960_, new_n38959_ );
xor  ( new_n38962_, new_n38961_, new_n5597_ );
nor  ( new_n38963_, new_n38962_, new_n38958_ );
nor  ( new_n38964_, new_n38963_, new_n38957_ );
or   ( new_n38965_, new_n38964_, new_n38948_ );
and  ( new_n38966_, new_n38965_, new_n38947_ );
or   ( new_n38967_, new_n2425_, new_n31654_ );
or   ( new_n38968_, new_n2427_, new_n31333_ );
and  ( new_n38969_, new_n38968_, new_n38967_ );
xor  ( new_n38970_, new_n38969_, new_n2120_ );
and  ( new_n38971_, new_n2000_, RIbb33378_192 );
or   ( new_n38972_, new_n38971_, new_n1843_ );
nand ( new_n38973_, new_n38971_, new_n1840_ );
and  ( new_n38974_, new_n38973_, new_n38972_ );
nand ( new_n38975_, new_n38974_, new_n38970_ );
or   ( new_n38976_, new_n38974_, new_n38970_ );
xor  ( new_n38977_, new_n38812_, new_n38808_ );
xnor ( new_n38978_, new_n38977_, new_n38818_ );
nand ( new_n38979_, new_n38978_, new_n38976_ );
and  ( new_n38980_, new_n38979_, new_n38975_ );
nor  ( new_n38981_, new_n38980_, new_n38966_ );
nand ( new_n38982_, new_n38980_, new_n38966_ );
or   ( new_n38983_, new_n4302_, new_n29263_ );
or   ( new_n38984_, new_n4304_, new_n28531_ );
and  ( new_n38985_, new_n38984_, new_n38983_ );
xor  ( new_n38986_, new_n38985_, new_n3895_ );
or   ( new_n38987_, new_n3896_, new_n29474_ );
or   ( new_n38988_, new_n3898_, new_n29261_ );
and  ( new_n38989_, new_n38988_, new_n38987_ );
xor  ( new_n38990_, new_n38989_, new_n3460_ );
or   ( new_n38991_, new_n38990_, new_n38986_ );
and  ( new_n38992_, new_n38990_, new_n38986_ );
or   ( new_n38993_, new_n3461_, new_n30120_ );
or   ( new_n38994_, new_n3463_, new_n29619_ );
and  ( new_n38995_, new_n38994_, new_n38993_ );
xor  ( new_n38996_, new_n38995_, new_n3116_ );
or   ( new_n38997_, new_n38996_, new_n38992_ );
and  ( new_n38998_, new_n38997_, new_n38991_ );
or   ( new_n38999_, new_n3117_, new_n30800_ );
or   ( new_n39000_, new_n3119_, new_n30227_ );
and  ( new_n39001_, new_n39000_, new_n38999_ );
xor  ( new_n39002_, new_n39001_, new_n2800_ );
or   ( new_n39003_, new_n2807_, new_n31333_ );
or   ( new_n39004_, new_n2809_, new_n30798_ );
and  ( new_n39005_, new_n39004_, new_n39003_ );
xor  ( new_n39006_, new_n39005_, new_n2424_ );
or   ( new_n39007_, new_n39006_, new_n39002_ );
and  ( new_n39008_, new_n39006_, new_n39002_ );
or   ( new_n39009_, new_n2425_, new_n31952_ );
or   ( new_n39010_, new_n2427_, new_n31654_ );
and  ( new_n39011_, new_n39010_, new_n39009_ );
xor  ( new_n39012_, new_n39011_, new_n2121_ );
or   ( new_n39013_, new_n39012_, new_n39008_ );
and  ( new_n39014_, new_n39013_, new_n39007_ );
nor  ( new_n39015_, new_n39014_, new_n38998_ );
nand ( new_n39016_, new_n39014_, new_n38998_ );
or   ( new_n39017_, new_n5604_, new_n27396_ );
or   ( new_n39018_, new_n5606_, new_n27085_ );
and  ( new_n39019_, new_n39018_, new_n39017_ );
xor  ( new_n39020_, new_n39019_, new_n5206_ );
or   ( new_n39021_, new_n5207_, new_n27763_ );
or   ( new_n39022_, new_n5209_, new_n27602_ );
and  ( new_n39023_, new_n39022_, new_n39021_ );
xor  ( new_n39024_, new_n39023_, new_n4708_ );
nor  ( new_n39025_, new_n39024_, new_n39020_ );
nand ( new_n39026_, new_n39024_, new_n39020_ );
or   ( new_n39027_, new_n4709_, new_n28314_ );
or   ( new_n39028_, new_n4711_, new_n28108_ );
and  ( new_n39029_, new_n39028_, new_n39027_ );
xor  ( new_n39030_, new_n39029_, new_n4295_ );
not  ( new_n39031_, new_n39030_ );
and  ( new_n39032_, new_n39031_, new_n39026_ );
or   ( new_n39033_, new_n39032_, new_n39025_ );
and  ( new_n39034_, new_n39033_, new_n39016_ );
or   ( new_n39035_, new_n39034_, new_n39015_ );
and  ( new_n39036_, new_n39035_, new_n38982_ );
or   ( new_n39037_, new_n39036_, new_n38981_ );
xor  ( new_n39038_, new_n38774_, new_n38770_ );
xnor ( new_n39039_, new_n39038_, new_n38780_ );
xor  ( new_n39040_, new_n38762_, new_n38756_ );
xor  ( new_n39041_, new_n39040_, new_n1843_ );
or   ( new_n39042_, new_n39041_, new_n39039_ );
xnor ( new_n39043_, new_n38744_, new_n38740_ );
xor  ( new_n39044_, new_n39043_, new_n38750_ );
xnor ( new_n39045_, new_n38796_, new_n38792_ );
xor  ( new_n39046_, new_n39045_, new_n38802_ );
or   ( new_n39047_, new_n39046_, new_n39044_ );
and  ( new_n39048_, new_n39046_, new_n39044_ );
xnor ( new_n39049_, new_n38830_, new_n38826_ );
xor  ( new_n39050_, new_n39049_, new_n38836_ );
or   ( new_n39051_, new_n39050_, new_n39048_ );
and  ( new_n39052_, new_n39051_, new_n39047_ );
or   ( new_n39053_, new_n39052_, new_n39042_ );
and  ( new_n39054_, new_n39052_, new_n39042_ );
xor  ( new_n39055_, new_n38579_, new_n38573_ );
xnor ( new_n39056_, new_n39055_, new_n38585_ );
or   ( new_n39057_, new_n39056_, new_n39054_ );
and  ( new_n39058_, new_n39057_, new_n39053_ );
nand ( new_n39059_, new_n39058_, new_n39037_ );
or   ( new_n39060_, new_n39058_, new_n39037_ );
xor  ( new_n39061_, new_n38820_, new_n38804_ );
xor  ( new_n39062_, new_n39061_, new_n38838_ );
xnor ( new_n39063_, new_n38848_, new_n38846_ );
xor  ( new_n39064_, new_n39063_, new_n38852_ );
and  ( new_n39065_, new_n39064_, new_n39062_ );
nor  ( new_n39066_, new_n39064_, new_n39062_ );
xor  ( new_n39067_, new_n38730_, new_n38728_ );
xor  ( new_n39068_, new_n39067_, new_n38734_ );
nor  ( new_n39069_, new_n39068_, new_n39066_ );
nor  ( new_n39070_, new_n39069_, new_n39065_ );
nand ( new_n39071_, new_n39070_, new_n39060_ );
and  ( new_n39072_, new_n39071_, new_n39059_ );
nor  ( new_n39073_, new_n39072_, new_n38912_ );
nand ( new_n39074_, new_n39072_, new_n38912_ );
xor  ( new_n39075_, new_n38854_, new_n38844_ );
xor  ( new_n39076_, new_n39075_, new_n38858_ );
xor  ( new_n39077_, new_n38786_, new_n38736_ );
xor  ( new_n39078_, new_n39077_, new_n38840_ );
nor  ( new_n39079_, new_n39078_, new_n39076_ );
and  ( new_n39080_, new_n39078_, new_n39076_ );
xor  ( new_n39081_, new_n38866_, new_n38864_ );
xor  ( new_n39082_, new_n39081_, new_n38871_ );
nor  ( new_n39083_, new_n39082_, new_n39080_ );
nor  ( new_n39084_, new_n39083_, new_n39079_ );
and  ( new_n39085_, new_n39084_, new_n39074_ );
or   ( new_n39086_, new_n39085_, new_n39073_ );
xor  ( new_n39087_, new_n38885_, new_n38875_ );
xor  ( new_n39088_, new_n39087_, new_n38889_ );
or   ( new_n39089_, new_n39088_, new_n39086_ );
and  ( new_n39090_, new_n39088_, new_n39086_ );
xor  ( new_n39091_, new_n38718_, new_n38716_ );
xor  ( new_n39092_, new_n39091_, new_n38722_ );
or   ( new_n39093_, new_n39092_, new_n39090_ );
and  ( new_n39094_, new_n39093_, new_n39089_ );
or   ( new_n39095_, new_n39094_, new_n38910_ );
and  ( new_n39096_, new_n39094_, new_n38910_ );
xor  ( new_n39097_, new_n38682_, new_n38680_ );
xor  ( new_n39098_, new_n39097_, new_n38695_ );
or   ( new_n39099_, new_n39098_, new_n39096_ );
and  ( new_n39100_, new_n39099_, new_n39095_ );
nor  ( new_n39101_, new_n39100_, new_n38908_ );
xor  ( new_n39102_, new_n39088_, new_n39086_ );
xor  ( new_n39103_, new_n39102_, new_n39092_ );
xor  ( new_n39104_, new_n38860_, new_n38842_ );
xor  ( new_n39105_, new_n39104_, new_n38873_ );
xnor ( new_n39106_, new_n38946_, new_n38928_ );
xor  ( new_n39107_, new_n39106_, new_n38964_ );
xor  ( new_n39108_, new_n39014_, new_n38998_ );
xor  ( new_n39109_, new_n39108_, new_n39033_ );
nor  ( new_n39110_, new_n39109_, new_n39107_ );
and  ( new_n39111_, new_n39109_, new_n39107_ );
xor  ( new_n39112_, new_n38974_, new_n38970_ );
xor  ( new_n39113_, new_n39112_, new_n38978_ );
nor  ( new_n39114_, new_n39113_, new_n39111_ );
nor  ( new_n39115_, new_n39114_, new_n39110_ );
or   ( new_n39116_, new_n4709_, new_n28531_ );
or   ( new_n39117_, new_n4711_, new_n28314_ );
and  ( new_n39118_, new_n39117_, new_n39116_ );
xor  ( new_n39119_, new_n39118_, new_n4295_ );
or   ( new_n39120_, new_n4302_, new_n29261_ );
or   ( new_n39121_, new_n4304_, new_n29263_ );
and  ( new_n39122_, new_n39121_, new_n39120_ );
xor  ( new_n39123_, new_n39122_, new_n3895_ );
or   ( new_n39124_, new_n39123_, new_n39119_ );
and  ( new_n39125_, new_n39123_, new_n39119_ );
or   ( new_n39126_, new_n3896_, new_n29619_ );
or   ( new_n39127_, new_n3898_, new_n29474_ );
and  ( new_n39128_, new_n39127_, new_n39126_ );
xor  ( new_n39129_, new_n39128_, new_n3460_ );
or   ( new_n39130_, new_n39129_, new_n39125_ );
and  ( new_n39131_, new_n39130_, new_n39124_ );
or   ( new_n39132_, new_n6173_, new_n27085_ );
or   ( new_n39133_, new_n6175_, new_n26762_ );
and  ( new_n39134_, new_n39133_, new_n39132_ );
xor  ( new_n39135_, new_n39134_, new_n5597_ );
or   ( new_n39136_, new_n5604_, new_n27602_ );
or   ( new_n39137_, new_n5606_, new_n27396_ );
and  ( new_n39138_, new_n39137_, new_n39136_ );
xor  ( new_n39139_, new_n39138_, new_n5206_ );
or   ( new_n39140_, new_n39139_, new_n39135_ );
and  ( new_n39141_, new_n39139_, new_n39135_ );
or   ( new_n39142_, new_n5207_, new_n28108_ );
or   ( new_n39143_, new_n5209_, new_n27763_ );
and  ( new_n39144_, new_n39143_, new_n39142_ );
xor  ( new_n39145_, new_n39144_, new_n4708_ );
or   ( new_n39146_, new_n39145_, new_n39141_ );
and  ( new_n39147_, new_n39146_, new_n39140_ );
nor  ( new_n39148_, new_n39147_, new_n39131_ );
and  ( new_n39149_, new_n39147_, new_n39131_ );
or   ( new_n39150_, new_n3461_, new_n30227_ );
or   ( new_n39151_, new_n3463_, new_n30120_ );
and  ( new_n39152_, new_n39151_, new_n39150_ );
xor  ( new_n39153_, new_n39152_, new_n3116_ );
or   ( new_n39154_, new_n3117_, new_n30798_ );
or   ( new_n39155_, new_n3119_, new_n30800_ );
and  ( new_n39156_, new_n39155_, new_n39154_ );
xor  ( new_n39157_, new_n39156_, new_n2800_ );
nor  ( new_n39158_, new_n39157_, new_n39153_ );
and  ( new_n39159_, new_n39157_, new_n39153_ );
or   ( new_n39160_, new_n2807_, new_n31654_ );
or   ( new_n39161_, new_n2809_, new_n31333_ );
and  ( new_n39162_, new_n39161_, new_n39160_ );
xor  ( new_n39163_, new_n39162_, new_n2424_ );
nor  ( new_n39164_, new_n39163_, new_n39159_ );
nor  ( new_n39165_, new_n39164_, new_n39158_ );
nor  ( new_n39166_, new_n39165_, new_n39149_ );
nor  ( new_n39167_, new_n39166_, new_n39148_ );
or   ( new_n39168_, new_n10059_, new_n24227_ );
or   ( new_n39169_, new_n10061_, new_n24006_ );
and  ( new_n39170_, new_n39169_, new_n39168_ );
xor  ( new_n39171_, new_n39170_, new_n9421_ );
and  ( new_n39172_, RIbb32388_158, RIbb2d888_64 );
or   ( new_n39173_, new_n23895_, RIbb2d888_64 );
and  ( new_n39174_, new_n39173_, RIbb2d900_63 );
or   ( new_n39175_, new_n39174_, new_n39172_ );
or   ( new_n39176_, new_n10770_, new_n23733_ );
and  ( new_n39177_, new_n39176_, new_n39175_ );
or   ( new_n39178_, new_n39177_, new_n39171_ );
and  ( new_n39179_, new_n39177_, new_n39171_ );
or   ( new_n39180_, new_n39179_, new_n2120_ );
and  ( new_n39181_, new_n39180_, new_n39178_ );
or   ( new_n39182_, new_n9422_, new_n24543_ );
or   ( new_n39183_, new_n9424_, new_n24418_ );
and  ( new_n39184_, new_n39183_, new_n39182_ );
xor  ( new_n39185_, new_n39184_, new_n8873_ );
or   ( new_n39186_, new_n8874_, new_n24925_ );
or   ( new_n39187_, new_n8876_, new_n24927_ );
and  ( new_n39188_, new_n39187_, new_n39186_ );
xor  ( new_n39189_, new_n39188_, new_n8257_ );
or   ( new_n39190_, new_n39189_, new_n39185_ );
and  ( new_n39191_, new_n39189_, new_n39185_ );
or   ( new_n39192_, new_n8264_, new_n25288_ );
or   ( new_n39193_, new_n8266_, new_n25048_ );
and  ( new_n39194_, new_n39193_, new_n39192_ );
xor  ( new_n39195_, new_n39194_, new_n7725_ );
or   ( new_n39196_, new_n39195_, new_n39191_ );
and  ( new_n39197_, new_n39196_, new_n39190_ );
nor  ( new_n39198_, new_n39197_, new_n39181_ );
and  ( new_n39199_, new_n39197_, new_n39181_ );
or   ( new_n39200_, new_n7732_, new_n25813_ );
or   ( new_n39201_, new_n7734_, new_n25486_ );
and  ( new_n39202_, new_n39201_, new_n39200_ );
xor  ( new_n39203_, new_n39202_, new_n7177_ );
or   ( new_n39204_, new_n7184_, new_n26063_ );
or   ( new_n39205_, new_n7186_, new_n26196_ );
and  ( new_n39206_, new_n39205_, new_n39204_ );
xor  ( new_n39207_, new_n39206_, new_n6638_ );
nor  ( new_n39208_, new_n39207_, new_n39203_ );
and  ( new_n39209_, new_n39207_, new_n39203_ );
or   ( new_n39210_, new_n6645_, new_n26620_ );
or   ( new_n39211_, new_n6647_, new_n26372_ );
and  ( new_n39212_, new_n39211_, new_n39210_ );
xor  ( new_n39213_, new_n39212_, new_n6166_ );
nor  ( new_n39214_, new_n39213_, new_n39209_ );
nor  ( new_n39215_, new_n39214_, new_n39208_ );
nor  ( new_n39216_, new_n39215_, new_n39199_ );
nor  ( new_n39217_, new_n39216_, new_n39198_ );
and  ( new_n39218_, new_n39217_, new_n39167_ );
nor  ( new_n39219_, new_n39217_, new_n39167_ );
xnor ( new_n39220_, new_n39006_, new_n39002_ );
xor  ( new_n39221_, new_n39220_, new_n39012_ );
xnor ( new_n39222_, new_n38990_, new_n38986_ );
xor  ( new_n39223_, new_n39222_, new_n38996_ );
nor  ( new_n39224_, new_n39223_, new_n39221_ );
and  ( new_n39225_, new_n39223_, new_n39221_ );
xor  ( new_n39226_, new_n39024_, new_n39020_ );
xor  ( new_n39227_, new_n39226_, new_n39031_ );
nor  ( new_n39228_, new_n39227_, new_n39225_ );
nor  ( new_n39229_, new_n39228_, new_n39224_ );
nor  ( new_n39230_, new_n39229_, new_n39219_ );
nor  ( new_n39231_, new_n39230_, new_n39218_ );
and  ( new_n39232_, new_n39231_, new_n39115_ );
xor  ( new_n39233_, new_n39046_, new_n39044_ );
xor  ( new_n39234_, new_n39233_, new_n39050_ );
xnor ( new_n39235_, new_n38938_, new_n38932_ );
xor  ( new_n39236_, new_n39235_, new_n38944_ );
xnor ( new_n39237_, new_n38920_, new_n38916_ );
xor  ( new_n39238_, new_n39237_, new_n38926_ );
or   ( new_n39239_, new_n39238_, new_n39236_ );
and  ( new_n39240_, new_n39238_, new_n39236_ );
xor  ( new_n39241_, new_n38956_, new_n38952_ );
xnor ( new_n39242_, new_n39241_, new_n38962_ );
or   ( new_n39243_, new_n39242_, new_n39240_ );
and  ( new_n39244_, new_n39243_, new_n39239_ );
nor  ( new_n39245_, new_n39244_, new_n39234_ );
and  ( new_n39246_, new_n39244_, new_n39234_ );
xor  ( new_n39247_, new_n39041_, new_n39039_ );
not  ( new_n39248_, new_n39247_ );
nor  ( new_n39249_, new_n39248_, new_n39246_ );
nor  ( new_n39250_, new_n39249_, new_n39245_ );
nor  ( new_n39251_, new_n39250_, new_n39232_ );
nor  ( new_n39252_, new_n39231_, new_n39115_ );
or   ( new_n39253_, new_n39252_, new_n39251_ );
xor  ( new_n39254_, new_n38782_, new_n38766_ );
xor  ( new_n39255_, new_n39254_, new_n38752_ );
xnor ( new_n39256_, new_n39052_, new_n39042_ );
xor  ( new_n39257_, new_n39256_, new_n39056_ );
or   ( new_n39258_, new_n39257_, new_n39255_ );
and  ( new_n39259_, new_n39257_, new_n39255_ );
xor  ( new_n39260_, new_n39064_, new_n39062_ );
xnor ( new_n39261_, new_n39260_, new_n39068_ );
or   ( new_n39262_, new_n39261_, new_n39259_ );
and  ( new_n39263_, new_n39262_, new_n39258_ );
nand ( new_n39264_, new_n39263_, new_n39253_ );
nor  ( new_n39265_, new_n39263_, new_n39253_ );
xor  ( new_n39266_, new_n39078_, new_n39076_ );
xor  ( new_n39267_, new_n39266_, new_n39082_ );
or   ( new_n39268_, new_n39267_, new_n39265_ );
and  ( new_n39269_, new_n39268_, new_n39264_ );
or   ( new_n39270_, new_n39269_, new_n39105_ );
and  ( new_n39271_, new_n39269_, new_n39105_ );
xor  ( new_n39272_, new_n39072_, new_n38912_ );
xor  ( new_n39273_, new_n39272_, new_n39084_ );
or   ( new_n39274_, new_n39273_, new_n39271_ );
and  ( new_n39275_, new_n39274_, new_n39270_ );
nor  ( new_n39276_, new_n39275_, new_n39103_ );
xnor ( new_n39277_, new_n39094_, new_n38910_ );
xor  ( new_n39278_, new_n39277_, new_n39098_ );
and  ( new_n39279_, new_n39278_, new_n39276_ );
not  ( new_n39280_, new_n39250_ );
xor  ( new_n39281_, new_n39231_, new_n39115_ );
nor  ( new_n39282_, new_n39281_, new_n39280_ );
not  ( new_n39283_, new_n39252_ );
and  ( new_n39284_, new_n39283_, new_n39251_ );
nor  ( new_n39285_, new_n39284_, new_n39282_ );
not  ( new_n39286_, new_n39285_ );
xnor ( new_n39287_, new_n39257_, new_n39255_ );
xor  ( new_n39288_, new_n39287_, new_n39261_ );
or   ( new_n39289_, new_n39288_, new_n39286_ );
xnor ( new_n39290_, new_n39217_, new_n39167_ );
xor  ( new_n39291_, new_n39290_, new_n39229_ );
xnor ( new_n39292_, new_n39109_, new_n39107_ );
xor  ( new_n39293_, new_n39292_, new_n39113_ );
nand ( new_n39294_, new_n39293_, new_n39291_ );
or   ( new_n39295_, new_n39293_, new_n39291_ );
xor  ( new_n39296_, new_n39244_, new_n39234_ );
xor  ( new_n39297_, new_n39296_, new_n39247_ );
nand ( new_n39298_, new_n39297_, new_n39295_ );
and  ( new_n39299_, new_n39298_, new_n39294_ );
xor  ( new_n39300_, new_n38980_, new_n38966_ );
xor  ( new_n39301_, new_n39300_, new_n39035_ );
or   ( new_n39302_, new_n39301_, new_n39299_ );
and  ( new_n39303_, new_n39301_, new_n39299_ );
xor  ( new_n39304_, new_n39197_, new_n39181_ );
xnor ( new_n39305_, new_n39304_, new_n39215_ );
xnor ( new_n39306_, new_n39147_, new_n39131_ );
xor  ( new_n39307_, new_n39306_, new_n39165_ );
nor  ( new_n39308_, new_n39307_, new_n39305_ );
and  ( new_n39309_, new_n2242_, RIbb33378_192 );
or   ( new_n39310_, new_n39309_, new_n2121_ );
nand ( new_n39311_, new_n39309_, new_n2118_ );
and  ( new_n39312_, new_n39311_, new_n39310_ );
xnor ( new_n39313_, new_n39157_, new_n39153_ );
xor  ( new_n39314_, new_n39313_, new_n39163_ );
nor  ( new_n39315_, new_n39314_, new_n39312_ );
nand ( new_n39316_, new_n39314_, new_n39312_ );
xor  ( new_n39317_, new_n39123_, new_n39119_ );
xnor ( new_n39318_, new_n39317_, new_n39129_ );
not  ( new_n39319_, new_n39318_ );
and  ( new_n39320_, new_n39319_, new_n39316_ );
or   ( new_n39321_, new_n39320_, new_n39315_ );
or   ( new_n39322_, new_n10059_, new_n24418_ );
or   ( new_n39323_, new_n10061_, new_n24227_ );
and  ( new_n39324_, new_n39323_, new_n39322_ );
xor  ( new_n39325_, new_n39324_, new_n9421_ );
and  ( new_n39326_, RIbb32400_159, RIbb2d888_64 );
or   ( new_n39327_, new_n24006_, RIbb2d888_64 );
and  ( new_n39328_, new_n39327_, RIbb2d900_63 );
or   ( new_n39329_, new_n39328_, new_n39326_ );
or   ( new_n39330_, new_n10770_, new_n23895_ );
and  ( new_n39331_, new_n39330_, new_n39329_ );
or   ( new_n39332_, new_n39331_, new_n39325_ );
and  ( new_n39333_, new_n39331_, new_n39325_ );
or   ( new_n39334_, new_n9422_, new_n24927_ );
or   ( new_n39335_, new_n9424_, new_n24543_ );
and  ( new_n39336_, new_n39335_, new_n39334_ );
xor  ( new_n39337_, new_n39336_, new_n8873_ );
or   ( new_n39338_, new_n39337_, new_n39333_ );
and  ( new_n39339_, new_n39338_, new_n39332_ );
or   ( new_n39340_, new_n7184_, new_n26372_ );
or   ( new_n39341_, new_n7186_, new_n26063_ );
and  ( new_n39342_, new_n39341_, new_n39340_ );
xor  ( new_n39343_, new_n39342_, new_n6638_ );
or   ( new_n39344_, new_n6645_, new_n26762_ );
or   ( new_n39345_, new_n6647_, new_n26620_ );
and  ( new_n39346_, new_n39345_, new_n39344_ );
xor  ( new_n39347_, new_n39346_, new_n6166_ );
or   ( new_n39348_, new_n39347_, new_n39343_ );
and  ( new_n39349_, new_n39347_, new_n39343_ );
or   ( new_n39350_, new_n6173_, new_n27396_ );
or   ( new_n39351_, new_n6175_, new_n27085_ );
and  ( new_n39352_, new_n39351_, new_n39350_ );
xor  ( new_n39353_, new_n39352_, new_n5597_ );
or   ( new_n39354_, new_n39353_, new_n39349_ );
and  ( new_n39355_, new_n39354_, new_n39348_ );
or   ( new_n39356_, new_n39355_, new_n39339_ );
and  ( new_n39357_, new_n39355_, new_n39339_ );
or   ( new_n39358_, new_n8874_, new_n25048_ );
or   ( new_n39359_, new_n8876_, new_n24925_ );
and  ( new_n39360_, new_n39359_, new_n39358_ );
xor  ( new_n39361_, new_n39360_, new_n8257_ );
or   ( new_n39362_, new_n8264_, new_n25486_ );
or   ( new_n39363_, new_n8266_, new_n25288_ );
and  ( new_n39364_, new_n39363_, new_n39362_ );
xor  ( new_n39365_, new_n39364_, new_n7725_ );
or   ( new_n39366_, new_n39365_, new_n39361_ );
and  ( new_n39367_, new_n39365_, new_n39361_ );
or   ( new_n39368_, new_n7732_, new_n26196_ );
or   ( new_n39369_, new_n7734_, new_n25813_ );
and  ( new_n39370_, new_n39369_, new_n39368_ );
xor  ( new_n39371_, new_n39370_, new_n7177_ );
or   ( new_n39372_, new_n39371_, new_n39367_ );
and  ( new_n39373_, new_n39372_, new_n39366_ );
or   ( new_n39374_, new_n39373_, new_n39357_ );
and  ( new_n39375_, new_n39374_, new_n39356_ );
or   ( new_n39376_, new_n39375_, new_n39321_ );
and  ( new_n39377_, new_n39375_, new_n39321_ );
or   ( new_n39378_, new_n4302_, new_n29474_ );
or   ( new_n39379_, new_n4304_, new_n29261_ );
and  ( new_n39380_, new_n39379_, new_n39378_ );
xor  ( new_n39381_, new_n39380_, new_n3895_ );
or   ( new_n39382_, new_n3896_, new_n30120_ );
or   ( new_n39383_, new_n3898_, new_n29619_ );
and  ( new_n39384_, new_n39383_, new_n39382_ );
xor  ( new_n39385_, new_n39384_, new_n3460_ );
nor  ( new_n39386_, new_n39385_, new_n39381_ );
and  ( new_n39387_, new_n39385_, new_n39381_ );
or   ( new_n39388_, new_n3461_, new_n30800_ );
or   ( new_n39389_, new_n3463_, new_n30227_ );
and  ( new_n39390_, new_n39389_, new_n39388_ );
xor  ( new_n39391_, new_n39390_, new_n3116_ );
nor  ( new_n39392_, new_n39391_, new_n39387_ );
nor  ( new_n39393_, new_n39392_, new_n39386_ );
or   ( new_n39394_, new_n3117_, new_n31333_ );
or   ( new_n39395_, new_n3119_, new_n30798_ );
and  ( new_n39396_, new_n39395_, new_n39394_ );
xor  ( new_n39397_, new_n39396_, new_n2800_ );
or   ( new_n39398_, new_n2807_, new_n31952_ );
or   ( new_n39399_, new_n2809_, new_n31654_ );
and  ( new_n39400_, new_n39399_, new_n39398_ );
xor  ( new_n39401_, new_n39400_, new_n2424_ );
and  ( new_n39402_, new_n39401_, new_n39397_ );
or   ( new_n39403_, new_n5604_, new_n27763_ );
or   ( new_n39404_, new_n5606_, new_n27602_ );
and  ( new_n39405_, new_n39404_, new_n39403_ );
xor  ( new_n39406_, new_n39405_, new_n5206_ );
or   ( new_n39407_, new_n5207_, new_n28314_ );
or   ( new_n39408_, new_n5209_, new_n28108_ );
and  ( new_n39409_, new_n39408_, new_n39407_ );
xor  ( new_n39410_, new_n39409_, new_n4708_ );
nor  ( new_n39411_, new_n39410_, new_n39406_ );
and  ( new_n39412_, new_n39410_, new_n39406_ );
or   ( new_n39413_, new_n4709_, new_n29263_ );
or   ( new_n39414_, new_n4711_, new_n28531_ );
and  ( new_n39415_, new_n39414_, new_n39413_ );
xor  ( new_n39416_, new_n39415_, new_n4295_ );
nor  ( new_n39417_, new_n39416_, new_n39412_ );
nor  ( new_n39418_, new_n39417_, new_n39411_ );
and  ( new_n39419_, new_n39418_, new_n39402_ );
nor  ( new_n39420_, new_n39419_, new_n39393_ );
nor  ( new_n39421_, new_n39418_, new_n39402_ );
nor  ( new_n39422_, new_n39421_, new_n39420_ );
or   ( new_n39423_, new_n39422_, new_n39377_ );
and  ( new_n39424_, new_n39423_, new_n39376_ );
and  ( new_n39425_, new_n39424_, new_n39308_ );
nor  ( new_n39426_, new_n39424_, new_n39308_ );
xor  ( new_n39427_, new_n39223_, new_n39221_ );
xor  ( new_n39428_, new_n39427_, new_n39227_ );
xnor ( new_n39429_, new_n39189_, new_n39185_ );
xor  ( new_n39430_, new_n39429_, new_n39195_ );
xnor ( new_n39431_, new_n39139_, new_n39135_ );
xor  ( new_n39432_, new_n39431_, new_n39145_ );
or   ( new_n39433_, new_n39432_, new_n39430_ );
and  ( new_n39434_, new_n39432_, new_n39430_ );
xor  ( new_n39435_, new_n39207_, new_n39203_ );
xnor ( new_n39436_, new_n39435_, new_n39213_ );
or   ( new_n39437_, new_n39436_, new_n39434_ );
and  ( new_n39438_, new_n39437_, new_n39433_ );
nor  ( new_n39439_, new_n39438_, new_n39428_ );
and  ( new_n39440_, new_n39438_, new_n39428_ );
xor  ( new_n39441_, new_n39238_, new_n39236_ );
xnor ( new_n39442_, new_n39441_, new_n39242_ );
not  ( new_n39443_, new_n39442_ );
nor  ( new_n39444_, new_n39443_, new_n39440_ );
nor  ( new_n39445_, new_n39444_, new_n39439_ );
nor  ( new_n39446_, new_n39445_, new_n39426_ );
nor  ( new_n39447_, new_n39446_, new_n39425_ );
or   ( new_n39448_, new_n39447_, new_n39303_ );
and  ( new_n39449_, new_n39448_, new_n39302_ );
nor  ( new_n39450_, new_n39449_, new_n39289_ );
and  ( new_n39451_, new_n39449_, new_n39289_ );
xor  ( new_n39452_, new_n39058_, new_n39037_ );
xor  ( new_n39453_, new_n39452_, new_n39070_ );
nor  ( new_n39454_, new_n39453_, new_n39451_ );
or   ( new_n39455_, new_n39454_, new_n39450_ );
xnor ( new_n39456_, new_n39269_, new_n39105_ );
xor  ( new_n39457_, new_n39456_, new_n39273_ );
and  ( new_n39458_, new_n39457_, new_n39455_ );
xor  ( new_n39459_, new_n39275_, new_n39103_ );
and  ( new_n39460_, new_n39459_, new_n39458_ );
xor  ( new_n39461_, new_n39449_, new_n39289_ );
xor  ( new_n39462_, new_n39461_, new_n39453_ );
xor  ( new_n39463_, new_n39263_, new_n39253_ );
xor  ( new_n39464_, new_n39463_, new_n39267_ );
nor  ( new_n39465_, new_n39464_, new_n39462_ );
xor  ( new_n39466_, new_n39457_, new_n39455_ );
and  ( new_n39467_, new_n39466_, new_n39465_ );
xor  ( new_n39468_, new_n39464_, new_n39462_ );
xor  ( new_n39469_, new_n39177_, new_n39171_ );
xor  ( new_n39470_, new_n39469_, new_n2121_ );
xnor ( new_n39471_, new_n39347_, new_n39343_ );
xor  ( new_n39472_, new_n39471_, new_n39353_ );
xnor ( new_n39473_, new_n39331_, new_n39325_ );
xor  ( new_n39474_, new_n39473_, new_n39337_ );
or   ( new_n39475_, new_n39474_, new_n39472_ );
and  ( new_n39476_, new_n39474_, new_n39472_ );
xor  ( new_n39477_, new_n39365_, new_n39361_ );
xnor ( new_n39478_, new_n39477_, new_n39371_ );
or   ( new_n39479_, new_n39478_, new_n39476_ );
and  ( new_n39480_, new_n39479_, new_n39475_ );
nor  ( new_n39481_, new_n39480_, new_n39470_ );
and  ( new_n39482_, new_n39480_, new_n39470_ );
xor  ( new_n39483_, new_n39432_, new_n39430_ );
xnor ( new_n39484_, new_n39483_, new_n39436_ );
not  ( new_n39485_, new_n39484_ );
nor  ( new_n39486_, new_n39485_, new_n39482_ );
nor  ( new_n39487_, new_n39486_, new_n39481_ );
or   ( new_n39488_, new_n7732_, new_n26063_ );
or   ( new_n39489_, new_n7734_, new_n26196_ );
and  ( new_n39490_, new_n39489_, new_n39488_ );
xor  ( new_n39491_, new_n39490_, new_n7177_ );
or   ( new_n39492_, new_n7184_, new_n26620_ );
or   ( new_n39493_, new_n7186_, new_n26372_ );
and  ( new_n39494_, new_n39493_, new_n39492_ );
xor  ( new_n39495_, new_n39494_, new_n6638_ );
nor  ( new_n39496_, new_n39495_, new_n39491_ );
nand ( new_n39497_, new_n39495_, new_n39491_ );
or   ( new_n39498_, new_n6645_, new_n27085_ );
or   ( new_n39499_, new_n6647_, new_n26762_ );
and  ( new_n39500_, new_n39499_, new_n39498_ );
xor  ( new_n39501_, new_n39500_, new_n6165_ );
and  ( new_n39502_, new_n39501_, new_n39497_ );
or   ( new_n39503_, new_n39502_, new_n39496_ );
or   ( new_n39504_, new_n10059_, new_n24543_ );
or   ( new_n39505_, new_n10061_, new_n24418_ );
and  ( new_n39506_, new_n39505_, new_n39504_ );
xor  ( new_n39507_, new_n39506_, new_n9421_ );
and  ( new_n39508_, RIbb32478_160, RIbb2d888_64 );
or   ( new_n39509_, new_n24227_, RIbb2d888_64 );
and  ( new_n39510_, new_n39509_, RIbb2d900_63 );
or   ( new_n39511_, new_n39510_, new_n39508_ );
or   ( new_n39512_, new_n10770_, new_n24006_ );
and  ( new_n39513_, new_n39512_, new_n39511_ );
nor  ( new_n39514_, new_n39513_, new_n39507_ );
nand ( new_n39515_, new_n39513_, new_n39507_ );
and  ( new_n39516_, new_n39515_, new_n2424_ );
or   ( new_n39517_, new_n39516_, new_n39514_ );
or   ( new_n39518_, new_n9422_, new_n24925_ );
or   ( new_n39519_, new_n9424_, new_n24927_ );
and  ( new_n39520_, new_n39519_, new_n39518_ );
xor  ( new_n39521_, new_n39520_, new_n8873_ );
or   ( new_n39522_, new_n8874_, new_n25288_ );
or   ( new_n39523_, new_n8876_, new_n25048_ );
and  ( new_n39524_, new_n39523_, new_n39522_ );
xor  ( new_n39525_, new_n39524_, new_n8257_ );
nor  ( new_n39526_, new_n39525_, new_n39521_ );
and  ( new_n39527_, new_n39525_, new_n39521_ );
or   ( new_n39528_, new_n8264_, new_n25813_ );
or   ( new_n39529_, new_n8266_, new_n25486_ );
and  ( new_n39530_, new_n39529_, new_n39528_ );
xor  ( new_n39531_, new_n39530_, new_n7725_ );
nor  ( new_n39532_, new_n39531_, new_n39527_ );
nor  ( new_n39533_, new_n39532_, new_n39526_ );
not  ( new_n39534_, new_n39533_ );
or   ( new_n39535_, new_n39534_, new_n39517_ );
and  ( new_n39536_, new_n39535_, new_n39503_ );
and  ( new_n39537_, new_n39534_, new_n39517_ );
or   ( new_n39538_, new_n39537_, new_n39536_ );
or   ( new_n39539_, new_n6173_, new_n27602_ );
or   ( new_n39540_, new_n6175_, new_n27396_ );
and  ( new_n39541_, new_n39540_, new_n39539_ );
xor  ( new_n39542_, new_n39541_, new_n5597_ );
or   ( new_n39543_, new_n5604_, new_n28108_ );
or   ( new_n39544_, new_n5606_, new_n27763_ );
and  ( new_n39545_, new_n39544_, new_n39543_ );
xor  ( new_n39546_, new_n39545_, new_n5206_ );
nor  ( new_n39547_, new_n39546_, new_n39542_ );
nand ( new_n39548_, new_n39546_, new_n39542_ );
or   ( new_n39549_, new_n5207_, new_n28531_ );
or   ( new_n39550_, new_n5209_, new_n28314_ );
and  ( new_n39551_, new_n39550_, new_n39549_ );
xor  ( new_n39552_, new_n39551_, new_n4708_ );
not  ( new_n39553_, new_n39552_ );
and  ( new_n39554_, new_n39553_, new_n39548_ );
or   ( new_n39555_, new_n39554_, new_n39547_ );
or   ( new_n39556_, new_n4709_, new_n29261_ );
or   ( new_n39557_, new_n4711_, new_n29263_ );
and  ( new_n39558_, new_n39557_, new_n39556_ );
xor  ( new_n39559_, new_n39558_, new_n4295_ );
or   ( new_n39560_, new_n4302_, new_n29619_ );
or   ( new_n39561_, new_n4304_, new_n29474_ );
and  ( new_n39562_, new_n39561_, new_n39560_ );
xor  ( new_n39563_, new_n39562_, new_n3895_ );
nor  ( new_n39564_, new_n39563_, new_n39559_ );
and  ( new_n39565_, new_n39563_, new_n39559_ );
or   ( new_n39566_, new_n3896_, new_n30227_ );
or   ( new_n39567_, new_n3898_, new_n30120_ );
and  ( new_n39568_, new_n39567_, new_n39566_ );
xor  ( new_n39569_, new_n39568_, new_n3460_ );
nor  ( new_n39570_, new_n39569_, new_n39565_ );
nor  ( new_n39571_, new_n39570_, new_n39564_ );
not  ( new_n39572_, new_n39571_ );
or   ( new_n39573_, new_n39572_, new_n39555_ );
and  ( new_n39574_, new_n39572_, new_n39555_ );
or   ( new_n39575_, new_n3461_, new_n30798_ );
or   ( new_n39576_, new_n3463_, new_n30800_ );
and  ( new_n39577_, new_n39576_, new_n39575_ );
xor  ( new_n39578_, new_n39577_, new_n3116_ );
or   ( new_n39579_, new_n3117_, new_n31654_ );
or   ( new_n39580_, new_n3119_, new_n31333_ );
and  ( new_n39581_, new_n39580_, new_n39579_ );
xor  ( new_n39582_, new_n39581_, new_n2800_ );
nand ( new_n39583_, new_n39582_, new_n39578_ );
nor  ( new_n39584_, new_n39582_, new_n39578_ );
and  ( new_n39585_, new_n2613_, RIbb33378_192 );
nor  ( new_n39586_, new_n39585_, new_n2424_ );
and  ( new_n39587_, new_n39585_, new_n2421_ );
nor  ( new_n39588_, new_n39587_, new_n39586_ );
or   ( new_n39589_, new_n39588_, new_n39584_ );
and  ( new_n39590_, new_n39589_, new_n39583_ );
or   ( new_n39591_, new_n39590_, new_n39574_ );
and  ( new_n39592_, new_n39591_, new_n39573_ );
nor  ( new_n39593_, new_n39592_, new_n39538_ );
and  ( new_n39594_, new_n39592_, new_n39538_ );
xnor ( new_n39595_, new_n39385_, new_n39381_ );
xor  ( new_n39596_, new_n39595_, new_n39391_ );
xnor ( new_n39597_, new_n39410_, new_n39406_ );
xor  ( new_n39598_, new_n39597_, new_n39416_ );
nor  ( new_n39599_, new_n39598_, new_n39596_ );
and  ( new_n39600_, new_n39598_, new_n39596_ );
xor  ( new_n39601_, new_n39401_, new_n39397_ );
not  ( new_n39602_, new_n39601_ );
nor  ( new_n39603_, new_n39602_, new_n39600_ );
nor  ( new_n39604_, new_n39603_, new_n39599_ );
nor  ( new_n39605_, new_n39604_, new_n39594_ );
nor  ( new_n39606_, new_n39605_, new_n39593_ );
and  ( new_n39607_, new_n39606_, new_n39487_ );
xor  ( new_n39608_, new_n39355_, new_n39339_ );
xor  ( new_n39609_, new_n39608_, new_n39373_ );
xor  ( new_n39610_, new_n39418_, new_n39402_ );
xor  ( new_n39611_, new_n39610_, new_n39393_ );
and  ( new_n39612_, new_n39611_, new_n39609_ );
nor  ( new_n39613_, new_n39611_, new_n39609_ );
not  ( new_n39614_, new_n39613_ );
xor  ( new_n39615_, new_n39314_, new_n39312_ );
xor  ( new_n39616_, new_n39615_, new_n39319_ );
and  ( new_n39617_, new_n39616_, new_n39614_ );
nor  ( new_n39618_, new_n39617_, new_n39612_ );
nor  ( new_n39619_, new_n39618_, new_n39607_ );
nor  ( new_n39620_, new_n39606_, new_n39487_ );
or   ( new_n39621_, new_n39620_, new_n39619_ );
xor  ( new_n39622_, new_n39293_, new_n39291_ );
xor  ( new_n39623_, new_n39622_, new_n39297_ );
or   ( new_n39624_, new_n39623_, new_n39621_ );
nand ( new_n39625_, new_n39623_, new_n39621_ );
xor  ( new_n39626_, new_n39438_, new_n39428_ );
xor  ( new_n39627_, new_n39626_, new_n39443_ );
xnor ( new_n39628_, new_n39375_, new_n39321_ );
xor  ( new_n39629_, new_n39628_, new_n39422_ );
nor  ( new_n39630_, new_n39629_, new_n39627_ );
and  ( new_n39631_, new_n39629_, new_n39627_ );
xor  ( new_n39632_, new_n39307_, new_n39305_ );
not  ( new_n39633_, new_n39632_ );
nor  ( new_n39634_, new_n39633_, new_n39631_ );
nor  ( new_n39635_, new_n39634_, new_n39630_ );
nand ( new_n39636_, new_n39635_, new_n39625_ );
and  ( new_n39637_, new_n39636_, new_n39624_ );
xnor ( new_n39638_, new_n39301_, new_n39299_ );
xor  ( new_n39639_, new_n39638_, new_n39447_ );
or   ( new_n39640_, new_n39639_, new_n39637_ );
and  ( new_n39641_, new_n39639_, new_n39637_ );
xor  ( new_n39642_, new_n39288_, new_n39286_ );
or   ( new_n39643_, new_n39642_, new_n39641_ );
and  ( new_n39644_, new_n39643_, new_n39640_ );
and  ( new_n39645_, new_n39644_, new_n39468_ );
xnor ( new_n39646_, new_n39639_, new_n39637_ );
xor  ( new_n39647_, new_n39646_, new_n39642_ );
xnor ( new_n39648_, new_n39606_, new_n39487_ );
and  ( new_n39649_, new_n39648_, new_n39618_ );
not  ( new_n39650_, new_n39619_ );
nor  ( new_n39651_, new_n39620_, new_n39650_ );
or   ( new_n39652_, new_n39651_, new_n39649_ );
xor  ( new_n39653_, new_n39571_, new_n39555_ );
xor  ( new_n39654_, new_n39653_, new_n39590_ );
xnor ( new_n39655_, new_n39474_, new_n39472_ );
xor  ( new_n39656_, new_n39655_, new_n39478_ );
or   ( new_n39657_, new_n39656_, new_n39654_ );
and  ( new_n39658_, new_n39656_, new_n39654_ );
xor  ( new_n39659_, new_n39598_, new_n39596_ );
xor  ( new_n39660_, new_n39659_, new_n39601_ );
or   ( new_n39661_, new_n39660_, new_n39658_ );
and  ( new_n39662_, new_n39661_, new_n39657_ );
xor  ( new_n39663_, new_n39611_, new_n39609_ );
xor  ( new_n39664_, new_n39663_, new_n39616_ );
nand ( new_n39665_, new_n39664_, new_n39662_ );
nor  ( new_n39666_, new_n39664_, new_n39662_ );
or   ( new_n39667_, new_n10059_, new_n24927_ );
or   ( new_n39668_, new_n10061_, new_n24543_ );
and  ( new_n39669_, new_n39668_, new_n39667_ );
xor  ( new_n39670_, new_n39669_, new_n9421_ );
and  ( new_n39671_, RIbb324f0_161, RIbb2d888_64 );
or   ( new_n39672_, new_n24418_, RIbb2d888_64 );
and  ( new_n39673_, new_n39672_, RIbb2d900_63 );
or   ( new_n39674_, new_n39673_, new_n39671_ );
or   ( new_n39675_, new_n10770_, new_n24227_ );
and  ( new_n39676_, new_n39675_, new_n39674_ );
or   ( new_n39677_, new_n39676_, new_n39670_ );
and  ( new_n39678_, new_n39676_, new_n39670_ );
or   ( new_n39679_, new_n9422_, new_n25048_ );
or   ( new_n39680_, new_n9424_, new_n24925_ );
and  ( new_n39681_, new_n39680_, new_n39679_ );
xor  ( new_n39682_, new_n39681_, new_n8873_ );
or   ( new_n39683_, new_n39682_, new_n39678_ );
and  ( new_n39684_, new_n39683_, new_n39677_ );
or   ( new_n39685_, new_n8874_, new_n25486_ );
or   ( new_n39686_, new_n8876_, new_n25288_ );
and  ( new_n39687_, new_n39686_, new_n39685_ );
xor  ( new_n39688_, new_n39687_, new_n8257_ );
or   ( new_n39689_, new_n8264_, new_n26196_ );
or   ( new_n39690_, new_n8266_, new_n25813_ );
and  ( new_n39691_, new_n39690_, new_n39689_ );
xor  ( new_n39692_, new_n39691_, new_n7725_ );
or   ( new_n39693_, new_n39692_, new_n39688_ );
and  ( new_n39694_, new_n39692_, new_n39688_ );
or   ( new_n39695_, new_n7732_, new_n26372_ );
or   ( new_n39696_, new_n7734_, new_n26063_ );
and  ( new_n39697_, new_n39696_, new_n39695_ );
xor  ( new_n39698_, new_n39697_, new_n7177_ );
or   ( new_n39699_, new_n39698_, new_n39694_ );
and  ( new_n39700_, new_n39699_, new_n39693_ );
or   ( new_n39701_, new_n39700_, new_n39684_ );
and  ( new_n39702_, new_n39700_, new_n39684_ );
or   ( new_n39703_, new_n7184_, new_n26762_ );
or   ( new_n39704_, new_n7186_, new_n26620_ );
and  ( new_n39705_, new_n39704_, new_n39703_ );
xor  ( new_n39706_, new_n39705_, new_n6638_ );
or   ( new_n39707_, new_n6645_, new_n27396_ );
or   ( new_n39708_, new_n6647_, new_n27085_ );
and  ( new_n39709_, new_n39708_, new_n39707_ );
xor  ( new_n39710_, new_n39709_, new_n6166_ );
nor  ( new_n39711_, new_n39710_, new_n39706_ );
and  ( new_n39712_, new_n39710_, new_n39706_ );
or   ( new_n39713_, new_n6173_, new_n27763_ );
or   ( new_n39714_, new_n6175_, new_n27602_ );
and  ( new_n39715_, new_n39714_, new_n39713_ );
xor  ( new_n39716_, new_n39715_, new_n5597_ );
nor  ( new_n39717_, new_n39716_, new_n39712_ );
nor  ( new_n39718_, new_n39717_, new_n39711_ );
or   ( new_n39719_, new_n39718_, new_n39702_ );
and  ( new_n39720_, new_n39719_, new_n39701_ );
xnor ( new_n39721_, new_n39582_, new_n39578_ );
xor  ( new_n39722_, new_n39721_, new_n39588_ );
or   ( new_n39723_, new_n5604_, new_n28314_ );
or   ( new_n39724_, new_n5606_, new_n28108_ );
and  ( new_n39725_, new_n39724_, new_n39723_ );
xor  ( new_n39726_, new_n39725_, new_n5206_ );
or   ( new_n39727_, new_n5207_, new_n29263_ );
or   ( new_n39728_, new_n5209_, new_n28531_ );
and  ( new_n39729_, new_n39728_, new_n39727_ );
xor  ( new_n39730_, new_n39729_, new_n4708_ );
or   ( new_n39731_, new_n39730_, new_n39726_ );
and  ( new_n39732_, new_n39730_, new_n39726_ );
or   ( new_n39733_, new_n4709_, new_n29474_ );
or   ( new_n39734_, new_n4711_, new_n29261_ );
and  ( new_n39735_, new_n39734_, new_n39733_ );
xor  ( new_n39736_, new_n39735_, new_n4295_ );
or   ( new_n39737_, new_n39736_, new_n39732_ );
and  ( new_n39738_, new_n39737_, new_n39731_ );
or   ( new_n39739_, new_n39738_, new_n39722_ );
and  ( new_n39740_, new_n39738_, new_n39722_ );
or   ( new_n39741_, new_n4302_, new_n30120_ );
or   ( new_n39742_, new_n4304_, new_n29619_ );
and  ( new_n39743_, new_n39742_, new_n39741_ );
xor  ( new_n39744_, new_n39743_, new_n3895_ );
or   ( new_n39745_, new_n3896_, new_n30800_ );
or   ( new_n39746_, new_n3898_, new_n30227_ );
and  ( new_n39747_, new_n39746_, new_n39745_ );
xor  ( new_n39748_, new_n39747_, new_n3460_ );
nor  ( new_n39749_, new_n39748_, new_n39744_ );
and  ( new_n39750_, new_n39748_, new_n39744_ );
or   ( new_n39751_, new_n3461_, new_n31333_ );
or   ( new_n39752_, new_n3463_, new_n30798_ );
and  ( new_n39753_, new_n39752_, new_n39751_ );
xor  ( new_n39754_, new_n39753_, new_n3116_ );
nor  ( new_n39755_, new_n39754_, new_n39750_ );
nor  ( new_n39756_, new_n39755_, new_n39749_ );
or   ( new_n39757_, new_n39756_, new_n39740_ );
and  ( new_n39758_, new_n39757_, new_n39739_ );
and  ( new_n39759_, new_n39758_, new_n39720_ );
nor  ( new_n39760_, new_n39758_, new_n39720_ );
xnor ( new_n39761_, new_n39563_, new_n39559_ );
xor  ( new_n39762_, new_n39761_, new_n39569_ );
xor  ( new_n39763_, new_n39495_, new_n39491_ );
xor  ( new_n39764_, new_n39763_, new_n39501_ );
nor  ( new_n39765_, new_n39764_, new_n39762_ );
and  ( new_n39766_, new_n39764_, new_n39762_ );
xor  ( new_n39767_, new_n39546_, new_n39542_ );
xor  ( new_n39768_, new_n39767_, new_n39553_ );
nor  ( new_n39769_, new_n39768_, new_n39766_ );
nor  ( new_n39770_, new_n39769_, new_n39765_ );
nor  ( new_n39771_, new_n39770_, new_n39760_ );
nor  ( new_n39772_, new_n39771_, new_n39759_ );
or   ( new_n39773_, new_n39772_, new_n39666_ );
and  ( new_n39774_, new_n39773_, new_n39665_ );
nor  ( new_n39775_, new_n39774_, new_n39652_ );
and  ( new_n39776_, new_n39774_, new_n39652_ );
xor  ( new_n39777_, new_n39629_, new_n39627_ );
xor  ( new_n39778_, new_n39777_, new_n39633_ );
nor  ( new_n39779_, new_n39778_, new_n39776_ );
or   ( new_n39780_, new_n39779_, new_n39775_ );
xnor ( new_n39781_, new_n39424_, new_n39308_ );
xor  ( new_n39782_, new_n39781_, new_n39445_ );
nand ( new_n39783_, new_n39782_, new_n39780_ );
nor  ( new_n39784_, new_n39782_, new_n39780_ );
xor  ( new_n39785_, new_n39623_, new_n39621_ );
xor  ( new_n39786_, new_n39785_, new_n39635_ );
or   ( new_n39787_, new_n39786_, new_n39784_ );
and  ( new_n39788_, new_n39787_, new_n39783_ );
nor  ( new_n39789_, new_n39788_, new_n39647_ );
xor  ( new_n39790_, new_n39782_, new_n39780_ );
xor  ( new_n39791_, new_n39790_, new_n39786_ );
xor  ( new_n39792_, new_n39592_, new_n39538_ );
xor  ( new_n39793_, new_n39792_, new_n39604_ );
xnor ( new_n39794_, new_n39664_, new_n39662_ );
xnor ( new_n39795_, new_n39794_, new_n39772_ );
or   ( new_n39796_, new_n39795_, new_n39793_ );
xor  ( new_n39797_, new_n39480_, new_n39470_ );
xor  ( new_n39798_, new_n39797_, new_n39485_ );
xor  ( new_n39799_, new_n39533_, new_n39517_ );
xor  ( new_n39800_, new_n39799_, new_n39503_ );
xnor ( new_n39801_, new_n39758_, new_n39720_ );
xor  ( new_n39802_, new_n39801_, new_n39770_ );
nand ( new_n39803_, new_n39802_, new_n39800_ );
nor  ( new_n39804_, new_n39802_, new_n39800_ );
xor  ( new_n39805_, new_n39656_, new_n39654_ );
xnor ( new_n39806_, new_n39805_, new_n39660_ );
or   ( new_n39807_, new_n39806_, new_n39804_ );
and  ( new_n39808_, new_n39807_, new_n39803_ );
or   ( new_n39809_, new_n39808_, new_n39798_ );
and  ( new_n39810_, new_n39808_, new_n39798_ );
xor  ( new_n39811_, new_n39700_, new_n39684_ );
xnor ( new_n39812_, new_n39811_, new_n39718_ );
xnor ( new_n39813_, new_n39738_, new_n39722_ );
xor  ( new_n39814_, new_n39813_, new_n39756_ );
or   ( new_n39815_, new_n39814_, new_n39812_ );
or   ( new_n39816_, new_n3117_, new_n31952_ );
or   ( new_n39817_, new_n3119_, new_n31654_ );
and  ( new_n39818_, new_n39817_, new_n39816_ );
xor  ( new_n39819_, new_n39818_, new_n2800_ );
or   ( new_n39820_, new_n4709_, new_n29619_ );
or   ( new_n39821_, new_n4711_, new_n29474_ );
and  ( new_n39822_, new_n39821_, new_n39820_ );
xor  ( new_n39823_, new_n39822_, new_n4295_ );
or   ( new_n39824_, new_n4302_, new_n30227_ );
or   ( new_n39825_, new_n4304_, new_n30120_ );
and  ( new_n39826_, new_n39825_, new_n39824_ );
xor  ( new_n39827_, new_n39826_, new_n3895_ );
or   ( new_n39828_, new_n39827_, new_n39823_ );
and  ( new_n39829_, new_n39827_, new_n39823_ );
or   ( new_n39830_, new_n3896_, new_n30798_ );
or   ( new_n39831_, new_n3898_, new_n30800_ );
and  ( new_n39832_, new_n39831_, new_n39830_ );
xor  ( new_n39833_, new_n39832_, new_n3460_ );
or   ( new_n39834_, new_n39833_, new_n39829_ );
and  ( new_n39835_, new_n39834_, new_n39828_ );
or   ( new_n39836_, new_n39835_, new_n39819_ );
and  ( new_n39837_, new_n39835_, new_n39819_ );
or   ( new_n39838_, new_n6173_, new_n28108_ );
or   ( new_n39839_, new_n6175_, new_n27763_ );
and  ( new_n39840_, new_n39839_, new_n39838_ );
xor  ( new_n39841_, new_n39840_, new_n5597_ );
or   ( new_n39842_, new_n5604_, new_n28531_ );
or   ( new_n39843_, new_n5606_, new_n28314_ );
and  ( new_n39844_, new_n39843_, new_n39842_ );
xor  ( new_n39845_, new_n39844_, new_n5206_ );
nor  ( new_n39846_, new_n39845_, new_n39841_ );
and  ( new_n39847_, new_n39845_, new_n39841_ );
or   ( new_n39848_, new_n5207_, new_n29261_ );
or   ( new_n39849_, new_n5209_, new_n29263_ );
and  ( new_n39850_, new_n39849_, new_n39848_ );
xor  ( new_n39851_, new_n39850_, new_n4708_ );
nor  ( new_n39852_, new_n39851_, new_n39847_ );
nor  ( new_n39853_, new_n39852_, new_n39846_ );
or   ( new_n39854_, new_n39853_, new_n39837_ );
and  ( new_n39855_, new_n39854_, new_n39836_ );
or   ( new_n39856_, new_n9422_, new_n25288_ );
or   ( new_n39857_, new_n9424_, new_n25048_ );
and  ( new_n39858_, new_n39857_, new_n39856_ );
xor  ( new_n39859_, new_n39858_, new_n8873_ );
or   ( new_n39860_, new_n8874_, new_n25813_ );
or   ( new_n39861_, new_n8876_, new_n25486_ );
and  ( new_n39862_, new_n39861_, new_n39860_ );
xor  ( new_n39863_, new_n39862_, new_n8257_ );
nor  ( new_n39864_, new_n39863_, new_n39859_ );
and  ( new_n39865_, new_n39863_, new_n39859_ );
or   ( new_n39866_, new_n8264_, new_n26063_ );
or   ( new_n39867_, new_n8266_, new_n26196_ );
and  ( new_n39868_, new_n39867_, new_n39866_ );
xor  ( new_n39869_, new_n39868_, new_n7725_ );
nor  ( new_n39870_, new_n39869_, new_n39865_ );
nor  ( new_n39871_, new_n39870_, new_n39864_ );
or   ( new_n39872_, new_n10059_, new_n24925_ );
or   ( new_n39873_, new_n10061_, new_n24927_ );
and  ( new_n39874_, new_n39873_, new_n39872_ );
xor  ( new_n39875_, new_n39874_, new_n9421_ );
and  ( new_n39876_, RIbb32568_162, RIbb2d888_64 );
or   ( new_n39877_, new_n24543_, RIbb2d888_64 );
and  ( new_n39878_, new_n39877_, RIbb2d900_63 );
or   ( new_n39879_, new_n39878_, new_n39876_ );
or   ( new_n39880_, new_n10770_, new_n24418_ );
and  ( new_n39881_, new_n39880_, new_n39879_ );
nor  ( new_n39882_, new_n39881_, new_n39875_ );
and  ( new_n39883_, new_n39881_, new_n39875_ );
nor  ( new_n39884_, new_n39883_, new_n2799_ );
nor  ( new_n39885_, new_n39884_, new_n39882_ );
or   ( new_n39886_, new_n7732_, new_n26620_ );
or   ( new_n39887_, new_n7734_, new_n26372_ );
and  ( new_n39888_, new_n39887_, new_n39886_ );
xor  ( new_n39889_, new_n39888_, new_n7177_ );
or   ( new_n39890_, new_n7184_, new_n27085_ );
or   ( new_n39891_, new_n7186_, new_n26762_ );
and  ( new_n39892_, new_n39891_, new_n39890_ );
xor  ( new_n39893_, new_n39892_, new_n6638_ );
or   ( new_n39894_, new_n39893_, new_n39889_ );
and  ( new_n39895_, new_n39893_, new_n39889_ );
or   ( new_n39896_, new_n6645_, new_n27602_ );
or   ( new_n39897_, new_n6647_, new_n27396_ );
and  ( new_n39898_, new_n39897_, new_n39896_ );
xor  ( new_n39899_, new_n39898_, new_n6166_ );
or   ( new_n39900_, new_n39899_, new_n39895_ );
and  ( new_n39901_, new_n39900_, new_n39894_ );
and  ( new_n39902_, new_n39901_, new_n39885_ );
or   ( new_n39903_, new_n39902_, new_n39871_ );
or   ( new_n39904_, new_n39901_, new_n39885_ );
and  ( new_n39905_, new_n39904_, new_n39903_ );
nand ( new_n39906_, new_n39905_, new_n39855_ );
nor  ( new_n39907_, new_n39905_, new_n39855_ );
xnor ( new_n39908_, new_n39730_, new_n39726_ );
xor  ( new_n39909_, new_n39908_, new_n39736_ );
xnor ( new_n39910_, new_n39748_, new_n39744_ );
xor  ( new_n39911_, new_n39910_, new_n39754_ );
nor  ( new_n39912_, new_n39911_, new_n39909_ );
and  ( new_n39913_, new_n39911_, new_n39909_ );
xor  ( new_n39914_, new_n39710_, new_n39706_ );
xnor ( new_n39915_, new_n39914_, new_n39716_ );
nor  ( new_n39916_, new_n39915_, new_n39913_ );
nor  ( new_n39917_, new_n39916_, new_n39912_ );
or   ( new_n39918_, new_n39917_, new_n39907_ );
and  ( new_n39919_, new_n39918_, new_n39906_ );
nor  ( new_n39920_, new_n39919_, new_n39815_ );
and  ( new_n39921_, new_n39919_, new_n39815_ );
xor  ( new_n39922_, new_n39513_, new_n39507_ );
xor  ( new_n39923_, new_n39922_, new_n2424_ );
xnor ( new_n39924_, new_n39525_, new_n39521_ );
xor  ( new_n39925_, new_n39924_, new_n39531_ );
nor  ( new_n39926_, new_n39925_, new_n39923_ );
and  ( new_n39927_, new_n39925_, new_n39923_ );
not  ( new_n39928_, new_n39927_ );
xor  ( new_n39929_, new_n39764_, new_n39762_ );
xnor ( new_n39930_, new_n39929_, new_n39768_ );
and  ( new_n39931_, new_n39930_, new_n39928_ );
nor  ( new_n39932_, new_n39931_, new_n39926_ );
nor  ( new_n39933_, new_n39932_, new_n39921_ );
nor  ( new_n39934_, new_n39933_, new_n39920_ );
or   ( new_n39935_, new_n39934_, new_n39810_ );
and  ( new_n39936_, new_n39935_, new_n39809_ );
or   ( new_n39937_, new_n39936_, new_n39796_ );
and  ( new_n39938_, new_n39936_, new_n39796_ );
xor  ( new_n39939_, new_n39774_, new_n39652_ );
xor  ( new_n39940_, new_n39939_, new_n39778_ );
or   ( new_n39941_, new_n39940_, new_n39938_ );
and  ( new_n39942_, new_n39941_, new_n39937_ );
nor  ( new_n39943_, new_n39942_, new_n39791_ );
xnor ( new_n39944_, new_n39802_, new_n39800_ );
xor  ( new_n39945_, new_n39944_, new_n39806_ );
or   ( new_n39946_, new_n8874_, new_n26196_ );
or   ( new_n39947_, new_n8876_, new_n25813_ );
and  ( new_n39948_, new_n39947_, new_n39946_ );
xor  ( new_n39949_, new_n39948_, new_n8257_ );
or   ( new_n39950_, new_n8264_, new_n26372_ );
or   ( new_n39951_, new_n8266_, new_n26063_ );
and  ( new_n39952_, new_n39951_, new_n39950_ );
xor  ( new_n39953_, new_n39952_, new_n7725_ );
or   ( new_n39954_, new_n39953_, new_n39949_ );
and  ( new_n39955_, new_n39953_, new_n39949_ );
or   ( new_n39956_, new_n7732_, new_n26762_ );
or   ( new_n39957_, new_n7734_, new_n26620_ );
and  ( new_n39958_, new_n39957_, new_n39956_ );
xor  ( new_n39959_, new_n39958_, new_n7177_ );
or   ( new_n39960_, new_n39959_, new_n39955_ );
and  ( new_n39961_, new_n39960_, new_n39954_ );
or   ( new_n39962_, new_n7184_, new_n27396_ );
or   ( new_n39963_, new_n7186_, new_n27085_ );
and  ( new_n39964_, new_n39963_, new_n39962_ );
xor  ( new_n39965_, new_n39964_, new_n6638_ );
or   ( new_n39966_, new_n6645_, new_n27763_ );
or   ( new_n39967_, new_n6647_, new_n27602_ );
and  ( new_n39968_, new_n39967_, new_n39966_ );
xor  ( new_n39969_, new_n39968_, new_n6166_ );
or   ( new_n39970_, new_n39969_, new_n39965_ );
and  ( new_n39971_, new_n39969_, new_n39965_ );
or   ( new_n39972_, new_n6173_, new_n28314_ );
or   ( new_n39973_, new_n6175_, new_n28108_ );
and  ( new_n39974_, new_n39973_, new_n39972_ );
xor  ( new_n39975_, new_n39974_, new_n5597_ );
or   ( new_n39976_, new_n39975_, new_n39971_ );
and  ( new_n39977_, new_n39976_, new_n39970_ );
or   ( new_n39978_, new_n39977_, new_n39961_ );
and  ( new_n39979_, new_n39977_, new_n39961_ );
or   ( new_n39980_, new_n10059_, new_n25048_ );
or   ( new_n39981_, new_n10061_, new_n24925_ );
and  ( new_n39982_, new_n39981_, new_n39980_ );
xor  ( new_n39983_, new_n39982_, new_n9421_ );
and  ( new_n39984_, RIbb325e0_163, RIbb2d888_64 );
or   ( new_n39985_, new_n24927_, RIbb2d888_64 );
and  ( new_n39986_, new_n39985_, RIbb2d900_63 );
or   ( new_n39987_, new_n39986_, new_n39984_ );
or   ( new_n39988_, new_n10770_, new_n24543_ );
and  ( new_n39989_, new_n39988_, new_n39987_ );
nor  ( new_n39990_, new_n39989_, new_n39983_ );
and  ( new_n39991_, new_n39989_, new_n39983_ );
or   ( new_n39992_, new_n9422_, new_n25486_ );
or   ( new_n39993_, new_n9424_, new_n25288_ );
and  ( new_n39994_, new_n39993_, new_n39992_ );
xor  ( new_n39995_, new_n39994_, new_n8873_ );
nor  ( new_n39996_, new_n39995_, new_n39991_ );
nor  ( new_n39997_, new_n39996_, new_n39990_ );
or   ( new_n39998_, new_n39997_, new_n39979_ );
and  ( new_n39999_, new_n39998_, new_n39978_ );
or   ( new_n40000_, new_n3461_, new_n31654_ );
or   ( new_n40001_, new_n3463_, new_n31333_ );
and  ( new_n40002_, new_n40001_, new_n40000_ );
xor  ( new_n40003_, new_n40002_, new_n3116_ );
or   ( new_n40004_, new_n4302_, new_n30800_ );
or   ( new_n40005_, new_n4304_, new_n30227_ );
and  ( new_n40006_, new_n40005_, new_n40004_ );
xor  ( new_n40007_, new_n40006_, new_n3895_ );
or   ( new_n40008_, new_n3896_, new_n31333_ );
or   ( new_n40009_, new_n3898_, new_n30798_ );
and  ( new_n40010_, new_n40009_, new_n40008_ );
xor  ( new_n40011_, new_n40010_, new_n3460_ );
or   ( new_n40012_, new_n40011_, new_n40007_ );
and  ( new_n40013_, new_n40011_, new_n40007_ );
or   ( new_n40014_, new_n3461_, new_n31952_ );
or   ( new_n40015_, new_n3463_, new_n31654_ );
and  ( new_n40016_, new_n40015_, new_n40014_ );
xor  ( new_n40017_, new_n40016_, new_n3116_ );
or   ( new_n40018_, new_n40017_, new_n40013_ );
and  ( new_n40019_, new_n40018_, new_n40012_ );
or   ( new_n40020_, new_n40019_, new_n40003_ );
and  ( new_n40021_, new_n40019_, new_n40003_ );
or   ( new_n40022_, new_n5604_, new_n29263_ );
or   ( new_n40023_, new_n5606_, new_n28531_ );
and  ( new_n40024_, new_n40023_, new_n40022_ );
xor  ( new_n40025_, new_n40024_, new_n5206_ );
or   ( new_n40026_, new_n5207_, new_n29474_ );
or   ( new_n40027_, new_n5209_, new_n29261_ );
and  ( new_n40028_, new_n40027_, new_n40026_ );
xor  ( new_n40029_, new_n40028_, new_n4708_ );
nor  ( new_n40030_, new_n40029_, new_n40025_ );
and  ( new_n40031_, new_n40029_, new_n40025_ );
or   ( new_n40032_, new_n4709_, new_n30120_ );
or   ( new_n40033_, new_n4711_, new_n29619_ );
and  ( new_n40034_, new_n40033_, new_n40032_ );
xor  ( new_n40035_, new_n40034_, new_n4295_ );
nor  ( new_n40036_, new_n40035_, new_n40031_ );
nor  ( new_n40037_, new_n40036_, new_n40030_ );
or   ( new_n40038_, new_n40037_, new_n40021_ );
and  ( new_n40039_, new_n40038_, new_n40020_ );
nor  ( new_n40040_, new_n40039_, new_n39999_ );
nand ( new_n40041_, new_n40039_, new_n39999_ );
and  ( new_n40042_, new_n2928_, RIbb33378_192 );
or   ( new_n40043_, new_n40042_, new_n2800_ );
nand ( new_n40044_, new_n40042_, new_n2797_ );
and  ( new_n40045_, new_n40044_, new_n40043_ );
xnor ( new_n40046_, new_n39845_, new_n39841_ );
xor  ( new_n40047_, new_n40046_, new_n39851_ );
nor  ( new_n40048_, new_n40047_, new_n40045_ );
and  ( new_n40049_, new_n40047_, new_n40045_ );
xor  ( new_n40050_, new_n39827_, new_n39823_ );
xnor ( new_n40051_, new_n40050_, new_n39833_ );
nor  ( new_n40052_, new_n40051_, new_n40049_ );
nor  ( new_n40053_, new_n40052_, new_n40048_ );
and  ( new_n40054_, new_n40053_, new_n40041_ );
or   ( new_n40055_, new_n40054_, new_n40040_ );
xor  ( new_n40056_, new_n39911_, new_n39909_ );
xor  ( new_n40057_, new_n40056_, new_n39915_ );
xnor ( new_n40058_, new_n39835_, new_n39819_ );
xor  ( new_n40059_, new_n40058_, new_n39853_ );
or   ( new_n40060_, new_n40059_, new_n40057_ );
and  ( new_n40061_, new_n40059_, new_n40057_ );
xnor ( new_n40062_, new_n39901_, new_n39885_ );
xnor ( new_n40063_, new_n40062_, new_n39871_ );
not  ( new_n40064_, new_n40063_ );
or   ( new_n40065_, new_n40064_, new_n40061_ );
and  ( new_n40066_, new_n40065_, new_n40060_ );
nand ( new_n40067_, new_n40066_, new_n40055_ );
or   ( new_n40068_, new_n40066_, new_n40055_ );
xnor ( new_n40069_, new_n39692_, new_n39688_ );
xor  ( new_n40070_, new_n40069_, new_n39698_ );
xnor ( new_n40071_, new_n39863_, new_n39859_ );
xor  ( new_n40072_, new_n40071_, new_n39869_ );
xnor ( new_n40073_, new_n39893_, new_n39889_ );
xor  ( new_n40074_, new_n40073_, new_n39899_ );
or   ( new_n40075_, new_n40074_, new_n40072_ );
and  ( new_n40076_, new_n40074_, new_n40072_ );
xor  ( new_n40077_, new_n39881_, new_n39875_ );
xor  ( new_n40078_, new_n40077_, new_n2800_ );
or   ( new_n40079_, new_n40078_, new_n40076_ );
and  ( new_n40080_, new_n40079_, new_n40075_ );
nor  ( new_n40081_, new_n40080_, new_n40070_ );
and  ( new_n40082_, new_n40080_, new_n40070_ );
xor  ( new_n40083_, new_n39676_, new_n39670_ );
xnor ( new_n40084_, new_n40083_, new_n39682_ );
nor  ( new_n40085_, new_n40084_, new_n40082_ );
nor  ( new_n40086_, new_n40085_, new_n40081_ );
nand ( new_n40087_, new_n40086_, new_n40068_ );
and  ( new_n40088_, new_n40087_, new_n40067_ );
or   ( new_n40089_, new_n40088_, new_n39945_ );
nand ( new_n40090_, new_n40088_, new_n39945_ );
xor  ( new_n40091_, new_n39925_, new_n39923_ );
xor  ( new_n40092_, new_n40091_, new_n39930_ );
xnor ( new_n40093_, new_n39905_, new_n39855_ );
xor  ( new_n40094_, new_n40093_, new_n39917_ );
and  ( new_n40095_, new_n40094_, new_n40092_ );
nor  ( new_n40096_, new_n40094_, new_n40092_ );
xor  ( new_n40097_, new_n39814_, new_n39812_ );
not  ( new_n40098_, new_n40097_ );
nor  ( new_n40099_, new_n40098_, new_n40096_ );
nor  ( new_n40100_, new_n40099_, new_n40095_ );
nand ( new_n40101_, new_n40100_, new_n40090_ );
and  ( new_n40102_, new_n40101_, new_n40089_ );
xnor ( new_n40103_, new_n39808_, new_n39798_ );
xor  ( new_n40104_, new_n40103_, new_n39934_ );
nor  ( new_n40105_, new_n40104_, new_n40102_ );
nand ( new_n40106_, new_n40104_, new_n40102_ );
xnor ( new_n40107_, new_n39795_, new_n39793_ );
and  ( new_n40108_, new_n40107_, new_n40106_ );
or   ( new_n40109_, new_n40108_, new_n40105_ );
xor  ( new_n40110_, new_n39936_, new_n39796_ );
xor  ( new_n40111_, new_n40110_, new_n39940_ );
nor  ( new_n40112_, new_n40111_, new_n40109_ );
xor  ( new_n40113_, new_n40104_, new_n40102_ );
xor  ( new_n40114_, new_n40113_, new_n40107_ );
xor  ( new_n40115_, new_n40039_, new_n39999_ );
xnor ( new_n40116_, new_n40115_, new_n40053_ );
xnor ( new_n40117_, new_n40080_, new_n40070_ );
xor  ( new_n40118_, new_n40117_, new_n40084_ );
nand ( new_n40119_, new_n40118_, new_n40116_ );
xor  ( new_n40120_, new_n40074_, new_n40072_ );
xor  ( new_n40121_, new_n40120_, new_n40078_ );
xnor ( new_n40122_, new_n40019_, new_n40003_ );
xor  ( new_n40123_, new_n40122_, new_n40037_ );
or   ( new_n40124_, new_n40123_, new_n40121_ );
nand ( new_n40125_, new_n40123_, new_n40121_ );
xor  ( new_n40126_, new_n40047_, new_n40045_ );
xnor ( new_n40127_, new_n40126_, new_n40051_ );
nand ( new_n40128_, new_n40127_, new_n40125_ );
and  ( new_n40129_, new_n40128_, new_n40124_ );
xor  ( new_n40130_, new_n40011_, new_n40007_ );
xor  ( new_n40131_, new_n40130_, new_n40017_ );
or   ( new_n40132_, new_n6173_, new_n28531_ );
or   ( new_n40133_, new_n6175_, new_n28314_ );
and  ( new_n40134_, new_n40133_, new_n40132_ );
xor  ( new_n40135_, new_n40134_, new_n5597_ );
or   ( new_n40136_, new_n5604_, new_n29261_ );
or   ( new_n40137_, new_n5606_, new_n29263_ );
and  ( new_n40138_, new_n40137_, new_n40136_ );
xor  ( new_n40139_, new_n40138_, new_n5206_ );
or   ( new_n40140_, new_n40139_, new_n40135_ );
and  ( new_n40141_, new_n40139_, new_n40135_ );
or   ( new_n40142_, new_n5207_, new_n29619_ );
or   ( new_n40143_, new_n5209_, new_n29474_ );
and  ( new_n40144_, new_n40143_, new_n40142_ );
xor  ( new_n40145_, new_n40144_, new_n4708_ );
or   ( new_n40146_, new_n40145_, new_n40141_ );
and  ( new_n40147_, new_n40146_, new_n40140_ );
or   ( new_n40148_, new_n40147_, new_n40131_ );
and  ( new_n40149_, new_n40147_, new_n40131_ );
or   ( new_n40150_, new_n4709_, new_n30227_ );
or   ( new_n40151_, new_n4711_, new_n30120_ );
and  ( new_n40152_, new_n40151_, new_n40150_ );
xor  ( new_n40153_, new_n40152_, new_n4295_ );
or   ( new_n40154_, new_n4302_, new_n30798_ );
or   ( new_n40155_, new_n4304_, new_n30800_ );
and  ( new_n40156_, new_n40155_, new_n40154_ );
xor  ( new_n40157_, new_n40156_, new_n3895_ );
nor  ( new_n40158_, new_n40157_, new_n40153_ );
and  ( new_n40159_, new_n40157_, new_n40153_ );
or   ( new_n40160_, new_n3896_, new_n31654_ );
or   ( new_n40161_, new_n3898_, new_n31333_ );
and  ( new_n40162_, new_n40161_, new_n40160_ );
xor  ( new_n40163_, new_n40162_, new_n3460_ );
nor  ( new_n40164_, new_n40163_, new_n40159_ );
nor  ( new_n40165_, new_n40164_, new_n40158_ );
or   ( new_n40166_, new_n40165_, new_n40149_ );
and  ( new_n40167_, new_n40166_, new_n40148_ );
or   ( new_n40168_, new_n7732_, new_n27085_ );
or   ( new_n40169_, new_n7734_, new_n26762_ );
and  ( new_n40170_, new_n40169_, new_n40168_ );
xor  ( new_n40171_, new_n40170_, new_n7177_ );
or   ( new_n40172_, new_n7184_, new_n27602_ );
or   ( new_n40173_, new_n7186_, new_n27396_ );
and  ( new_n40174_, new_n40173_, new_n40172_ );
xor  ( new_n40175_, new_n40174_, new_n6638_ );
nor  ( new_n40176_, new_n40175_, new_n40171_ );
and  ( new_n40177_, new_n40175_, new_n40171_ );
or   ( new_n40178_, new_n6645_, new_n28108_ );
or   ( new_n40179_, new_n6647_, new_n27763_ );
and  ( new_n40180_, new_n40179_, new_n40178_ );
xor  ( new_n40181_, new_n40180_, new_n6166_ );
nor  ( new_n40182_, new_n40181_, new_n40177_ );
nor  ( new_n40183_, new_n40182_, new_n40176_ );
or   ( new_n40184_, new_n10059_, new_n25288_ );
or   ( new_n40185_, new_n10061_, new_n25048_ );
and  ( new_n40186_, new_n40185_, new_n40184_ );
xor  ( new_n40187_, new_n40186_, new_n9421_ );
and  ( new_n40188_, RIbb32658_164, RIbb2d888_64 );
or   ( new_n40189_, new_n24925_, RIbb2d888_64 );
and  ( new_n40190_, new_n40189_, RIbb2d900_63 );
or   ( new_n40191_, new_n40190_, new_n40188_ );
or   ( new_n40192_, new_n10770_, new_n24927_ );
and  ( new_n40193_, new_n40192_, new_n40191_ );
nor  ( new_n40194_, new_n40193_, new_n40187_ );
and  ( new_n40195_, new_n40193_, new_n40187_ );
nor  ( new_n40196_, new_n40195_, new_n3115_ );
nor  ( new_n40197_, new_n40196_, new_n40194_ );
or   ( new_n40198_, new_n9422_, new_n25813_ );
or   ( new_n40199_, new_n9424_, new_n25486_ );
and  ( new_n40200_, new_n40199_, new_n40198_ );
xor  ( new_n40201_, new_n40200_, new_n8873_ );
or   ( new_n40202_, new_n8874_, new_n26063_ );
or   ( new_n40203_, new_n8876_, new_n26196_ );
and  ( new_n40204_, new_n40203_, new_n40202_ );
xor  ( new_n40205_, new_n40204_, new_n8257_ );
or   ( new_n40206_, new_n40205_, new_n40201_ );
and  ( new_n40207_, new_n40205_, new_n40201_ );
or   ( new_n40208_, new_n8264_, new_n26620_ );
or   ( new_n40209_, new_n8266_, new_n26372_ );
and  ( new_n40210_, new_n40209_, new_n40208_ );
xor  ( new_n40211_, new_n40210_, new_n7725_ );
or   ( new_n40212_, new_n40211_, new_n40207_ );
and  ( new_n40213_, new_n40212_, new_n40206_ );
and  ( new_n40214_, new_n40213_, new_n40197_ );
or   ( new_n40215_, new_n40214_, new_n40183_ );
or   ( new_n40216_, new_n40213_, new_n40197_ );
and  ( new_n40217_, new_n40216_, new_n40215_ );
nand ( new_n40218_, new_n40217_, new_n40167_ );
nor  ( new_n40219_, new_n40217_, new_n40167_ );
xnor ( new_n40220_, new_n39969_, new_n39965_ );
xor  ( new_n40221_, new_n40220_, new_n39975_ );
xnor ( new_n40222_, new_n39953_, new_n39949_ );
xor  ( new_n40223_, new_n40222_, new_n39959_ );
nor  ( new_n40224_, new_n40223_, new_n40221_ );
and  ( new_n40225_, new_n40223_, new_n40221_ );
xor  ( new_n40226_, new_n40029_, new_n40025_ );
xnor ( new_n40227_, new_n40226_, new_n40035_ );
nor  ( new_n40228_, new_n40227_, new_n40225_ );
nor  ( new_n40229_, new_n40228_, new_n40224_ );
or   ( new_n40230_, new_n40229_, new_n40219_ );
and  ( new_n40231_, new_n40230_, new_n40218_ );
or   ( new_n40232_, new_n40231_, new_n40129_ );
and  ( new_n40233_, new_n40231_, new_n40129_ );
xor  ( new_n40234_, new_n40059_, new_n40057_ );
xor  ( new_n40235_, new_n40234_, new_n40064_ );
or   ( new_n40236_, new_n40235_, new_n40233_ );
and  ( new_n40237_, new_n40236_, new_n40232_ );
nor  ( new_n40238_, new_n40237_, new_n40119_ );
nand ( new_n40239_, new_n40237_, new_n40119_ );
xor  ( new_n40240_, new_n40094_, new_n40092_ );
xor  ( new_n40241_, new_n40240_, new_n40097_ );
and  ( new_n40242_, new_n40241_, new_n40239_ );
or   ( new_n40243_, new_n40242_, new_n40238_ );
xnor ( new_n40244_, new_n39919_, new_n39815_ );
xor  ( new_n40245_, new_n40244_, new_n39932_ );
nand ( new_n40246_, new_n40245_, new_n40243_ );
nor  ( new_n40247_, new_n40245_, new_n40243_ );
xor  ( new_n40248_, new_n40088_, new_n39945_ );
xor  ( new_n40249_, new_n40248_, new_n40100_ );
or   ( new_n40250_, new_n40249_, new_n40247_ );
and  ( new_n40251_, new_n40250_, new_n40246_ );
nor  ( new_n40252_, new_n40251_, new_n40114_ );
xor  ( new_n40253_, new_n40245_, new_n40243_ );
xor  ( new_n40254_, new_n40253_, new_n40249_ );
or   ( new_n40255_, new_n7184_, new_n27763_ );
or   ( new_n40256_, new_n7186_, new_n27602_ );
and  ( new_n40257_, new_n40256_, new_n40255_ );
xor  ( new_n40258_, new_n40257_, new_n6638_ );
or   ( new_n40259_, new_n6645_, new_n28314_ );
or   ( new_n40260_, new_n6647_, new_n28108_ );
and  ( new_n40261_, new_n40260_, new_n40259_ );
xor  ( new_n40262_, new_n40261_, new_n6166_ );
or   ( new_n40263_, new_n40262_, new_n40258_ );
and  ( new_n40264_, new_n40262_, new_n40258_ );
or   ( new_n40265_, new_n6173_, new_n29263_ );
or   ( new_n40266_, new_n6175_, new_n28531_ );
and  ( new_n40267_, new_n40266_, new_n40265_ );
xor  ( new_n40268_, new_n40267_, new_n5597_ );
or   ( new_n40269_, new_n40268_, new_n40264_ );
and  ( new_n40270_, new_n40269_, new_n40263_ );
or   ( new_n40271_, new_n10059_, new_n25486_ );
or   ( new_n40272_, new_n10061_, new_n25288_ );
and  ( new_n40273_, new_n40272_, new_n40271_ );
xor  ( new_n40274_, new_n40273_, new_n9421_ );
and  ( new_n40275_, RIbb326d0_165, RIbb2d888_64 );
or   ( new_n40276_, new_n25048_, RIbb2d888_64 );
and  ( new_n40277_, new_n40276_, RIbb2d900_63 );
or   ( new_n40278_, new_n40277_, new_n40275_ );
or   ( new_n40279_, new_n10770_, new_n24925_ );
and  ( new_n40280_, new_n40279_, new_n40278_ );
or   ( new_n40281_, new_n40280_, new_n40274_ );
and  ( new_n40282_, new_n40280_, new_n40274_ );
or   ( new_n40283_, new_n9422_, new_n26196_ );
or   ( new_n40284_, new_n9424_, new_n25813_ );
and  ( new_n40285_, new_n40284_, new_n40283_ );
xor  ( new_n40286_, new_n40285_, new_n8873_ );
or   ( new_n40287_, new_n40286_, new_n40282_ );
and  ( new_n40288_, new_n40287_, new_n40281_ );
nor  ( new_n40289_, new_n40288_, new_n40270_ );
nand ( new_n40290_, new_n40288_, new_n40270_ );
or   ( new_n40291_, new_n8874_, new_n26372_ );
or   ( new_n40292_, new_n8876_, new_n26063_ );
and  ( new_n40293_, new_n40292_, new_n40291_ );
xor  ( new_n40294_, new_n40293_, new_n8257_ );
or   ( new_n40295_, new_n8264_, new_n26762_ );
or   ( new_n40296_, new_n8266_, new_n26620_ );
and  ( new_n40297_, new_n40296_, new_n40295_ );
xor  ( new_n40298_, new_n40297_, new_n7725_ );
nor  ( new_n40299_, new_n40298_, new_n40294_ );
nand ( new_n40300_, new_n40298_, new_n40294_ );
or   ( new_n40301_, new_n7732_, new_n27396_ );
or   ( new_n40302_, new_n7734_, new_n27085_ );
and  ( new_n40303_, new_n40302_, new_n40301_ );
xor  ( new_n40304_, new_n40303_, new_n7176_ );
and  ( new_n40305_, new_n40304_, new_n40300_ );
or   ( new_n40306_, new_n40305_, new_n40299_ );
and  ( new_n40307_, new_n40306_, new_n40290_ );
or   ( new_n40308_, new_n40307_, new_n40289_ );
and  ( new_n40309_, new_n3291_, RIbb33378_192 );
or   ( new_n40310_, new_n40309_, new_n3116_ );
nand ( new_n40311_, new_n40309_, new_n3113_ );
and  ( new_n40312_, new_n40311_, new_n40310_ );
xnor ( new_n40313_, new_n40157_, new_n40153_ );
xor  ( new_n40314_, new_n40313_, new_n40163_ );
or   ( new_n40315_, new_n40314_, new_n40312_ );
and  ( new_n40316_, new_n40314_, new_n40312_ );
or   ( new_n40317_, new_n5604_, new_n29474_ );
or   ( new_n40318_, new_n5606_, new_n29261_ );
and  ( new_n40319_, new_n40318_, new_n40317_ );
xor  ( new_n40320_, new_n40319_, new_n5206_ );
or   ( new_n40321_, new_n5207_, new_n30120_ );
or   ( new_n40322_, new_n5209_, new_n29619_ );
and  ( new_n40323_, new_n40322_, new_n40321_ );
xor  ( new_n40324_, new_n40323_, new_n4708_ );
nor  ( new_n40325_, new_n40324_, new_n40320_ );
and  ( new_n40326_, new_n40324_, new_n40320_ );
or   ( new_n40327_, new_n4709_, new_n30800_ );
or   ( new_n40328_, new_n4711_, new_n30227_ );
and  ( new_n40329_, new_n40328_, new_n40327_ );
xor  ( new_n40330_, new_n40329_, new_n4295_ );
nor  ( new_n40331_, new_n40330_, new_n40326_ );
nor  ( new_n40332_, new_n40331_, new_n40325_ );
not  ( new_n40333_, new_n40332_ );
or   ( new_n40334_, new_n40333_, new_n40316_ );
and  ( new_n40335_, new_n40334_, new_n40315_ );
and  ( new_n40336_, new_n40335_, new_n40308_ );
xnor ( new_n40337_, new_n40175_, new_n40171_ );
xor  ( new_n40338_, new_n40337_, new_n40181_ );
xnor ( new_n40339_, new_n40205_, new_n40201_ );
xor  ( new_n40340_, new_n40339_, new_n40211_ );
nor  ( new_n40341_, new_n40340_, new_n40338_ );
and  ( new_n40342_, new_n40340_, new_n40338_ );
xor  ( new_n40343_, new_n40139_, new_n40135_ );
xnor ( new_n40344_, new_n40343_, new_n40145_ );
nor  ( new_n40345_, new_n40344_, new_n40342_ );
nor  ( new_n40346_, new_n40345_, new_n40341_ );
or   ( new_n40347_, new_n40346_, new_n40336_ );
or   ( new_n40348_, new_n40335_, new_n40308_ );
and  ( new_n40349_, new_n40348_, new_n40347_ );
xnor ( new_n40350_, new_n39977_, new_n39961_ );
xor  ( new_n40351_, new_n40350_, new_n39997_ );
and  ( new_n40352_, new_n40351_, new_n40349_ );
xor  ( new_n40353_, new_n40223_, new_n40221_ );
xor  ( new_n40354_, new_n40353_, new_n40227_ );
xnor ( new_n40355_, new_n40147_, new_n40131_ );
xor  ( new_n40356_, new_n40355_, new_n40165_ );
nor  ( new_n40357_, new_n40356_, new_n40354_ );
and  ( new_n40358_, new_n40356_, new_n40354_ );
xor  ( new_n40359_, new_n39989_, new_n39983_ );
xnor ( new_n40360_, new_n40359_, new_n39995_ );
nor  ( new_n40361_, new_n40360_, new_n40358_ );
nor  ( new_n40362_, new_n40361_, new_n40357_ );
nor  ( new_n40363_, new_n40362_, new_n40352_ );
nor  ( new_n40364_, new_n40351_, new_n40349_ );
or   ( new_n40365_, new_n40364_, new_n40363_ );
xnor ( new_n40366_, new_n40231_, new_n40129_ );
xor  ( new_n40367_, new_n40366_, new_n40235_ );
nor  ( new_n40368_, new_n40367_, new_n40365_ );
nand ( new_n40369_, new_n40367_, new_n40365_ );
xnor ( new_n40370_, new_n40118_, new_n40116_ );
and  ( new_n40371_, new_n40370_, new_n40369_ );
or   ( new_n40372_, new_n40371_, new_n40368_ );
xor  ( new_n40373_, new_n40066_, new_n40055_ );
xor  ( new_n40374_, new_n40373_, new_n40086_ );
or   ( new_n40375_, new_n40374_, new_n40372_ );
and  ( new_n40376_, new_n40374_, new_n40372_ );
xnor ( new_n40377_, new_n40237_, new_n40119_ );
xor  ( new_n40378_, new_n40377_, new_n40241_ );
or   ( new_n40379_, new_n40378_, new_n40376_ );
and  ( new_n40380_, new_n40379_, new_n40375_ );
nor  ( new_n40381_, new_n40380_, new_n40254_ );
xor  ( new_n40382_, new_n40374_, new_n40372_ );
xor  ( new_n40383_, new_n40382_, new_n40378_ );
xor  ( new_n40384_, new_n40351_, new_n40349_ );
xor  ( new_n40385_, new_n40384_, new_n40362_ );
xnor ( new_n40386_, new_n40217_, new_n40167_ );
xnor ( new_n40387_, new_n40386_, new_n40229_ );
nor  ( new_n40388_, new_n40387_, new_n40385_ );
xor  ( new_n40389_, new_n40335_, new_n40308_ );
xor  ( new_n40390_, new_n40389_, new_n40346_ );
xnor ( new_n40391_, new_n40356_, new_n40354_ );
xnor ( new_n40392_, new_n40391_, new_n40360_ );
nor  ( new_n40393_, new_n40392_, new_n40390_ );
xor  ( new_n40394_, new_n40123_, new_n40121_ );
xor  ( new_n40395_, new_n40394_, new_n40127_ );
or   ( new_n40396_, new_n40395_, new_n40393_ );
and  ( new_n40397_, new_n40395_, new_n40393_ );
or   ( new_n40398_, new_n4302_, new_n31333_ );
or   ( new_n40399_, new_n4304_, new_n30798_ );
and  ( new_n40400_, new_n40399_, new_n40398_ );
xor  ( new_n40401_, new_n40400_, new_n3895_ );
or   ( new_n40402_, new_n6173_, new_n29261_ );
or   ( new_n40403_, new_n6175_, new_n29263_ );
and  ( new_n40404_, new_n40403_, new_n40402_ );
xor  ( new_n40405_, new_n40404_, new_n5597_ );
or   ( new_n40406_, new_n5604_, new_n29619_ );
or   ( new_n40407_, new_n5606_, new_n29474_ );
and  ( new_n40408_, new_n40407_, new_n40406_ );
xor  ( new_n40409_, new_n40408_, new_n5206_ );
or   ( new_n40410_, new_n40409_, new_n40405_ );
and  ( new_n40411_, new_n40409_, new_n40405_ );
or   ( new_n40412_, new_n5207_, new_n30227_ );
or   ( new_n40413_, new_n5209_, new_n30120_ );
and  ( new_n40414_, new_n40413_, new_n40412_ );
xor  ( new_n40415_, new_n40414_, new_n4708_ );
or   ( new_n40416_, new_n40415_, new_n40411_ );
and  ( new_n40417_, new_n40416_, new_n40410_ );
or   ( new_n40418_, new_n40417_, new_n40401_ );
nand ( new_n40419_, new_n40417_, new_n40401_ );
or   ( new_n40420_, new_n4709_, new_n30798_ );
or   ( new_n40421_, new_n4711_, new_n30800_ );
and  ( new_n40422_, new_n40421_, new_n40420_ );
xor  ( new_n40423_, new_n40422_, new_n4295_ );
or   ( new_n40424_, new_n4302_, new_n31654_ );
or   ( new_n40425_, new_n4304_, new_n31333_ );
and  ( new_n40426_, new_n40425_, new_n40424_ );
xor  ( new_n40427_, new_n40426_, new_n3895_ );
and  ( new_n40428_, new_n40427_, new_n40423_ );
nor  ( new_n40429_, new_n40427_, new_n40423_ );
and  ( new_n40430_, new_n3731_, RIbb33378_192 );
nor  ( new_n40431_, new_n40430_, new_n3460_ );
and  ( new_n40432_, new_n40430_, new_n3457_ );
nor  ( new_n40433_, new_n40432_, new_n40431_ );
nor  ( new_n40434_, new_n40433_, new_n40429_ );
nor  ( new_n40435_, new_n40434_, new_n40428_ );
nand ( new_n40436_, new_n40435_, new_n40419_ );
and  ( new_n40437_, new_n40436_, new_n40418_ );
or   ( new_n40438_, new_n7732_, new_n27602_ );
or   ( new_n40439_, new_n7734_, new_n27396_ );
and  ( new_n40440_, new_n40439_, new_n40438_ );
xor  ( new_n40441_, new_n40440_, new_n7177_ );
or   ( new_n40442_, new_n7184_, new_n28108_ );
or   ( new_n40443_, new_n7186_, new_n27763_ );
and  ( new_n40444_, new_n40443_, new_n40442_ );
xor  ( new_n40445_, new_n40444_, new_n6638_ );
nor  ( new_n40446_, new_n40445_, new_n40441_ );
and  ( new_n40447_, new_n40445_, new_n40441_ );
or   ( new_n40448_, new_n6645_, new_n28531_ );
or   ( new_n40449_, new_n6647_, new_n28314_ );
and  ( new_n40450_, new_n40449_, new_n40448_ );
xor  ( new_n40451_, new_n40450_, new_n6166_ );
nor  ( new_n40452_, new_n40451_, new_n40447_ );
nor  ( new_n40453_, new_n40452_, new_n40446_ );
or   ( new_n40454_, new_n10059_, new_n25813_ );
or   ( new_n40455_, new_n10061_, new_n25486_ );
and  ( new_n40456_, new_n40455_, new_n40454_ );
xor  ( new_n40457_, new_n40456_, new_n9421_ );
and  ( new_n40458_, RIbb32748_166, RIbb2d888_64 );
or   ( new_n40459_, new_n25288_, RIbb2d888_64 );
and  ( new_n40460_, new_n40459_, RIbb2d900_63 );
or   ( new_n40461_, new_n40460_, new_n40458_ );
or   ( new_n40462_, new_n10770_, new_n25048_ );
and  ( new_n40463_, new_n40462_, new_n40461_ );
nor  ( new_n40464_, new_n40463_, new_n40457_ );
and  ( new_n40465_, new_n40463_, new_n40457_ );
nor  ( new_n40466_, new_n40465_, new_n3459_ );
nor  ( new_n40467_, new_n40466_, new_n40464_ );
or   ( new_n40468_, new_n9422_, new_n26063_ );
or   ( new_n40469_, new_n9424_, new_n26196_ );
and  ( new_n40470_, new_n40469_, new_n40468_ );
xor  ( new_n40471_, new_n40470_, new_n8873_ );
or   ( new_n40472_, new_n8874_, new_n26620_ );
or   ( new_n40473_, new_n8876_, new_n26372_ );
and  ( new_n40474_, new_n40473_, new_n40472_ );
xor  ( new_n40475_, new_n40474_, new_n8257_ );
or   ( new_n40476_, new_n40475_, new_n40471_ );
and  ( new_n40477_, new_n40475_, new_n40471_ );
or   ( new_n40478_, new_n8264_, new_n27085_ );
or   ( new_n40479_, new_n8266_, new_n26762_ );
and  ( new_n40480_, new_n40479_, new_n40478_ );
xor  ( new_n40481_, new_n40480_, new_n7725_ );
or   ( new_n40482_, new_n40481_, new_n40477_ );
and  ( new_n40483_, new_n40482_, new_n40476_ );
and  ( new_n40484_, new_n40483_, new_n40467_ );
or   ( new_n40485_, new_n40484_, new_n40453_ );
or   ( new_n40486_, new_n40483_, new_n40467_ );
and  ( new_n40487_, new_n40486_, new_n40485_ );
nor  ( new_n40488_, new_n40487_, new_n40437_ );
nand ( new_n40489_, new_n40487_, new_n40437_ );
or   ( new_n40490_, new_n3896_, new_n31952_ );
or   ( new_n40491_, new_n3898_, new_n31654_ );
and  ( new_n40492_, new_n40491_, new_n40490_ );
xor  ( new_n40493_, new_n40492_, new_n3459_ );
xnor ( new_n40494_, new_n40324_, new_n40320_ );
xor  ( new_n40495_, new_n40494_, new_n40330_ );
and  ( new_n40496_, new_n40495_, new_n40493_ );
or   ( new_n40497_, new_n40495_, new_n40493_ );
xor  ( new_n40498_, new_n40262_, new_n40258_ );
xnor ( new_n40499_, new_n40498_, new_n40268_ );
and  ( new_n40500_, new_n40499_, new_n40497_ );
or   ( new_n40501_, new_n40500_, new_n40496_ );
and  ( new_n40502_, new_n40501_, new_n40489_ );
or   ( new_n40503_, new_n40502_, new_n40488_ );
xor  ( new_n40504_, new_n40193_, new_n40187_ );
xnor ( new_n40505_, new_n40504_, new_n3116_ );
xnor ( new_n40506_, new_n40340_, new_n40338_ );
xor  ( new_n40507_, new_n40506_, new_n40344_ );
nand ( new_n40508_, new_n40507_, new_n40505_ );
nor  ( new_n40509_, new_n40507_, new_n40505_ );
xor  ( new_n40510_, new_n40314_, new_n40312_ );
xor  ( new_n40511_, new_n40510_, new_n40333_ );
or   ( new_n40512_, new_n40511_, new_n40509_ );
and  ( new_n40513_, new_n40512_, new_n40508_ );
and  ( new_n40514_, new_n40513_, new_n40503_ );
nor  ( new_n40515_, new_n40513_, new_n40503_ );
xnor ( new_n40516_, new_n40213_, new_n40197_ );
xnor ( new_n40517_, new_n40516_, new_n40183_ );
nor  ( new_n40518_, new_n40517_, new_n40515_ );
nor  ( new_n40519_, new_n40518_, new_n40514_ );
or   ( new_n40520_, new_n40519_, new_n40397_ );
and  ( new_n40521_, new_n40520_, new_n40396_ );
nand ( new_n40522_, new_n40521_, new_n40388_ );
nor  ( new_n40523_, new_n40521_, new_n40388_ );
xor  ( new_n40524_, new_n40367_, new_n40365_ );
xor  ( new_n40525_, new_n40524_, new_n40370_ );
or   ( new_n40526_, new_n40525_, new_n40523_ );
and  ( new_n40527_, new_n40526_, new_n40522_ );
nor  ( new_n40528_, new_n40527_, new_n40383_ );
xor  ( new_n40529_, new_n40521_, new_n40388_ );
xor  ( new_n40530_, new_n40529_, new_n40525_ );
xor  ( new_n40531_, new_n40288_, new_n40270_ );
xor  ( new_n40532_, new_n40531_, new_n40306_ );
xnor ( new_n40533_, new_n40280_, new_n40274_ );
xor  ( new_n40534_, new_n40533_, new_n40286_ );
xor  ( new_n40535_, new_n40298_, new_n40294_ );
xor  ( new_n40536_, new_n40535_, new_n40304_ );
or   ( new_n40537_, new_n40536_, new_n40534_ );
and  ( new_n40538_, new_n40536_, new_n40534_ );
xor  ( new_n40539_, new_n40495_, new_n40493_ );
xor  ( new_n40540_, new_n40539_, new_n40499_ );
or   ( new_n40541_, new_n40540_, new_n40538_ );
and  ( new_n40542_, new_n40541_, new_n40537_ );
or   ( new_n40543_, new_n40542_, new_n40532_ );
and  ( new_n40544_, new_n40542_, new_n40532_ );
or   ( new_n40545_, new_n10059_, new_n26196_ );
or   ( new_n40546_, new_n10061_, new_n25813_ );
and  ( new_n40547_, new_n40546_, new_n40545_ );
xor  ( new_n40548_, new_n40547_, new_n9421_ );
and  ( new_n40549_, RIbb327c0_167, RIbb2d888_64 );
or   ( new_n40550_, new_n25486_, RIbb2d888_64 );
and  ( new_n40551_, new_n40550_, RIbb2d900_63 );
or   ( new_n40552_, new_n40551_, new_n40549_ );
or   ( new_n40553_, new_n10770_, new_n25288_ );
and  ( new_n40554_, new_n40553_, new_n40552_ );
or   ( new_n40555_, new_n40554_, new_n40548_ );
and  ( new_n40556_, new_n40554_, new_n40548_ );
or   ( new_n40557_, new_n9422_, new_n26372_ );
or   ( new_n40558_, new_n9424_, new_n26063_ );
and  ( new_n40559_, new_n40558_, new_n40557_ );
xor  ( new_n40560_, new_n40559_, new_n8873_ );
or   ( new_n40561_, new_n40560_, new_n40556_ );
and  ( new_n40562_, new_n40561_, new_n40555_ );
or   ( new_n40563_, new_n8874_, new_n26762_ );
or   ( new_n40564_, new_n8876_, new_n26620_ );
and  ( new_n40565_, new_n40564_, new_n40563_ );
xor  ( new_n40566_, new_n40565_, new_n8257_ );
or   ( new_n40567_, new_n8264_, new_n27396_ );
or   ( new_n40568_, new_n8266_, new_n27085_ );
and  ( new_n40569_, new_n40568_, new_n40567_ );
xor  ( new_n40570_, new_n40569_, new_n7725_ );
or   ( new_n40571_, new_n40570_, new_n40566_ );
and  ( new_n40572_, new_n40570_, new_n40566_ );
or   ( new_n40573_, new_n7732_, new_n27763_ );
or   ( new_n40574_, new_n7734_, new_n27602_ );
and  ( new_n40575_, new_n40574_, new_n40573_ );
xor  ( new_n40576_, new_n40575_, new_n7177_ );
or   ( new_n40577_, new_n40576_, new_n40572_ );
and  ( new_n40578_, new_n40577_, new_n40571_ );
or   ( new_n40579_, new_n40578_, new_n40562_ );
and  ( new_n40580_, new_n40578_, new_n40562_ );
or   ( new_n40581_, new_n7184_, new_n28314_ );
or   ( new_n40582_, new_n7186_, new_n28108_ );
and  ( new_n40583_, new_n40582_, new_n40581_ );
xor  ( new_n40584_, new_n40583_, new_n6638_ );
or   ( new_n40585_, new_n6645_, new_n29263_ );
or   ( new_n40586_, new_n6647_, new_n28531_ );
and  ( new_n40587_, new_n40586_, new_n40585_ );
xor  ( new_n40588_, new_n40587_, new_n6166_ );
or   ( new_n40589_, new_n40588_, new_n40584_ );
and  ( new_n40590_, new_n40588_, new_n40584_ );
or   ( new_n40591_, new_n6173_, new_n29474_ );
or   ( new_n40592_, new_n6175_, new_n29261_ );
and  ( new_n40593_, new_n40592_, new_n40591_ );
xor  ( new_n40594_, new_n40593_, new_n5597_ );
or   ( new_n40595_, new_n40594_, new_n40590_ );
and  ( new_n40596_, new_n40595_, new_n40589_ );
or   ( new_n40597_, new_n40596_, new_n40580_ );
and  ( new_n40598_, new_n40597_, new_n40579_ );
xnor ( new_n40599_, new_n40427_, new_n40423_ );
xor  ( new_n40600_, new_n40599_, new_n40433_ );
or   ( new_n40601_, new_n5604_, new_n30120_ );
or   ( new_n40602_, new_n5606_, new_n29619_ );
and  ( new_n40603_, new_n40602_, new_n40601_ );
xor  ( new_n40604_, new_n40603_, new_n5206_ );
or   ( new_n40605_, new_n5207_, new_n30800_ );
or   ( new_n40606_, new_n5209_, new_n30227_ );
and  ( new_n40607_, new_n40606_, new_n40605_ );
xor  ( new_n40608_, new_n40607_, new_n4708_ );
or   ( new_n40609_, new_n40608_, new_n40604_ );
and  ( new_n40610_, new_n40608_, new_n40604_ );
or   ( new_n40611_, new_n4709_, new_n31333_ );
or   ( new_n40612_, new_n4711_, new_n30798_ );
and  ( new_n40613_, new_n40612_, new_n40611_ );
xor  ( new_n40614_, new_n40613_, new_n4295_ );
or   ( new_n40615_, new_n40614_, new_n40610_ );
and  ( new_n40616_, new_n40615_, new_n40609_ );
or   ( new_n40617_, new_n40616_, new_n40600_ );
nand ( new_n40618_, new_n40616_, new_n40600_ );
xor  ( new_n40619_, new_n40409_, new_n40405_ );
xnor ( new_n40620_, new_n40619_, new_n40415_ );
nand ( new_n40621_, new_n40620_, new_n40618_ );
and  ( new_n40622_, new_n40621_, new_n40617_ );
and  ( new_n40623_, new_n40622_, new_n40598_ );
nor  ( new_n40624_, new_n40622_, new_n40598_ );
xnor ( new_n40625_, new_n40445_, new_n40441_ );
xor  ( new_n40626_, new_n40625_, new_n40451_ );
xor  ( new_n40627_, new_n40463_, new_n40457_ );
xor  ( new_n40628_, new_n40627_, new_n3460_ );
nor  ( new_n40629_, new_n40628_, new_n40626_ );
and  ( new_n40630_, new_n40628_, new_n40626_ );
xor  ( new_n40631_, new_n40475_, new_n40471_ );
xnor ( new_n40632_, new_n40631_, new_n40481_ );
nor  ( new_n40633_, new_n40632_, new_n40630_ );
nor  ( new_n40634_, new_n40633_, new_n40629_ );
nor  ( new_n40635_, new_n40634_, new_n40624_ );
nor  ( new_n40636_, new_n40635_, new_n40623_ );
or   ( new_n40637_, new_n40636_, new_n40544_ );
and  ( new_n40638_, new_n40637_, new_n40543_ );
xnor ( new_n40639_, new_n40513_, new_n40503_ );
xor  ( new_n40640_, new_n40639_, new_n40517_ );
or   ( new_n40641_, new_n40640_, new_n40638_ );
and  ( new_n40642_, new_n40640_, new_n40638_ );
xnor ( new_n40643_, new_n40392_, new_n40390_ );
or   ( new_n40644_, new_n40643_, new_n40642_ );
and  ( new_n40645_, new_n40644_, new_n40641_ );
xnor ( new_n40646_, new_n40395_, new_n40393_ );
xor  ( new_n40647_, new_n40646_, new_n40519_ );
or   ( new_n40648_, new_n40647_, new_n40645_ );
and  ( new_n40649_, new_n40647_, new_n40645_ );
xnor ( new_n40650_, new_n40387_, new_n40385_ );
or   ( new_n40651_, new_n40650_, new_n40649_ );
and  ( new_n40652_, new_n40651_, new_n40648_ );
nor  ( new_n40653_, new_n40652_, new_n40530_ );
xor  ( new_n40654_, new_n40647_, new_n40645_ );
xor  ( new_n40655_, new_n40654_, new_n40650_ );
xor  ( new_n40656_, new_n40542_, new_n40532_ );
xnor ( new_n40657_, new_n40656_, new_n40636_ );
not  ( new_n40658_, new_n40657_ );
xor  ( new_n40659_, new_n40487_, new_n40437_ );
xor  ( new_n40660_, new_n40659_, new_n40501_ );
or   ( new_n40661_, new_n40660_, new_n40658_ );
xor  ( new_n40662_, new_n40483_, new_n40467_ );
xor  ( new_n40663_, new_n40662_, new_n40453_ );
xnor ( new_n40664_, new_n40622_, new_n40598_ );
xor  ( new_n40665_, new_n40664_, new_n40634_ );
or   ( new_n40666_, new_n40665_, new_n40663_ );
and  ( new_n40667_, new_n40665_, new_n40663_ );
xor  ( new_n40668_, new_n40536_, new_n40534_ );
xnor ( new_n40669_, new_n40668_, new_n40540_ );
or   ( new_n40670_, new_n40669_, new_n40667_ );
and  ( new_n40671_, new_n40670_, new_n40666_ );
xnor ( new_n40672_, new_n40507_, new_n40505_ );
xor  ( new_n40673_, new_n40672_, new_n40511_ );
nand ( new_n40674_, new_n40673_, new_n40671_ );
nor  ( new_n40675_, new_n40673_, new_n40671_ );
xor  ( new_n40676_, new_n40417_, new_n40401_ );
xor  ( new_n40677_, new_n40676_, new_n40435_ );
or   ( new_n40678_, new_n4709_, new_n31654_ );
or   ( new_n40679_, new_n4711_, new_n31333_ );
and  ( new_n40680_, new_n40679_, new_n40678_ );
xor  ( new_n40681_, new_n40680_, new_n4295_ );
not  ( new_n40682_, new_n40681_ );
and  ( new_n40683_, new_n4032_, RIbb33378_192 );
or   ( new_n40684_, new_n40683_, new_n3895_ );
nand ( new_n40685_, new_n40683_, new_n3892_ );
and  ( new_n40686_, new_n40685_, new_n40684_ );
nor  ( new_n40687_, new_n40686_, new_n40682_ );
or   ( new_n40688_, new_n4302_, new_n31952_ );
or   ( new_n40689_, new_n4304_, new_n31654_ );
and  ( new_n40690_, new_n40689_, new_n40688_ );
xor  ( new_n40691_, new_n40690_, new_n3895_ );
or   ( new_n40692_, new_n40691_, new_n40687_ );
and  ( new_n40693_, new_n40691_, new_n40687_ );
or   ( new_n40694_, new_n6173_, new_n29619_ );
or   ( new_n40695_, new_n6175_, new_n29474_ );
and  ( new_n40696_, new_n40695_, new_n40694_ );
xor  ( new_n40697_, new_n40696_, new_n5597_ );
or   ( new_n40698_, new_n5604_, new_n30227_ );
or   ( new_n40699_, new_n5606_, new_n30120_ );
and  ( new_n40700_, new_n40699_, new_n40698_ );
xor  ( new_n40701_, new_n40700_, new_n5206_ );
nor  ( new_n40702_, new_n40701_, new_n40697_ );
and  ( new_n40703_, new_n40701_, new_n40697_ );
or   ( new_n40704_, new_n5207_, new_n30798_ );
or   ( new_n40705_, new_n5209_, new_n30800_ );
and  ( new_n40706_, new_n40705_, new_n40704_ );
xor  ( new_n40707_, new_n40706_, new_n4708_ );
nor  ( new_n40708_, new_n40707_, new_n40703_ );
nor  ( new_n40709_, new_n40708_, new_n40702_ );
or   ( new_n40710_, new_n40709_, new_n40693_ );
and  ( new_n40711_, new_n40710_, new_n40692_ );
or   ( new_n40712_, new_n9422_, new_n26620_ );
or   ( new_n40713_, new_n9424_, new_n26372_ );
and  ( new_n40714_, new_n40713_, new_n40712_ );
xor  ( new_n40715_, new_n40714_, new_n8873_ );
or   ( new_n40716_, new_n8874_, new_n27085_ );
or   ( new_n40717_, new_n8876_, new_n26762_ );
and  ( new_n40718_, new_n40717_, new_n40716_ );
xor  ( new_n40719_, new_n40718_, new_n8257_ );
or   ( new_n40720_, new_n40719_, new_n40715_ );
and  ( new_n40721_, new_n40719_, new_n40715_ );
or   ( new_n40722_, new_n8264_, new_n27602_ );
or   ( new_n40723_, new_n8266_, new_n27396_ );
and  ( new_n40724_, new_n40723_, new_n40722_ );
xor  ( new_n40725_, new_n40724_, new_n7725_ );
or   ( new_n40726_, new_n40725_, new_n40721_ );
and  ( new_n40727_, new_n40726_, new_n40720_ );
or   ( new_n40728_, new_n10059_, new_n26063_ );
or   ( new_n40729_, new_n10061_, new_n26196_ );
and  ( new_n40730_, new_n40729_, new_n40728_ );
xor  ( new_n40731_, new_n40730_, new_n9421_ );
and  ( new_n40732_, RIbb32838_168, RIbb2d888_64 );
or   ( new_n40733_, new_n25813_, RIbb2d888_64 );
and  ( new_n40734_, new_n40733_, RIbb2d900_63 );
or   ( new_n40735_, new_n40734_, new_n40732_ );
or   ( new_n40736_, new_n10770_, new_n25486_ );
and  ( new_n40737_, new_n40736_, new_n40735_ );
nor  ( new_n40738_, new_n40737_, new_n40731_ );
and  ( new_n40739_, new_n40737_, new_n40731_ );
nor  ( new_n40740_, new_n40739_, new_n3894_ );
nor  ( new_n40741_, new_n40740_, new_n40738_ );
or   ( new_n40742_, new_n7732_, new_n28108_ );
or   ( new_n40743_, new_n7734_, new_n27763_ );
and  ( new_n40744_, new_n40743_, new_n40742_ );
xor  ( new_n40745_, new_n40744_, new_n7177_ );
or   ( new_n40746_, new_n7184_, new_n28531_ );
or   ( new_n40747_, new_n7186_, new_n28314_ );
and  ( new_n40748_, new_n40747_, new_n40746_ );
xor  ( new_n40749_, new_n40748_, new_n6638_ );
or   ( new_n40750_, new_n40749_, new_n40745_ );
and  ( new_n40751_, new_n40749_, new_n40745_ );
or   ( new_n40752_, new_n6645_, new_n29261_ );
or   ( new_n40753_, new_n6647_, new_n29263_ );
and  ( new_n40754_, new_n40753_, new_n40752_ );
xor  ( new_n40755_, new_n40754_, new_n6166_ );
or   ( new_n40756_, new_n40755_, new_n40751_ );
and  ( new_n40757_, new_n40756_, new_n40750_ );
and  ( new_n40758_, new_n40757_, new_n40741_ );
or   ( new_n40759_, new_n40758_, new_n40727_ );
or   ( new_n40760_, new_n40757_, new_n40741_ );
and  ( new_n40761_, new_n40760_, new_n40759_ );
nand ( new_n40762_, new_n40761_, new_n40711_ );
nor  ( new_n40763_, new_n40761_, new_n40711_ );
xnor ( new_n40764_, new_n40570_, new_n40566_ );
xor  ( new_n40765_, new_n40764_, new_n40576_ );
xnor ( new_n40766_, new_n40608_, new_n40604_ );
xor  ( new_n40767_, new_n40766_, new_n40614_ );
nor  ( new_n40768_, new_n40767_, new_n40765_ );
and  ( new_n40769_, new_n40767_, new_n40765_ );
xor  ( new_n40770_, new_n40588_, new_n40584_ );
xnor ( new_n40771_, new_n40770_, new_n40594_ );
nor  ( new_n40772_, new_n40771_, new_n40769_ );
nor  ( new_n40773_, new_n40772_, new_n40768_ );
or   ( new_n40774_, new_n40773_, new_n40763_ );
and  ( new_n40775_, new_n40774_, new_n40762_ );
or   ( new_n40776_, new_n40775_, new_n40677_ );
and  ( new_n40777_, new_n40775_, new_n40677_ );
xor  ( new_n40778_, new_n40578_, new_n40562_ );
xor  ( new_n40779_, new_n40778_, new_n40596_ );
xnor ( new_n40780_, new_n40628_, new_n40626_ );
xor  ( new_n40781_, new_n40780_, new_n40632_ );
and  ( new_n40782_, new_n40781_, new_n40779_ );
nor  ( new_n40783_, new_n40781_, new_n40779_ );
xor  ( new_n40784_, new_n40616_, new_n40600_ );
xor  ( new_n40785_, new_n40784_, new_n40620_ );
nor  ( new_n40786_, new_n40785_, new_n40783_ );
nor  ( new_n40787_, new_n40786_, new_n40782_ );
or   ( new_n40788_, new_n40787_, new_n40777_ );
and  ( new_n40789_, new_n40788_, new_n40776_ );
or   ( new_n40790_, new_n40789_, new_n40675_ );
and  ( new_n40791_, new_n40790_, new_n40674_ );
or   ( new_n40792_, new_n40791_, new_n40661_ );
and  ( new_n40793_, new_n40791_, new_n40661_ );
xor  ( new_n40794_, new_n40640_, new_n40638_ );
xor  ( new_n40795_, new_n40794_, new_n40643_ );
or   ( new_n40796_, new_n40795_, new_n40793_ );
and  ( new_n40797_, new_n40796_, new_n40792_ );
nor  ( new_n40798_, new_n40797_, new_n40655_ );
xor  ( new_n40799_, new_n40791_, new_n40661_ );
xor  ( new_n40800_, new_n40799_, new_n40795_ );
xor  ( new_n40801_, new_n40673_, new_n40671_ );
xor  ( new_n40802_, new_n40801_, new_n40789_ );
xor  ( new_n40803_, new_n40781_, new_n40779_ );
xor  ( new_n40804_, new_n40803_, new_n40785_ );
xor  ( new_n40805_, new_n40767_, new_n40765_ );
xor  ( new_n40806_, new_n40805_, new_n40771_ );
xnor ( new_n40807_, new_n40691_, new_n40687_ );
xor  ( new_n40808_, new_n40807_, new_n40709_ );
or   ( new_n40809_, new_n40808_, new_n40806_ );
and  ( new_n40810_, new_n40808_, new_n40806_ );
xor  ( new_n40811_, new_n40554_, new_n40548_ );
xnor ( new_n40812_, new_n40811_, new_n40560_ );
or   ( new_n40813_, new_n40812_, new_n40810_ );
and  ( new_n40814_, new_n40813_, new_n40809_ );
nor  ( new_n40815_, new_n40814_, new_n40804_ );
nand ( new_n40816_, new_n40814_, new_n40804_ );
or   ( new_n40817_, new_n7184_, new_n29263_ );
or   ( new_n40818_, new_n7186_, new_n28531_ );
and  ( new_n40819_, new_n40818_, new_n40817_ );
xor  ( new_n40820_, new_n40819_, new_n6638_ );
or   ( new_n40821_, new_n6645_, new_n29474_ );
or   ( new_n40822_, new_n6647_, new_n29261_ );
and  ( new_n40823_, new_n40822_, new_n40821_ );
xor  ( new_n40824_, new_n40823_, new_n6166_ );
or   ( new_n40825_, new_n40824_, new_n40820_ );
and  ( new_n40826_, new_n40824_, new_n40820_ );
or   ( new_n40827_, new_n6173_, new_n30120_ );
or   ( new_n40828_, new_n6175_, new_n29619_ );
and  ( new_n40829_, new_n40828_, new_n40827_ );
xor  ( new_n40830_, new_n40829_, new_n5597_ );
or   ( new_n40831_, new_n40830_, new_n40826_ );
and  ( new_n40832_, new_n40831_, new_n40825_ );
or   ( new_n40833_, new_n8874_, new_n27396_ );
or   ( new_n40834_, new_n8876_, new_n27085_ );
and  ( new_n40835_, new_n40834_, new_n40833_ );
xor  ( new_n40836_, new_n40835_, new_n8257_ );
or   ( new_n40837_, new_n8264_, new_n27763_ );
or   ( new_n40838_, new_n8266_, new_n27602_ );
and  ( new_n40839_, new_n40838_, new_n40837_ );
xor  ( new_n40840_, new_n40839_, new_n7725_ );
or   ( new_n40841_, new_n40840_, new_n40836_ );
and  ( new_n40842_, new_n40840_, new_n40836_ );
or   ( new_n40843_, new_n7732_, new_n28314_ );
or   ( new_n40844_, new_n7734_, new_n28108_ );
and  ( new_n40845_, new_n40844_, new_n40843_ );
xor  ( new_n40846_, new_n40845_, new_n7177_ );
or   ( new_n40847_, new_n40846_, new_n40842_ );
and  ( new_n40848_, new_n40847_, new_n40841_ );
or   ( new_n40849_, new_n40848_, new_n40832_ );
and  ( new_n40850_, new_n40848_, new_n40832_ );
or   ( new_n40851_, new_n10059_, new_n26372_ );
or   ( new_n40852_, new_n10061_, new_n26063_ );
and  ( new_n40853_, new_n40852_, new_n40851_ );
xor  ( new_n40854_, new_n40853_, new_n9421_ );
and  ( new_n40855_, RIbb328b0_169, RIbb2d888_64 );
or   ( new_n40856_, new_n26196_, RIbb2d888_64 );
and  ( new_n40857_, new_n40856_, RIbb2d900_63 );
or   ( new_n40858_, new_n40857_, new_n40855_ );
or   ( new_n40859_, new_n10770_, new_n25813_ );
and  ( new_n40860_, new_n40859_, new_n40858_ );
or   ( new_n40861_, new_n40860_, new_n40854_ );
and  ( new_n40862_, new_n40860_, new_n40854_ );
or   ( new_n40863_, new_n9422_, new_n26762_ );
or   ( new_n40864_, new_n9424_, new_n26620_ );
and  ( new_n40865_, new_n40864_, new_n40863_ );
xor  ( new_n40866_, new_n40865_, new_n8873_ );
or   ( new_n40867_, new_n40866_, new_n40862_ );
and  ( new_n40868_, new_n40867_, new_n40861_ );
or   ( new_n40869_, new_n40868_, new_n40850_ );
and  ( new_n40870_, new_n40869_, new_n40849_ );
xor  ( new_n40871_, new_n40701_, new_n40697_ );
xor  ( new_n40872_, new_n40871_, new_n40707_ );
or   ( new_n40873_, new_n5604_, new_n30800_ );
or   ( new_n40874_, new_n5606_, new_n30227_ );
and  ( new_n40875_, new_n40874_, new_n40873_ );
xor  ( new_n40876_, new_n40875_, new_n5206_ );
or   ( new_n40877_, new_n5207_, new_n31333_ );
or   ( new_n40878_, new_n5209_, new_n30798_ );
and  ( new_n40879_, new_n40878_, new_n40877_ );
xor  ( new_n40880_, new_n40879_, new_n4708_ );
or   ( new_n40881_, new_n40880_, new_n40876_ );
and  ( new_n40882_, new_n40880_, new_n40876_ );
or   ( new_n40883_, new_n4709_, new_n31952_ );
or   ( new_n40884_, new_n4711_, new_n31654_ );
and  ( new_n40885_, new_n40884_, new_n40883_ );
xor  ( new_n40886_, new_n40885_, new_n4295_ );
or   ( new_n40887_, new_n40886_, new_n40882_ );
and  ( new_n40888_, new_n40887_, new_n40881_ );
or   ( new_n40889_, new_n40888_, new_n40872_ );
and  ( new_n40890_, new_n40888_, new_n40872_ );
xor  ( new_n40891_, new_n40686_, new_n40682_ );
or   ( new_n40892_, new_n40891_, new_n40890_ );
and  ( new_n40893_, new_n40892_, new_n40889_ );
and  ( new_n40894_, new_n40893_, new_n40870_ );
or   ( new_n40895_, new_n40893_, new_n40870_ );
xnor ( new_n40896_, new_n40719_, new_n40715_ );
xor  ( new_n40897_, new_n40896_, new_n40725_ );
xor  ( new_n40898_, new_n40737_, new_n40731_ );
xor  ( new_n40899_, new_n40898_, new_n3895_ );
nor  ( new_n40900_, new_n40899_, new_n40897_ );
and  ( new_n40901_, new_n40899_, new_n40897_ );
xor  ( new_n40902_, new_n40749_, new_n40745_ );
xnor ( new_n40903_, new_n40902_, new_n40755_ );
nor  ( new_n40904_, new_n40903_, new_n40901_ );
nor  ( new_n40905_, new_n40904_, new_n40900_ );
not  ( new_n40906_, new_n40905_ );
and  ( new_n40907_, new_n40906_, new_n40895_ );
or   ( new_n40908_, new_n40907_, new_n40894_ );
and  ( new_n40909_, new_n40908_, new_n40816_ );
or   ( new_n40910_, new_n40909_, new_n40815_ );
xnor ( new_n40911_, new_n40775_, new_n40677_ );
xor  ( new_n40912_, new_n40911_, new_n40787_ );
nand ( new_n40913_, new_n40912_, new_n40910_ );
nor  ( new_n40914_, new_n40912_, new_n40910_ );
xor  ( new_n40915_, new_n40665_, new_n40663_ );
xnor ( new_n40916_, new_n40915_, new_n40669_ );
or   ( new_n40917_, new_n40916_, new_n40914_ );
and  ( new_n40918_, new_n40917_, new_n40913_ );
or   ( new_n40919_, new_n40918_, new_n40802_ );
nand ( new_n40920_, new_n40918_, new_n40802_ );
xor  ( new_n40921_, new_n40660_, new_n40658_ );
nand ( new_n40922_, new_n40921_, new_n40920_ );
and  ( new_n40923_, new_n40922_, new_n40919_ );
nor  ( new_n40924_, new_n40923_, new_n40800_ );
xor  ( new_n40925_, new_n40893_, new_n40870_ );
xor  ( new_n40926_, new_n40925_, new_n40906_ );
xnor ( new_n40927_, new_n40808_, new_n40806_ );
xor  ( new_n40928_, new_n40927_, new_n40812_ );
nand ( new_n40929_, new_n40928_, new_n40926_ );
xnor ( new_n40930_, new_n40757_, new_n40741_ );
xor  ( new_n40931_, new_n40930_, new_n40727_ );
xor  ( new_n40932_, new_n40848_, new_n40832_ );
xor  ( new_n40933_, new_n40932_, new_n40868_ );
xnor ( new_n40934_, new_n40899_, new_n40897_ );
xor  ( new_n40935_, new_n40934_, new_n40903_ );
nand ( new_n40936_, new_n40935_, new_n40933_ );
nor  ( new_n40937_, new_n40935_, new_n40933_ );
xnor ( new_n40938_, new_n40888_, new_n40872_ );
xor  ( new_n40939_, new_n40938_, new_n40891_ );
or   ( new_n40940_, new_n40939_, new_n40937_ );
and  ( new_n40941_, new_n40940_, new_n40936_ );
or   ( new_n40942_, new_n40941_, new_n40931_ );
nand ( new_n40943_, new_n40941_, new_n40931_ );
xor  ( new_n40944_, new_n40840_, new_n40836_ );
xnor ( new_n40945_, new_n40944_, new_n40846_ );
xnor ( new_n40946_, new_n40860_, new_n40854_ );
xor  ( new_n40947_, new_n40946_, new_n40866_ );
nor  ( new_n40948_, new_n40947_, new_n40945_ );
or   ( new_n40949_, new_n9422_, new_n27085_ );
or   ( new_n40950_, new_n9424_, new_n26762_ );
and  ( new_n40951_, new_n40950_, new_n40949_ );
xor  ( new_n40952_, new_n40951_, new_n8873_ );
or   ( new_n40953_, new_n8874_, new_n27602_ );
or   ( new_n40954_, new_n8876_, new_n27396_ );
and  ( new_n40955_, new_n40954_, new_n40953_ );
xor  ( new_n40956_, new_n40955_, new_n8257_ );
or   ( new_n40957_, new_n40956_, new_n40952_ );
and  ( new_n40958_, new_n40956_, new_n40952_ );
or   ( new_n40959_, new_n8264_, new_n28108_ );
or   ( new_n40960_, new_n8266_, new_n27763_ );
and  ( new_n40961_, new_n40960_, new_n40959_ );
xor  ( new_n40962_, new_n40961_, new_n7725_ );
or   ( new_n40963_, new_n40962_, new_n40958_ );
and  ( new_n40964_, new_n40963_, new_n40957_ );
or   ( new_n40965_, new_n10059_, new_n26620_ );
or   ( new_n40966_, new_n10061_, new_n26372_ );
and  ( new_n40967_, new_n40966_, new_n40965_ );
xor  ( new_n40968_, new_n40967_, new_n9421_ );
and  ( new_n40969_, RIbb32928_170, RIbb2d888_64 );
or   ( new_n40970_, new_n26063_, RIbb2d888_64 );
and  ( new_n40971_, new_n40970_, RIbb2d900_63 );
or   ( new_n40972_, new_n40971_, new_n40969_ );
or   ( new_n40973_, new_n10770_, new_n26196_ );
and  ( new_n40974_, new_n40973_, new_n40972_ );
nor  ( new_n40975_, new_n40974_, new_n40968_ );
and  ( new_n40976_, new_n40974_, new_n40968_ );
nor  ( new_n40977_, new_n40976_, new_n4294_ );
nor  ( new_n40978_, new_n40977_, new_n40975_ );
or   ( new_n40979_, new_n7732_, new_n28531_ );
or   ( new_n40980_, new_n7734_, new_n28314_ );
and  ( new_n40981_, new_n40980_, new_n40979_ );
xor  ( new_n40982_, new_n40981_, new_n7177_ );
or   ( new_n40983_, new_n7184_, new_n29261_ );
or   ( new_n40984_, new_n7186_, new_n29263_ );
and  ( new_n40985_, new_n40984_, new_n40983_ );
xor  ( new_n40986_, new_n40985_, new_n6638_ );
or   ( new_n40987_, new_n40986_, new_n40982_ );
and  ( new_n40988_, new_n40986_, new_n40982_ );
or   ( new_n40989_, new_n6645_, new_n29619_ );
or   ( new_n40990_, new_n6647_, new_n29474_ );
and  ( new_n40991_, new_n40990_, new_n40989_ );
xor  ( new_n40992_, new_n40991_, new_n6166_ );
or   ( new_n40993_, new_n40992_, new_n40988_ );
and  ( new_n40994_, new_n40993_, new_n40987_ );
and  ( new_n40995_, new_n40994_, new_n40978_ );
or   ( new_n40996_, new_n40995_, new_n40964_ );
or   ( new_n40997_, new_n40994_, new_n40978_ );
and  ( new_n40998_, new_n40997_, new_n40996_ );
nor  ( new_n40999_, new_n40998_, new_n40948_ );
and  ( new_n41000_, new_n40998_, new_n40948_ );
xor  ( new_n41001_, new_n40880_, new_n40876_ );
xor  ( new_n41002_, new_n41001_, new_n40886_ );
or   ( new_n41003_, new_n6173_, new_n30227_ );
or   ( new_n41004_, new_n6175_, new_n30120_ );
and  ( new_n41005_, new_n41004_, new_n41003_ );
xor  ( new_n41006_, new_n41005_, new_n5597_ );
or   ( new_n41007_, new_n5604_, new_n30798_ );
or   ( new_n41008_, new_n5606_, new_n30800_ );
and  ( new_n41009_, new_n41008_, new_n41007_ );
xor  ( new_n41010_, new_n41009_, new_n5206_ );
or   ( new_n41011_, new_n41010_, new_n41006_ );
and  ( new_n41012_, new_n41010_, new_n41006_ );
or   ( new_n41013_, new_n5207_, new_n31654_ );
or   ( new_n41014_, new_n5209_, new_n31333_ );
and  ( new_n41015_, new_n41014_, new_n41013_ );
xor  ( new_n41016_, new_n41015_, new_n4708_ );
or   ( new_n41017_, new_n41016_, new_n41012_ );
and  ( new_n41018_, new_n41017_, new_n41011_ );
nor  ( new_n41019_, new_n41018_, new_n41002_ );
and  ( new_n41020_, new_n41018_, new_n41002_ );
not  ( new_n41021_, new_n41020_ );
xor  ( new_n41022_, new_n40824_, new_n40820_ );
xnor ( new_n41023_, new_n41022_, new_n40830_ );
and  ( new_n41024_, new_n41023_, new_n41021_ );
nor  ( new_n41025_, new_n41024_, new_n41019_ );
nor  ( new_n41026_, new_n41025_, new_n41000_ );
nor  ( new_n41027_, new_n41026_, new_n40999_ );
nand ( new_n41028_, new_n41027_, new_n40943_ );
and  ( new_n41029_, new_n41028_, new_n40942_ );
nor  ( new_n41030_, new_n41029_, new_n40929_ );
nand ( new_n41031_, new_n41029_, new_n40929_ );
xor  ( new_n41032_, new_n40761_, new_n40711_ );
xnor ( new_n41033_, new_n41032_, new_n40773_ );
and  ( new_n41034_, new_n41033_, new_n41031_ );
or   ( new_n41035_, new_n41034_, new_n41030_ );
xnor ( new_n41036_, new_n40912_, new_n40910_ );
xor  ( new_n41037_, new_n41036_, new_n40916_ );
and  ( new_n41038_, new_n41037_, new_n41035_ );
xor  ( new_n41039_, new_n40918_, new_n40802_ );
xor  ( new_n41040_, new_n41039_, new_n40921_ );
and  ( new_n41041_, new_n41040_, new_n41038_ );
xor  ( new_n41042_, new_n41029_, new_n40929_ );
xnor ( new_n41043_, new_n41042_, new_n41033_ );
xor  ( new_n41044_, new_n40814_, new_n40804_ );
xnor ( new_n41045_, new_n41044_, new_n40908_ );
nor  ( new_n41046_, new_n41045_, new_n41043_ );
xor  ( new_n41047_, new_n41037_, new_n41035_ );
and  ( new_n41048_, new_n41047_, new_n41046_ );
xnor ( new_n41049_, new_n41045_, new_n41043_ );
xor  ( new_n41050_, new_n40935_, new_n40933_ );
xor  ( new_n41051_, new_n41050_, new_n40939_ );
xnor ( new_n41052_, new_n40994_, new_n40978_ );
xor  ( new_n41053_, new_n41052_, new_n40964_ );
xor  ( new_n41054_, new_n41018_, new_n41002_ );
xor  ( new_n41055_, new_n41054_, new_n41023_ );
or   ( new_n41056_, new_n41055_, new_n41053_ );
and  ( new_n41057_, new_n41055_, new_n41053_ );
xnor ( new_n41058_, new_n40947_, new_n40945_ );
or   ( new_n41059_, new_n41058_, new_n41057_ );
and  ( new_n41060_, new_n41059_, new_n41056_ );
nor  ( new_n41061_, new_n41060_, new_n41051_ );
and  ( new_n41062_, new_n41060_, new_n41051_ );
xor  ( new_n41063_, new_n40956_, new_n40952_ );
xnor ( new_n41064_, new_n41063_, new_n40962_ );
xor  ( new_n41065_, new_n40974_, new_n40968_ );
xor  ( new_n41066_, new_n41065_, new_n4295_ );
nor  ( new_n41067_, new_n41066_, new_n41064_ );
or   ( new_n41068_, new_n7184_, new_n29474_ );
or   ( new_n41069_, new_n7186_, new_n29261_ );
and  ( new_n41070_, new_n41069_, new_n41068_ );
xor  ( new_n41071_, new_n41070_, new_n6638_ );
or   ( new_n41072_, new_n6645_, new_n30120_ );
or   ( new_n41073_, new_n6647_, new_n29619_ );
and  ( new_n41074_, new_n41073_, new_n41072_ );
xor  ( new_n41075_, new_n41074_, new_n6166_ );
or   ( new_n41076_, new_n41075_, new_n41071_ );
and  ( new_n41077_, new_n41075_, new_n41071_ );
or   ( new_n41078_, new_n6173_, new_n30800_ );
or   ( new_n41079_, new_n6175_, new_n30227_ );
and  ( new_n41080_, new_n41079_, new_n41078_ );
xor  ( new_n41081_, new_n41080_, new_n5597_ );
or   ( new_n41082_, new_n41081_, new_n41077_ );
and  ( new_n41083_, new_n41082_, new_n41076_ );
or   ( new_n41084_, new_n10059_, new_n26762_ );
or   ( new_n41085_, new_n10061_, new_n26620_ );
and  ( new_n41086_, new_n41085_, new_n41084_ );
xor  ( new_n41087_, new_n41086_, new_n9421_ );
and  ( new_n41088_, RIbb329a0_171, RIbb2d888_64 );
or   ( new_n41089_, new_n26372_, RIbb2d888_64 );
and  ( new_n41090_, new_n41089_, RIbb2d900_63 );
or   ( new_n41091_, new_n41090_, new_n41088_ );
or   ( new_n41092_, new_n10770_, new_n26063_ );
and  ( new_n41093_, new_n41092_, new_n41091_ );
or   ( new_n41094_, new_n41093_, new_n41087_ );
and  ( new_n41095_, new_n41093_, new_n41087_ );
or   ( new_n41096_, new_n9422_, new_n27396_ );
or   ( new_n41097_, new_n9424_, new_n27085_ );
and  ( new_n41098_, new_n41097_, new_n41096_ );
xor  ( new_n41099_, new_n41098_, new_n8873_ );
or   ( new_n41100_, new_n41099_, new_n41095_ );
and  ( new_n41101_, new_n41100_, new_n41094_ );
or   ( new_n41102_, new_n41101_, new_n41083_ );
and  ( new_n41103_, new_n41101_, new_n41083_ );
or   ( new_n41104_, new_n8874_, new_n27763_ );
or   ( new_n41105_, new_n8876_, new_n27602_ );
and  ( new_n41106_, new_n41105_, new_n41104_ );
xor  ( new_n41107_, new_n41106_, new_n8257_ );
or   ( new_n41108_, new_n8264_, new_n28314_ );
or   ( new_n41109_, new_n8266_, new_n28108_ );
and  ( new_n41110_, new_n41109_, new_n41108_ );
xor  ( new_n41111_, new_n41110_, new_n7725_ );
or   ( new_n41112_, new_n41111_, new_n41107_ );
and  ( new_n41113_, new_n41111_, new_n41107_ );
or   ( new_n41114_, new_n7732_, new_n29263_ );
or   ( new_n41115_, new_n7734_, new_n28531_ );
and  ( new_n41116_, new_n41115_, new_n41114_ );
xor  ( new_n41117_, new_n41116_, new_n7177_ );
or   ( new_n41118_, new_n41117_, new_n41113_ );
and  ( new_n41119_, new_n41118_, new_n41112_ );
or   ( new_n41120_, new_n41119_, new_n41103_ );
and  ( new_n41121_, new_n41120_, new_n41102_ );
and  ( new_n41122_, new_n41121_, new_n41067_ );
nor  ( new_n41123_, new_n41121_, new_n41067_ );
and  ( new_n41124_, new_n4541_, RIbb33378_192 );
or   ( new_n41125_, new_n41124_, new_n4295_ );
nand ( new_n41126_, new_n41124_, new_n4292_ );
and  ( new_n41127_, new_n41126_, new_n41125_ );
xnor ( new_n41128_, new_n41010_, new_n41006_ );
xor  ( new_n41129_, new_n41128_, new_n41016_ );
nor  ( new_n41130_, new_n41129_, new_n41127_ );
and  ( new_n41131_, new_n41129_, new_n41127_ );
xor  ( new_n41132_, new_n40986_, new_n40982_ );
xnor ( new_n41133_, new_n41132_, new_n40992_ );
nor  ( new_n41134_, new_n41133_, new_n41131_ );
nor  ( new_n41135_, new_n41134_, new_n41130_ );
nor  ( new_n41136_, new_n41135_, new_n41123_ );
nor  ( new_n41137_, new_n41136_, new_n41122_ );
nor  ( new_n41138_, new_n41137_, new_n41062_ );
or   ( new_n41139_, new_n41138_, new_n41061_ );
xor  ( new_n41140_, new_n40941_, new_n40931_ );
xor  ( new_n41141_, new_n41140_, new_n41027_ );
nand ( new_n41142_, new_n41141_, new_n41139_ );
nor  ( new_n41143_, new_n41141_, new_n41139_ );
xnor ( new_n41144_, new_n40928_, new_n40926_ );
or   ( new_n41145_, new_n41144_, new_n41143_ );
and  ( new_n41146_, new_n41145_, new_n41142_ );
nor  ( new_n41147_, new_n41146_, new_n41049_ );
xor  ( new_n41148_, new_n41141_, new_n41139_ );
xor  ( new_n41149_, new_n41148_, new_n41144_ );
xor  ( new_n41150_, new_n41060_, new_n41051_ );
xor  ( new_n41151_, new_n41150_, new_n41137_ );
xnor ( new_n41152_, new_n40998_, new_n40948_ );
xor  ( new_n41153_, new_n41152_, new_n41025_ );
or   ( new_n41154_, new_n41153_, new_n41151_ );
and  ( new_n41155_, new_n41153_, new_n41151_ );
xor  ( new_n41156_, new_n41055_, new_n41053_ );
xor  ( new_n41157_, new_n41156_, new_n41058_ );
xor  ( new_n41158_, new_n41101_, new_n41083_ );
xor  ( new_n41159_, new_n41158_, new_n41119_ );
xnor ( new_n41160_, new_n41129_, new_n41127_ );
xor  ( new_n41161_, new_n41160_, new_n41133_ );
nand ( new_n41162_, new_n41161_, new_n41159_ );
or   ( new_n41163_, new_n41161_, new_n41159_ );
xor  ( new_n41164_, new_n41066_, new_n41064_ );
nand ( new_n41165_, new_n41164_, new_n41163_ );
and  ( new_n41166_, new_n41165_, new_n41162_ );
nor  ( new_n41167_, new_n41166_, new_n41157_ );
and  ( new_n41168_, new_n41166_, new_n41157_ );
or   ( new_n41169_, new_n10059_, new_n27085_ );
or   ( new_n41170_, new_n10061_, new_n26762_ );
and  ( new_n41171_, new_n41170_, new_n41169_ );
xor  ( new_n41172_, new_n41171_, new_n9421_ );
and  ( new_n41173_, RIbb32a18_172, RIbb2d888_64 );
or   ( new_n41174_, new_n26620_, RIbb2d888_64 );
and  ( new_n41175_, new_n41174_, RIbb2d900_63 );
or   ( new_n41176_, new_n41175_, new_n41173_ );
or   ( new_n41177_, new_n10770_, new_n26372_ );
and  ( new_n41178_, new_n41177_, new_n41176_ );
or   ( new_n41179_, new_n41178_, new_n41172_ );
and  ( new_n41180_, new_n41178_, new_n41172_ );
or   ( new_n41181_, new_n41180_, new_n4707_ );
and  ( new_n41182_, new_n41181_, new_n41179_ );
or   ( new_n41183_, new_n9422_, new_n27602_ );
or   ( new_n41184_, new_n9424_, new_n27396_ );
and  ( new_n41185_, new_n41184_, new_n41183_ );
xor  ( new_n41186_, new_n41185_, new_n8873_ );
or   ( new_n41187_, new_n8874_, new_n28108_ );
or   ( new_n41188_, new_n8876_, new_n27763_ );
and  ( new_n41189_, new_n41188_, new_n41187_ );
xor  ( new_n41190_, new_n41189_, new_n8257_ );
or   ( new_n41191_, new_n41190_, new_n41186_ );
and  ( new_n41192_, new_n41190_, new_n41186_ );
or   ( new_n41193_, new_n8264_, new_n28531_ );
or   ( new_n41194_, new_n8266_, new_n28314_ );
and  ( new_n41195_, new_n41194_, new_n41193_ );
xor  ( new_n41196_, new_n41195_, new_n7725_ );
or   ( new_n41197_, new_n41196_, new_n41192_ );
and  ( new_n41198_, new_n41197_, new_n41191_ );
nor  ( new_n41199_, new_n41198_, new_n41182_ );
nand ( new_n41200_, new_n41198_, new_n41182_ );
or   ( new_n41201_, new_n7732_, new_n29261_ );
or   ( new_n41202_, new_n7734_, new_n29263_ );
and  ( new_n41203_, new_n41202_, new_n41201_ );
xor  ( new_n41204_, new_n41203_, new_n7177_ );
or   ( new_n41205_, new_n7184_, new_n29619_ );
or   ( new_n41206_, new_n7186_, new_n29474_ );
and  ( new_n41207_, new_n41206_, new_n41205_ );
xor  ( new_n41208_, new_n41207_, new_n6638_ );
nor  ( new_n41209_, new_n41208_, new_n41204_ );
and  ( new_n41210_, new_n41208_, new_n41204_ );
or   ( new_n41211_, new_n6645_, new_n30227_ );
or   ( new_n41212_, new_n6647_, new_n30120_ );
and  ( new_n41213_, new_n41212_, new_n41211_ );
xor  ( new_n41214_, new_n41213_, new_n6166_ );
nor  ( new_n41215_, new_n41214_, new_n41210_ );
nor  ( new_n41216_, new_n41215_, new_n41209_ );
not  ( new_n41217_, new_n41216_ );
and  ( new_n41218_, new_n41217_, new_n41200_ );
or   ( new_n41219_, new_n41218_, new_n41199_ );
xnor ( new_n41220_, new_n41093_, new_n41087_ );
xor  ( new_n41221_, new_n41220_, new_n41099_ );
xnor ( new_n41222_, new_n41075_, new_n41071_ );
xor  ( new_n41223_, new_n41222_, new_n41081_ );
or   ( new_n41224_, new_n41223_, new_n41221_ );
and  ( new_n41225_, new_n41223_, new_n41221_ );
xor  ( new_n41226_, new_n41111_, new_n41107_ );
xnor ( new_n41227_, new_n41226_, new_n41117_ );
or   ( new_n41228_, new_n41227_, new_n41225_ );
and  ( new_n41229_, new_n41228_, new_n41224_ );
nor  ( new_n41230_, new_n41229_, new_n41219_ );
and  ( new_n41231_, new_n41229_, new_n41219_ );
or   ( new_n41232_, new_n5604_, new_n31333_ );
or   ( new_n41233_, new_n5606_, new_n30798_ );
and  ( new_n41234_, new_n41233_, new_n41232_ );
xor  ( new_n41235_, new_n41234_, new_n5205_ );
or   ( new_n41236_, new_n6173_, new_n30798_ );
or   ( new_n41237_, new_n6175_, new_n30800_ );
and  ( new_n41238_, new_n41237_, new_n41236_ );
xor  ( new_n41239_, new_n41238_, new_n5597_ );
or   ( new_n41240_, new_n5604_, new_n31654_ );
or   ( new_n41241_, new_n5606_, new_n31333_ );
and  ( new_n41242_, new_n41241_, new_n41240_ );
xor  ( new_n41243_, new_n41242_, new_n5206_ );
nand ( new_n41244_, new_n41243_, new_n41239_ );
nor  ( new_n41245_, new_n41243_, new_n41239_ );
and  ( new_n41246_, new_n4958_, RIbb33378_192 );
nor  ( new_n41247_, new_n41246_, new_n4708_ );
and  ( new_n41248_, new_n41246_, new_n4705_ );
nor  ( new_n41249_, new_n41248_, new_n41247_ );
or   ( new_n41250_, new_n41249_, new_n41245_ );
and  ( new_n41251_, new_n41250_, new_n41244_ );
nor  ( new_n41252_, new_n41251_, new_n41235_ );
and  ( new_n41253_, new_n41251_, new_n41235_ );
or   ( new_n41254_, new_n5207_, new_n31952_ );
or   ( new_n41255_, new_n5209_, new_n31654_ );
and  ( new_n41256_, new_n41255_, new_n41254_ );
xor  ( new_n41257_, new_n41256_, new_n4708_ );
not  ( new_n41258_, new_n41257_ );
nor  ( new_n41259_, new_n41258_, new_n41253_ );
nor  ( new_n41260_, new_n41259_, new_n41252_ );
nor  ( new_n41261_, new_n41260_, new_n41231_ );
nor  ( new_n41262_, new_n41261_, new_n41230_ );
nor  ( new_n41263_, new_n41262_, new_n41168_ );
nor  ( new_n41264_, new_n41263_, new_n41167_ );
or   ( new_n41265_, new_n41264_, new_n41155_ );
and  ( new_n41266_, new_n41265_, new_n41154_ );
nor  ( new_n41267_, new_n41266_, new_n41149_ );
xnor ( new_n41268_, new_n41166_, new_n41157_ );
xor  ( new_n41269_, new_n41268_, new_n41262_ );
xnor ( new_n41270_, new_n41121_, new_n41067_ );
xor  ( new_n41271_, new_n41270_, new_n41135_ );
and  ( new_n41272_, new_n41271_, new_n41269_ );
nor  ( new_n41273_, new_n41271_, new_n41269_ );
or   ( new_n41274_, new_n10059_, new_n27396_ );
or   ( new_n41275_, new_n10061_, new_n27085_ );
and  ( new_n41276_, new_n41275_, new_n41274_ );
xor  ( new_n41277_, new_n41276_, new_n9421_ );
and  ( new_n41278_, RIbb32a90_173, RIbb2d888_64 );
or   ( new_n41279_, new_n26762_, RIbb2d888_64 );
and  ( new_n41280_, new_n41279_, RIbb2d900_63 );
or   ( new_n41281_, new_n41280_, new_n41278_ );
or   ( new_n41282_, new_n10770_, new_n26620_ );
and  ( new_n41283_, new_n41282_, new_n41281_ );
or   ( new_n41284_, new_n41283_, new_n41277_ );
and  ( new_n41285_, new_n41283_, new_n41277_ );
or   ( new_n41286_, new_n9422_, new_n27763_ );
or   ( new_n41287_, new_n9424_, new_n27602_ );
and  ( new_n41288_, new_n41287_, new_n41286_ );
xor  ( new_n41289_, new_n41288_, new_n8873_ );
or   ( new_n41290_, new_n41289_, new_n41285_ );
and  ( new_n41291_, new_n41290_, new_n41284_ );
or   ( new_n41292_, new_n7184_, new_n30120_ );
or   ( new_n41293_, new_n7186_, new_n29619_ );
and  ( new_n41294_, new_n41293_, new_n41292_ );
xor  ( new_n41295_, new_n41294_, new_n6638_ );
or   ( new_n41296_, new_n6645_, new_n30800_ );
or   ( new_n41297_, new_n6647_, new_n30227_ );
and  ( new_n41298_, new_n41297_, new_n41296_ );
xor  ( new_n41299_, new_n41298_, new_n6166_ );
or   ( new_n41300_, new_n41299_, new_n41295_ );
and  ( new_n41301_, new_n41299_, new_n41295_ );
or   ( new_n41302_, new_n6173_, new_n31333_ );
or   ( new_n41303_, new_n6175_, new_n30798_ );
and  ( new_n41304_, new_n41303_, new_n41302_ );
xor  ( new_n41305_, new_n41304_, new_n5597_ );
or   ( new_n41306_, new_n41305_, new_n41301_ );
and  ( new_n41307_, new_n41306_, new_n41300_ );
or   ( new_n41308_, new_n41307_, new_n41291_ );
and  ( new_n41309_, new_n41307_, new_n41291_ );
or   ( new_n41310_, new_n8874_, new_n28314_ );
or   ( new_n41311_, new_n8876_, new_n28108_ );
and  ( new_n41312_, new_n41311_, new_n41310_ );
xor  ( new_n41313_, new_n41312_, new_n8257_ );
or   ( new_n41314_, new_n8264_, new_n29263_ );
or   ( new_n41315_, new_n8266_, new_n28531_ );
and  ( new_n41316_, new_n41315_, new_n41314_ );
xor  ( new_n41317_, new_n41316_, new_n7725_ );
nor  ( new_n41318_, new_n41317_, new_n41313_ );
and  ( new_n41319_, new_n41317_, new_n41313_ );
or   ( new_n41320_, new_n7732_, new_n29474_ );
or   ( new_n41321_, new_n7734_, new_n29261_ );
and  ( new_n41322_, new_n41321_, new_n41320_ );
xor  ( new_n41323_, new_n41322_, new_n7177_ );
nor  ( new_n41324_, new_n41323_, new_n41319_ );
nor  ( new_n41325_, new_n41324_, new_n41318_ );
or   ( new_n41326_, new_n41325_, new_n41309_ );
and  ( new_n41327_, new_n41326_, new_n41308_ );
xnor ( new_n41328_, new_n41223_, new_n41221_ );
xor  ( new_n41329_, new_n41328_, new_n41227_ );
or   ( new_n41330_, new_n41329_, new_n41327_ );
nand ( new_n41331_, new_n41329_, new_n41327_ );
xor  ( new_n41332_, new_n41190_, new_n41186_ );
xor  ( new_n41333_, new_n41332_, new_n41196_ );
xnor ( new_n41334_, new_n41243_, new_n41239_ );
xor  ( new_n41335_, new_n41334_, new_n41249_ );
and  ( new_n41336_, new_n41335_, new_n41333_ );
nor  ( new_n41337_, new_n41335_, new_n41333_ );
xor  ( new_n41338_, new_n41208_, new_n41204_ );
xnor ( new_n41339_, new_n41338_, new_n41214_ );
nor  ( new_n41340_, new_n41339_, new_n41337_ );
nor  ( new_n41341_, new_n41340_, new_n41336_ );
nand ( new_n41342_, new_n41341_, new_n41331_ );
and  ( new_n41343_, new_n41342_, new_n41330_ );
xnor ( new_n41344_, new_n41229_, new_n41219_ );
xor  ( new_n41345_, new_n41344_, new_n41260_ );
and  ( new_n41346_, new_n41345_, new_n41343_ );
nor  ( new_n41347_, new_n41345_, new_n41343_ );
xor  ( new_n41348_, new_n41161_, new_n41159_ );
xor  ( new_n41349_, new_n41348_, new_n41164_ );
not  ( new_n41350_, new_n41349_ );
nor  ( new_n41351_, new_n41350_, new_n41347_ );
nor  ( new_n41352_, new_n41351_, new_n41346_ );
nor  ( new_n41353_, new_n41352_, new_n41273_ );
or   ( new_n41354_, new_n41353_, new_n41272_ );
xnor ( new_n41355_, new_n41153_, new_n41151_ );
xor  ( new_n41356_, new_n41355_, new_n41264_ );
and  ( new_n41357_, new_n41356_, new_n41354_ );
xor  ( new_n41358_, new_n41271_, new_n41269_ );
xor  ( new_n41359_, new_n41358_, new_n41352_ );
xor  ( new_n41360_, new_n41198_, new_n41182_ );
xor  ( new_n41361_, new_n41360_, new_n41217_ );
xor  ( new_n41362_, new_n41329_, new_n41327_ );
xor  ( new_n41363_, new_n41362_, new_n41341_ );
or   ( new_n41364_, new_n41363_, new_n41361_ );
xor  ( new_n41365_, new_n41307_, new_n41291_ );
xnor ( new_n41366_, new_n41365_, new_n41325_ );
xnor ( new_n41367_, new_n41335_, new_n41333_ );
xnor ( new_n41368_, new_n41367_, new_n41339_ );
nor  ( new_n41369_, new_n41368_, new_n41366_ );
xor  ( new_n41370_, new_n41178_, new_n41172_ );
xor  ( new_n41371_, new_n41370_, new_n4707_ );
or   ( new_n41372_, new_n5604_, new_n31952_ );
or   ( new_n41373_, new_n5606_, new_n31654_ );
and  ( new_n41374_, new_n41373_, new_n41372_ );
xor  ( new_n41375_, new_n41374_, new_n5205_ );
xnor ( new_n41376_, new_n41299_, new_n41295_ );
xor  ( new_n41377_, new_n41376_, new_n41305_ );
nand ( new_n41378_, new_n41377_, new_n41375_ );
nor  ( new_n41379_, new_n41377_, new_n41375_ );
xor  ( new_n41380_, new_n41317_, new_n41313_ );
xor  ( new_n41381_, new_n41380_, new_n41323_ );
or   ( new_n41382_, new_n41381_, new_n41379_ );
and  ( new_n41383_, new_n41382_, new_n41378_ );
or   ( new_n41384_, new_n41383_, new_n41371_ );
and  ( new_n41385_, new_n41383_, new_n41371_ );
or   ( new_n41386_, new_n10059_, new_n27602_ );
or   ( new_n41387_, new_n10061_, new_n27396_ );
and  ( new_n41388_, new_n41387_, new_n41386_ );
xor  ( new_n41389_, new_n41388_, new_n9421_ );
and  ( new_n41390_, RIbb32b08_174, RIbb2d888_64 );
or   ( new_n41391_, new_n27085_, RIbb2d888_64 );
and  ( new_n41392_, new_n41391_, RIbb2d900_63 );
or   ( new_n41393_, new_n41392_, new_n41390_ );
or   ( new_n41394_, new_n10770_, new_n26762_ );
and  ( new_n41395_, new_n41394_, new_n41393_ );
or   ( new_n41396_, new_n41395_, new_n41389_ );
and  ( new_n41397_, new_n41395_, new_n41389_ );
or   ( new_n41398_, new_n41397_, new_n5205_ );
and  ( new_n41399_, new_n41398_, new_n41396_ );
or   ( new_n41400_, new_n7732_, new_n29619_ );
or   ( new_n41401_, new_n7734_, new_n29474_ );
and  ( new_n41402_, new_n41401_, new_n41400_ );
xor  ( new_n41403_, new_n41402_, new_n7177_ );
or   ( new_n41404_, new_n7184_, new_n30227_ );
or   ( new_n41405_, new_n7186_, new_n30120_ );
and  ( new_n41406_, new_n41405_, new_n41404_ );
xor  ( new_n41407_, new_n41406_, new_n6638_ );
or   ( new_n41408_, new_n41407_, new_n41403_ );
and  ( new_n41409_, new_n41407_, new_n41403_ );
or   ( new_n41410_, new_n6645_, new_n30798_ );
or   ( new_n41411_, new_n6647_, new_n30800_ );
and  ( new_n41412_, new_n41411_, new_n41410_ );
xor  ( new_n41413_, new_n41412_, new_n6166_ );
or   ( new_n41414_, new_n41413_, new_n41409_ );
and  ( new_n41415_, new_n41414_, new_n41408_ );
nor  ( new_n41416_, new_n41415_, new_n41399_ );
and  ( new_n41417_, new_n41415_, new_n41399_ );
or   ( new_n41418_, new_n9422_, new_n28108_ );
or   ( new_n41419_, new_n9424_, new_n27763_ );
and  ( new_n41420_, new_n41419_, new_n41418_ );
xor  ( new_n41421_, new_n41420_, new_n8873_ );
or   ( new_n41422_, new_n8874_, new_n28531_ );
or   ( new_n41423_, new_n8876_, new_n28314_ );
and  ( new_n41424_, new_n41423_, new_n41422_ );
xor  ( new_n41425_, new_n41424_, new_n8257_ );
nor  ( new_n41426_, new_n41425_, new_n41421_ );
and  ( new_n41427_, new_n41425_, new_n41421_ );
or   ( new_n41428_, new_n8264_, new_n29261_ );
or   ( new_n41429_, new_n8266_, new_n29263_ );
and  ( new_n41430_, new_n41429_, new_n41428_ );
xor  ( new_n41431_, new_n41430_, new_n7725_ );
nor  ( new_n41432_, new_n41431_, new_n41427_ );
nor  ( new_n41433_, new_n41432_, new_n41426_ );
nor  ( new_n41434_, new_n41433_, new_n41417_ );
nor  ( new_n41435_, new_n41434_, new_n41416_ );
or   ( new_n41436_, new_n41435_, new_n41385_ );
and  ( new_n41437_, new_n41436_, new_n41384_ );
nand ( new_n41438_, new_n41437_, new_n41369_ );
nor  ( new_n41439_, new_n41437_, new_n41369_ );
xor  ( new_n41440_, new_n41251_, new_n41235_ );
xor  ( new_n41441_, new_n41440_, new_n41258_ );
or   ( new_n41442_, new_n41441_, new_n41439_ );
and  ( new_n41443_, new_n41442_, new_n41438_ );
or   ( new_n41444_, new_n41443_, new_n41364_ );
and  ( new_n41445_, new_n41443_, new_n41364_ );
xor  ( new_n41446_, new_n41345_, new_n41343_ );
xor  ( new_n41447_, new_n41446_, new_n41350_ );
or   ( new_n41448_, new_n41447_, new_n41445_ );
and  ( new_n41449_, new_n41448_, new_n41444_ );
nor  ( new_n41450_, new_n41449_, new_n41359_ );
xor  ( new_n41451_, new_n41443_, new_n41364_ );
xor  ( new_n41452_, new_n41451_, new_n41447_ );
xor  ( new_n41453_, new_n41437_, new_n41369_ );
xor  ( new_n41454_, new_n41453_, new_n41441_ );
xor  ( new_n41455_, new_n41283_, new_n41277_ );
xor  ( new_n41456_, new_n41455_, new_n41289_ );
or   ( new_n41457_, new_n6173_, new_n31654_ );
or   ( new_n41458_, new_n6175_, new_n31333_ );
and  ( new_n41459_, new_n41458_, new_n41457_ );
xor  ( new_n41460_, new_n41459_, new_n5596_ );
and  ( new_n41461_, new_n5371_, RIbb33378_192 );
or   ( new_n41462_, new_n41461_, new_n5206_ );
nand ( new_n41463_, new_n41461_, new_n5203_ );
and  ( new_n41464_, new_n41463_, new_n41462_ );
nand ( new_n41465_, new_n41464_, new_n41460_ );
or   ( new_n41466_, new_n41464_, new_n41460_ );
xor  ( new_n41467_, new_n41407_, new_n41403_ );
xnor ( new_n41468_, new_n41467_, new_n41413_ );
nand ( new_n41469_, new_n41468_, new_n41466_ );
and  ( new_n41470_, new_n41469_, new_n41465_ );
nor  ( new_n41471_, new_n41470_, new_n41456_ );
nand ( new_n41472_, new_n41470_, new_n41456_ );
or   ( new_n41473_, new_n10059_, new_n27763_ );
or   ( new_n41474_, new_n10061_, new_n27602_ );
and  ( new_n41475_, new_n41474_, new_n41473_ );
xor  ( new_n41476_, new_n41475_, new_n9421_ );
and  ( new_n41477_, RIbb32b80_175, RIbb2d888_64 );
or   ( new_n41478_, new_n27396_, RIbb2d888_64 );
and  ( new_n41479_, new_n41478_, RIbb2d900_63 );
or   ( new_n41480_, new_n41479_, new_n41477_ );
or   ( new_n41481_, new_n10770_, new_n27085_ );
and  ( new_n41482_, new_n41481_, new_n41480_ );
or   ( new_n41483_, new_n41482_, new_n41476_ );
and  ( new_n41484_, new_n41482_, new_n41476_ );
or   ( new_n41485_, new_n9422_, new_n28314_ );
or   ( new_n41486_, new_n9424_, new_n28108_ );
and  ( new_n41487_, new_n41486_, new_n41485_ );
xor  ( new_n41488_, new_n41487_, new_n8873_ );
or   ( new_n41489_, new_n41488_, new_n41484_ );
and  ( new_n41490_, new_n41489_, new_n41483_ );
or   ( new_n41491_, new_n8874_, new_n29263_ );
or   ( new_n41492_, new_n8876_, new_n28531_ );
and  ( new_n41493_, new_n41492_, new_n41491_ );
xor  ( new_n41494_, new_n41493_, new_n8257_ );
or   ( new_n41495_, new_n8264_, new_n29474_ );
or   ( new_n41496_, new_n8266_, new_n29261_ );
and  ( new_n41497_, new_n41496_, new_n41495_ );
xor  ( new_n41498_, new_n41497_, new_n7725_ );
or   ( new_n41499_, new_n41498_, new_n41494_ );
and  ( new_n41500_, new_n41498_, new_n41494_ );
or   ( new_n41501_, new_n7732_, new_n30120_ );
or   ( new_n41502_, new_n7734_, new_n29619_ );
and  ( new_n41503_, new_n41502_, new_n41501_ );
xor  ( new_n41504_, new_n41503_, new_n7177_ );
or   ( new_n41505_, new_n41504_, new_n41500_ );
and  ( new_n41506_, new_n41505_, new_n41499_ );
nor  ( new_n41507_, new_n41506_, new_n41490_ );
nand ( new_n41508_, new_n41506_, new_n41490_ );
or   ( new_n41509_, new_n7184_, new_n30800_ );
or   ( new_n41510_, new_n7186_, new_n30227_ );
and  ( new_n41511_, new_n41510_, new_n41509_ );
xor  ( new_n41512_, new_n41511_, new_n6638_ );
or   ( new_n41513_, new_n6645_, new_n31333_ );
or   ( new_n41514_, new_n6647_, new_n30798_ );
and  ( new_n41515_, new_n41514_, new_n41513_ );
xor  ( new_n41516_, new_n41515_, new_n6166_ );
nor  ( new_n41517_, new_n41516_, new_n41512_ );
nand ( new_n41518_, new_n41516_, new_n41512_ );
or   ( new_n41519_, new_n6173_, new_n31952_ );
or   ( new_n41520_, new_n6175_, new_n31654_ );
and  ( new_n41521_, new_n41520_, new_n41519_ );
xor  ( new_n41522_, new_n41521_, new_n5597_ );
not  ( new_n41523_, new_n41522_ );
and  ( new_n41524_, new_n41523_, new_n41518_ );
or   ( new_n41525_, new_n41524_, new_n41517_ );
and  ( new_n41526_, new_n41525_, new_n41508_ );
or   ( new_n41527_, new_n41526_, new_n41507_ );
and  ( new_n41528_, new_n41527_, new_n41472_ );
or   ( new_n41529_, new_n41528_, new_n41471_ );
xnor ( new_n41530_, new_n41383_, new_n41371_ );
xor  ( new_n41531_, new_n41530_, new_n41435_ );
or   ( new_n41532_, new_n41531_, new_n41529_ );
and  ( new_n41533_, new_n41531_, new_n41529_ );
xnor ( new_n41534_, new_n41368_, new_n41366_ );
or   ( new_n41535_, new_n41534_, new_n41533_ );
and  ( new_n41536_, new_n41535_, new_n41532_ );
or   ( new_n41537_, new_n41536_, new_n41454_ );
and  ( new_n41538_, new_n41536_, new_n41454_ );
xnor ( new_n41539_, new_n41363_, new_n41361_ );
or   ( new_n41540_, new_n41539_, new_n41538_ );
and  ( new_n41541_, new_n41540_, new_n41537_ );
nor  ( new_n41542_, new_n41541_, new_n41452_ );
xor  ( new_n41543_, new_n41536_, new_n41454_ );
xor  ( new_n41544_, new_n41543_, new_n41539_ );
xor  ( new_n41545_, new_n41415_, new_n41399_ );
xnor ( new_n41546_, new_n41545_, new_n41433_ );
xor  ( new_n41547_, new_n41470_, new_n41456_ );
xor  ( new_n41548_, new_n41547_, new_n41527_ );
nor  ( new_n41549_, new_n41548_, new_n41546_ );
xor  ( new_n41550_, new_n41377_, new_n41375_ );
xor  ( new_n41551_, new_n41550_, new_n41381_ );
xor  ( new_n41552_, new_n41425_, new_n41421_ );
xor  ( new_n41553_, new_n41552_, new_n41431_ );
or   ( new_n41554_, new_n9422_, new_n28531_ );
or   ( new_n41555_, new_n9424_, new_n28314_ );
and  ( new_n41556_, new_n41555_, new_n41554_ );
xor  ( new_n41557_, new_n41556_, new_n8873_ );
or   ( new_n41558_, new_n8874_, new_n29261_ );
or   ( new_n41559_, new_n8876_, new_n29263_ );
and  ( new_n41560_, new_n41559_, new_n41558_ );
xor  ( new_n41561_, new_n41560_, new_n8257_ );
nor  ( new_n41562_, new_n41561_, new_n41557_ );
and  ( new_n41563_, new_n41561_, new_n41557_ );
or   ( new_n41564_, new_n8264_, new_n29619_ );
or   ( new_n41565_, new_n8266_, new_n29474_ );
and  ( new_n41566_, new_n41565_, new_n41564_ );
xor  ( new_n41567_, new_n41566_, new_n7725_ );
nor  ( new_n41568_, new_n41567_, new_n41563_ );
nor  ( new_n41569_, new_n41568_, new_n41562_ );
or   ( new_n41570_, new_n10059_, new_n28108_ );
or   ( new_n41571_, new_n10061_, new_n27763_ );
and  ( new_n41572_, new_n41571_, new_n41570_ );
xor  ( new_n41573_, new_n41572_, new_n9421_ );
and  ( new_n41574_, RIbb32bf8_176, RIbb2d888_64 );
or   ( new_n41575_, new_n27602_, RIbb2d888_64 );
and  ( new_n41576_, new_n41575_, RIbb2d900_63 );
or   ( new_n41577_, new_n41576_, new_n41574_ );
or   ( new_n41578_, new_n10770_, new_n27396_ );
and  ( new_n41579_, new_n41578_, new_n41577_ );
nor  ( new_n41580_, new_n41579_, new_n41573_ );
and  ( new_n41581_, new_n41579_, new_n41573_ );
nor  ( new_n41582_, new_n41581_, new_n5596_ );
nor  ( new_n41583_, new_n41582_, new_n41580_ );
or   ( new_n41584_, new_n7732_, new_n30227_ );
or   ( new_n41585_, new_n7734_, new_n30120_ );
and  ( new_n41586_, new_n41585_, new_n41584_ );
xor  ( new_n41587_, new_n41586_, new_n7177_ );
or   ( new_n41588_, new_n7184_, new_n30798_ );
or   ( new_n41589_, new_n7186_, new_n30800_ );
and  ( new_n41590_, new_n41589_, new_n41588_ );
xor  ( new_n41591_, new_n41590_, new_n6638_ );
or   ( new_n41592_, new_n41591_, new_n41587_ );
and  ( new_n41593_, new_n41591_, new_n41587_ );
or   ( new_n41594_, new_n6645_, new_n31654_ );
or   ( new_n41595_, new_n6647_, new_n31333_ );
and  ( new_n41596_, new_n41595_, new_n41594_ );
xor  ( new_n41597_, new_n41596_, new_n6166_ );
or   ( new_n41598_, new_n41597_, new_n41593_ );
and  ( new_n41599_, new_n41598_, new_n41592_ );
and  ( new_n41600_, new_n41599_, new_n41583_ );
or   ( new_n41601_, new_n41600_, new_n41569_ );
or   ( new_n41602_, new_n41599_, new_n41583_ );
and  ( new_n41603_, new_n41602_, new_n41601_ );
or   ( new_n41604_, new_n41603_, new_n41553_ );
nand ( new_n41605_, new_n41603_, new_n41553_ );
xnor ( new_n41606_, new_n41498_, new_n41494_ );
xor  ( new_n41607_, new_n41606_, new_n41504_ );
xnor ( new_n41608_, new_n41482_, new_n41476_ );
xor  ( new_n41609_, new_n41608_, new_n41488_ );
nor  ( new_n41610_, new_n41609_, new_n41607_ );
and  ( new_n41611_, new_n41609_, new_n41607_ );
xor  ( new_n41612_, new_n41516_, new_n41512_ );
xor  ( new_n41613_, new_n41612_, new_n41523_ );
nor  ( new_n41614_, new_n41613_, new_n41611_ );
nor  ( new_n41615_, new_n41614_, new_n41610_ );
nand ( new_n41616_, new_n41615_, new_n41605_ );
and  ( new_n41617_, new_n41616_, new_n41604_ );
or   ( new_n41618_, new_n41617_, new_n41551_ );
nand ( new_n41619_, new_n41617_, new_n41551_ );
xor  ( new_n41620_, new_n41395_, new_n41389_ );
xor  ( new_n41621_, new_n41620_, new_n5206_ );
xor  ( new_n41622_, new_n41506_, new_n41490_ );
xor  ( new_n41623_, new_n41622_, new_n41525_ );
nor  ( new_n41624_, new_n41623_, new_n41621_ );
and  ( new_n41625_, new_n41623_, new_n41621_ );
xor  ( new_n41626_, new_n41464_, new_n41460_ );
xor  ( new_n41627_, new_n41626_, new_n41468_ );
nor  ( new_n41628_, new_n41627_, new_n41625_ );
nor  ( new_n41629_, new_n41628_, new_n41624_ );
nand ( new_n41630_, new_n41629_, new_n41619_ );
and  ( new_n41631_, new_n41630_, new_n41618_ );
nand ( new_n41632_, new_n41631_, new_n41549_ );
nor  ( new_n41633_, new_n41631_, new_n41549_ );
xor  ( new_n41634_, new_n41531_, new_n41529_ );
xor  ( new_n41635_, new_n41634_, new_n41534_ );
or   ( new_n41636_, new_n41635_, new_n41633_ );
and  ( new_n41637_, new_n41636_, new_n41632_ );
nor  ( new_n41638_, new_n41637_, new_n41544_ );
xor  ( new_n41639_, new_n41631_, new_n41549_ );
xor  ( new_n41640_, new_n41639_, new_n41635_ );
xor  ( new_n41641_, new_n41617_, new_n41551_ );
xor  ( new_n41642_, new_n41641_, new_n41629_ );
and  ( new_n41643_, new_n5915_, RIbb33378_192 );
or   ( new_n41644_, new_n41643_, new_n5597_ );
nand ( new_n41645_, new_n41643_, new_n5594_ );
and  ( new_n41646_, new_n41645_, new_n41644_ );
xnor ( new_n41647_, new_n41591_, new_n41587_ );
xor  ( new_n41648_, new_n41647_, new_n41597_ );
nor  ( new_n41649_, new_n41648_, new_n41646_ );
nand ( new_n41650_, new_n41648_, new_n41646_ );
xor  ( new_n41651_, new_n41561_, new_n41557_ );
xor  ( new_n41652_, new_n41651_, new_n41567_ );
and  ( new_n41653_, new_n41652_, new_n41650_ );
or   ( new_n41654_, new_n41653_, new_n41649_ );
xnor ( new_n41655_, new_n41609_, new_n41607_ );
xor  ( new_n41656_, new_n41655_, new_n41613_ );
nor  ( new_n41657_, new_n41656_, new_n41654_ );
nand ( new_n41658_, new_n41656_, new_n41654_ );
or   ( new_n41659_, new_n10059_, new_n28314_ );
or   ( new_n41660_, new_n10061_, new_n28108_ );
and  ( new_n41661_, new_n41660_, new_n41659_ );
xor  ( new_n41662_, new_n41661_, new_n9421_ );
and  ( new_n41663_, RIbb32c70_177, RIbb2d888_64 );
or   ( new_n41664_, new_n27763_, RIbb2d888_64 );
and  ( new_n41665_, new_n41664_, RIbb2d900_63 );
or   ( new_n41666_, new_n41665_, new_n41663_ );
or   ( new_n41667_, new_n10770_, new_n27602_ );
and  ( new_n41668_, new_n41667_, new_n41666_ );
nor  ( new_n41669_, new_n41668_, new_n41662_ );
nand ( new_n41670_, new_n41668_, new_n41662_ );
or   ( new_n41671_, new_n9422_, new_n29263_ );
or   ( new_n41672_, new_n9424_, new_n28531_ );
and  ( new_n41673_, new_n41672_, new_n41671_ );
xor  ( new_n41674_, new_n41673_, new_n8872_ );
and  ( new_n41675_, new_n41674_, new_n41670_ );
or   ( new_n41676_, new_n41675_, new_n41669_ );
or   ( new_n41677_, new_n7184_, new_n31333_ );
or   ( new_n41678_, new_n7186_, new_n30798_ );
and  ( new_n41679_, new_n41678_, new_n41677_ );
xor  ( new_n41680_, new_n41679_, new_n6638_ );
or   ( new_n41681_, new_n6645_, new_n31952_ );
or   ( new_n41682_, new_n6647_, new_n31654_ );
and  ( new_n41683_, new_n41682_, new_n41681_ );
xor  ( new_n41684_, new_n41683_, new_n6166_ );
and  ( new_n41685_, new_n41684_, new_n41680_ );
not  ( new_n41686_, new_n41685_ );
or   ( new_n41687_, new_n8874_, new_n29474_ );
or   ( new_n41688_, new_n8876_, new_n29261_ );
and  ( new_n41689_, new_n41688_, new_n41687_ );
xor  ( new_n41690_, new_n41689_, new_n8257_ );
or   ( new_n41691_, new_n8264_, new_n30120_ );
or   ( new_n41692_, new_n8266_, new_n29619_ );
and  ( new_n41693_, new_n41692_, new_n41691_ );
xor  ( new_n41694_, new_n41693_, new_n7725_ );
nor  ( new_n41695_, new_n41694_, new_n41690_ );
and  ( new_n41696_, new_n41694_, new_n41690_ );
or   ( new_n41697_, new_n7732_, new_n30800_ );
or   ( new_n41698_, new_n7734_, new_n30227_ );
and  ( new_n41699_, new_n41698_, new_n41697_ );
xor  ( new_n41700_, new_n41699_, new_n7177_ );
nor  ( new_n41701_, new_n41700_, new_n41696_ );
nor  ( new_n41702_, new_n41701_, new_n41695_ );
not  ( new_n41703_, new_n41702_ );
or   ( new_n41704_, new_n41703_, new_n41686_ );
and  ( new_n41705_, new_n41704_, new_n41676_ );
and  ( new_n41706_, new_n41703_, new_n41686_ );
or   ( new_n41707_, new_n41706_, new_n41705_ );
and  ( new_n41708_, new_n41707_, new_n41658_ );
or   ( new_n41709_, new_n41708_, new_n41657_ );
xor  ( new_n41710_, new_n41603_, new_n41553_ );
xor  ( new_n41711_, new_n41710_, new_n41615_ );
or   ( new_n41712_, new_n41711_, new_n41709_ );
and  ( new_n41713_, new_n41711_, new_n41709_ );
xor  ( new_n41714_, new_n41623_, new_n41621_ );
xor  ( new_n41715_, new_n41714_, new_n41627_ );
or   ( new_n41716_, new_n41715_, new_n41713_ );
and  ( new_n41717_, new_n41716_, new_n41712_ );
or   ( new_n41718_, new_n41717_, new_n41642_ );
nand ( new_n41719_, new_n41717_, new_n41642_ );
xor  ( new_n41720_, new_n41548_, new_n41546_ );
nand ( new_n41721_, new_n41720_, new_n41719_ );
and  ( new_n41722_, new_n41721_, new_n41718_ );
nor  ( new_n41723_, new_n41722_, new_n41640_ );
xor  ( new_n41724_, new_n41685_, new_n41676_ );
xor  ( new_n41725_, new_n41724_, new_n41702_ );
not  ( new_n41726_, new_n41725_ );
xor  ( new_n41727_, new_n41648_, new_n41646_ );
xor  ( new_n41728_, new_n41727_, new_n41652_ );
nand ( new_n41729_, new_n41728_, new_n41726_ );
xor  ( new_n41730_, new_n41579_, new_n41573_ );
xor  ( new_n41731_, new_n41730_, new_n5597_ );
xor  ( new_n41732_, new_n41668_, new_n41662_ );
xor  ( new_n41733_, new_n41732_, new_n41674_ );
xnor ( new_n41734_, new_n41694_, new_n41690_ );
xor  ( new_n41735_, new_n41734_, new_n41700_ );
or   ( new_n41736_, new_n41735_, new_n41733_ );
nand ( new_n41737_, new_n41735_, new_n41733_ );
xor  ( new_n41738_, new_n41684_, new_n41680_ );
nand ( new_n41739_, new_n41738_, new_n41737_ );
and  ( new_n41740_, new_n41739_, new_n41736_ );
or   ( new_n41741_, new_n41740_, new_n41731_ );
and  ( new_n41742_, new_n41740_, new_n41731_ );
or   ( new_n41743_, new_n10059_, new_n28531_ );
or   ( new_n41744_, new_n10061_, new_n28314_ );
and  ( new_n41745_, new_n41744_, new_n41743_ );
xor  ( new_n41746_, new_n41745_, new_n9421_ );
and  ( new_n41747_, RIbb32ce8_178, RIbb2d888_64 );
or   ( new_n41748_, new_n28108_, RIbb2d888_64 );
and  ( new_n41749_, new_n41748_, RIbb2d900_63 );
or   ( new_n41750_, new_n41749_, new_n41747_ );
or   ( new_n41751_, new_n10770_, new_n27763_ );
and  ( new_n41752_, new_n41751_, new_n41750_ );
or   ( new_n41753_, new_n41752_, new_n41746_ );
and  ( new_n41754_, new_n41752_, new_n41746_ );
or   ( new_n41755_, new_n41754_, new_n6165_ );
and  ( new_n41756_, new_n41755_, new_n41753_ );
or   ( new_n41757_, new_n9422_, new_n29261_ );
or   ( new_n41758_, new_n9424_, new_n29263_ );
and  ( new_n41759_, new_n41758_, new_n41757_ );
xor  ( new_n41760_, new_n41759_, new_n8873_ );
or   ( new_n41761_, new_n8874_, new_n29619_ );
or   ( new_n41762_, new_n8876_, new_n29474_ );
and  ( new_n41763_, new_n41762_, new_n41761_ );
xor  ( new_n41764_, new_n41763_, new_n8257_ );
or   ( new_n41765_, new_n41764_, new_n41760_ );
and  ( new_n41766_, new_n41764_, new_n41760_ );
or   ( new_n41767_, new_n8264_, new_n30227_ );
or   ( new_n41768_, new_n8266_, new_n30120_ );
and  ( new_n41769_, new_n41768_, new_n41767_ );
xor  ( new_n41770_, new_n41769_, new_n7725_ );
or   ( new_n41771_, new_n41770_, new_n41766_ );
and  ( new_n41772_, new_n41771_, new_n41765_ );
and  ( new_n41773_, new_n41772_, new_n41756_ );
nor  ( new_n41774_, new_n41772_, new_n41756_ );
or   ( new_n41775_, new_n7732_, new_n30798_ );
or   ( new_n41776_, new_n7734_, new_n30800_ );
and  ( new_n41777_, new_n41776_, new_n41775_ );
xor  ( new_n41778_, new_n41777_, new_n7177_ );
or   ( new_n41779_, new_n7184_, new_n31654_ );
or   ( new_n41780_, new_n7186_, new_n31333_ );
and  ( new_n41781_, new_n41780_, new_n41779_ );
xor  ( new_n41782_, new_n41781_, new_n6638_ );
and  ( new_n41783_, new_n41782_, new_n41778_ );
nor  ( new_n41784_, new_n41782_, new_n41778_ );
and  ( new_n41785_, new_n6508_, RIbb33378_192 );
nor  ( new_n41786_, new_n41785_, new_n6166_ );
and  ( new_n41787_, new_n41785_, new_n6163_ );
nor  ( new_n41788_, new_n41787_, new_n41786_ );
nor  ( new_n41789_, new_n41788_, new_n41784_ );
nor  ( new_n41790_, new_n41789_, new_n41783_ );
nor  ( new_n41791_, new_n41790_, new_n41774_ );
nor  ( new_n41792_, new_n41791_, new_n41773_ );
or   ( new_n41793_, new_n41792_, new_n41742_ );
and  ( new_n41794_, new_n41793_, new_n41741_ );
or   ( new_n41795_, new_n41794_, new_n41729_ );
and  ( new_n41796_, new_n41794_, new_n41729_ );
xnor ( new_n41797_, new_n41599_, new_n41583_ );
xnor ( new_n41798_, new_n41797_, new_n41569_ );
not  ( new_n41799_, new_n41798_ );
or   ( new_n41800_, new_n41799_, new_n41796_ );
and  ( new_n41801_, new_n41800_, new_n41795_ );
xor  ( new_n41802_, new_n41711_, new_n41709_ );
xor  ( new_n41803_, new_n41802_, new_n41715_ );
nor  ( new_n41804_, new_n41803_, new_n41801_ );
xor  ( new_n41805_, new_n41717_, new_n41642_ );
xor  ( new_n41806_, new_n41805_, new_n41720_ );
and  ( new_n41807_, new_n41806_, new_n41804_ );
xor  ( new_n41808_, new_n41794_, new_n41729_ );
xor  ( new_n41809_, new_n41808_, new_n41799_ );
xor  ( new_n41810_, new_n41656_, new_n41654_ );
xor  ( new_n41811_, new_n41810_, new_n41707_ );
nor  ( new_n41812_, new_n41811_, new_n41809_ );
xor  ( new_n41813_, new_n41803_, new_n41801_ );
and  ( new_n41814_, new_n41813_, new_n41812_ );
xnor ( new_n41815_, new_n41811_, new_n41809_ );
xor  ( new_n41816_, new_n41752_, new_n41746_ );
xor  ( new_n41817_, new_n41816_, new_n6166_ );
xnor ( new_n41818_, new_n41764_, new_n41760_ );
xor  ( new_n41819_, new_n41818_, new_n41770_ );
nor  ( new_n41820_, new_n41819_, new_n41817_ );
xor  ( new_n41821_, new_n41735_, new_n41733_ );
xor  ( new_n41822_, new_n41821_, new_n41738_ );
or   ( new_n41823_, new_n41822_, new_n41820_ );
and  ( new_n41824_, new_n41822_, new_n41820_ );
xnor ( new_n41825_, new_n41782_, new_n41778_ );
xor  ( new_n41826_, new_n41825_, new_n41788_ );
or   ( new_n41827_, new_n10059_, new_n29263_ );
or   ( new_n41828_, new_n10061_, new_n28531_ );
and  ( new_n41829_, new_n41828_, new_n41827_ );
xor  ( new_n41830_, new_n41829_, new_n9421_ );
and  ( new_n41831_, RIbb32d60_179, RIbb2d888_64 );
or   ( new_n41832_, new_n28314_, RIbb2d888_64 );
and  ( new_n41833_, new_n41832_, RIbb2d900_63 );
or   ( new_n41834_, new_n41833_, new_n41831_ );
or   ( new_n41835_, new_n10770_, new_n28108_ );
and  ( new_n41836_, new_n41835_, new_n41834_ );
or   ( new_n41837_, new_n41836_, new_n41830_ );
and  ( new_n41838_, new_n41836_, new_n41830_ );
or   ( new_n41839_, new_n9422_, new_n29474_ );
or   ( new_n41840_, new_n9424_, new_n29261_ );
and  ( new_n41841_, new_n41840_, new_n41839_ );
xor  ( new_n41842_, new_n41841_, new_n8873_ );
or   ( new_n41843_, new_n41842_, new_n41838_ );
and  ( new_n41844_, new_n41843_, new_n41837_ );
nor  ( new_n41845_, new_n41844_, new_n41826_ );
and  ( new_n41846_, new_n41844_, new_n41826_ );
or   ( new_n41847_, new_n8874_, new_n30120_ );
or   ( new_n41848_, new_n8876_, new_n29619_ );
and  ( new_n41849_, new_n41848_, new_n41847_ );
xor  ( new_n41850_, new_n41849_, new_n8257_ );
or   ( new_n41851_, new_n8264_, new_n30800_ );
or   ( new_n41852_, new_n8266_, new_n30227_ );
and  ( new_n41853_, new_n41852_, new_n41851_ );
xor  ( new_n41854_, new_n41853_, new_n7725_ );
nor  ( new_n41855_, new_n41854_, new_n41850_ );
and  ( new_n41856_, new_n41854_, new_n41850_ );
or   ( new_n41857_, new_n7732_, new_n31333_ );
or   ( new_n41858_, new_n7734_, new_n30798_ );
and  ( new_n41859_, new_n41858_, new_n41857_ );
xor  ( new_n41860_, new_n41859_, new_n7177_ );
nor  ( new_n41861_, new_n41860_, new_n41856_ );
nor  ( new_n41862_, new_n41861_, new_n41855_ );
nor  ( new_n41863_, new_n41862_, new_n41846_ );
nor  ( new_n41864_, new_n41863_, new_n41845_ );
or   ( new_n41865_, new_n41864_, new_n41824_ );
and  ( new_n41866_, new_n41865_, new_n41823_ );
xnor ( new_n41867_, new_n41740_, new_n41731_ );
xor  ( new_n41868_, new_n41867_, new_n41792_ );
nand ( new_n41869_, new_n41868_, new_n41866_ );
or   ( new_n41870_, new_n41868_, new_n41866_ );
xor  ( new_n41871_, new_n41728_, new_n41726_ );
nand ( new_n41872_, new_n41871_, new_n41870_ );
and  ( new_n41873_, new_n41872_, new_n41869_ );
nor  ( new_n41874_, new_n41873_, new_n41815_ );
xor  ( new_n41875_, new_n41868_, new_n41866_ );
xor  ( new_n41876_, new_n41875_, new_n41871_ );
xnor ( new_n41877_, new_n41772_, new_n41756_ );
xor  ( new_n41878_, new_n41877_, new_n41790_ );
or   ( new_n41879_, new_n7184_, new_n31952_ );
or   ( new_n41880_, new_n7186_, new_n31654_ );
and  ( new_n41881_, new_n41880_, new_n41879_ );
xor  ( new_n41882_, new_n41881_, new_n6638_ );
or   ( new_n41883_, new_n10059_, new_n29261_ );
or   ( new_n41884_, new_n10061_, new_n29263_ );
and  ( new_n41885_, new_n41884_, new_n41883_ );
xor  ( new_n41886_, new_n41885_, new_n9421_ );
and  ( new_n41887_, RIbb32dd8_180, RIbb2d888_64 );
or   ( new_n41888_, new_n28531_, RIbb2d888_64 );
and  ( new_n41889_, new_n41888_, RIbb2d900_63 );
or   ( new_n41890_, new_n41889_, new_n41887_ );
or   ( new_n41891_, new_n10770_, new_n28314_ );
and  ( new_n41892_, new_n41891_, new_n41890_ );
or   ( new_n41893_, new_n41892_, new_n41886_ );
and  ( new_n41894_, new_n41892_, new_n41886_ );
or   ( new_n41895_, new_n41894_, new_n6637_ );
and  ( new_n41896_, new_n41895_, new_n41893_ );
nor  ( new_n41897_, new_n41896_, new_n41882_ );
nand ( new_n41898_, new_n41896_, new_n41882_ );
or   ( new_n41899_, new_n9422_, new_n29619_ );
or   ( new_n41900_, new_n9424_, new_n29474_ );
and  ( new_n41901_, new_n41900_, new_n41899_ );
xor  ( new_n41902_, new_n41901_, new_n8873_ );
or   ( new_n41903_, new_n8874_, new_n30227_ );
or   ( new_n41904_, new_n8876_, new_n30120_ );
and  ( new_n41905_, new_n41904_, new_n41903_ );
xor  ( new_n41906_, new_n41905_, new_n8257_ );
nor  ( new_n41907_, new_n41906_, new_n41902_ );
nand ( new_n41908_, new_n41906_, new_n41902_ );
or   ( new_n41909_, new_n8264_, new_n30798_ );
or   ( new_n41910_, new_n8266_, new_n30800_ );
and  ( new_n41911_, new_n41910_, new_n41909_ );
xor  ( new_n41912_, new_n41911_, new_n7724_ );
and  ( new_n41913_, new_n41912_, new_n41908_ );
or   ( new_n41914_, new_n41913_, new_n41907_ );
and  ( new_n41915_, new_n41914_, new_n41898_ );
or   ( new_n41916_, new_n41915_, new_n41897_ );
xnor ( new_n41917_, new_n41844_, new_n41826_ );
xor  ( new_n41918_, new_n41917_, new_n41862_ );
nand ( new_n41919_, new_n41918_, new_n41916_ );
nor  ( new_n41920_, new_n41918_, new_n41916_ );
xor  ( new_n41921_, new_n41819_, new_n41817_ );
or   ( new_n41922_, new_n41921_, new_n41920_ );
and  ( new_n41923_, new_n41922_, new_n41919_ );
or   ( new_n41924_, new_n41923_, new_n41878_ );
nand ( new_n41925_, new_n41923_, new_n41878_ );
xor  ( new_n41926_, new_n41822_, new_n41820_ );
xnor ( new_n41927_, new_n41926_, new_n41864_ );
nand ( new_n41928_, new_n41927_, new_n41925_ );
and  ( new_n41929_, new_n41928_, new_n41924_ );
and  ( new_n41930_, new_n41929_, new_n41876_ );
xor  ( new_n41931_, new_n41836_, new_n41830_ );
xnor ( new_n41932_, new_n41931_, new_n41842_ );
xor  ( new_n41933_, new_n41896_, new_n41882_ );
xor  ( new_n41934_, new_n41933_, new_n41914_ );
or   ( new_n41935_, new_n41934_, new_n41932_ );
xnor ( new_n41936_, new_n41918_, new_n41916_ );
xor  ( new_n41937_, new_n41936_, new_n41921_ );
or   ( new_n41938_, new_n41937_, new_n41935_ );
nand ( new_n41939_, new_n41937_, new_n41935_ );
xor  ( new_n41940_, new_n41854_, new_n41850_ );
xor  ( new_n41941_, new_n41940_, new_n41860_ );
or   ( new_n41942_, new_n7732_, new_n31654_ );
or   ( new_n41943_, new_n7734_, new_n31333_ );
and  ( new_n41944_, new_n41943_, new_n41942_ );
xor  ( new_n41945_, new_n41944_, new_n7177_ );
or   ( new_n41946_, new_n8874_, new_n30800_ );
or   ( new_n41947_, new_n8876_, new_n30227_ );
and  ( new_n41948_, new_n41947_, new_n41946_ );
xor  ( new_n41949_, new_n41948_, new_n8257_ );
or   ( new_n41950_, new_n8264_, new_n31333_ );
or   ( new_n41951_, new_n8266_, new_n30798_ );
and  ( new_n41952_, new_n41951_, new_n41950_ );
xor  ( new_n41953_, new_n41952_, new_n7725_ );
or   ( new_n41954_, new_n41953_, new_n41949_ );
and  ( new_n41955_, new_n41953_, new_n41949_ );
or   ( new_n41956_, new_n7732_, new_n31952_ );
or   ( new_n41957_, new_n7734_, new_n31654_ );
and  ( new_n41958_, new_n41957_, new_n41956_ );
xor  ( new_n41959_, new_n41958_, new_n7177_ );
or   ( new_n41960_, new_n41959_, new_n41955_ );
and  ( new_n41961_, new_n41960_, new_n41954_ );
or   ( new_n41962_, new_n41961_, new_n41945_ );
and  ( new_n41963_, new_n41961_, new_n41945_ );
or   ( new_n41964_, new_n10059_, new_n29474_ );
or   ( new_n41965_, new_n10061_, new_n29261_ );
and  ( new_n41966_, new_n41965_, new_n41964_ );
xor  ( new_n41967_, new_n41966_, new_n9421_ );
and  ( new_n41968_, RIbb32e50_181, RIbb2d888_64 );
or   ( new_n41969_, new_n29263_, RIbb2d888_64 );
and  ( new_n41970_, new_n41969_, RIbb2d900_63 );
or   ( new_n41971_, new_n41970_, new_n41968_ );
or   ( new_n41972_, new_n10770_, new_n28531_ );
and  ( new_n41973_, new_n41972_, new_n41971_ );
nor  ( new_n41974_, new_n41973_, new_n41967_ );
and  ( new_n41975_, new_n41973_, new_n41967_ );
or   ( new_n41976_, new_n9422_, new_n30120_ );
or   ( new_n41977_, new_n9424_, new_n29619_ );
and  ( new_n41978_, new_n41977_, new_n41976_ );
xor  ( new_n41979_, new_n41978_, new_n8873_ );
nor  ( new_n41980_, new_n41979_, new_n41975_ );
nor  ( new_n41981_, new_n41980_, new_n41974_ );
or   ( new_n41982_, new_n41981_, new_n41963_ );
and  ( new_n41983_, new_n41982_, new_n41962_ );
nor  ( new_n41984_, new_n41983_, new_n41941_ );
and  ( new_n41985_, new_n41983_, new_n41941_ );
not  ( new_n41986_, new_n41985_ );
and  ( new_n41987_, new_n6908_, RIbb33378_192 );
or   ( new_n41988_, new_n41987_, new_n6638_ );
nand ( new_n41989_, new_n41987_, new_n6635_ );
and  ( new_n41990_, new_n41989_, new_n41988_ );
xor  ( new_n41991_, new_n41906_, new_n41902_ );
xor  ( new_n41992_, new_n41991_, new_n41912_ );
nor  ( new_n41993_, new_n41992_, new_n41990_ );
and  ( new_n41994_, new_n41992_, new_n41990_ );
xor  ( new_n41995_, new_n41892_, new_n41886_ );
xor  ( new_n41996_, new_n41995_, new_n6638_ );
nor  ( new_n41997_, new_n41996_, new_n41994_ );
nor  ( new_n41998_, new_n41997_, new_n41993_ );
and  ( new_n41999_, new_n41998_, new_n41986_ );
nor  ( new_n42000_, new_n41999_, new_n41984_ );
nand ( new_n42001_, new_n42000_, new_n41939_ );
and  ( new_n42002_, new_n42001_, new_n41938_ );
xor  ( new_n42003_, new_n41923_, new_n41878_ );
xor  ( new_n42004_, new_n42003_, new_n41927_ );
nor  ( new_n42005_, new_n42004_, new_n42002_ );
xor  ( new_n42006_, new_n41937_, new_n41935_ );
xor  ( new_n42007_, new_n42006_, new_n42000_ );
xnor ( new_n42008_, new_n41992_, new_n41990_ );
xor  ( new_n42009_, new_n42008_, new_n41996_ );
xor  ( new_n42010_, new_n41953_, new_n41949_ );
xor  ( new_n42011_, new_n42010_, new_n41959_ );
or   ( new_n42012_, new_n9422_, new_n30227_ );
or   ( new_n42013_, new_n9424_, new_n30120_ );
and  ( new_n42014_, new_n42013_, new_n42012_ );
xor  ( new_n42015_, new_n42014_, new_n8873_ );
or   ( new_n42016_, new_n8874_, new_n30798_ );
or   ( new_n42017_, new_n8876_, new_n30800_ );
and  ( new_n42018_, new_n42017_, new_n42016_ );
xor  ( new_n42019_, new_n42018_, new_n8257_ );
or   ( new_n42020_, new_n42019_, new_n42015_ );
and  ( new_n42021_, new_n42019_, new_n42015_ );
or   ( new_n42022_, new_n8264_, new_n31654_ );
or   ( new_n42023_, new_n8266_, new_n31333_ );
and  ( new_n42024_, new_n42023_, new_n42022_ );
xor  ( new_n42025_, new_n42024_, new_n7725_ );
or   ( new_n42026_, new_n42025_, new_n42021_ );
and  ( new_n42027_, new_n42026_, new_n42020_ );
or   ( new_n42028_, new_n42027_, new_n42011_ );
and  ( new_n42029_, new_n42027_, new_n42011_ );
or   ( new_n42030_, new_n10059_, new_n29619_ );
or   ( new_n42031_, new_n10061_, new_n29474_ );
and  ( new_n42032_, new_n42031_, new_n42030_ );
xor  ( new_n42033_, new_n42032_, new_n9421_ );
and  ( new_n42034_, RIbb32ec8_182, RIbb2d888_64 );
or   ( new_n42035_, new_n29261_, RIbb2d888_64 );
and  ( new_n42036_, new_n42035_, RIbb2d900_63 );
or   ( new_n42037_, new_n42036_, new_n42034_ );
or   ( new_n42038_, new_n10770_, new_n29263_ );
and  ( new_n42039_, new_n42038_, new_n42037_ );
nor  ( new_n42040_, new_n42039_, new_n42033_ );
and  ( new_n42041_, new_n42039_, new_n42033_ );
nor  ( new_n42042_, new_n42041_, new_n7176_ );
nor  ( new_n42043_, new_n42042_, new_n42040_ );
or   ( new_n42044_, new_n42043_, new_n42029_ );
and  ( new_n42045_, new_n42044_, new_n42028_ );
nor  ( new_n42046_, new_n42045_, new_n42009_ );
nand ( new_n42047_, new_n42045_, new_n42009_ );
xor  ( new_n42048_, new_n41961_, new_n41945_ );
xnor ( new_n42049_, new_n42048_, new_n41981_ );
and  ( new_n42050_, new_n42049_, new_n42047_ );
or   ( new_n42051_, new_n42050_, new_n42046_ );
xor  ( new_n42052_, new_n41983_, new_n41941_ );
xor  ( new_n42053_, new_n42052_, new_n41998_ );
nand ( new_n42054_, new_n42053_, new_n42051_ );
nor  ( new_n42055_, new_n42053_, new_n42051_ );
xor  ( new_n42056_, new_n41934_, new_n41932_ );
or   ( new_n42057_, new_n42056_, new_n42055_ );
and  ( new_n42058_, new_n42057_, new_n42054_ );
and  ( new_n42059_, new_n42058_, new_n42007_ );
and  ( new_n42060_, new_n7487_, RIbb33378_192 );
or   ( new_n42061_, new_n42060_, new_n7177_ );
nand ( new_n42062_, new_n42060_, new_n7174_ );
and  ( new_n42063_, new_n42062_, new_n42061_ );
xnor ( new_n42064_, new_n42019_, new_n42015_ );
xor  ( new_n42065_, new_n42064_, new_n42025_ );
or   ( new_n42066_, new_n42065_, new_n42063_ );
nand ( new_n42067_, new_n42065_, new_n42063_ );
or   ( new_n42068_, new_n10059_, new_n30120_ );
or   ( new_n42069_, new_n10061_, new_n29619_ );
and  ( new_n42070_, new_n42069_, new_n42068_ );
xor  ( new_n42071_, new_n42070_, new_n9421_ );
and  ( new_n42072_, RIbb32f40_183, RIbb2d888_64 );
or   ( new_n42073_, new_n29474_, RIbb2d888_64 );
and  ( new_n42074_, new_n42073_, RIbb2d900_63 );
or   ( new_n42075_, new_n42074_, new_n42072_ );
or   ( new_n42076_, new_n10770_, new_n29261_ );
and  ( new_n42077_, new_n42076_, new_n42075_ );
nor  ( new_n42078_, new_n42077_, new_n42071_ );
and  ( new_n42079_, new_n42077_, new_n42071_ );
or   ( new_n42080_, new_n9422_, new_n30800_ );
or   ( new_n42081_, new_n9424_, new_n30227_ );
and  ( new_n42082_, new_n42081_, new_n42080_ );
xor  ( new_n42083_, new_n42082_, new_n8873_ );
nor  ( new_n42084_, new_n42083_, new_n42079_ );
nor  ( new_n42085_, new_n42084_, new_n42078_ );
nand ( new_n42086_, new_n42085_, new_n42067_ );
and  ( new_n42087_, new_n42086_, new_n42066_ );
xnor ( new_n42088_, new_n41973_, new_n41967_ );
xor  ( new_n42089_, new_n42088_, new_n41979_ );
nor  ( new_n42090_, new_n42089_, new_n42087_ );
and  ( new_n42091_, new_n42089_, new_n42087_ );
xor  ( new_n42092_, new_n42027_, new_n42011_ );
xnor ( new_n42093_, new_n42092_, new_n42043_ );
nor  ( new_n42094_, new_n42093_, new_n42091_ );
or   ( new_n42095_, new_n42094_, new_n42090_ );
xnor ( new_n42096_, new_n42045_, new_n42009_ );
xor  ( new_n42097_, new_n42096_, new_n42049_ );
nand ( new_n42098_, new_n42097_, new_n42095_ );
xnor ( new_n42099_, new_n42053_, new_n42051_ );
xor  ( new_n42100_, new_n42099_, new_n42056_ );
nor  ( new_n42101_, new_n42100_, new_n42098_ );
xor  ( new_n42102_, new_n42089_, new_n42087_ );
xor  ( new_n42103_, new_n42102_, new_n42093_ );
or   ( new_n42104_, new_n8264_, new_n31952_ );
or   ( new_n42105_, new_n8266_, new_n31654_ );
and  ( new_n42106_, new_n42105_, new_n42104_ );
xor  ( new_n42107_, new_n42106_, new_n7724_ );
xnor ( new_n42108_, new_n42077_, new_n42071_ );
xor  ( new_n42109_, new_n42108_, new_n42083_ );
or   ( new_n42110_, new_n42109_, new_n42107_ );
xor  ( new_n42111_, new_n42039_, new_n42033_ );
xor  ( new_n42112_, new_n42111_, new_n7177_ );
or   ( new_n42113_, new_n42112_, new_n42110_ );
and  ( new_n42114_, new_n42112_, new_n42110_ );
or   ( new_n42115_, new_n8874_, new_n31333_ );
or   ( new_n42116_, new_n8876_, new_n30798_ );
and  ( new_n42117_, new_n42116_, new_n42115_ );
xor  ( new_n42118_, new_n42117_, new_n8256_ );
or   ( new_n42119_, new_n9422_, new_n30798_ );
or   ( new_n42120_, new_n9424_, new_n30800_ );
and  ( new_n42121_, new_n42120_, new_n42119_ );
xor  ( new_n42122_, new_n42121_, new_n8873_ );
or   ( new_n42123_, new_n8874_, new_n31654_ );
or   ( new_n42124_, new_n8876_, new_n31333_ );
and  ( new_n42125_, new_n42124_, new_n42123_ );
xor  ( new_n42126_, new_n42125_, new_n8257_ );
nand ( new_n42127_, new_n42126_, new_n42122_ );
nor  ( new_n42128_, new_n42126_, new_n42122_ );
and  ( new_n42129_, new_n8040_, RIbb33378_192 );
nor  ( new_n42130_, new_n42129_, new_n7725_ );
and  ( new_n42131_, new_n42129_, new_n7722_ );
nor  ( new_n42132_, new_n42131_, new_n42130_ );
or   ( new_n42133_, new_n42132_, new_n42128_ );
and  ( new_n42134_, new_n42133_, new_n42127_ );
nor  ( new_n42135_, new_n42134_, new_n42118_ );
and  ( new_n42136_, new_n42134_, new_n42118_ );
or   ( new_n42137_, new_n10059_, new_n30227_ );
or   ( new_n42138_, new_n10061_, new_n30120_ );
and  ( new_n42139_, new_n42138_, new_n42137_ );
xor  ( new_n42140_, new_n42139_, new_n9421_ );
and  ( new_n42141_, RIbb32fb8_184, RIbb2d888_64 );
or   ( new_n42142_, new_n29619_, RIbb2d888_64 );
and  ( new_n42143_, new_n42142_, RIbb2d900_63 );
or   ( new_n42144_, new_n42143_, new_n42141_ );
or   ( new_n42145_, new_n10770_, new_n29474_ );
and  ( new_n42146_, new_n42145_, new_n42144_ );
nor  ( new_n42147_, new_n42146_, new_n42140_ );
and  ( new_n42148_, new_n42146_, new_n42140_ );
nor  ( new_n42149_, new_n42148_, new_n7724_ );
nor  ( new_n42150_, new_n42149_, new_n42147_ );
not  ( new_n42151_, new_n42150_ );
nor  ( new_n42152_, new_n42151_, new_n42136_ );
nor  ( new_n42153_, new_n42152_, new_n42135_ );
or   ( new_n42154_, new_n42153_, new_n42114_ );
and  ( new_n42155_, new_n42154_, new_n42113_ );
nor  ( new_n42156_, new_n42155_, new_n42103_ );
xor  ( new_n42157_, new_n42097_, new_n42095_ );
and  ( new_n42158_, new_n42157_, new_n42156_ );
xor  ( new_n42159_, new_n42065_, new_n42063_ );
xor  ( new_n42160_, new_n42159_, new_n42085_ );
xnor ( new_n42161_, new_n42112_, new_n42110_ );
xor  ( new_n42162_, new_n42161_, new_n42153_ );
and  ( new_n42163_, new_n42162_, new_n42160_ );
xor  ( new_n42164_, new_n42155_, new_n42103_ );
and  ( new_n42165_, new_n42164_, new_n42163_ );
xor  ( new_n42166_, new_n42162_, new_n42160_ );
xor  ( new_n42167_, new_n42109_, new_n42107_ );
xor  ( new_n42168_, new_n42146_, new_n42140_ );
xor  ( new_n42169_, new_n42168_, new_n7724_ );
or   ( new_n42170_, new_n10059_, new_n30800_ );
or   ( new_n42171_, new_n10061_, new_n30227_ );
and  ( new_n42172_, new_n42171_, new_n42170_ );
xor  ( new_n42173_, new_n42172_, new_n9421_ );
and  ( new_n42174_, RIbb33030_185, RIbb2d888_64 );
or   ( new_n42175_, new_n30120_, RIbb2d888_64 );
and  ( new_n42176_, new_n42175_, RIbb2d900_63 );
or   ( new_n42177_, new_n42176_, new_n42174_ );
or   ( new_n42178_, new_n10770_, new_n29619_ );
and  ( new_n42179_, new_n42178_, new_n42177_ );
or   ( new_n42180_, new_n42179_, new_n42173_ );
and  ( new_n42181_, new_n42179_, new_n42173_ );
or   ( new_n42182_, new_n9422_, new_n31333_ );
or   ( new_n42183_, new_n9424_, new_n30798_ );
and  ( new_n42184_, new_n42183_, new_n42182_ );
xor  ( new_n42185_, new_n42184_, new_n8873_ );
or   ( new_n42186_, new_n42185_, new_n42181_ );
and  ( new_n42187_, new_n42186_, new_n42180_ );
or   ( new_n42188_, new_n42187_, new_n42169_ );
and  ( new_n42189_, new_n42187_, new_n42169_ );
xor  ( new_n42190_, new_n42126_, new_n42122_ );
xnor ( new_n42191_, new_n42190_, new_n42132_ );
or   ( new_n42192_, new_n42191_, new_n42189_ );
and  ( new_n42193_, new_n42192_, new_n42188_ );
or   ( new_n42194_, new_n42193_, new_n42167_ );
and  ( new_n42195_, new_n42193_, new_n42167_ );
xor  ( new_n42196_, new_n42134_, new_n42118_ );
xor  ( new_n42197_, new_n42196_, new_n42150_ );
or   ( new_n42198_, new_n42197_, new_n42195_ );
and  ( new_n42199_, new_n42198_, new_n42194_ );
and  ( new_n42200_, new_n42199_, new_n42166_ );
or   ( new_n42201_, new_n9422_, new_n31654_ );
or   ( new_n42202_, new_n9424_, new_n31333_ );
and  ( new_n42203_, new_n42202_, new_n42201_ );
xor  ( new_n42204_, new_n42203_, new_n8873_ );
not  ( new_n42205_, new_n42204_ );
and  ( new_n42206_, new_n8649_, RIbb33378_192 );
or   ( new_n42207_, new_n42206_, new_n8257_ );
nand ( new_n42208_, new_n42206_, new_n8254_ );
and  ( new_n42209_, new_n42208_, new_n42207_ );
nor  ( new_n42210_, new_n42209_, new_n42205_ );
or   ( new_n42211_, new_n8874_, new_n31952_ );
or   ( new_n42212_, new_n8876_, new_n31654_ );
and  ( new_n42213_, new_n42212_, new_n42211_ );
xor  ( new_n42214_, new_n42213_, new_n8257_ );
nor  ( new_n42215_, new_n42214_, new_n42210_ );
or   ( new_n42216_, new_n10059_, new_n30798_ );
or   ( new_n42217_, new_n10061_, new_n30800_ );
and  ( new_n42218_, new_n42217_, new_n42216_ );
xor  ( new_n42219_, new_n42218_, new_n9421_ );
and  ( new_n42220_, RIbb330a8_186, RIbb2d888_64 );
or   ( new_n42221_, new_n30227_, RIbb2d888_64 );
and  ( new_n42222_, new_n42221_, RIbb2d900_63 );
or   ( new_n42223_, new_n42222_, new_n42220_ );
or   ( new_n42224_, new_n10770_, new_n30120_ );
and  ( new_n42225_, new_n42224_, new_n42223_ );
nor  ( new_n42226_, new_n42225_, new_n42219_ );
and  ( new_n42227_, new_n42225_, new_n42219_ );
nor  ( new_n42228_, new_n42227_, new_n8256_ );
nor  ( new_n42229_, new_n42228_, new_n42226_ );
and  ( new_n42230_, new_n42214_, new_n42210_ );
nor  ( new_n42231_, new_n42230_, new_n42229_ );
or   ( new_n42232_, new_n42231_, new_n42215_ );
xnor ( new_n42233_, new_n42187_, new_n42169_ );
xor  ( new_n42234_, new_n42233_, new_n42191_ );
or   ( new_n42235_, new_n42234_, new_n42232_ );
xnor ( new_n42236_, new_n42193_, new_n42167_ );
xor  ( new_n42237_, new_n42236_, new_n42197_ );
nor  ( new_n42238_, new_n42237_, new_n42235_ );
xor  ( new_n42239_, new_n42179_, new_n42173_ );
xor  ( new_n42240_, new_n42239_, new_n42185_ );
xor  ( new_n42241_, new_n42214_, new_n42210_ );
xor  ( new_n42242_, new_n42241_, new_n42229_ );
and  ( new_n42243_, new_n42242_, new_n42240_ );
xor  ( new_n42244_, new_n42234_, new_n42232_ );
and  ( new_n42245_, new_n42244_, new_n42243_ );
xor  ( new_n42246_, new_n42242_, new_n42240_ );
xor  ( new_n42247_, new_n42225_, new_n42219_ );
xor  ( new_n42248_, new_n42247_, new_n8256_ );
or   ( new_n42249_, new_n10059_, new_n31333_ );
or   ( new_n42250_, new_n10061_, new_n30798_ );
and  ( new_n42251_, new_n42250_, new_n42249_ );
xor  ( new_n42252_, new_n42251_, new_n9421_ );
and  ( new_n42253_, RIbb33120_187, RIbb2d888_64 );
or   ( new_n42254_, new_n30800_, RIbb2d888_64 );
and  ( new_n42255_, new_n42254_, RIbb2d900_63 );
or   ( new_n42256_, new_n42255_, new_n42253_ );
or   ( new_n42257_, new_n10770_, new_n30227_ );
and  ( new_n42258_, new_n42257_, new_n42256_ );
or   ( new_n42259_, new_n42258_, new_n42252_ );
and  ( new_n42260_, new_n42258_, new_n42252_ );
or   ( new_n42261_, new_n9422_, new_n31952_ );
or   ( new_n42262_, new_n9424_, new_n31654_ );
and  ( new_n42263_, new_n42262_, new_n42261_ );
xor  ( new_n42264_, new_n42263_, new_n8873_ );
or   ( new_n42265_, new_n42264_, new_n42260_ );
and  ( new_n42266_, new_n42265_, new_n42259_ );
or   ( new_n42267_, new_n42266_, new_n42248_ );
and  ( new_n42268_, new_n42266_, new_n42248_ );
xor  ( new_n42269_, new_n42209_, new_n42205_ );
or   ( new_n42270_, new_n42269_, new_n42268_ );
and  ( new_n42271_, new_n42270_, new_n42267_ );
and  ( new_n42272_, new_n42271_, new_n42246_ );
or   ( new_n42273_, new_n10059_, new_n31654_ );
or   ( new_n42274_, new_n10061_, new_n31333_ );
and  ( new_n42275_, new_n42274_, new_n42273_ );
xor  ( new_n42276_, new_n42275_, new_n9421_ );
and  ( new_n42277_, RIbb33198_188, RIbb2d888_64 );
or   ( new_n42278_, new_n30798_, RIbb2d888_64 );
and  ( new_n42279_, new_n42278_, RIbb2d900_63 );
or   ( new_n42280_, new_n42279_, new_n42277_ );
or   ( new_n42281_, new_n10770_, new_n30800_ );
and  ( new_n42282_, new_n42281_, new_n42280_ );
nor  ( new_n42283_, new_n42282_, new_n42276_ );
nand ( new_n42284_, new_n42282_, new_n42276_ );
and  ( new_n42285_, new_n42284_, new_n8873_ );
or   ( new_n42286_, new_n42285_, new_n42283_ );
xnor ( new_n42287_, new_n42258_, new_n42252_ );
xor  ( new_n42288_, new_n42287_, new_n42264_ );
or   ( new_n42289_, new_n42288_, new_n42286_ );
xnor ( new_n42290_, new_n42266_, new_n42248_ );
xor  ( new_n42291_, new_n42290_, new_n42269_ );
nor  ( new_n42292_, new_n42291_, new_n42289_ );
and  ( new_n42293_, new_n9185_, RIbb33378_192 );
or   ( new_n42294_, new_n42293_, new_n8873_ );
nand ( new_n42295_, new_n42293_, new_n8870_ );
and  ( new_n42296_, new_n42295_, new_n42294_ );
xor  ( new_n42297_, new_n42282_, new_n42276_ );
xor  ( new_n42298_, new_n42297_, new_n8873_ );
nor  ( new_n42299_, new_n42298_, new_n42296_ );
xor  ( new_n42300_, new_n42288_, new_n42286_ );
and  ( new_n42301_, new_n42300_, new_n42299_ );
or   ( new_n42302_, new_n10059_, new_n31952_ );
or   ( new_n42303_, new_n10061_, new_n31654_ );
and  ( new_n42304_, new_n42303_, new_n42302_ );
xor  ( new_n42305_, new_n42304_, new_n9421_ );
and  ( new_n42306_, RIbb33210_189, RIbb2d888_64 );
or   ( new_n42307_, new_n31333_, RIbb2d888_64 );
and  ( new_n42308_, new_n42307_, RIbb2d900_63 );
or   ( new_n42309_, new_n42308_, new_n42306_ );
or   ( new_n42310_, new_n10770_, new_n30798_ );
and  ( new_n42311_, new_n42310_, new_n42309_ );
and  ( new_n42312_, new_n42311_, new_n42305_ );
xor  ( new_n42313_, new_n42298_, new_n42296_ );
and  ( new_n42314_, new_n42313_, new_n42312_ );
and  ( new_n42315_, RIbb33288_190, RIbb2d888_64 );
or   ( new_n42316_, new_n31654_, RIbb2d888_64 );
and  ( new_n42317_, new_n42316_, RIbb2d900_63 );
or   ( new_n42318_, new_n42317_, new_n42315_ );
or   ( new_n42319_, new_n10770_, new_n31333_ );
and  ( new_n42320_, new_n42319_, new_n42318_ );
and  ( new_n42321_, new_n42320_, new_n9420_ );
xor  ( new_n42322_, new_n42311_, new_n42305_ );
and  ( new_n42323_, new_n42322_, new_n42321_ );
xor  ( new_n42324_, new_n42320_, new_n9421_ );
and  ( new_n42325_, new_n9738_, RIbb33378_192 );
or   ( new_n42326_, new_n42325_, new_n9421_ );
nand ( new_n42327_, new_n42325_, new_n9418_ );
and  ( new_n42328_, new_n42327_, new_n42326_ );
nor  ( new_n42329_, new_n42328_, new_n42324_ );
and  ( new_n42330_, RIbb33378_192, RIbb2d888_64 );
nor  ( new_n42331_, new_n42330_, new_n10052_ );
and  ( new_n42332_, RIbb33300_191, RIbb2d888_64 );
or   ( new_n42333_, new_n31952_, RIbb2d888_64 );
and  ( new_n42334_, new_n42333_, RIbb2d900_63 );
or   ( new_n42335_, new_n42334_, new_n42332_ );
or   ( new_n42336_, new_n10770_, new_n31654_ );
and  ( new_n42337_, new_n42336_, new_n42335_ );
and  ( new_n42338_, new_n42337_, new_n42331_ );
xor  ( new_n42339_, new_n42328_, new_n42324_ );
and  ( new_n42340_, new_n42339_, new_n42338_ );
nor  ( new_n42341_, new_n42340_, new_n42329_ );
not  ( new_n42342_, new_n42341_ );
xor  ( new_n42343_, new_n42322_, new_n42321_ );
and  ( new_n42344_, new_n42343_, new_n42342_ );
nor  ( new_n42345_, new_n42344_, new_n42323_ );
not  ( new_n42346_, new_n42345_ );
xor  ( new_n42347_, new_n42313_, new_n42312_ );
and  ( new_n42348_, new_n42347_, new_n42346_ );
nor  ( new_n42349_, new_n42348_, new_n42314_ );
not  ( new_n42350_, new_n42349_ );
xor  ( new_n42351_, new_n42300_, new_n42299_ );
and  ( new_n42352_, new_n42351_, new_n42350_ );
nor  ( new_n42353_, new_n42352_, new_n42301_ );
not  ( new_n42354_, new_n42353_ );
xor  ( new_n42355_, new_n42291_, new_n42289_ );
and  ( new_n42356_, new_n42355_, new_n42354_ );
nor  ( new_n42357_, new_n42356_, new_n42292_ );
not  ( new_n42358_, new_n42357_ );
xor  ( new_n42359_, new_n42271_, new_n42246_ );
and  ( new_n42360_, new_n42359_, new_n42358_ );
nor  ( new_n42361_, new_n42360_, new_n42272_ );
not  ( new_n42362_, new_n42361_ );
xor  ( new_n42363_, new_n42244_, new_n42243_ );
and  ( new_n42364_, new_n42363_, new_n42362_ );
nor  ( new_n42365_, new_n42364_, new_n42245_ );
not  ( new_n42366_, new_n42365_ );
xor  ( new_n42367_, new_n42237_, new_n42235_ );
and  ( new_n42368_, new_n42367_, new_n42366_ );
or   ( new_n42369_, new_n42368_, new_n42238_ );
xor  ( new_n42370_, new_n42199_, new_n42166_ );
and  ( new_n42371_, new_n42370_, new_n42369_ );
or   ( new_n42372_, new_n42371_, new_n42200_ );
xor  ( new_n42373_, new_n42164_, new_n42163_ );
and  ( new_n42374_, new_n42373_, new_n42372_ );
or   ( new_n42375_, new_n42374_, new_n42165_ );
xor  ( new_n42376_, new_n42157_, new_n42156_ );
and  ( new_n42377_, new_n42376_, new_n42375_ );
or   ( new_n42378_, new_n42377_, new_n42158_ );
xor  ( new_n42379_, new_n42100_, new_n42098_ );
and  ( new_n42380_, new_n42379_, new_n42378_ );
or   ( new_n42381_, new_n42380_, new_n42101_ );
xor  ( new_n42382_, new_n42058_, new_n42007_ );
and  ( new_n42383_, new_n42382_, new_n42381_ );
or   ( new_n42384_, new_n42383_, new_n42059_ );
xor  ( new_n42385_, new_n42004_, new_n42002_ );
and  ( new_n42386_, new_n42385_, new_n42384_ );
or   ( new_n42387_, new_n42386_, new_n42005_ );
xor  ( new_n42388_, new_n41929_, new_n41876_ );
and  ( new_n42389_, new_n42388_, new_n42387_ );
or   ( new_n42390_, new_n42389_, new_n41930_ );
xor  ( new_n42391_, new_n41873_, new_n41815_ );
and  ( new_n42392_, new_n42391_, new_n42390_ );
or   ( new_n42393_, new_n42392_, new_n41874_ );
xor  ( new_n42394_, new_n41813_, new_n41812_ );
and  ( new_n42395_, new_n42394_, new_n42393_ );
or   ( new_n42396_, new_n42395_, new_n41814_ );
xor  ( new_n42397_, new_n41806_, new_n41804_ );
and  ( new_n42398_, new_n42397_, new_n42396_ );
or   ( new_n42399_, new_n42398_, new_n41807_ );
xor  ( new_n42400_, new_n41722_, new_n41640_ );
and  ( new_n42401_, new_n42400_, new_n42399_ );
or   ( new_n42402_, new_n42401_, new_n41723_ );
xor  ( new_n42403_, new_n41637_, new_n41544_ );
and  ( new_n42404_, new_n42403_, new_n42402_ );
or   ( new_n42405_, new_n42404_, new_n41638_ );
xor  ( new_n42406_, new_n41541_, new_n41452_ );
and  ( new_n42407_, new_n42406_, new_n42405_ );
or   ( new_n42408_, new_n42407_, new_n41542_ );
xor  ( new_n42409_, new_n41449_, new_n41359_ );
and  ( new_n42410_, new_n42409_, new_n42408_ );
or   ( new_n42411_, new_n42410_, new_n41450_ );
xor  ( new_n42412_, new_n41356_, new_n41354_ );
and  ( new_n42413_, new_n42412_, new_n42411_ );
or   ( new_n42414_, new_n42413_, new_n41357_ );
xor  ( new_n42415_, new_n41266_, new_n41149_ );
and  ( new_n42416_, new_n42415_, new_n42414_ );
or   ( new_n42417_, new_n42416_, new_n41267_ );
xor  ( new_n42418_, new_n41146_, new_n41049_ );
and  ( new_n42419_, new_n42418_, new_n42417_ );
or   ( new_n42420_, new_n42419_, new_n41147_ );
xor  ( new_n42421_, new_n41047_, new_n41046_ );
and  ( new_n42422_, new_n42421_, new_n42420_ );
or   ( new_n42423_, new_n42422_, new_n41048_ );
xor  ( new_n42424_, new_n41040_, new_n41038_ );
and  ( new_n42425_, new_n42424_, new_n42423_ );
or   ( new_n42426_, new_n42425_, new_n41041_ );
xor  ( new_n42427_, new_n40923_, new_n40800_ );
and  ( new_n42428_, new_n42427_, new_n42426_ );
or   ( new_n42429_, new_n42428_, new_n40924_ );
xor  ( new_n42430_, new_n40797_, new_n40655_ );
and  ( new_n42431_, new_n42430_, new_n42429_ );
or   ( new_n42432_, new_n42431_, new_n40798_ );
xor  ( new_n42433_, new_n40652_, new_n40530_ );
and  ( new_n42434_, new_n42433_, new_n42432_ );
or   ( new_n42435_, new_n42434_, new_n40653_ );
xor  ( new_n42436_, new_n40527_, new_n40383_ );
and  ( new_n42437_, new_n42436_, new_n42435_ );
or   ( new_n42438_, new_n42437_, new_n40528_ );
xor  ( new_n42439_, new_n40380_, new_n40254_ );
and  ( new_n42440_, new_n42439_, new_n42438_ );
or   ( new_n42441_, new_n42440_, new_n40381_ );
xor  ( new_n42442_, new_n40251_, new_n40114_ );
and  ( new_n42443_, new_n42442_, new_n42441_ );
or   ( new_n42444_, new_n42443_, new_n40252_ );
xor  ( new_n42445_, new_n40111_, new_n40109_ );
and  ( new_n42446_, new_n42445_, new_n42444_ );
or   ( new_n42447_, new_n42446_, new_n40112_ );
xor  ( new_n42448_, new_n39942_, new_n39791_ );
and  ( new_n42449_, new_n42448_, new_n42447_ );
or   ( new_n42450_, new_n42449_, new_n39943_ );
xor  ( new_n42451_, new_n39788_, new_n39647_ );
and  ( new_n42452_, new_n42451_, new_n42450_ );
or   ( new_n42453_, new_n42452_, new_n39789_ );
xor  ( new_n42454_, new_n39644_, new_n39468_ );
and  ( new_n42455_, new_n42454_, new_n42453_ );
or   ( new_n42456_, new_n42455_, new_n39645_ );
xor  ( new_n42457_, new_n39466_, new_n39465_ );
and  ( new_n42458_, new_n42457_, new_n42456_ );
or   ( new_n42459_, new_n42458_, new_n39467_ );
xor  ( new_n42460_, new_n39459_, new_n39458_ );
and  ( new_n42461_, new_n42460_, new_n42459_ );
or   ( new_n42462_, new_n42461_, new_n39460_ );
xor  ( new_n42463_, new_n39278_, new_n39276_ );
and  ( new_n42464_, new_n42463_, new_n42462_ );
or   ( new_n42465_, new_n42464_, new_n39279_ );
xor  ( new_n42466_, new_n39100_, new_n38908_ );
and  ( new_n42467_, new_n42466_, new_n42465_ );
or   ( new_n42468_, new_n42467_, new_n39101_ );
xor  ( new_n42469_, new_n38906_, new_n38904_ );
and  ( new_n42470_, new_n42469_, new_n42468_ );
or   ( new_n42471_, new_n42470_, new_n38907_ );
xor  ( new_n42472_, new_n38710_, new_n38523_ );
and  ( new_n42473_, new_n42472_, new_n42471_ );
or   ( new_n42474_, new_n42473_, new_n38711_ );
xor  ( new_n42475_, new_n38520_, new_n38308_ );
and  ( new_n42476_, new_n42475_, new_n42474_ );
or   ( new_n42477_, new_n42476_, new_n38521_ );
xor  ( new_n42478_, new_n38305_, new_n38106_ );
and  ( new_n42479_, new_n42478_, new_n42477_ );
or   ( new_n42480_, new_n42479_, new_n38306_ );
xor  ( new_n42481_, new_n38103_, new_n37907_ );
and  ( new_n42482_, new_n42481_, new_n42480_ );
or   ( new_n42483_, new_n42482_, new_n38104_ );
xor  ( new_n42484_, new_n37904_, new_n37693_ );
and  ( new_n42485_, new_n42484_, new_n42483_ );
or   ( new_n42486_, new_n42485_, new_n37905_ );
xor  ( new_n42487_, new_n37690_, new_n37477_ );
and  ( new_n42488_, new_n42487_, new_n42486_ );
or   ( new_n42489_, new_n42488_, new_n37691_ );
xor  ( new_n42490_, new_n37474_, new_n37472_ );
and  ( new_n42491_, new_n42490_, new_n42489_ );
or   ( new_n42492_, new_n42491_, new_n37475_ );
xor  ( new_n42493_, new_n37240_, new_n37004_ );
and  ( new_n42494_, new_n42493_, new_n42492_ );
or   ( new_n42495_, new_n42494_, new_n37241_ );
xor  ( new_n42496_, new_n37001_, new_n36778_ );
and  ( new_n42497_, new_n42496_, new_n42495_ );
or   ( new_n42498_, new_n42497_, new_n37002_ );
xor  ( new_n42499_, new_n36775_, new_n36551_ );
and  ( new_n42500_, new_n42499_, new_n42498_ );
or   ( new_n42501_, new_n42500_, new_n36776_ );
xor  ( new_n42502_, new_n36548_, new_n36297_ );
and  ( new_n42503_, new_n42502_, new_n42501_ );
or   ( new_n42504_, new_n42503_, new_n36549_ );
xor  ( new_n42505_, new_n36294_, new_n36063_ );
and  ( new_n42506_, new_n42505_, new_n42504_ );
or   ( new_n42507_, new_n42506_, new_n36295_ );
xor  ( new_n42508_, new_n36060_, new_n35813_ );
and  ( new_n42509_, new_n42508_, new_n42507_ );
or   ( new_n42510_, new_n42509_, new_n36061_ );
xor  ( new_n42511_, new_n35811_, new_n35810_ );
and  ( new_n42512_, new_n42511_, new_n42510_ );
or   ( new_n42513_, new_n42512_, new_n35812_ );
xor  ( new_n42514_, new_n35804_, new_n35803_ );
and  ( new_n42515_, new_n42514_, new_n42513_ );
or   ( new_n42516_, new_n42515_, new_n35805_ );
xor  ( new_n42517_, new_n35535_, new_n35534_ );
and  ( new_n42518_, new_n42517_, new_n42516_ );
or   ( new_n42519_, new_n42518_, new_n35536_ );
xor  ( new_n42520_, new_n35267_, new_n35265_ );
and  ( new_n42521_, new_n42520_, new_n42519_ );
or   ( new_n42522_, new_n42521_, new_n35268_ );
xor  ( new_n42523_, new_n34996_, new_n34718_ );
and  ( new_n42524_, new_n42523_, new_n42522_ );
nor  ( new_n42525_, new_n42524_, new_n34997_ );
not  ( new_n42526_, new_n42525_ );
xor  ( new_n42527_, new_n34716_, new_n34715_ );
and  ( new_n42528_, new_n42527_, new_n42526_ );
or   ( new_n42529_, new_n42528_, new_n34717_ );
xor  ( new_n42530_, new_n34438_, new_n34436_ );
and  ( new_n42531_, new_n42530_, new_n42529_ );
or   ( new_n42532_, new_n42531_, new_n34439_ );
xor  ( new_n42533_, new_n34164_, new_n33859_ );
and  ( new_n42534_, new_n42533_, new_n42532_ );
or   ( new_n42535_, new_n42534_, new_n34165_ );
xor  ( new_n42536_, new_n33857_, new_n33855_ );
and  ( new_n42537_, new_n42536_, new_n42535_ );
or   ( new_n42538_, new_n42537_, new_n33858_ );
xor  ( new_n42539_, new_n33574_, new_n33288_ );
and  ( new_n42540_, new_n42539_, new_n42538_ );
or   ( new_n42541_, new_n42540_, new_n33575_ );
xor  ( new_n42542_, new_n33285_, new_n32969_ );
and  ( new_n42543_, new_n42542_, new_n42541_ );
nor  ( new_n42544_, new_n42543_, new_n33286_ );
not  ( new_n42545_, new_n42544_ );
xor  ( new_n42546_, new_n32966_, new_n32664_ );
and  ( new_n42547_, new_n42546_, new_n42545_ );
or   ( new_n42548_, new_n42547_, new_n32967_ );
xor  ( new_n42549_, new_n32661_, new_n32344_ );
and  ( new_n42550_, new_n42549_, new_n42548_ );
nor  ( new_n42551_, new_n42550_, new_n32662_ );
not  ( new_n42552_, new_n42551_ );
xor  ( new_n42553_, new_n32341_, new_n32021_ );
and  ( new_n42554_, new_n42553_, new_n42552_ );
or   ( new_n42555_, new_n42554_, new_n32342_ );
xor  ( new_n42556_, new_n32018_, new_n31708_ );
and  ( new_n42557_, new_n42556_, new_n42555_ );
or   ( new_n42558_, new_n42557_, new_n32019_ );
xor  ( new_n42559_, new_n31705_, new_n31398_ );
and  ( new_n42560_, new_n42559_, new_n42558_ );
or   ( new_n42561_, new_n42560_, new_n31706_ );
xor  ( new_n42562_, new_n31396_, new_n31394_ );
and  ( new_n42563_, new_n42562_, new_n42561_ );
or   ( new_n42564_, new_n42563_, new_n31397_ );
xor  ( new_n42565_, new_n31079_, new_n30767_ );
and  ( new_n42566_, new_n42565_, new_n42564_ );
or   ( new_n42567_, new_n42566_, new_n31080_ );
xor  ( new_n42568_, new_n30765_, new_n30764_ );
and  ( new_n42569_, new_n42568_, new_n42567_ );
nor  ( new_n42570_, new_n42569_, new_n30766_ );
not  ( new_n42571_, new_n42570_ );
xor  ( new_n42572_, new_n30459_, new_n30457_ );
and  ( new_n42573_, new_n42572_, new_n42571_ );
nor  ( new_n42574_, new_n42573_, new_n30460_ );
not  ( new_n42575_, new_n42574_ );
xor  ( new_n42576_, new_n30170_, new_n29875_ );
and  ( new_n42577_, new_n42576_, new_n42575_ );
nor  ( new_n42578_, new_n42577_, new_n30171_ );
not  ( new_n42579_, new_n42578_ );
xor  ( new_n42580_, new_n29873_, new_n29872_ );
and  ( new_n42581_, new_n42580_, new_n42579_ );
or   ( new_n42582_, new_n42581_, new_n29874_ );
xor  ( new_n42583_, new_n29588_, new_n29587_ );
and  ( new_n42584_, new_n42583_, new_n42582_ );
or   ( new_n42585_, new_n42584_, new_n29589_ );
xor  ( new_n42586_, new_n29310_, new_n29309_ );
and  ( new_n42587_, new_n42586_, new_n42585_ );
or   ( new_n42588_, new_n42587_, new_n29311_ );
xor  ( new_n42589_, new_n29021_, new_n29020_ );
and  ( new_n42590_, new_n42589_, new_n42588_ );
or   ( new_n42591_, new_n42590_, new_n29022_ );
xor  ( new_n42592_, new_n28761_, new_n28760_ );
and  ( new_n42593_, new_n42592_, new_n42591_ );
nor  ( new_n42594_, new_n42593_, new_n28762_ );
not  ( new_n42595_, new_n42594_ );
xor  ( new_n42596_, new_n28500_, new_n28499_ );
and  ( new_n42597_, new_n42596_, new_n42595_ );
or   ( new_n42598_, new_n42597_, new_n28501_ );
xor  ( new_n42599_, new_n28244_, new_n28243_ );
and  ( new_n42600_, new_n42599_, new_n42598_ );
or   ( new_n42601_, new_n42600_, new_n28245_ );
xor  ( new_n42602_, new_n27983_, new_n27982_ );
and  ( new_n42603_, new_n42602_, new_n42601_ );
nor  ( new_n42604_, new_n42603_, new_n27984_ );
not  ( new_n42605_, new_n42604_ );
xor  ( new_n42606_, new_n27727_, new_n27726_ );
and  ( new_n42607_, new_n42606_, new_n42605_ );
or   ( new_n42608_, new_n42607_, new_n27728_ );
xor  ( new_n42609_, new_n27474_, new_n27473_ );
and  ( new_n42610_, new_n42609_, new_n42608_ );
or   ( new_n42611_, new_n42610_, new_n27475_ );
xor  ( new_n42612_, new_n27222_, new_n27221_ );
and  ( new_n42613_, new_n42612_, new_n42611_ );
or   ( new_n42614_, new_n42613_, new_n27223_ );
xor  ( new_n42615_, new_n26974_, new_n26973_ );
and  ( new_n42616_, new_n42615_, new_n42614_ );
nor  ( new_n42617_, new_n42616_, new_n26975_ );
not  ( new_n42618_, new_n42617_ );
xor  ( new_n42619_, new_n26730_, new_n26729_ );
and  ( new_n42620_, new_n42619_, new_n42618_ );
or   ( new_n42621_, new_n42620_, new_n26731_ );
xor  ( new_n42622_, new_n26503_, new_n26501_ );
and  ( new_n42623_, new_n42622_, new_n42621_ );
or   ( new_n42624_, new_n42623_, new_n26504_ );
xor  ( new_n42625_, new_n26264_, new_n25846_ );
and  ( new_n42626_, new_n42625_, new_n42624_ );
nor  ( new_n42627_, new_n42626_, new_n26265_ );
not  ( new_n42628_, new_n42627_ );
xor  ( new_n42629_, new_n25843_, new_n25644_ );
and  ( new_n42630_, new_n42629_, new_n42628_ );
or   ( new_n42631_, new_n42630_, new_n25844_ );
xor  ( new_n42632_, new_n25641_, new_n25437_ );
and  ( new_n42633_, new_n42632_, new_n42631_ );
nor  ( new_n42634_, new_n42633_, new_n25642_ );
not  ( new_n42635_, new_n42634_ );
xor  ( new_n42636_, new_n25435_, new_n25434_ );
and  ( new_n42637_, new_n42636_, new_n42635_ );
nor  ( new_n42638_, new_n42637_, new_n25436_ );
not  ( new_n42639_, new_n42638_ );
xor  ( new_n42640_, new_n25229_, new_n25228_ );
and  ( new_n42641_, new_n42640_, new_n42639_ );
or   ( new_n42642_, new_n42641_, new_n25230_ );
xor  ( new_n42643_, new_n25033_, new_n25032_ );
and  ( new_n42644_, new_n42643_, new_n42642_ );
nor  ( new_n42645_, new_n42644_, new_n25034_ );
not  ( new_n42646_, new_n42645_ );
xor  ( new_n42647_, new_n24840_, new_n24839_ );
and  ( new_n42648_, new_n42647_, new_n42646_ );
or   ( new_n42649_, new_n42648_, new_n24841_ );
xor  ( new_n42650_, new_n24666_, new_n24665_ );
and  ( new_n42651_, new_n42650_, new_n42649_ );
or   ( new_n42652_, new_n42651_, new_n24667_ );
xor  ( new_n42653_, new_n24489_, new_n24488_ );
and  ( new_n42654_, new_n42653_, new_n42652_ );
nor  ( new_n42655_, new_n42654_, new_n24490_ );
not  ( new_n42656_, new_n42655_ );
xor  ( new_n42657_, new_n24323_, new_n24322_ );
and  ( new_n42658_, new_n42657_, new_n42656_ );
nor  ( new_n42659_, new_n42658_, new_n24324_ );
not  ( new_n42660_, new_n42659_ );
xor  ( new_n42661_, new_n24153_, new_n24152_ );
and  ( new_n42662_, new_n42661_, new_n42660_ );
or   ( new_n42663_, new_n42662_, new_n24154_ );
xor  ( new_n42664_, new_n23987_, new_n23986_ );
and  ( new_n42665_, new_n42664_, new_n42663_ );
nor  ( new_n42666_, new_n42665_, new_n23988_ );
not  ( new_n42667_, new_n42666_ );
xor  ( new_n42668_, new_n23823_, new_n23822_ );
and  ( new_n42669_, new_n42668_, new_n42667_ );
nor  ( new_n42670_, new_n42669_, new_n23824_ );
not  ( new_n42671_, new_n42670_ );
xor  ( new_n42672_, new_n23663_, new_n23661_ );
and  ( new_n42673_, new_n42672_, new_n42671_ );
nor  ( new_n42674_, new_n42673_, new_n23664_ );
not  ( new_n42675_, new_n42674_ );
xor  ( new_n42676_, new_n23494_, new_n23227_ );
and  ( new_n42677_, new_n42676_, new_n42675_ );
nor  ( new_n42678_, new_n42677_, new_n23495_ );
not  ( new_n42679_, new_n42678_ );
xor  ( new_n42680_, new_n23224_, new_n23096_ );
and  ( new_n42681_, new_n42680_, new_n42679_ );
nor  ( new_n42682_, new_n42681_, new_n23225_ );
not  ( new_n42683_, new_n42682_ );
xor  ( new_n42684_, new_n23094_, new_n23093_ );
and  ( new_n42685_, new_n42684_, new_n42683_ );
nor  ( new_n42686_, new_n42685_, new_n23095_ );
not  ( new_n42687_, new_n42686_ );
xor  ( new_n42688_, new_n22966_, new_n22965_ );
and  ( new_n42689_, new_n42688_, new_n42687_ );
nor  ( new_n42690_, new_n42689_, new_n22967_ );
not  ( new_n42691_, new_n42690_ );
xor  ( new_n42692_, new_n22850_, new_n22849_ );
and  ( new_n42693_, new_n42692_, new_n42691_ );
or   ( new_n42694_, new_n42693_, new_n22851_ );
xor  ( new_n42695_, new_n22734_, new_n22733_ );
and  ( new_n42696_, new_n42695_, new_n42694_ );
nor  ( new_n42697_, new_n42696_, new_n22735_ );
not  ( new_n42698_, new_n42697_ );
xor  ( new_n42699_, new_n22622_, new_n22621_ );
and  ( new_n42700_, new_n42699_, new_n42698_ );
or   ( new_n42701_, new_n42700_, new_n22623_ );
xor  ( new_n42702_, new_n22509_, new_n22508_ );
and  ( new_n42703_, new_n42702_, new_n42701_ );
nor  ( new_n42704_, new_n42703_, new_n22510_ );
not  ( new_n42705_, new_n42704_ );
xor  ( new_n42706_, new_n22401_, new_n22399_ );
and  ( new_n42707_, new_n42706_, new_n42705_ );
nor  ( new_n42708_, new_n42707_, new_n22402_ );
not  ( new_n42709_, new_n42708_ );
xor  ( new_n42710_, new_n22294_, new_n22124_ );
and  ( new_n42711_, new_n42710_, new_n42709_ );
or   ( new_n42712_, new_n42711_, new_n22295_ );
xor  ( new_n42713_, new_n22122_, new_n22121_ );
and  ( new_n42714_, new_n42713_, new_n42712_ );
or   ( new_n42715_, new_n42714_, new_n22123_ );
xor  ( new_n42716_, new_n22049_, new_n22023_ );
and  ( new_n42717_, new_n42716_, new_n42715_ );
or   ( new_n42718_, new_n42717_, new_n22050_ );
nor  ( new_n42719_, new_n22048_, new_n22044_ );
and  ( new_n42720_, new_n22037_, new_n22035_ );
or   ( new_n42721_, new_n22037_, new_n22035_ );
and  ( new_n42722_, new_n22043_, new_n42721_ );
or   ( new_n42723_, new_n42722_, new_n42720_ );
xnor ( new_n42724_, new_n21724_, new_n21711_ );
xor  ( new_n42725_, new_n21772_, new_n21761_ );
xor  ( new_n42726_, new_n42725_, new_n21786_ );
xor  ( new_n42727_, new_n42726_, new_n42724_ );
or   ( new_n42728_, new_n22029_, new_n22025_ );
and  ( new_n42729_, new_n22029_, new_n22025_ );
or   ( new_n42730_, new_n22034_, new_n42729_ );
and  ( new_n42731_, new_n42730_, new_n42728_ );
xor  ( new_n42732_, new_n42731_, new_n42727_ );
xor  ( new_n42733_, new_n42732_, new_n42723_ );
xor  ( new_n42734_, new_n42733_, new_n42719_ );
xor  ( new_n42735_, new_n42734_, new_n42718_ );
xor  ( new_n42736_, new_n42716_, new_n42715_ );
xor  ( new_n42737_, new_n21608_, new_n21607_ );
xor  ( new_n42738_, new_n42713_, new_n42712_ );
or   ( new_n42739_, new_n42738_, new_n42737_ );
and  ( new_n42740_, new_n42738_, new_n42737_ );
xor  ( new_n42741_, new_n42706_, new_n42705_ );
xor  ( new_n42742_, new_n21597_, new_n21596_ );
xor  ( new_n42743_, new_n42702_, new_n42701_ );
nor  ( new_n42744_, new_n42743_, new_n42742_ );
and  ( new_n42745_, new_n42743_, new_n42742_ );
xor  ( new_n42746_, new_n42699_, new_n42698_ );
xor  ( new_n42747_, new_n21590_, new_n21589_ );
xor  ( new_n42748_, new_n42695_, new_n42694_ );
nor  ( new_n42749_, new_n42748_, new_n42747_ );
and  ( new_n42750_, new_n42748_, new_n42747_ );
xor  ( new_n42751_, new_n42668_, new_n42667_ );
xor  ( new_n42752_, new_n21559_, new_n21558_ );
xor  ( new_n42753_, new_n42664_, new_n42663_ );
nor  ( new_n42754_, new_n42753_, new_n42752_ );
and  ( new_n42755_, new_n42753_, new_n42752_ );
xor  ( new_n42756_, new_n42657_, new_n42656_ );
xor  ( new_n42757_, new_n21548_, new_n21547_ );
xor  ( new_n42758_, new_n42653_, new_n42652_ );
nor  ( new_n42759_, new_n42758_, new_n42757_ );
xor  ( new_n42760_, new_n21545_, new_n21544_ );
xor  ( new_n42761_, new_n42650_, new_n42649_ );
nor  ( new_n42762_, new_n42761_, new_n42760_ );
and  ( new_n42763_, new_n42761_, new_n42760_ );
xor  ( new_n42764_, new_n42647_, new_n42646_ );
xor  ( new_n42765_, new_n21538_, new_n21537_ );
xor  ( new_n42766_, new_n42643_, new_n42642_ );
nor  ( new_n42767_, new_n42766_, new_n42765_ );
and  ( new_n42768_, new_n42766_, new_n42765_ );
xor  ( new_n42769_, new_n42636_, new_n42635_ );
xor  ( new_n42770_, new_n21527_, new_n21526_ );
xor  ( new_n42771_, new_n42632_, new_n42631_ );
nor  ( new_n42772_, new_n42771_, new_n42770_ );
xor  ( new_n42773_, new_n21524_, new_n21523_ );
xor  ( new_n42774_, new_n42629_, new_n42628_ );
nor  ( new_n42775_, new_n42774_, new_n42773_ );
and  ( new_n42776_, new_n42774_, new_n42773_ );
xor  ( new_n42777_, new_n42625_, new_n42624_ );
xor  ( new_n42778_, new_n21516_, new_n21515_ );
xor  ( new_n42779_, new_n42622_, new_n42621_ );
or   ( new_n42780_, new_n42779_, new_n42778_ );
and  ( new_n42781_, new_n42779_, new_n42778_ );
xor  ( new_n42782_, new_n42619_, new_n42618_ );
xor  ( new_n42783_, new_n21509_, new_n21508_ );
xor  ( new_n42784_, new_n42615_, new_n42614_ );
nor  ( new_n42785_, new_n42784_, new_n42783_ );
xor  ( new_n42786_, new_n21506_, new_n21505_ );
xor  ( new_n42787_, new_n42612_, new_n42611_ );
nor  ( new_n42788_, new_n42787_, new_n42786_ );
xor  ( new_n42789_, new_n21503_, new_n21502_ );
xor  ( new_n42790_, new_n42609_, new_n42608_ );
nor  ( new_n42791_, new_n42790_, new_n42789_ );
and  ( new_n42792_, new_n42790_, new_n42789_ );
xor  ( new_n42793_, new_n42606_, new_n42605_ );
xor  ( new_n42794_, new_n21496_, new_n21495_ );
xor  ( new_n42795_, new_n42602_, new_n42601_ );
nor  ( new_n42796_, new_n42795_, new_n42794_ );
xor  ( new_n42797_, new_n21493_, new_n21492_ );
xor  ( new_n42798_, new_n42599_, new_n42598_ );
nor  ( new_n42799_, new_n42798_, new_n42797_ );
and  ( new_n42800_, new_n42798_, new_n42797_ );
xor  ( new_n42801_, new_n42596_, new_n42595_ );
xor  ( new_n42802_, new_n21486_, new_n21485_ );
xor  ( new_n42803_, new_n42592_, new_n42591_ );
nor  ( new_n42804_, new_n42803_, new_n42802_ );
xor  ( new_n42805_, new_n21483_, new_n21482_ );
xor  ( new_n42806_, new_n42589_, new_n42588_ );
nor  ( new_n42807_, new_n42806_, new_n42805_ );
xor  ( new_n42808_, new_n21480_, new_n21479_ );
xor  ( new_n42809_, new_n42586_, new_n42585_ );
nor  ( new_n42810_, new_n42809_, new_n42808_ );
xor  ( new_n42811_, new_n21477_, new_n21476_ );
xor  ( new_n42812_, new_n42583_, new_n42582_ );
nor  ( new_n42813_, new_n42812_, new_n42811_ );
and  ( new_n42814_, new_n42812_, new_n42811_ );
xor  ( new_n42815_, new_n42572_, new_n42571_ );
xor  ( new_n42816_, new_n21462_, new_n21461_ );
xor  ( new_n42817_, new_n42568_, new_n42567_ );
nor  ( new_n42818_, new_n42817_, new_n42816_ );
xor  ( new_n42819_, new_n21459_, new_n21458_ );
xor  ( new_n42820_, new_n42565_, new_n42564_ );
nor  ( new_n42821_, new_n42820_, new_n42819_ );
xor  ( new_n42822_, new_n21456_, new_n21455_ );
xor  ( new_n42823_, new_n42562_, new_n42561_ );
nor  ( new_n42824_, new_n42823_, new_n42822_ );
xor  ( new_n42825_, new_n21453_, new_n21452_ );
xor  ( new_n42826_, new_n42559_, new_n42558_ );
nor  ( new_n42827_, new_n42826_, new_n42825_ );
xor  ( new_n42828_, new_n21450_, new_n21449_ );
xor  ( new_n42829_, new_n42556_, new_n42555_ );
nor  ( new_n42830_, new_n42829_, new_n42828_ );
and  ( new_n42831_, new_n42829_, new_n42828_ );
xor  ( new_n42832_, new_n42553_, new_n42552_ );
xor  ( new_n42833_, new_n21443_, new_n21442_ );
xor  ( new_n42834_, new_n42549_, new_n42548_ );
nor  ( new_n42835_, new_n42834_, new_n42833_ );
and  ( new_n42836_, new_n42834_, new_n42833_ );
xor  ( new_n42837_, new_n42546_, new_n42545_ );
xor  ( new_n42838_, new_n21436_, new_n21435_ );
xor  ( new_n42839_, new_n42542_, new_n42541_ );
nor  ( new_n42840_, new_n42839_, new_n42838_ );
xor  ( new_n42841_, new_n21433_, new_n21432_ );
xor  ( new_n42842_, new_n42539_, new_n42538_ );
nor  ( new_n42843_, new_n42842_, new_n42841_ );
xor  ( new_n42844_, new_n21430_, new_n21429_ );
xor  ( new_n42845_, new_n42536_, new_n42535_ );
nor  ( new_n42846_, new_n42845_, new_n42844_ );
xor  ( new_n42847_, new_n21427_, new_n21426_ );
xor  ( new_n42848_, new_n42533_, new_n42532_ );
nor  ( new_n42849_, new_n42848_, new_n42847_ );
xor  ( new_n42850_, new_n21424_, new_n21423_ );
xor  ( new_n42851_, new_n42530_, new_n42529_ );
nor  ( new_n42852_, new_n42851_, new_n42850_ );
and  ( new_n42853_, new_n42851_, new_n42850_ );
xor  ( new_n42854_, new_n42527_, new_n42526_ );
xor  ( new_n42855_, new_n21417_, new_n21416_ );
xor  ( new_n42856_, new_n42523_, new_n42522_ );
nor  ( new_n42857_, new_n42856_, new_n42855_ );
xor  ( new_n42858_, new_n21414_, new_n21413_ );
xor  ( new_n42859_, new_n42520_, new_n42519_ );
nor  ( new_n42860_, new_n42859_, new_n42858_ );
xor  ( new_n42861_, new_n21411_, new_n21410_ );
xor  ( new_n42862_, new_n42517_, new_n42516_ );
nor  ( new_n42863_, new_n42862_, new_n42861_ );
xor  ( new_n42864_, new_n21408_, new_n21407_ );
xor  ( new_n42865_, new_n42514_, new_n42513_ );
nor  ( new_n42866_, new_n42865_, new_n42864_ );
xor  ( new_n42867_, new_n21405_, new_n21404_ );
xor  ( new_n42868_, new_n42511_, new_n42510_ );
nor  ( new_n42869_, new_n42868_, new_n42867_ );
xor  ( new_n42870_, new_n21402_, new_n21401_ );
xor  ( new_n42871_, new_n42508_, new_n42507_ );
nor  ( new_n42872_, new_n42871_, new_n42870_ );
xor  ( new_n42873_, new_n21399_, new_n21398_ );
xor  ( new_n42874_, new_n42505_, new_n42504_ );
nor  ( new_n42875_, new_n42874_, new_n42873_ );
xor  ( new_n42876_, new_n21396_, new_n21395_ );
xor  ( new_n42877_, new_n42502_, new_n42501_ );
nor  ( new_n42878_, new_n42877_, new_n42876_ );
xor  ( new_n42879_, new_n21393_, new_n21392_ );
xor  ( new_n42880_, new_n42499_, new_n42498_ );
nor  ( new_n42881_, new_n42880_, new_n42879_ );
xor  ( new_n42882_, new_n21390_, new_n21389_ );
xor  ( new_n42883_, new_n42496_, new_n42495_ );
nor  ( new_n42884_, new_n42883_, new_n42882_ );
xor  ( new_n42885_, new_n21387_, new_n21386_ );
xor  ( new_n42886_, new_n42493_, new_n42492_ );
nor  ( new_n42887_, new_n42886_, new_n42885_ );
xor  ( new_n42888_, new_n21384_, new_n21383_ );
xor  ( new_n42889_, new_n42490_, new_n42489_ );
nor  ( new_n42890_, new_n42889_, new_n42888_ );
xor  ( new_n42891_, new_n21381_, new_n21380_ );
xor  ( new_n42892_, new_n42487_, new_n42486_ );
nor  ( new_n42893_, new_n42892_, new_n42891_ );
xor  ( new_n42894_, new_n21378_, new_n21377_ );
xor  ( new_n42895_, new_n42484_, new_n42483_ );
nor  ( new_n42896_, new_n42895_, new_n42894_ );
xor  ( new_n42897_, new_n21375_, new_n21374_ );
xor  ( new_n42898_, new_n42481_, new_n42480_ );
nor  ( new_n42899_, new_n42898_, new_n42897_ );
xor  ( new_n42900_, new_n21372_, new_n21371_ );
xor  ( new_n42901_, new_n42478_, new_n42477_ );
nor  ( new_n42902_, new_n42901_, new_n42900_ );
xor  ( new_n42903_, new_n21369_, new_n21368_ );
xor  ( new_n42904_, new_n42475_, new_n42474_ );
nor  ( new_n42905_, new_n42904_, new_n42903_ );
xor  ( new_n42906_, new_n21366_, new_n21365_ );
xor  ( new_n42907_, new_n42472_, new_n42471_ );
nor  ( new_n42908_, new_n42907_, new_n42906_ );
xor  ( new_n42909_, new_n21363_, new_n21362_ );
xor  ( new_n42910_, new_n42469_, new_n42468_ );
nor  ( new_n42911_, new_n42910_, new_n42909_ );
xor  ( new_n42912_, new_n21360_, new_n21359_ );
xor  ( new_n42913_, new_n42466_, new_n42465_ );
nor  ( new_n42914_, new_n42913_, new_n42912_ );
xor  ( new_n42915_, new_n21357_, new_n21356_ );
xor  ( new_n42916_, new_n42463_, new_n42462_ );
nor  ( new_n42917_, new_n42916_, new_n42915_ );
xor  ( new_n42918_, new_n21354_, new_n21353_ );
xor  ( new_n42919_, new_n42460_, new_n42459_ );
nor  ( new_n42920_, new_n42919_, new_n42918_ );
xor  ( new_n42921_, new_n21351_, new_n21350_ );
xor  ( new_n42922_, new_n42457_, new_n42456_ );
nor  ( new_n42923_, new_n42922_, new_n42921_ );
xor  ( new_n42924_, new_n21348_, new_n21347_ );
xor  ( new_n42925_, new_n42454_, new_n42453_ );
nor  ( new_n42926_, new_n42925_, new_n42924_ );
xor  ( new_n42927_, new_n21345_, new_n21344_ );
xor  ( new_n42928_, new_n42451_, new_n42450_ );
nor  ( new_n42929_, new_n42928_, new_n42927_ );
xor  ( new_n42930_, new_n21342_, new_n21341_ );
xor  ( new_n42931_, new_n42448_, new_n42447_ );
nor  ( new_n42932_, new_n42931_, new_n42930_ );
xor  ( new_n42933_, new_n21339_, new_n21338_ );
xor  ( new_n42934_, new_n42445_, new_n42444_ );
nor  ( new_n42935_, new_n42934_, new_n42933_ );
xor  ( new_n42936_, new_n21336_, new_n21335_ );
xor  ( new_n42937_, new_n42442_, new_n42441_ );
nor  ( new_n42938_, new_n42937_, new_n42936_ );
xor  ( new_n42939_, new_n21333_, new_n21332_ );
xor  ( new_n42940_, new_n42439_, new_n42438_ );
nor  ( new_n42941_, new_n42940_, new_n42939_ );
xor  ( new_n42942_, new_n21330_, new_n21329_ );
xor  ( new_n42943_, new_n42436_, new_n42435_ );
nor  ( new_n42944_, new_n42943_, new_n42942_ );
and  ( new_n42945_, new_n42943_, new_n42942_ );
xor  ( new_n42946_, new_n42433_, new_n42432_ );
xor  ( new_n42947_, new_n21323_, new_n21322_ );
xor  ( new_n42948_, new_n42430_, new_n42429_ );
or   ( new_n42949_, new_n42948_, new_n42947_ );
and  ( new_n42950_, new_n42948_, new_n42947_ );
xor  ( new_n42951_, new_n21320_, new_n21319_ );
xor  ( new_n42952_, new_n42427_, new_n42426_ );
nor  ( new_n42953_, new_n42952_, new_n42951_ );
xor  ( new_n42954_, new_n21317_, new_n21316_ );
xor  ( new_n42955_, new_n42424_, new_n42423_ );
nor  ( new_n42956_, new_n42955_, new_n42954_ );
xor  ( new_n42957_, new_n21314_, new_n21313_ );
xor  ( new_n42958_, new_n42421_, new_n42420_ );
nor  ( new_n42959_, new_n42958_, new_n42957_ );
xor  ( new_n42960_, new_n21311_, new_n21310_ );
xor  ( new_n42961_, new_n42418_, new_n42417_ );
nor  ( new_n42962_, new_n42961_, new_n42960_ );
xor  ( new_n42963_, new_n21308_, new_n21307_ );
xor  ( new_n42964_, new_n42415_, new_n42414_ );
nor  ( new_n42965_, new_n42964_, new_n42963_ );
xor  ( new_n42966_, new_n21305_, new_n21304_ );
xor  ( new_n42967_, new_n42412_, new_n42411_ );
nor  ( new_n42968_, new_n42967_, new_n42966_ );
xor  ( new_n42969_, new_n21302_, new_n21301_ );
xor  ( new_n42970_, new_n42409_, new_n42408_ );
nor  ( new_n42971_, new_n42970_, new_n42969_ );
xor  ( new_n42972_, new_n21299_, new_n21298_ );
xor  ( new_n42973_, new_n42406_, new_n42405_ );
nor  ( new_n42974_, new_n42973_, new_n42972_ );
xor  ( new_n42975_, new_n21296_, new_n21295_ );
xor  ( new_n42976_, new_n42403_, new_n42402_ );
nor  ( new_n42977_, new_n42976_, new_n42975_ );
xor  ( new_n42978_, new_n21293_, new_n21292_ );
xor  ( new_n42979_, new_n42400_, new_n42399_ );
nor  ( new_n42980_, new_n42979_, new_n42978_ );
xor  ( new_n42981_, new_n21290_, new_n21289_ );
xor  ( new_n42982_, new_n42397_, new_n42396_ );
nor  ( new_n42983_, new_n42982_, new_n42981_ );
xor  ( new_n42984_, new_n21287_, new_n21286_ );
xor  ( new_n42985_, new_n42394_, new_n42393_ );
nor  ( new_n42986_, new_n42985_, new_n42984_ );
xor  ( new_n42987_, new_n21284_, new_n21283_ );
xor  ( new_n42988_, new_n42391_, new_n42390_ );
nor  ( new_n42989_, new_n42988_, new_n42987_ );
and  ( new_n42990_, new_n42988_, new_n42987_ );
xor  ( new_n42991_, new_n21281_, new_n21280_ );
xor  ( new_n42992_, new_n42388_, new_n42387_ );
nor  ( new_n42993_, new_n42992_, new_n42991_ );
and  ( new_n42994_, new_n42992_, new_n42991_ );
xor  ( new_n42995_, new_n21278_, new_n21277_ );
xor  ( new_n42996_, new_n42385_, new_n42384_ );
nor  ( new_n42997_, new_n42996_, new_n42995_ );
and  ( new_n42998_, new_n42996_, new_n42995_ );
xor  ( new_n42999_, new_n21275_, new_n21274_ );
xor  ( new_n43000_, new_n42382_, new_n42381_ );
nor  ( new_n43001_, new_n43000_, new_n42999_ );
xor  ( new_n43002_, new_n21272_, new_n21271_ );
xor  ( new_n43003_, new_n42379_, new_n42378_ );
nor  ( new_n43004_, new_n43003_, new_n43002_ );
xor  ( new_n43005_, new_n21269_, new_n21268_ );
xor  ( new_n43006_, new_n42376_, new_n42375_ );
nor  ( new_n43007_, new_n43006_, new_n43005_ );
xor  ( new_n43008_, new_n21266_, new_n21265_ );
xor  ( new_n43009_, new_n42373_, new_n42372_ );
nor  ( new_n43010_, new_n43009_, new_n43008_ );
xor  ( new_n43011_, new_n21263_, new_n21262_ );
xor  ( new_n43012_, new_n42370_, new_n42369_ );
nor  ( new_n43013_, new_n43012_, new_n43011_ );
and  ( new_n43014_, new_n43012_, new_n43011_ );
xor  ( new_n43015_, new_n42339_, new_n42338_ );
xor  ( new_n43016_, new_n21232_, new_n21231_ );
and  ( new_n43017_, new_n43016_, new_n43015_ );
not  ( new_n43018_, new_n43017_ );
and  ( new_n43019_, RIbb33378_192, RIbb31578_128 );
and  ( new_n43020_, new_n43019_, RIbb2d888_64 );
and  ( new_n43021_, new_n43020_, new_n42337_ );
xor  ( new_n43022_, new_n42337_, new_n42331_ );
nor  ( new_n43023_, new_n43022_, new_n43020_ );
not  ( new_n43024_, new_n43023_ );
xor  ( new_n43025_, new_n21230_, new_n21224_ );
and  ( new_n43026_, new_n43025_, new_n43024_ );
nor  ( new_n43027_, new_n43026_, new_n43021_ );
and  ( new_n43028_, new_n43027_, new_n43018_ );
nor  ( new_n43029_, new_n43016_, new_n43015_ );
nor  ( new_n43030_, new_n43029_, new_n43028_ );
xor  ( new_n43031_, new_n42343_, new_n42342_ );
xor  ( new_n43032_, new_n21236_, new_n21235_ );
and  ( new_n43033_, new_n43032_, new_n43031_ );
nor  ( new_n43034_, new_n43033_, new_n43030_ );
nor  ( new_n43035_, new_n43032_, new_n43031_ );
nor  ( new_n43036_, new_n43035_, new_n43034_ );
xor  ( new_n43037_, new_n42347_, new_n42346_ );
xor  ( new_n43038_, new_n21240_, new_n21239_ );
and  ( new_n43039_, new_n43038_, new_n43037_ );
nor  ( new_n43040_, new_n43039_, new_n43036_ );
nor  ( new_n43041_, new_n43038_, new_n43037_ );
nor  ( new_n43042_, new_n43041_, new_n43040_ );
xor  ( new_n43043_, new_n42351_, new_n42350_ );
xor  ( new_n43044_, new_n21244_, new_n21243_ );
and  ( new_n43045_, new_n43044_, new_n43043_ );
nor  ( new_n43046_, new_n43045_, new_n43042_ );
nor  ( new_n43047_, new_n43044_, new_n43043_ );
nor  ( new_n43048_, new_n43047_, new_n43046_ );
xor  ( new_n43049_, new_n42355_, new_n42354_ );
xor  ( new_n43050_, new_n21248_, new_n21247_ );
and  ( new_n43051_, new_n43050_, new_n43049_ );
nor  ( new_n43052_, new_n43051_, new_n43048_ );
nor  ( new_n43053_, new_n43050_, new_n43049_ );
nor  ( new_n43054_, new_n43053_, new_n43052_ );
xor  ( new_n43055_, new_n42359_, new_n42358_ );
xor  ( new_n43056_, new_n21252_, new_n21251_ );
and  ( new_n43057_, new_n43056_, new_n43055_ );
nor  ( new_n43058_, new_n43057_, new_n43054_ );
nor  ( new_n43059_, new_n43056_, new_n43055_ );
nor  ( new_n43060_, new_n43059_, new_n43058_ );
xor  ( new_n43061_, new_n42363_, new_n42362_ );
xor  ( new_n43062_, new_n21256_, new_n21255_ );
and  ( new_n43063_, new_n43062_, new_n43061_ );
nor  ( new_n43064_, new_n43063_, new_n43060_ );
nor  ( new_n43065_, new_n43062_, new_n43061_ );
nor  ( new_n43066_, new_n43065_, new_n43064_ );
xor  ( new_n43067_, new_n42367_, new_n42366_ );
xor  ( new_n43068_, new_n21260_, new_n21259_ );
and  ( new_n43069_, new_n43068_, new_n43067_ );
nor  ( new_n43070_, new_n43069_, new_n43066_ );
nor  ( new_n43071_, new_n43068_, new_n43067_ );
nor  ( new_n43072_, new_n43071_, new_n43070_ );
nor  ( new_n43073_, new_n43072_, new_n43014_ );
nor  ( new_n43074_, new_n43073_, new_n43013_ );
and  ( new_n43075_, new_n43009_, new_n43008_ );
nor  ( new_n43076_, new_n43075_, new_n43074_ );
nor  ( new_n43077_, new_n43076_, new_n43010_ );
and  ( new_n43078_, new_n43006_, new_n43005_ );
nor  ( new_n43079_, new_n43078_, new_n43077_ );
nor  ( new_n43080_, new_n43079_, new_n43007_ );
and  ( new_n43081_, new_n43003_, new_n43002_ );
nor  ( new_n43082_, new_n43081_, new_n43080_ );
nor  ( new_n43083_, new_n43082_, new_n43004_ );
and  ( new_n43084_, new_n43000_, new_n42999_ );
nor  ( new_n43085_, new_n43084_, new_n43083_ );
nor  ( new_n43086_, new_n43085_, new_n43001_ );
nor  ( new_n43087_, new_n43086_, new_n42998_ );
nor  ( new_n43088_, new_n43087_, new_n42997_ );
nor  ( new_n43089_, new_n43088_, new_n42994_ );
nor  ( new_n43090_, new_n43089_, new_n42993_ );
nor  ( new_n43091_, new_n43090_, new_n42990_ );
nor  ( new_n43092_, new_n43091_, new_n42989_ );
and  ( new_n43093_, new_n42985_, new_n42984_ );
nor  ( new_n43094_, new_n43093_, new_n43092_ );
nor  ( new_n43095_, new_n43094_, new_n42986_ );
and  ( new_n43096_, new_n42982_, new_n42981_ );
nor  ( new_n43097_, new_n43096_, new_n43095_ );
nor  ( new_n43098_, new_n43097_, new_n42983_ );
and  ( new_n43099_, new_n42979_, new_n42978_ );
nor  ( new_n43100_, new_n43099_, new_n43098_ );
nor  ( new_n43101_, new_n43100_, new_n42980_ );
and  ( new_n43102_, new_n42976_, new_n42975_ );
nor  ( new_n43103_, new_n43102_, new_n43101_ );
nor  ( new_n43104_, new_n43103_, new_n42977_ );
and  ( new_n43105_, new_n42973_, new_n42972_ );
nor  ( new_n43106_, new_n43105_, new_n43104_ );
nor  ( new_n43107_, new_n43106_, new_n42974_ );
and  ( new_n43108_, new_n42970_, new_n42969_ );
nor  ( new_n43109_, new_n43108_, new_n43107_ );
nor  ( new_n43110_, new_n43109_, new_n42971_ );
and  ( new_n43111_, new_n42967_, new_n42966_ );
nor  ( new_n43112_, new_n43111_, new_n43110_ );
nor  ( new_n43113_, new_n43112_, new_n42968_ );
and  ( new_n43114_, new_n42964_, new_n42963_ );
nor  ( new_n43115_, new_n43114_, new_n43113_ );
nor  ( new_n43116_, new_n43115_, new_n42965_ );
and  ( new_n43117_, new_n42961_, new_n42960_ );
nor  ( new_n43118_, new_n43117_, new_n43116_ );
nor  ( new_n43119_, new_n43118_, new_n42962_ );
and  ( new_n43120_, new_n42958_, new_n42957_ );
nor  ( new_n43121_, new_n43120_, new_n43119_ );
nor  ( new_n43122_, new_n43121_, new_n42959_ );
and  ( new_n43123_, new_n42955_, new_n42954_ );
nor  ( new_n43124_, new_n43123_, new_n43122_ );
nor  ( new_n43125_, new_n43124_, new_n42956_ );
and  ( new_n43126_, new_n42952_, new_n42951_ );
nor  ( new_n43127_, new_n43126_, new_n43125_ );
nor  ( new_n43128_, new_n43127_, new_n42953_ );
or   ( new_n43129_, new_n43128_, new_n42950_ );
and  ( new_n43130_, new_n43129_, new_n42949_ );
nor  ( new_n43131_, new_n43130_, new_n42946_ );
and  ( new_n43132_, new_n43130_, new_n42946_ );
xor  ( new_n43133_, new_n21327_, new_n21326_ );
nor  ( new_n43134_, new_n43133_, new_n43132_ );
nor  ( new_n43135_, new_n43134_, new_n43131_ );
nor  ( new_n43136_, new_n43135_, new_n42945_ );
nor  ( new_n43137_, new_n43136_, new_n42944_ );
and  ( new_n43138_, new_n42940_, new_n42939_ );
nor  ( new_n43139_, new_n43138_, new_n43137_ );
nor  ( new_n43140_, new_n43139_, new_n42941_ );
and  ( new_n43141_, new_n42937_, new_n42936_ );
nor  ( new_n43142_, new_n43141_, new_n43140_ );
nor  ( new_n43143_, new_n43142_, new_n42938_ );
and  ( new_n43144_, new_n42934_, new_n42933_ );
nor  ( new_n43145_, new_n43144_, new_n43143_ );
nor  ( new_n43146_, new_n43145_, new_n42935_ );
and  ( new_n43147_, new_n42931_, new_n42930_ );
nor  ( new_n43148_, new_n43147_, new_n43146_ );
nor  ( new_n43149_, new_n43148_, new_n42932_ );
and  ( new_n43150_, new_n42928_, new_n42927_ );
nor  ( new_n43151_, new_n43150_, new_n43149_ );
nor  ( new_n43152_, new_n43151_, new_n42929_ );
and  ( new_n43153_, new_n42925_, new_n42924_ );
nor  ( new_n43154_, new_n43153_, new_n43152_ );
nor  ( new_n43155_, new_n43154_, new_n42926_ );
and  ( new_n43156_, new_n42922_, new_n42921_ );
nor  ( new_n43157_, new_n43156_, new_n43155_ );
nor  ( new_n43158_, new_n43157_, new_n42923_ );
and  ( new_n43159_, new_n42919_, new_n42918_ );
nor  ( new_n43160_, new_n43159_, new_n43158_ );
nor  ( new_n43161_, new_n43160_, new_n42920_ );
and  ( new_n43162_, new_n42916_, new_n42915_ );
nor  ( new_n43163_, new_n43162_, new_n43161_ );
nor  ( new_n43164_, new_n43163_, new_n42917_ );
and  ( new_n43165_, new_n42913_, new_n42912_ );
nor  ( new_n43166_, new_n43165_, new_n43164_ );
nor  ( new_n43167_, new_n43166_, new_n42914_ );
and  ( new_n43168_, new_n42910_, new_n42909_ );
nor  ( new_n43169_, new_n43168_, new_n43167_ );
nor  ( new_n43170_, new_n43169_, new_n42911_ );
and  ( new_n43171_, new_n42907_, new_n42906_ );
nor  ( new_n43172_, new_n43171_, new_n43170_ );
nor  ( new_n43173_, new_n43172_, new_n42908_ );
and  ( new_n43174_, new_n42904_, new_n42903_ );
nor  ( new_n43175_, new_n43174_, new_n43173_ );
nor  ( new_n43176_, new_n43175_, new_n42905_ );
and  ( new_n43177_, new_n42901_, new_n42900_ );
nor  ( new_n43178_, new_n43177_, new_n43176_ );
nor  ( new_n43179_, new_n43178_, new_n42902_ );
and  ( new_n43180_, new_n42898_, new_n42897_ );
nor  ( new_n43181_, new_n43180_, new_n43179_ );
nor  ( new_n43182_, new_n43181_, new_n42899_ );
and  ( new_n43183_, new_n42895_, new_n42894_ );
nor  ( new_n43184_, new_n43183_, new_n43182_ );
nor  ( new_n43185_, new_n43184_, new_n42896_ );
and  ( new_n43186_, new_n42892_, new_n42891_ );
nor  ( new_n43187_, new_n43186_, new_n43185_ );
nor  ( new_n43188_, new_n43187_, new_n42893_ );
and  ( new_n43189_, new_n42889_, new_n42888_ );
nor  ( new_n43190_, new_n43189_, new_n43188_ );
nor  ( new_n43191_, new_n43190_, new_n42890_ );
and  ( new_n43192_, new_n42886_, new_n42885_ );
nor  ( new_n43193_, new_n43192_, new_n43191_ );
nor  ( new_n43194_, new_n43193_, new_n42887_ );
and  ( new_n43195_, new_n42883_, new_n42882_ );
nor  ( new_n43196_, new_n43195_, new_n43194_ );
nor  ( new_n43197_, new_n43196_, new_n42884_ );
and  ( new_n43198_, new_n42880_, new_n42879_ );
nor  ( new_n43199_, new_n43198_, new_n43197_ );
nor  ( new_n43200_, new_n43199_, new_n42881_ );
and  ( new_n43201_, new_n42877_, new_n42876_ );
nor  ( new_n43202_, new_n43201_, new_n43200_ );
nor  ( new_n43203_, new_n43202_, new_n42878_ );
and  ( new_n43204_, new_n42874_, new_n42873_ );
nor  ( new_n43205_, new_n43204_, new_n43203_ );
nor  ( new_n43206_, new_n43205_, new_n42875_ );
and  ( new_n43207_, new_n42871_, new_n42870_ );
nor  ( new_n43208_, new_n43207_, new_n43206_ );
nor  ( new_n43209_, new_n43208_, new_n42872_ );
and  ( new_n43210_, new_n42868_, new_n42867_ );
nor  ( new_n43211_, new_n43210_, new_n43209_ );
nor  ( new_n43212_, new_n43211_, new_n42869_ );
and  ( new_n43213_, new_n42865_, new_n42864_ );
nor  ( new_n43214_, new_n43213_, new_n43212_ );
nor  ( new_n43215_, new_n43214_, new_n42866_ );
and  ( new_n43216_, new_n42862_, new_n42861_ );
nor  ( new_n43217_, new_n43216_, new_n43215_ );
nor  ( new_n43218_, new_n43217_, new_n42863_ );
and  ( new_n43219_, new_n42859_, new_n42858_ );
nor  ( new_n43220_, new_n43219_, new_n43218_ );
nor  ( new_n43221_, new_n43220_, new_n42860_ );
and  ( new_n43222_, new_n42856_, new_n42855_ );
nor  ( new_n43223_, new_n43222_, new_n43221_ );
nor  ( new_n43224_, new_n43223_, new_n42857_ );
xor  ( new_n43225_, new_n21421_, new_n21420_ );
and  ( new_n43226_, new_n43225_, new_n43224_ );
nor  ( new_n43227_, new_n43226_, new_n42854_ );
nor  ( new_n43228_, new_n43225_, new_n43224_ );
nor  ( new_n43229_, new_n43228_, new_n43227_ );
nor  ( new_n43230_, new_n43229_, new_n42853_ );
nor  ( new_n43231_, new_n43230_, new_n42852_ );
and  ( new_n43232_, new_n42848_, new_n42847_ );
nor  ( new_n43233_, new_n43232_, new_n43231_ );
nor  ( new_n43234_, new_n43233_, new_n42849_ );
and  ( new_n43235_, new_n42845_, new_n42844_ );
nor  ( new_n43236_, new_n43235_, new_n43234_ );
nor  ( new_n43237_, new_n43236_, new_n42846_ );
and  ( new_n43238_, new_n42842_, new_n42841_ );
nor  ( new_n43239_, new_n43238_, new_n43237_ );
nor  ( new_n43240_, new_n43239_, new_n42843_ );
and  ( new_n43241_, new_n42839_, new_n42838_ );
nor  ( new_n43242_, new_n43241_, new_n43240_ );
nor  ( new_n43243_, new_n43242_, new_n42840_ );
xor  ( new_n43244_, new_n21440_, new_n21439_ );
and  ( new_n43245_, new_n43244_, new_n43243_ );
nor  ( new_n43246_, new_n43245_, new_n42837_ );
nor  ( new_n43247_, new_n43244_, new_n43243_ );
nor  ( new_n43248_, new_n43247_, new_n43246_ );
nor  ( new_n43249_, new_n43248_, new_n42836_ );
nor  ( new_n43250_, new_n43249_, new_n42835_ );
xor  ( new_n43251_, new_n21447_, new_n21446_ );
and  ( new_n43252_, new_n43251_, new_n43250_ );
nor  ( new_n43253_, new_n43252_, new_n42832_ );
nor  ( new_n43254_, new_n43251_, new_n43250_ );
nor  ( new_n43255_, new_n43254_, new_n43253_ );
nor  ( new_n43256_, new_n43255_, new_n42831_ );
nor  ( new_n43257_, new_n43256_, new_n42830_ );
and  ( new_n43258_, new_n42826_, new_n42825_ );
nor  ( new_n43259_, new_n43258_, new_n43257_ );
nor  ( new_n43260_, new_n43259_, new_n42827_ );
and  ( new_n43261_, new_n42823_, new_n42822_ );
nor  ( new_n43262_, new_n43261_, new_n43260_ );
nor  ( new_n43263_, new_n43262_, new_n42824_ );
and  ( new_n43264_, new_n42820_, new_n42819_ );
nor  ( new_n43265_, new_n43264_, new_n43263_ );
nor  ( new_n43266_, new_n43265_, new_n42821_ );
and  ( new_n43267_, new_n42817_, new_n42816_ );
nor  ( new_n43268_, new_n43267_, new_n43266_ );
nor  ( new_n43269_, new_n43268_, new_n42818_ );
xor  ( new_n43270_, new_n21466_, new_n21465_ );
and  ( new_n43271_, new_n43270_, new_n43269_ );
nor  ( new_n43272_, new_n43271_, new_n42815_ );
nor  ( new_n43273_, new_n43270_, new_n43269_ );
nor  ( new_n43274_, new_n43273_, new_n43272_ );
xor  ( new_n43275_, new_n42576_, new_n42575_ );
xor  ( new_n43276_, new_n21470_, new_n21469_ );
and  ( new_n43277_, new_n43276_, new_n43275_ );
nor  ( new_n43278_, new_n43277_, new_n43274_ );
nor  ( new_n43279_, new_n43276_, new_n43275_ );
nor  ( new_n43280_, new_n43279_, new_n43278_ );
xor  ( new_n43281_, new_n42580_, new_n42579_ );
xor  ( new_n43282_, new_n21474_, new_n21473_ );
and  ( new_n43283_, new_n43282_, new_n43281_ );
nor  ( new_n43284_, new_n43283_, new_n43280_ );
nor  ( new_n43285_, new_n43282_, new_n43281_ );
nor  ( new_n43286_, new_n43285_, new_n43284_ );
nor  ( new_n43287_, new_n43286_, new_n42814_ );
nor  ( new_n43288_, new_n43287_, new_n42813_ );
and  ( new_n43289_, new_n42809_, new_n42808_ );
nor  ( new_n43290_, new_n43289_, new_n43288_ );
nor  ( new_n43291_, new_n43290_, new_n42810_ );
and  ( new_n43292_, new_n42806_, new_n42805_ );
nor  ( new_n43293_, new_n43292_, new_n43291_ );
nor  ( new_n43294_, new_n43293_, new_n42807_ );
and  ( new_n43295_, new_n42803_, new_n42802_ );
nor  ( new_n43296_, new_n43295_, new_n43294_ );
nor  ( new_n43297_, new_n43296_, new_n42804_ );
xor  ( new_n43298_, new_n21490_, new_n21489_ );
and  ( new_n43299_, new_n43298_, new_n43297_ );
nor  ( new_n43300_, new_n43299_, new_n42801_ );
nor  ( new_n43301_, new_n43298_, new_n43297_ );
nor  ( new_n43302_, new_n43301_, new_n43300_ );
nor  ( new_n43303_, new_n43302_, new_n42800_ );
nor  ( new_n43304_, new_n43303_, new_n42799_ );
and  ( new_n43305_, new_n42795_, new_n42794_ );
nor  ( new_n43306_, new_n43305_, new_n43304_ );
nor  ( new_n43307_, new_n43306_, new_n42796_ );
xor  ( new_n43308_, new_n21500_, new_n21499_ );
and  ( new_n43309_, new_n43308_, new_n43307_ );
nor  ( new_n43310_, new_n43309_, new_n42793_ );
nor  ( new_n43311_, new_n43308_, new_n43307_ );
nor  ( new_n43312_, new_n43311_, new_n43310_ );
nor  ( new_n43313_, new_n43312_, new_n42792_ );
nor  ( new_n43314_, new_n43313_, new_n42791_ );
and  ( new_n43315_, new_n42787_, new_n42786_ );
nor  ( new_n43316_, new_n43315_, new_n43314_ );
nor  ( new_n43317_, new_n43316_, new_n42788_ );
and  ( new_n43318_, new_n42784_, new_n42783_ );
nor  ( new_n43319_, new_n43318_, new_n43317_ );
nor  ( new_n43320_, new_n43319_, new_n42785_ );
xor  ( new_n43321_, new_n21513_, new_n21512_ );
and  ( new_n43322_, new_n43321_, new_n43320_ );
nor  ( new_n43323_, new_n43322_, new_n42782_ );
nor  ( new_n43324_, new_n43321_, new_n43320_ );
nor  ( new_n43325_, new_n43324_, new_n43323_ );
or   ( new_n43326_, new_n43325_, new_n42781_ );
and  ( new_n43327_, new_n43326_, new_n42780_ );
nor  ( new_n43328_, new_n43327_, new_n42777_ );
and  ( new_n43329_, new_n43327_, new_n42777_ );
xor  ( new_n43330_, new_n21520_, new_n21519_ );
nor  ( new_n43331_, new_n43330_, new_n43329_ );
nor  ( new_n43332_, new_n43331_, new_n43328_ );
nor  ( new_n43333_, new_n43332_, new_n42776_ );
nor  ( new_n43334_, new_n43333_, new_n42775_ );
and  ( new_n43335_, new_n42771_, new_n42770_ );
nor  ( new_n43336_, new_n43335_, new_n43334_ );
nor  ( new_n43337_, new_n43336_, new_n42772_ );
xor  ( new_n43338_, new_n21531_, new_n21530_ );
and  ( new_n43339_, new_n43338_, new_n43337_ );
nor  ( new_n43340_, new_n43339_, new_n42769_ );
nor  ( new_n43341_, new_n43338_, new_n43337_ );
nor  ( new_n43342_, new_n43341_, new_n43340_ );
xor  ( new_n43343_, new_n42640_, new_n42639_ );
xor  ( new_n43344_, new_n21535_, new_n21534_ );
and  ( new_n43345_, new_n43344_, new_n43343_ );
nor  ( new_n43346_, new_n43345_, new_n43342_ );
nor  ( new_n43347_, new_n43344_, new_n43343_ );
nor  ( new_n43348_, new_n43347_, new_n43346_ );
nor  ( new_n43349_, new_n43348_, new_n42768_ );
nor  ( new_n43350_, new_n43349_, new_n42767_ );
xor  ( new_n43351_, new_n21542_, new_n21541_ );
and  ( new_n43352_, new_n43351_, new_n43350_ );
nor  ( new_n43353_, new_n43352_, new_n42764_ );
nor  ( new_n43354_, new_n43351_, new_n43350_ );
nor  ( new_n43355_, new_n43354_, new_n43353_ );
nor  ( new_n43356_, new_n43355_, new_n42763_ );
nor  ( new_n43357_, new_n43356_, new_n42762_ );
and  ( new_n43358_, new_n42758_, new_n42757_ );
nor  ( new_n43359_, new_n43358_, new_n43357_ );
nor  ( new_n43360_, new_n43359_, new_n42759_ );
xor  ( new_n43361_, new_n21552_, new_n21551_ );
and  ( new_n43362_, new_n43361_, new_n43360_ );
nor  ( new_n43363_, new_n43362_, new_n42756_ );
nor  ( new_n43364_, new_n43361_, new_n43360_ );
nor  ( new_n43365_, new_n43364_, new_n43363_ );
xor  ( new_n43366_, new_n42661_, new_n42660_ );
xor  ( new_n43367_, new_n21556_, new_n21555_ );
and  ( new_n43368_, new_n43367_, new_n43366_ );
nor  ( new_n43369_, new_n43368_, new_n43365_ );
nor  ( new_n43370_, new_n43367_, new_n43366_ );
nor  ( new_n43371_, new_n43370_, new_n43369_ );
nor  ( new_n43372_, new_n43371_, new_n42755_ );
nor  ( new_n43373_, new_n43372_, new_n42754_ );
xor  ( new_n43374_, new_n21563_, new_n21562_ );
and  ( new_n43375_, new_n43374_, new_n43373_ );
nor  ( new_n43376_, new_n43375_, new_n42751_ );
nor  ( new_n43377_, new_n43374_, new_n43373_ );
nor  ( new_n43378_, new_n43377_, new_n43376_ );
xor  ( new_n43379_, new_n42672_, new_n42671_ );
xor  ( new_n43380_, new_n21567_, new_n21566_ );
and  ( new_n43381_, new_n43380_, new_n43379_ );
nor  ( new_n43382_, new_n43381_, new_n43378_ );
nor  ( new_n43383_, new_n43380_, new_n43379_ );
nor  ( new_n43384_, new_n43383_, new_n43382_ );
xor  ( new_n43385_, new_n42676_, new_n42675_ );
xor  ( new_n43386_, new_n21571_, new_n21570_ );
and  ( new_n43387_, new_n43386_, new_n43385_ );
nor  ( new_n43388_, new_n43387_, new_n43384_ );
nor  ( new_n43389_, new_n43386_, new_n43385_ );
nor  ( new_n43390_, new_n43389_, new_n43388_ );
xor  ( new_n43391_, new_n42680_, new_n42679_ );
xor  ( new_n43392_, new_n21575_, new_n21574_ );
and  ( new_n43393_, new_n43392_, new_n43391_ );
nor  ( new_n43394_, new_n43393_, new_n43390_ );
nor  ( new_n43395_, new_n43392_, new_n43391_ );
nor  ( new_n43396_, new_n43395_, new_n43394_ );
xor  ( new_n43397_, new_n42684_, new_n42683_ );
xor  ( new_n43398_, new_n21579_, new_n21578_ );
and  ( new_n43399_, new_n43398_, new_n43397_ );
nor  ( new_n43400_, new_n43399_, new_n43396_ );
nor  ( new_n43401_, new_n43398_, new_n43397_ );
nor  ( new_n43402_, new_n43401_, new_n43400_ );
xor  ( new_n43403_, new_n42688_, new_n42687_ );
xor  ( new_n43404_, new_n21583_, new_n21582_ );
and  ( new_n43405_, new_n43404_, new_n43403_ );
nor  ( new_n43406_, new_n43405_, new_n43402_ );
nor  ( new_n43407_, new_n43404_, new_n43403_ );
nor  ( new_n43408_, new_n43407_, new_n43406_ );
xor  ( new_n43409_, new_n42692_, new_n42691_ );
xor  ( new_n43410_, new_n21587_, new_n21586_ );
and  ( new_n43411_, new_n43410_, new_n43409_ );
nor  ( new_n43412_, new_n43411_, new_n43408_ );
nor  ( new_n43413_, new_n43410_, new_n43409_ );
nor  ( new_n43414_, new_n43413_, new_n43412_ );
nor  ( new_n43415_, new_n43414_, new_n42750_ );
nor  ( new_n43416_, new_n43415_, new_n42749_ );
xor  ( new_n43417_, new_n21594_, new_n21593_ );
and  ( new_n43418_, new_n43417_, new_n43416_ );
nor  ( new_n43419_, new_n43418_, new_n42746_ );
nor  ( new_n43420_, new_n43417_, new_n43416_ );
nor  ( new_n43421_, new_n43420_, new_n43419_ );
nor  ( new_n43422_, new_n43421_, new_n42745_ );
nor  ( new_n43423_, new_n43422_, new_n42744_ );
xor  ( new_n43424_, new_n21601_, new_n21600_ );
and  ( new_n43425_, new_n43424_, new_n43423_ );
nor  ( new_n43426_, new_n43425_, new_n42741_ );
nor  ( new_n43427_, new_n43424_, new_n43423_ );
nor  ( new_n43428_, new_n43427_, new_n43426_ );
xor  ( new_n43429_, new_n42710_, new_n42709_ );
xor  ( new_n43430_, new_n21605_, new_n21604_ );
and  ( new_n43431_, new_n43430_, new_n43429_ );
nor  ( new_n43432_, new_n43431_, new_n43428_ );
nor  ( new_n43433_, new_n43430_, new_n43429_ );
nor  ( new_n43434_, new_n43433_, new_n43432_ );
or   ( new_n43435_, new_n43434_, new_n42740_ );
and  ( new_n43436_, new_n43435_, new_n42739_ );
xor  ( new_n43437_, new_n21611_, new_n21610_ );
and  ( new_n43438_, new_n43437_, new_n43436_ );
or   ( new_n43439_, new_n43438_, new_n42736_ );
or   ( new_n43440_, new_n43437_, new_n43436_ );
and  ( new_n43441_, new_n43440_, new_n43439_ );
nor  ( new_n43442_, new_n43441_, new_n42735_ );
and  ( new_n43443_, new_n43441_, new_n42735_ );
xor  ( new_n43444_, new_n21615_, new_n21614_ );
nor  ( new_n43445_, new_n43444_, new_n43443_ );
nor  ( new_n43446_, new_n43445_, new_n43442_ );
xor  ( new_n43447_, RIbb315f0_129, RIbb2d810_65 );
and  ( new_n43448_, RIbb31668_130, RIbb2d798_66 );
and  ( new_n43449_, new_n21694_, new_n333_ );
and  ( new_n43450_, RIbb316e0_131, RIbb2d720_67 );
and  ( new_n43451_, new_n21703_, new_n319_ );
and  ( new_n43452_, RIbb31758_132, RIbb2d6a8_68 );
and  ( new_n43453_, new_n21701_, new_n313_ );
and  ( new_n43454_, RIbb317d0_133, RIbb2d630_69 );
and  ( new_n43455_, RIbb31848_134, RIbb2d5b8_70 );
and  ( new_n43456_, new_n21672_, new_n279_ );
and  ( new_n43457_, RIbb318c0_135, RIbb2d540_71 );
and  ( new_n43458_, RIbb31938_136, RIbb2d4c8_72 );
and  ( new_n43459_, new_n21678_, new_n294_ );
and  ( new_n43460_, RIbb319b0_137, RIbb2d450_73 );
and  ( new_n43461_, new_n21687_, new_n270_ );
and  ( new_n43462_, RIbb31a28_138, RIbb2d3d8_74 );
and  ( new_n43463_, new_n21685_, new_n264_ );
and  ( new_n43464_, RIbb31aa0_139, RIbb2d360_75 );
and  ( new_n43465_, new_n21751_, new_n348_ );
and  ( new_n43466_, RIbb31b18_140, RIbb2d2e8_76 );
and  ( new_n43467_, new_n21792_, new_n419_ );
and  ( new_n43468_, RIbb31b90_141, RIbb2d270_77 );
and  ( new_n43469_, new_n21842_, new_n443_ );
and  ( new_n43470_, RIbb31c08_142, RIbb2d1f8_78 );
and  ( new_n43471_, new_n21840_, new_n509_ );
and  ( new_n43472_, RIbb31c80_143, RIbb2d180_79 );
and  ( new_n43473_, new_n21847_, new_n515_ );
and  ( new_n43474_, RIbb31cf8_144, RIbb2d108_80 );
and  ( new_n43475_, new_n22098_, new_n775_ );
and  ( new_n43476_, new_n22129_, new_n805_ );
not  ( new_n43477_, new_n43476_ );
and  ( new_n43478_, new_n22423_, new_n1168_ );
not  ( new_n43479_, new_n43478_ );
and  ( new_n43480_, new_n22207_, new_n886_ );
and  ( new_n43481_, new_n22304_, new_n986_ );
nor  ( new_n43482_, new_n43481_, new_n43480_ );
and  ( new_n43483_, new_n43482_, new_n43479_ );
and  ( new_n43484_, new_n43483_, new_n43477_ );
and  ( new_n43485_, new_n22829_, new_n1525_ );
not  ( new_n43486_, new_n43485_ );
and  ( new_n43487_, new_n22975_, new_n1523_ );
and  ( new_n43488_, new_n23733_, new_n2475_ );
and  ( new_n43489_, new_n23554_, new_n2291_ );
nor  ( new_n43490_, new_n43489_, new_n43488_ );
and  ( new_n43491_, new_n23895_, new_n2646_ );
not  ( new_n43492_, new_n43491_ );
and  ( new_n43493_, new_n24006_, new_n2751_ );
and  ( new_n43494_, new_n27602_, new_n6425_ );
not  ( new_n43495_, new_n43494_ );
and  ( new_n43496_, new_n28314_, new_n7149_ );
not  ( new_n43497_, new_n43496_ );
and  ( new_n43498_, new_n43497_, new_n43495_ );
and  ( new_n43499_, new_n28108_, new_n6943_ );
not  ( new_n43500_, new_n43499_ );
and  ( new_n43501_, new_n27763_, new_n6589_ );
not  ( new_n43502_, new_n43501_ );
and  ( new_n43503_, new_n43502_, new_n43500_ );
and  ( new_n43504_, new_n43503_, new_n43498_ );
not  ( new_n43505_, new_n43504_ );
and  ( new_n43506_, new_n29263_, new_n8117_ );
and  ( new_n43507_, new_n29261_, new_n8115_ );
nor  ( new_n43508_, new_n43507_, new_n43506_ );
and  ( new_n43509_, new_n28531_, new_n7373_ );
and  ( new_n43510_, new_n29474_, new_n8352_ );
nor  ( new_n43511_, new_n43510_, new_n43509_ );
and  ( new_n43512_, new_n43511_, new_n43508_ );
and  ( new_n43513_, new_n30120_, new_n8995_ );
and  ( new_n43514_, new_n29619_, new_n8481_ );
nor  ( new_n43515_, new_n43514_, new_n43513_ );
and  ( new_n43516_, new_n30227_, new_n9099_ );
not  ( new_n43517_, new_n43516_ );
and  ( new_n43518_, new_n30800_, new_n9681_ );
and  ( new_n43519_, new_n30798_, new_n9679_ );
and  ( new_n43520_, RIbb33210_189, RIbb2bbf0_125 );
and  ( new_n43521_, new_n31333_, new_n10220_ );
and  ( new_n43522_, RIbb33288_190, RIbb2bb78_126 );
and  ( new_n43523_, new_n31654_, new_n10541_ );
and  ( new_n43524_, RIbb33300_191, RIbb31500_127 );
nor  ( new_n43525_, new_n43524_, new_n43019_ );
nor  ( new_n43526_, new_n43525_, new_n43523_ );
nor  ( new_n43527_, new_n43526_, new_n43522_ );
nor  ( new_n43528_, new_n43527_, new_n43521_ );
nor  ( new_n43529_, new_n43528_, new_n43520_ );
nor  ( new_n43530_, new_n43529_, new_n43519_ );
not  ( new_n43531_, new_n43530_ );
nor  ( new_n43532_, new_n43531_, new_n43518_ );
and  ( new_n43533_, new_n43532_, new_n43517_ );
and  ( new_n43534_, new_n43533_, new_n43515_ );
and  ( new_n43535_, new_n43534_, new_n43512_ );
and  ( new_n43536_, RIbb32f40_183, RIbb2bec0_119 );
and  ( new_n43537_, RIbb32fb8_184, RIbb2be48_120 );
nor  ( new_n43538_, new_n43537_, new_n43536_ );
not  ( new_n43539_, new_n43538_ );
and  ( new_n43540_, new_n43539_, new_n43508_ );
not  ( new_n43541_, new_n43540_ );
and  ( new_n43542_, RIbb32ec8_182, RIbb2bf38_118 );
and  ( new_n43543_, RIbb32e50_181, RIbb2bfb0_117 );
nor  ( new_n43544_, new_n43543_, new_n43542_ );
and  ( new_n43545_, new_n43544_, new_n43541_ );
nor  ( new_n43546_, new_n43545_, new_n43509_ );
nor  ( new_n43547_, new_n43546_, new_n43535_ );
nor  ( new_n43548_, new_n43547_, new_n43505_ );
and  ( new_n43549_, new_n26762_, new_n5570_ );
and  ( new_n43550_, new_n26620_, new_n5428_ );
nor  ( new_n43551_, new_n43550_, new_n43549_ );
and  ( new_n43552_, new_n27085_, new_n5899_ );
not  ( new_n43553_, new_n43552_ );
and  ( new_n43554_, new_n27396_, new_n6219_ );
not  ( new_n43555_, new_n43554_ );
and  ( new_n43556_, new_n43555_, new_n43553_ );
and  ( new_n43557_, new_n43556_, new_n43551_ );
and  ( new_n43558_, new_n25813_, new_n4603_ );
not  ( new_n43559_, new_n43558_ );
and  ( new_n43560_, new_n26372_, new_n5171_ );
not  ( new_n43561_, new_n43560_ );
and  ( new_n43562_, new_n43561_, new_n43559_ );
and  ( new_n43563_, new_n26063_, new_n4859_ );
not  ( new_n43564_, new_n43563_ );
and  ( new_n43565_, new_n26196_, new_n4995_ );
not  ( new_n43566_, new_n43565_ );
and  ( new_n43567_, new_n43566_, new_n43564_ );
and  ( new_n43568_, new_n43567_, new_n43562_ );
and  ( new_n43569_, new_n24418_, new_n3178_ );
not  ( new_n43570_, new_n43569_ );
and  ( new_n43571_, new_n24927_, new_n3696_ );
not  ( new_n43572_, new_n43571_ );
and  ( new_n43573_, new_n43572_, new_n43570_ );
and  ( new_n43574_, new_n24543_, new_n3306_ );
not  ( new_n43575_, new_n43574_ );
and  ( new_n43576_, new_n24227_, new_n2981_ );
not  ( new_n43577_, new_n43576_ );
and  ( new_n43578_, new_n43577_, new_n43575_ );
and  ( new_n43579_, new_n43578_, new_n43573_ );
and  ( new_n43580_, new_n24925_, new_n3694_ );
not  ( new_n43581_, new_n43580_ );
and  ( new_n43582_, new_n25486_, new_n4267_ );
not  ( new_n43583_, new_n43582_ );
and  ( new_n43584_, new_n43583_, new_n43581_ );
and  ( new_n43585_, new_n25288_, new_n4069_ );
not  ( new_n43586_, new_n43585_ );
and  ( new_n43587_, new_n25048_, new_n3820_ );
not  ( new_n43588_, new_n43587_ );
and  ( new_n43589_, new_n43588_, new_n43586_ );
and  ( new_n43590_, new_n43589_, new_n43584_ );
and  ( new_n43591_, new_n43590_, new_n43579_ );
and  ( new_n43592_, new_n43591_, new_n43568_ );
and  ( new_n43593_, new_n43592_, new_n43557_ );
and  ( new_n43594_, new_n43593_, new_n43548_ );
not  ( new_n43595_, new_n43594_ );
and  ( new_n43596_, RIbb32a90_173, RIbb2c370_109 );
and  ( new_n43597_, RIbb32bf8_176, RIbb2c208_112 );
and  ( new_n43598_, new_n43597_, new_n43553_ );
not  ( new_n43599_, new_n43598_ );
and  ( new_n43600_, RIbb32b80_175, RIbb2c280_111 );
and  ( new_n43601_, RIbb32b08_174, RIbb2c2f8_110 );
nor  ( new_n43602_, new_n43601_, new_n43600_ );
and  ( new_n43603_, new_n43602_, new_n43599_ );
not  ( new_n43604_, new_n43603_ );
and  ( new_n43605_, new_n43604_, new_n43551_ );
nor  ( new_n43606_, new_n43605_, new_n43596_ );
not  ( new_n43607_, new_n43606_ );
and  ( new_n43608_, RIbb33030_185, RIbb2bdd0_121 );
and  ( new_n43609_, RIbb330a8_186, RIbb2bd58_122 );
and  ( new_n43610_, RIbb33120_187, RIbb2bce0_123 );
and  ( new_n43611_, RIbb33198_188, RIbb2bc68_124 );
nor  ( new_n43612_, new_n43611_, new_n43610_ );
nor  ( new_n43613_, new_n43612_, new_n43516_ );
nor  ( new_n43614_, new_n43613_, new_n43609_ );
not  ( new_n43615_, new_n43614_ );
and  ( new_n43616_, new_n43615_, new_n43515_ );
nor  ( new_n43617_, new_n43616_, new_n43608_ );
not  ( new_n43618_, new_n43617_ );
and  ( new_n43619_, new_n43512_, new_n43504_ );
and  ( new_n43620_, new_n43619_, new_n43618_ );
not  ( new_n43621_, new_n43620_ );
and  ( new_n43622_, RIbb32c70_177, RIbb2c190_113 );
and  ( new_n43623_, RIbb32ce8_178, RIbb2c118_114 );
and  ( new_n43624_, RIbb32d60_179, RIbb2c0a0_115 );
and  ( new_n43625_, RIbb32dd8_180, RIbb2c028_116 );
nor  ( new_n43626_, new_n43625_, new_n43624_ );
nor  ( new_n43627_, new_n43626_, new_n43499_ );
nor  ( new_n43628_, new_n43627_, new_n43623_ );
not  ( new_n43629_, new_n43628_ );
and  ( new_n43630_, new_n43502_, new_n43495_ );
and  ( new_n43631_, new_n43630_, new_n43629_ );
nor  ( new_n43632_, new_n43631_, new_n43622_ );
and  ( new_n43633_, new_n43632_, new_n43621_ );
not  ( new_n43634_, new_n43633_ );
and  ( new_n43635_, new_n43634_, new_n43557_ );
nor  ( new_n43636_, new_n43635_, new_n43607_ );
not  ( new_n43637_, new_n43636_ );
and  ( new_n43638_, new_n43637_, new_n43592_ );
not  ( new_n43639_, new_n43638_ );
and  ( new_n43640_, RIbb328b0_169, RIbb2c550_105 );
and  ( new_n43641_, RIbb32928_170, RIbb2c4d8_106 );
and  ( new_n43642_, RIbb329a0_171, RIbb2c460_107 );
and  ( new_n43643_, RIbb32a18_172, RIbb2c3e8_108 );
nor  ( new_n43644_, new_n43643_, new_n43642_ );
nor  ( new_n43645_, new_n43644_, new_n43563_ );
nor  ( new_n43646_, new_n43645_, new_n43641_ );
not  ( new_n43647_, new_n43646_ );
and  ( new_n43648_, new_n43566_, new_n43559_ );
and  ( new_n43649_, new_n43648_, new_n43647_ );
nor  ( new_n43650_, new_n43649_, new_n43640_ );
not  ( new_n43651_, new_n43650_ );
and  ( new_n43652_, new_n43651_, new_n43590_ );
and  ( new_n43653_, RIbb326d0_165, RIbb2c730_101 );
and  ( new_n43654_, RIbb32748_166, RIbb2c6b8_102 );
and  ( new_n43655_, RIbb327c0_167, RIbb2c640_103 );
and  ( new_n43656_, RIbb32838_168, RIbb2c5c8_104 );
nor  ( new_n43657_, new_n43656_, new_n43655_ );
nor  ( new_n43658_, new_n43657_, new_n43585_ );
nor  ( new_n43659_, new_n43658_, new_n43654_ );
not  ( new_n43660_, new_n43659_ );
and  ( new_n43661_, new_n43588_, new_n43581_ );
and  ( new_n43662_, new_n43661_, new_n43660_ );
nor  ( new_n43663_, new_n43662_, new_n43653_ );
not  ( new_n43664_, new_n43663_ );
nor  ( new_n43665_, new_n43664_, new_n43652_ );
not  ( new_n43666_, new_n43665_ );
and  ( new_n43667_, new_n43666_, new_n43579_ );
not  ( new_n43668_, new_n43667_ );
and  ( new_n43669_, RIbb32568_162, RIbb2c898_98 );
and  ( new_n43670_, RIbb325e0_163, RIbb2c820_99 );
and  ( new_n43671_, RIbb32658_164, RIbb2c7a8_100 );
nor  ( new_n43672_, new_n43671_, new_n43670_ );
nor  ( new_n43673_, new_n43672_, new_n43574_ );
nor  ( new_n43674_, new_n43673_, new_n43669_ );
not  ( new_n43675_, new_n43674_ );
and  ( new_n43676_, new_n43577_, new_n43570_ );
and  ( new_n43677_, new_n43676_, new_n43675_ );
and  ( new_n43678_, RIbb324f0_161, RIbb2c910_97 );
nor  ( new_n43679_, new_n43678_, new_n43677_ );
and  ( new_n43680_, new_n43679_, new_n43668_ );
and  ( new_n43681_, new_n43680_, new_n43639_ );
and  ( new_n43682_, new_n43681_, new_n43595_ );
nor  ( new_n43683_, new_n43682_, new_n43493_ );
and  ( new_n43684_, new_n43683_, new_n43492_ );
and  ( new_n43685_, new_n43684_, new_n43490_ );
and  ( new_n43686_, new_n23166_, new_n1899_ );
and  ( new_n43687_, new_n22973_, new_n1754_ );
nor  ( new_n43688_, new_n43687_, new_n43686_ );
and  ( new_n43689_, new_n23252_, new_n2057_ );
not  ( new_n43690_, new_n43689_ );
and  ( new_n43691_, new_n23370_, new_n2178_ );
not  ( new_n43692_, new_n43691_ );
and  ( new_n43693_, new_n43692_, new_n43690_ );
and  ( new_n43694_, new_n43693_, new_n43688_ );
and  ( new_n43695_, new_n43694_, new_n43685_ );
not  ( new_n43696_, new_n43695_ );
and  ( new_n43697_, RIbb32310_157, RIbb2caf0_93 );
and  ( new_n43698_, RIbb32388_158, RIbb2ca78_94 );
and  ( new_n43699_, RIbb32400_159, RIbb2ca00_95 );
and  ( new_n43700_, RIbb32478_160, RIbb2c988_96 );
nor  ( new_n43701_, new_n43700_, new_n43699_ );
nor  ( new_n43702_, new_n43701_, new_n43491_ );
nor  ( new_n43703_, new_n43702_, new_n43698_ );
not  ( new_n43704_, new_n43703_ );
and  ( new_n43705_, new_n43704_, new_n43490_ );
nor  ( new_n43706_, new_n43705_, new_n43697_ );
not  ( new_n43707_, new_n43706_ );
and  ( new_n43708_, new_n43707_, new_n43694_ );
not  ( new_n43709_, new_n43708_ );
and  ( new_n43710_, RIbb321a8_154, RIbb2cc58_90 );
and  ( new_n43711_, RIbb32220_155, RIbb2cbe0_91 );
and  ( new_n43712_, RIbb32298_156, RIbb2cb68_92 );
nor  ( new_n43713_, new_n43712_, new_n43711_ );
nor  ( new_n43714_, new_n43713_, new_n43689_ );
nor  ( new_n43715_, new_n43714_, new_n43710_ );
not  ( new_n43716_, new_n43715_ );
and  ( new_n43717_, new_n43716_, new_n43688_ );
and  ( new_n43718_, RIbb32130_153, RIbb2ccd0_89 );
nor  ( new_n43719_, new_n43718_, new_n43717_ );
and  ( new_n43720_, new_n43719_, new_n43709_ );
and  ( new_n43721_, new_n43720_, new_n43696_ );
nor  ( new_n43722_, new_n43721_, new_n43487_ );
and  ( new_n43723_, new_n43722_, new_n43486_ );
and  ( new_n43724_, new_n22641_, new_n1318_ );
and  ( new_n43725_, new_n22590_, new_n1213_ );
nor  ( new_n43726_, new_n43725_, new_n43724_ );
and  ( new_n43727_, new_n43726_, new_n43723_ );
and  ( new_n43728_, new_n43727_, new_n43484_ );
not  ( new_n43729_, new_n43728_ );
and  ( new_n43730_, RIbb31f50_149, RIbb2ceb0_85 );
and  ( new_n43731_, RIbb31fc8_150, RIbb2ce38_86 );
and  ( new_n43732_, RIbb32040_151, RIbb2cdc0_87 );
and  ( new_n43733_, RIbb320b8_152, RIbb2cd48_88 );
nor  ( new_n43734_, new_n43733_, new_n43732_ );
nor  ( new_n43735_, new_n43734_, new_n43485_ );
nor  ( new_n43736_, new_n43735_, new_n43731_ );
not  ( new_n43737_, new_n43736_ );
and  ( new_n43738_, new_n43737_, new_n43726_ );
nor  ( new_n43739_, new_n43738_, new_n43730_ );
not  ( new_n43740_, new_n43739_ );
and  ( new_n43741_, new_n43740_, new_n43484_ );
not  ( new_n43742_, new_n43741_ );
and  ( new_n43743_, RIbb31d70_145, RIbb2d090_81 );
and  ( new_n43744_, RIbb31de8_146, RIbb2d018_82 );
and  ( new_n43745_, RIbb31e60_147, RIbb2cfa0_83 );
and  ( new_n43746_, RIbb31ed8_148, RIbb2cf28_84 );
nor  ( new_n43747_, new_n43746_, new_n43745_ );
not  ( new_n43748_, new_n43747_ );
and  ( new_n43749_, new_n43748_, new_n43482_ );
nor  ( new_n43750_, new_n43749_, new_n43744_ );
nor  ( new_n43751_, new_n43750_, new_n43476_ );
nor  ( new_n43752_, new_n43751_, new_n43743_ );
and  ( new_n43753_, new_n43752_, new_n43742_ );
and  ( new_n43754_, new_n43753_, new_n43729_ );
nor  ( new_n43755_, new_n43754_, new_n43475_ );
nor  ( new_n43756_, new_n43755_, new_n43474_ );
nor  ( new_n43757_, new_n43756_, new_n43473_ );
nor  ( new_n43758_, new_n43757_, new_n43472_ );
nor  ( new_n43759_, new_n43758_, new_n43471_ );
nor  ( new_n43760_, new_n43759_, new_n43470_ );
nor  ( new_n43761_, new_n43760_, new_n43469_ );
nor  ( new_n43762_, new_n43761_, new_n43468_ );
nor  ( new_n43763_, new_n43762_, new_n43467_ );
nor  ( new_n43764_, new_n43763_, new_n43466_ );
nor  ( new_n43765_, new_n43764_, new_n43465_ );
nor  ( new_n43766_, new_n43765_, new_n43464_ );
nor  ( new_n43767_, new_n43766_, new_n43463_ );
nor  ( new_n43768_, new_n43767_, new_n43462_ );
nor  ( new_n43769_, new_n43768_, new_n43461_ );
nor  ( new_n43770_, new_n43769_, new_n43460_ );
nor  ( new_n43771_, new_n43770_, new_n43459_ );
nor  ( new_n43772_, new_n43771_, new_n43458_ );
and  ( new_n43773_, new_n21680_, new_n301_ );
nor  ( new_n43774_, new_n43773_, new_n43772_ );
nor  ( new_n43775_, new_n43774_, new_n43457_ );
nor  ( new_n43776_, new_n43775_, new_n43456_ );
nor  ( new_n43777_, new_n43776_, new_n43455_ );
and  ( new_n43778_, new_n21674_, new_n285_ );
nor  ( new_n43779_, new_n43778_, new_n43777_ );
nor  ( new_n43780_, new_n43779_, new_n43454_ );
nor  ( new_n43781_, new_n43780_, new_n43453_ );
nor  ( new_n43782_, new_n43781_, new_n43452_ );
nor  ( new_n43783_, new_n43782_, new_n43451_ );
nor  ( new_n43784_, new_n43783_, new_n43450_ );
nor  ( new_n43785_, new_n43784_, new_n43449_ );
nor  ( new_n43786_, new_n43785_, new_n43448_ );
xnor ( new_n43787_, new_n43786_, new_n43447_ );
xor  ( new_n43788_, new_n43787_, RIbb2f160_11 );
nand ( new_n43789_, new_n43788_, new_n373_ );
and  ( new_n43790_, RIbb315f0_129, RIbb2d810_65 );
and  ( new_n43791_, new_n21696_, new_n339_ );
nor  ( new_n43792_, new_n43786_, new_n43791_ );
nor  ( new_n43793_, new_n43792_, new_n43790_ );
xor  ( new_n43794_, new_n43793_, RIbb2f160_11 );
or   ( new_n43795_, new_n43794_, new_n411_ );
and  ( new_n43796_, new_n43795_, new_n43789_ );
nor  ( new_n43797_, new_n43796_, new_n402_ );
xor  ( new_n43798_, RIbb31758_132, new_n313_ );
xor  ( new_n43799_, new_n43798_, new_n43780_ );
xor  ( new_n43800_, new_n43799_, new_n309_ );
nor  ( new_n43801_, new_n43800_, new_n320_ );
xor  ( new_n43802_, RIbb317d0_133, RIbb2d630_69 );
xnor ( new_n43803_, new_n43802_, new_n43777_ );
xor  ( new_n43804_, new_n43803_, RIbb2f340_7 );
and  ( new_n43805_, new_n43804_, new_n316_ );
or   ( new_n43806_, new_n43805_, new_n43801_ );
xor  ( new_n43807_, new_n43796_, new_n402_ );
and  ( new_n43808_, new_n43807_, new_n43806_ );
nor  ( new_n43809_, new_n43808_, new_n43797_ );
not  ( new_n43810_, new_n43809_ );
xor  ( new_n43811_, RIbb31b18_140, RIbb2d2e8_76 );
xnor ( new_n43812_, new_n43811_, new_n43762_ );
and  ( new_n43813_, new_n1318_, new_n1213_ );
and  ( new_n43814_, new_n1523_, new_n1525_ );
and  ( new_n43815_, new_n43814_, new_n43813_ );
and  ( new_n43816_, new_n886_, new_n805_ );
and  ( new_n43817_, new_n1168_, new_n986_ );
and  ( new_n43818_, new_n43817_, new_n43816_ );
and  ( new_n43819_, new_n43818_, new_n43815_ );
and  ( new_n43820_, new_n2475_, new_n2291_ );
and  ( new_n43821_, new_n2751_, new_n2646_ );
and  ( new_n43822_, new_n43821_, new_n43820_ );
and  ( new_n43823_, new_n1899_, new_n1754_ );
and  ( new_n43824_, new_n2178_, new_n2057_ );
and  ( new_n43825_, new_n43824_, new_n43823_ );
and  ( new_n43826_, new_n43825_, new_n43822_ );
and  ( new_n43827_, new_n43826_, new_n43819_ );
and  ( new_n43828_, new_n285_, new_n279_ );
and  ( new_n43829_, new_n301_, new_n294_ );
and  ( new_n43830_, new_n43829_, new_n43828_ );
and  ( new_n43831_, new_n339_, new_n333_ );
and  ( new_n43832_, new_n319_, new_n313_ );
and  ( new_n43833_, new_n43832_, new_n43831_ );
and  ( new_n43834_, new_n43833_, new_n43830_ );
and  ( new_n43835_, new_n509_, new_n443_ );
and  ( new_n43836_, new_n775_, new_n515_ );
and  ( new_n43837_, new_n43836_, new_n43835_ );
and  ( new_n43838_, new_n270_, new_n264_ );
and  ( new_n43839_, new_n348_, new_n419_ );
and  ( new_n43840_, new_n43839_, new_n43838_ );
and  ( new_n43841_, new_n43840_, new_n43837_ );
and  ( new_n43842_, new_n43841_, new_n43834_ );
and  ( new_n43843_, new_n43842_, new_n43827_ );
and  ( new_n43844_, RIbb2bf38_118, new_n7373_ );
and  ( new_n43845_, RIbb2be48_120, RIbb2bec0_119 );
and  ( new_n43846_, new_n43845_, new_n43844_ );
and  ( new_n43847_, new_n6589_, new_n6425_ );
and  ( new_n43848_, new_n7149_, new_n6943_ );
and  ( new_n43849_, new_n43848_, new_n43847_ );
and  ( new_n43850_, new_n43849_, new_n43846_ );
and  ( new_n43851_, RIbb2bb78_126, new_n9679_ );
and  ( new_n43852_, new_n10841_, new_n10541_ );
and  ( new_n43853_, new_n43852_, new_n43851_ );
and  ( new_n43854_, RIbb2bd58_122, RIbb2bdd0_121 );
and  ( new_n43855_, new_n9681_, RIbb2bce0_123 );
and  ( new_n43856_, new_n43855_, new_n43854_ );
and  ( new_n43857_, new_n43856_, new_n43853_ );
and  ( new_n43858_, new_n43857_, new_n43850_ );
and  ( new_n43859_, new_n3820_, new_n3694_ );
and  ( new_n43860_, new_n4267_, new_n4069_ );
and  ( new_n43861_, new_n43860_, new_n43859_ );
and  ( new_n43862_, new_n3178_, new_n2981_ );
and  ( new_n43863_, new_n3696_, new_n3306_ );
and  ( new_n43864_, new_n43863_, new_n43862_ );
and  ( new_n43865_, new_n43864_, new_n43861_ );
and  ( new_n43866_, new_n5570_, new_n5428_ );
and  ( new_n43867_, new_n6219_, new_n5899_ );
and  ( new_n43868_, new_n43867_, new_n43866_ );
and  ( new_n43869_, new_n4995_, new_n4603_ );
and  ( new_n43870_, new_n5171_, new_n4859_ );
and  ( new_n43871_, new_n43870_, new_n43869_ );
and  ( new_n43872_, new_n43871_, new_n43868_ );
and  ( new_n43873_, new_n43872_, new_n43865_ );
and  ( new_n43874_, new_n43873_, new_n43858_ );
and  ( new_n43875_, new_n43874_, new_n43843_ );
not  ( new_n43876_, new_n43875_ );
and  ( new_n43877_, new_n43876_, RIbb2f610_1 );
and  ( new_n43878_, new_n43875_, RIbb2f598_2 );
nor  ( new_n43879_, new_n43878_, new_n43877_ );
not  ( new_n43880_, new_n43879_ );
and  ( new_n43881_, new_n43880_, new_n43812_ );
not  ( new_n43882_, new_n43881_ );
xor  ( new_n43883_, RIbb31848_134, RIbb2d5b8_70 );
xnor ( new_n43884_, new_n43883_, new_n43775_ );
xor  ( new_n43885_, new_n43884_, new_n275_ );
or   ( new_n43886_, new_n43885_, new_n286_ );
xor  ( new_n43887_, RIbb318c0_135, RIbb2d540_71 );
xnor ( new_n43888_, new_n43887_, new_n43772_ );
xor  ( new_n43889_, new_n43888_, new_n275_ );
or   ( new_n43890_, new_n43889_, new_n283_ );
and  ( new_n43891_, new_n43890_, new_n43886_ );
nor  ( new_n43892_, new_n43891_, new_n43882_ );
xor  ( new_n43893_, RIbb316e0_131, RIbb2d720_67 );
xnor ( new_n43894_, new_n43893_, new_n43782_ );
xor  ( new_n43895_, new_n43894_, RIbb2f250_9 );
and  ( new_n43896_, new_n43895_, new_n336_ );
xor  ( new_n43897_, RIbb31668_130, new_n333_ );
xor  ( new_n43898_, new_n43897_, new_n43784_ );
xor  ( new_n43899_, new_n43898_, new_n329_ );
nor  ( new_n43900_, new_n43899_, new_n340_ );
or   ( new_n43901_, new_n43900_, new_n43896_ );
xor  ( new_n43902_, new_n43891_, new_n43882_ );
and  ( new_n43903_, new_n43902_, new_n43901_ );
or   ( new_n43904_, new_n43903_, new_n43892_ );
not  ( new_n43905_, RIbb2f0e8_12 );
and  ( new_n43906_, new_n43905_, new_n400_ );
or   ( new_n43907_, new_n43906_, new_n328_ );
or   ( new_n43908_, new_n43794_, new_n409_ );
and  ( new_n43909_, new_n43908_, new_n43907_ );
xor  ( new_n43910_, new_n43909_, new_n43904_ );
xor  ( new_n43911_, new_n43910_, new_n43810_ );
not  ( new_n43912_, new_n43911_ );
xor  ( new_n43913_, RIbb31b90_141, RIbb2d270_77 );
xnor ( new_n43914_, new_n43913_, new_n43760_ );
and  ( new_n43915_, new_n43914_, new_n43880_ );
not  ( new_n43916_, new_n43915_ );
xor  ( new_n43917_, new_n43884_, new_n309_ );
or   ( new_n43918_, new_n43917_, new_n317_ );
nand ( new_n43919_, new_n43804_, new_n314_ );
and  ( new_n43920_, new_n43919_, new_n43918_ );
nor  ( new_n43921_, new_n43920_, new_n43916_ );
and  ( new_n43922_, new_n43788_, new_n371_ );
xor  ( new_n43923_, new_n43898_, new_n325_ );
nor  ( new_n43924_, new_n43923_, new_n409_ );
or   ( new_n43925_, new_n43924_, new_n43922_ );
xor  ( new_n43926_, new_n43920_, new_n43916_ );
and  ( new_n43927_, new_n43926_, new_n43925_ );
or   ( new_n43928_, new_n43927_, new_n43921_ );
xor  ( new_n43929_, new_n43807_, new_n43806_ );
nand ( new_n43930_, new_n43929_, new_n43928_ );
nor  ( new_n43931_, new_n43929_, new_n43928_ );
xor  ( new_n43932_, new_n43799_, new_n329_ );
or   ( new_n43933_, new_n43932_, new_n337_ );
nand ( new_n43934_, new_n43895_, new_n334_ );
and  ( new_n43935_, new_n43934_, new_n43933_ );
xor  ( new_n43936_, RIbb31938_136, RIbb2d4c8_72 );
xnor ( new_n43937_, new_n43936_, new_n43770_ );
xor  ( new_n43938_, new_n43937_, new_n275_ );
or   ( new_n43939_, new_n43938_, new_n283_ );
or   ( new_n43940_, new_n43889_, new_n286_ );
and  ( new_n43941_, new_n43940_, new_n43939_ );
or   ( new_n43942_, new_n43941_, new_n43935_ );
and  ( new_n43943_, new_n43876_, RIbb2f520_3 );
and  ( new_n43944_, new_n43875_, RIbb32fb8_184 );
nor  ( new_n43945_, new_n43944_, new_n43943_ );
and  ( new_n43946_, new_n43945_, new_n291_ );
nor  ( new_n43947_, RIbb2f4a8_4, RIbb2f430_5 );
nor  ( new_n43948_, new_n43945_, new_n43947_ );
nor  ( new_n43949_, new_n43948_, new_n43946_ );
not  ( new_n43950_, new_n43945_ );
xor  ( new_n43951_, RIbb31a28_138, RIbb2d3d8_74 );
xnor ( new_n43952_, new_n43951_, new_n43766_ );
xor  ( new_n43953_, new_n43952_, new_n43950_ );
and  ( new_n43954_, new_n43953_, new_n43949_ );
xor  ( new_n43955_, RIbb319b0_137, new_n270_ );
xor  ( new_n43956_, new_n43955_, new_n43768_ );
xor  ( new_n43957_, new_n43956_, new_n43945_ );
not  ( new_n43958_, new_n43957_ );
and  ( new_n43959_, new_n43958_, new_n295_ );
or   ( new_n43960_, new_n43959_, new_n43954_ );
xor  ( new_n43961_, new_n43941_, new_n43935_ );
nand ( new_n43962_, new_n43961_, new_n43960_ );
and  ( new_n43963_, new_n43962_, new_n43942_ );
or   ( new_n43964_, new_n43963_, new_n43931_ );
and  ( new_n43965_, new_n43964_, new_n43930_ );
nor  ( new_n43966_, new_n43965_, new_n43912_ );
xor  ( new_n43967_, new_n43965_, new_n43912_ );
nor  ( new_n43968_, RIbb2ef80_15, RIbb2eff8_14 );
not  ( new_n43969_, new_n43968_ );
and  ( new_n43970_, new_n43969_, new_n402_ );
xor  ( new_n43971_, new_n43793_, new_n400_ );
and  ( new_n43972_, new_n43971_, new_n456_ );
nor  ( new_n43973_, new_n43972_, new_n43970_ );
nand ( new_n43974_, new_n43876_, RIbb2f598_2 );
or   ( new_n43975_, new_n43876_, new_n296_ );
and  ( new_n43976_, new_n43975_, new_n43974_ );
xor  ( new_n43977_, new_n43976_, new_n43950_ );
not  ( new_n43978_, new_n43977_ );
xor  ( new_n43979_, new_n43952_, new_n43880_ );
nand ( new_n43980_, new_n43979_, new_n43978_ );
xor  ( new_n43981_, new_n43945_, new_n43880_ );
nor  ( new_n43982_, new_n43981_, new_n43978_ );
not  ( new_n43983_, new_n43982_ );
xor  ( new_n43984_, RIbb31aa0_139, RIbb2d360_75 );
xnor ( new_n43985_, new_n43984_, new_n43764_ );
xor  ( new_n43986_, new_n43985_, new_n43945_ );
not  ( new_n43987_, new_n43986_ );
or   ( new_n43988_, new_n43987_, new_n43983_ );
and  ( new_n43989_, new_n43988_, new_n43980_ );
nor  ( new_n43990_, new_n43989_, new_n43973_ );
and  ( new_n43991_, new_n43958_, new_n43949_ );
xor  ( new_n43992_, new_n43945_, new_n43937_ );
nor  ( new_n43993_, new_n43992_, new_n302_ );
nor  ( new_n43994_, new_n43993_, new_n43991_ );
not  ( new_n43995_, new_n43994_ );
xor  ( new_n43996_, new_n43989_, new_n43973_ );
and  ( new_n43997_, new_n43996_, new_n43995_ );
or   ( new_n43998_, new_n43997_, new_n43990_ );
nor  ( new_n43999_, new_n43899_, new_n337_ );
xor  ( new_n44000_, new_n43787_, RIbb2f250_9 );
and  ( new_n44001_, new_n44000_, new_n334_ );
or   ( new_n44002_, new_n44001_, new_n43999_ );
or   ( new_n44003_, new_n43885_, new_n283_ );
xor  ( new_n44004_, new_n43803_, new_n275_ );
or   ( new_n44005_, new_n44004_, new_n286_ );
and  ( new_n44006_, new_n44005_, new_n44003_ );
not  ( new_n44007_, new_n43949_ );
or   ( new_n44008_, new_n43992_, new_n44007_ );
xor  ( new_n44009_, new_n43945_, new_n43888_ );
or   ( new_n44010_, new_n44009_, new_n302_ );
and  ( new_n44011_, new_n44010_, new_n44008_ );
xor  ( new_n44012_, new_n44011_, new_n44006_ );
xor  ( new_n44013_, new_n44012_, new_n44002_ );
xor  ( new_n44014_, new_n44013_, new_n43998_ );
and  ( new_n44015_, new_n43982_, new_n43979_ );
xor  ( new_n44016_, new_n43956_, new_n43880_ );
and  ( new_n44017_, new_n44016_, new_n43978_ );
or   ( new_n44018_, new_n44017_, new_n44015_ );
and  ( new_n44019_, new_n43985_, new_n43880_ );
not  ( new_n44020_, new_n44019_ );
or   ( new_n44021_, new_n43800_, new_n317_ );
xor  ( new_n44022_, new_n43894_, RIbb2f340_7 );
nand ( new_n44023_, new_n44022_, new_n314_ );
and  ( new_n44024_, new_n44023_, new_n44021_ );
xor  ( new_n44025_, new_n44024_, new_n44020_ );
xor  ( new_n44026_, new_n44025_, new_n44018_ );
xor  ( new_n44027_, new_n44026_, new_n44014_ );
and  ( new_n44028_, new_n44027_, new_n43967_ );
nor  ( new_n44029_, new_n44028_, new_n43966_ );
not  ( new_n44030_, new_n44029_ );
or   ( new_n44031_, new_n44024_, new_n44020_ );
nand ( new_n44032_, new_n44025_, new_n44018_ );
nand ( new_n44033_, new_n44032_, new_n44031_ );
xor  ( new_n44034_, new_n43799_, new_n275_ );
or   ( new_n44035_, new_n44034_, new_n286_ );
or   ( new_n44036_, new_n44004_, new_n283_ );
and  ( new_n44037_, new_n44036_, new_n44035_ );
nand ( new_n44038_, new_n44000_, new_n336_ );
xor  ( new_n44039_, new_n43793_, RIbb2f250_9 );
or   ( new_n44040_, new_n44039_, new_n340_ );
and  ( new_n44041_, new_n44040_, new_n44038_ );
xor  ( new_n44042_, new_n44041_, new_n327_ );
xnor ( new_n44043_, new_n44042_, new_n44037_ );
xor  ( new_n44044_, new_n44043_, new_n44033_ );
nor  ( new_n44045_, new_n44009_, new_n44007_ );
xor  ( new_n44046_, new_n43945_, new_n43884_ );
nor  ( new_n44047_, new_n44046_, new_n302_ );
or   ( new_n44048_, new_n44047_, new_n44045_ );
xor  ( new_n44049_, new_n43937_, new_n43879_ );
nor  ( new_n44050_, new_n44049_, new_n43977_ );
and  ( new_n44051_, new_n44016_, new_n43982_ );
nor  ( new_n44052_, new_n44051_, new_n44050_ );
and  ( new_n44053_, new_n44022_, new_n316_ );
xor  ( new_n44054_, new_n43898_, new_n309_ );
nor  ( new_n44055_, new_n44054_, new_n320_ );
nor  ( new_n44056_, new_n44055_, new_n44053_ );
xor  ( new_n44057_, new_n44056_, new_n44052_ );
xor  ( new_n44058_, new_n44057_, new_n44048_ );
xor  ( new_n44059_, new_n44058_, new_n44044_ );
and  ( new_n44060_, new_n44059_, new_n44030_ );
xor  ( new_n44061_, new_n44059_, new_n44030_ );
and  ( new_n44062_, new_n44013_, new_n43998_ );
and  ( new_n44063_, new_n44026_, new_n44014_ );
nor  ( new_n44064_, new_n44063_, new_n44062_ );
and  ( new_n44065_, new_n43909_, new_n43904_ );
and  ( new_n44066_, new_n43910_, new_n43810_ );
or   ( new_n44067_, new_n44066_, new_n44065_ );
or   ( new_n44068_, new_n44011_, new_n44006_ );
nand ( new_n44069_, new_n44012_, new_n44002_ );
nand ( new_n44070_, new_n44069_, new_n44068_ );
and  ( new_n44071_, new_n43952_, new_n43880_ );
xnor ( new_n44072_, new_n44071_, new_n43909_ );
xor  ( new_n44073_, new_n44072_, new_n44070_ );
xor  ( new_n44074_, new_n44073_, new_n44067_ );
xnor ( new_n44075_, new_n44074_, new_n44064_ );
and  ( new_n44076_, new_n44075_, new_n44061_ );
nor  ( new_n44077_, new_n44076_, new_n44060_ );
or   ( new_n44078_, new_n44046_, new_n44007_ );
nor  ( new_n44079_, new_n43950_, new_n43803_ );
and  ( new_n44080_, new_n43950_, new_n43803_ );
or   ( new_n44081_, new_n44080_, new_n302_ );
or   ( new_n44082_, new_n44081_, new_n44079_ );
and  ( new_n44083_, new_n44082_, new_n44078_ );
or   ( new_n44084_, new_n44049_, new_n43983_ );
and  ( new_n44085_, new_n43888_, new_n43880_ );
nor  ( new_n44086_, new_n43888_, new_n43880_ );
or   ( new_n44087_, new_n44086_, new_n43977_ );
or   ( new_n44088_, new_n44087_, new_n44085_ );
and  ( new_n44089_, new_n44088_, new_n44084_ );
xor  ( new_n44090_, new_n44089_, new_n44083_ );
and  ( new_n44091_, new_n43956_, new_n43880_ );
or   ( new_n44092_, new_n44039_, new_n337_ );
and  ( new_n44093_, new_n44092_, new_n13845_ );
xor  ( new_n44094_, new_n44093_, new_n44091_ );
or   ( new_n44095_, new_n44041_, new_n327_ );
not  ( new_n44096_, new_n44037_ );
nand ( new_n44097_, new_n44042_, new_n44096_ );
and  ( new_n44098_, new_n44097_, new_n44095_ );
xor  ( new_n44099_, new_n44098_, new_n44094_ );
nor  ( new_n44100_, new_n44056_, new_n44052_ );
and  ( new_n44101_, new_n44057_, new_n44048_ );
or   ( new_n44102_, new_n44101_, new_n44100_ );
or   ( new_n44103_, new_n44034_, new_n283_ );
not  ( new_n44104_, new_n43894_ );
and  ( new_n44105_, new_n44104_, new_n275_ );
and  ( new_n44106_, new_n43894_, RIbb2f430_5 );
or   ( new_n44107_, new_n44106_, new_n286_ );
or   ( new_n44108_, new_n44107_, new_n44105_ );
and  ( new_n44109_, new_n44108_, new_n44103_ );
xor  ( new_n44110_, new_n44109_, new_n44102_ );
xor  ( new_n44111_, new_n44110_, new_n44099_ );
xor  ( new_n44112_, new_n44111_, new_n44090_ );
nand ( new_n44113_, new_n44043_, new_n44033_ );
nand ( new_n44114_, new_n44058_, new_n44044_ );
and  ( new_n44115_, new_n44114_, new_n44113_ );
or   ( new_n44116_, new_n44054_, new_n317_ );
nor  ( new_n44117_, new_n43787_, RIbb2f340_7 );
and  ( new_n44118_, new_n43787_, RIbb2f340_7 );
or   ( new_n44119_, new_n44118_, new_n320_ );
or   ( new_n44120_, new_n44119_, new_n44117_ );
and  ( new_n44121_, new_n44120_, new_n44116_ );
xor  ( new_n44122_, new_n44121_, new_n44115_ );
not  ( new_n44123_, new_n43909_ );
nand ( new_n44124_, new_n44071_, new_n44123_ );
nand ( new_n44125_, new_n44072_, new_n44070_ );
and  ( new_n44126_, new_n44125_, new_n44124_ );
xor  ( new_n44127_, new_n44126_, new_n44122_ );
xor  ( new_n44128_, new_n44127_, new_n44112_ );
xnor ( new_n44129_, new_n44128_, new_n44077_ );
and  ( new_n44130_, new_n44073_, new_n44067_ );
nor  ( new_n44131_, new_n44073_, new_n44067_ );
nor  ( new_n44132_, new_n44131_, new_n44064_ );
nor  ( new_n44133_, new_n44132_, new_n44130_ );
xnor ( new_n44134_, new_n44027_, new_n43967_ );
not  ( new_n44135_, new_n43973_ );
xor  ( new_n44136_, new_n43945_, new_n43812_ );
not  ( new_n44137_, new_n44136_ );
or   ( new_n44138_, new_n44137_, new_n43983_ );
not  ( new_n44139_, new_n43985_ );
and  ( new_n44140_, new_n44139_, new_n43879_ );
or   ( new_n44141_, new_n44019_, new_n43977_ );
or   ( new_n44142_, new_n44141_, new_n44140_ );
and  ( new_n44143_, new_n44142_, new_n44138_ );
nor  ( new_n44144_, new_n44143_, new_n44135_ );
xor  ( new_n44145_, new_n43787_, new_n400_ );
or   ( new_n44146_, new_n44145_, new_n524_ );
nand ( new_n44147_, new_n43971_, new_n454_ );
and  ( new_n44148_, new_n44147_, new_n44146_ );
nor  ( new_n44149_, new_n44148_, new_n522_ );
xor  ( new_n44150_, new_n43803_, RIbb2f250_9 );
and  ( new_n44151_, new_n44150_, new_n336_ );
nor  ( new_n44152_, new_n43932_, new_n340_ );
or   ( new_n44153_, new_n44152_, new_n44151_ );
xor  ( new_n44154_, new_n44148_, new_n522_ );
and  ( new_n44155_, new_n44154_, new_n44153_ );
or   ( new_n44156_, new_n44155_, new_n44149_ );
xor  ( new_n44157_, new_n44143_, new_n44135_ );
and  ( new_n44158_, new_n44157_, new_n44156_ );
or   ( new_n44159_, new_n44158_, new_n44144_ );
xor  ( new_n44160_, new_n43902_, new_n43901_ );
nand ( new_n44161_, new_n44160_, new_n44159_ );
or   ( new_n44162_, new_n44160_, new_n44159_ );
xor  ( new_n44163_, new_n43996_, new_n43995_ );
nand ( new_n44164_, new_n44163_, new_n44162_ );
and  ( new_n44165_, new_n44164_, new_n44161_ );
or   ( new_n44166_, new_n44165_, new_n44134_ );
or   ( new_n44167_, new_n43938_, new_n286_ );
xor  ( new_n44168_, new_n43956_, new_n275_ );
or   ( new_n44169_, new_n44168_, new_n283_ );
and  ( new_n44170_, new_n44169_, new_n44167_ );
xor  ( new_n44171_, new_n43894_, new_n325_ );
or   ( new_n44172_, new_n44171_, new_n409_ );
or   ( new_n44173_, new_n43923_, new_n411_ );
and  ( new_n44174_, new_n44173_, new_n44172_ );
or   ( new_n44175_, new_n44174_, new_n44170_ );
and  ( new_n44176_, new_n43953_, new_n295_ );
and  ( new_n44177_, new_n43987_, new_n43949_ );
or   ( new_n44178_, new_n44177_, new_n44176_ );
xor  ( new_n44179_, new_n44174_, new_n44170_ );
nand ( new_n44180_, new_n44179_, new_n44178_ );
and  ( new_n44181_, new_n44180_, new_n44175_ );
xor  ( new_n44182_, RIbb31c08_142, RIbb2d1f8_78 );
xnor ( new_n44183_, new_n44182_, new_n43758_ );
and  ( new_n44184_, new_n44183_, new_n43880_ );
xor  ( new_n44185_, new_n43888_, RIbb2f340_7 );
nand ( new_n44186_, new_n44185_, new_n316_ );
or   ( new_n44187_, new_n43917_, new_n320_ );
nand ( new_n44188_, new_n44187_, new_n44186_ );
nand ( new_n44189_, new_n44188_, new_n44184_ );
xnor ( new_n44190_, new_n44188_, new_n44184_ );
not  ( new_n44191_, new_n43914_ );
xor  ( new_n44192_, new_n43945_, new_n44191_ );
or   ( new_n44193_, new_n44192_, new_n43983_ );
nor  ( new_n44194_, new_n43880_, new_n43812_ );
or   ( new_n44195_, new_n43977_, new_n43881_ );
or   ( new_n44196_, new_n44195_, new_n44194_ );
and  ( new_n44197_, new_n44196_, new_n44193_ );
or   ( new_n44198_, new_n44197_, new_n44190_ );
and  ( new_n44199_, new_n44198_, new_n44189_ );
or   ( new_n44200_, new_n44199_, new_n44181_ );
xor  ( new_n44201_, new_n43961_, new_n43960_ );
xor  ( new_n44202_, new_n44199_, new_n44181_ );
nand ( new_n44203_, new_n44202_, new_n44201_ );
and  ( new_n44204_, new_n44203_, new_n44200_ );
xor  ( new_n44205_, new_n43929_, new_n43928_ );
xor  ( new_n44206_, new_n44205_, new_n43963_ );
nor  ( new_n44207_, new_n44206_, new_n44204_ );
xor  ( new_n44208_, new_n43926_, new_n43925_ );
xor  ( new_n44209_, new_n44157_, new_n44156_ );
and  ( new_n44210_, new_n44209_, new_n44208_ );
not  ( new_n44211_, RIbb2ef08_16 );
and  ( new_n44212_, new_n745_, new_n44211_ );
nor  ( new_n44213_, new_n44212_, new_n523_ );
xor  ( new_n44214_, new_n43793_, new_n520_ );
and  ( new_n44215_, new_n44214_, new_n662_ );
nor  ( new_n44216_, new_n44215_, new_n44213_ );
xor  ( new_n44217_, RIbb31c80_143, RIbb2d180_79 );
xnor ( new_n44218_, new_n44217_, new_n43756_ );
and  ( new_n44219_, new_n44218_, new_n43880_ );
xor  ( new_n44220_, new_n43884_, new_n329_ );
or   ( new_n44221_, new_n44220_, new_n337_ );
nand ( new_n44222_, new_n44150_, new_n334_ );
nand ( new_n44223_, new_n44222_, new_n44221_ );
nand ( new_n44224_, new_n44223_, new_n44219_ );
xnor ( new_n44225_, new_n44223_, new_n44219_ );
xor  ( new_n44226_, new_n44183_, new_n43950_ );
or   ( new_n44227_, new_n44226_, new_n43983_ );
and  ( new_n44228_, new_n44191_, new_n43879_ );
or   ( new_n44229_, new_n43977_, new_n43915_ );
or   ( new_n44230_, new_n44229_, new_n44228_ );
and  ( new_n44231_, new_n44230_, new_n44227_ );
or   ( new_n44232_, new_n44231_, new_n44225_ );
and  ( new_n44233_, new_n44232_, new_n44224_ );
nor  ( new_n44234_, new_n44233_, new_n44216_ );
xor  ( new_n44235_, new_n43898_, new_n400_ );
or   ( new_n44236_, new_n44235_, new_n524_ );
or   ( new_n44237_, new_n44145_, new_n526_ );
and  ( new_n44238_, new_n44237_, new_n44236_ );
or   ( new_n44239_, new_n44171_, new_n411_ );
xor  ( new_n44240_, new_n43799_, new_n325_ );
or   ( new_n44241_, new_n44240_, new_n409_ );
and  ( new_n44242_, new_n44241_, new_n44239_ );
nor  ( new_n44243_, new_n44242_, new_n44238_ );
xor  ( new_n44244_, new_n43937_, RIbb2f340_7 );
and  ( new_n44245_, new_n44244_, new_n316_ );
and  ( new_n44246_, new_n44185_, new_n314_ );
or   ( new_n44247_, new_n44246_, new_n44245_ );
xor  ( new_n44248_, new_n44242_, new_n44238_ );
and  ( new_n44249_, new_n44248_, new_n44247_ );
nor  ( new_n44250_, new_n44249_, new_n44243_ );
not  ( new_n44251_, new_n44250_ );
xor  ( new_n44252_, new_n44233_, new_n44216_ );
and  ( new_n44253_, new_n44252_, new_n44251_ );
or   ( new_n44254_, new_n44253_, new_n44234_ );
xor  ( new_n44255_, new_n44209_, new_n44208_ );
and  ( new_n44256_, new_n44255_, new_n44254_ );
or   ( new_n44257_, new_n44256_, new_n44210_ );
xor  ( new_n44258_, new_n44206_, new_n44204_ );
and  ( new_n44259_, new_n44258_, new_n44257_ );
nor  ( new_n44260_, new_n44259_, new_n44207_ );
not  ( new_n44261_, new_n44260_ );
xor  ( new_n44262_, new_n44165_, new_n44134_ );
nand ( new_n44263_, new_n44262_, new_n44261_ );
and  ( new_n44264_, new_n44263_, new_n44166_ );
xnor ( new_n44265_, new_n44075_, new_n44061_ );
or   ( new_n44266_, new_n44265_, new_n44264_ );
and  ( new_n44267_, new_n44265_, new_n44264_ );
xor  ( new_n44268_, new_n44258_, new_n44257_ );
xor  ( new_n44269_, new_n44160_, new_n44159_ );
xor  ( new_n44270_, new_n44269_, new_n44163_ );
and  ( new_n44271_, new_n44270_, new_n44268_ );
not  ( new_n44272_, new_n44216_ );
or   ( new_n44273_, new_n44136_, new_n44007_ );
or   ( new_n44274_, new_n43986_, new_n302_ );
and  ( new_n44275_, new_n44274_, new_n44273_ );
nor  ( new_n44276_, new_n44275_, new_n44272_ );
xor  ( new_n44277_, new_n43952_, new_n275_ );
nor  ( new_n44278_, new_n44277_, new_n283_ );
nor  ( new_n44279_, new_n44168_, new_n286_ );
or   ( new_n44280_, new_n44279_, new_n44278_ );
xor  ( new_n44281_, new_n44275_, new_n44272_ );
and  ( new_n44282_, new_n44281_, new_n44280_ );
or   ( new_n44283_, new_n44282_, new_n44276_ );
xor  ( new_n44284_, new_n44154_, new_n44153_ );
and  ( new_n44285_, new_n44284_, new_n44283_ );
xor  ( new_n44286_, new_n44179_, new_n44178_ );
xor  ( new_n44287_, new_n44284_, new_n44283_ );
and  ( new_n44288_, new_n44287_, new_n44286_ );
nor  ( new_n44289_, new_n44288_, new_n44285_ );
not  ( new_n44290_, new_n44289_ );
xor  ( new_n44291_, new_n44202_, new_n44201_ );
and  ( new_n44292_, new_n44291_, new_n44290_ );
xor  ( new_n44293_, new_n44291_, new_n44290_ );
xor  ( new_n44294_, new_n44255_, new_n44254_ );
and  ( new_n44295_, new_n44294_, new_n44293_ );
or   ( new_n44296_, new_n44295_, new_n44292_ );
xor  ( new_n44297_, new_n44270_, new_n44268_ );
and  ( new_n44298_, new_n44297_, new_n44296_ );
nor  ( new_n44299_, new_n44298_, new_n44271_ );
not  ( new_n44300_, new_n44299_ );
xor  ( new_n44301_, new_n44262_, new_n44261_ );
and  ( new_n44302_, new_n44301_, new_n44300_ );
nor  ( new_n44303_, new_n44301_, new_n44300_ );
xnor ( new_n44304_, new_n44294_, new_n44293_ );
xor  ( new_n44305_, new_n43787_, RIbb2ef80_15 );
nand ( new_n44306_, new_n44305_, new_n662_ );
nand ( new_n44307_, new_n44214_, new_n660_ );
and  ( new_n44308_, new_n44307_, new_n44306_ );
or   ( new_n44309_, new_n44308_, new_n747_ );
xor  ( new_n44310_, new_n43803_, RIbb2f160_11 );
and  ( new_n44311_, new_n44310_, new_n373_ );
nor  ( new_n44312_, new_n44240_, new_n411_ );
nor  ( new_n44313_, new_n44312_, new_n44311_ );
not  ( new_n44314_, new_n44313_ );
xor  ( new_n44315_, new_n44308_, new_n747_ );
nand ( new_n44316_, new_n44315_, new_n44314_ );
and  ( new_n44317_, new_n44316_, new_n44309_ );
xor  ( new_n44318_, RIbb31cf8_144, RIbb2d108_80 );
xnor ( new_n44319_, new_n44318_, new_n43754_ );
and  ( new_n44320_, new_n44319_, new_n43880_ );
not  ( new_n44321_, new_n44320_ );
xor  ( new_n44322_, new_n43894_, new_n400_ );
or   ( new_n44323_, new_n44322_, new_n524_ );
or   ( new_n44324_, new_n44235_, new_n526_ );
and  ( new_n44325_, new_n44324_, new_n44323_ );
or   ( new_n44326_, new_n44325_, new_n44321_ );
xor  ( new_n44327_, new_n43956_, new_n309_ );
nor  ( new_n44328_, new_n44327_, new_n317_ );
and  ( new_n44329_, new_n44244_, new_n314_ );
or   ( new_n44330_, new_n44329_, new_n44328_ );
xor  ( new_n44331_, new_n44325_, new_n44321_ );
nand ( new_n44332_, new_n44331_, new_n44330_ );
and  ( new_n44333_, new_n44332_, new_n44326_ );
nor  ( new_n44334_, new_n44333_, new_n44317_ );
or   ( new_n44335_, new_n44220_, new_n340_ );
xor  ( new_n44336_, new_n43888_, new_n329_ );
or   ( new_n44337_, new_n44336_, new_n337_ );
and  ( new_n44338_, new_n44337_, new_n44335_ );
xor  ( new_n44339_, new_n44218_, new_n43950_ );
or   ( new_n44340_, new_n44339_, new_n43983_ );
nor  ( new_n44341_, new_n44183_, new_n43880_ );
or   ( new_n44342_, new_n44184_, new_n43977_ );
or   ( new_n44343_, new_n44342_, new_n44341_ );
and  ( new_n44344_, new_n44343_, new_n44340_ );
nor  ( new_n44345_, new_n44344_, new_n44338_ );
and  ( new_n44346_, new_n44137_, new_n295_ );
and  ( new_n44347_, new_n44192_, new_n43949_ );
or   ( new_n44348_, new_n44347_, new_n44346_ );
xor  ( new_n44349_, new_n44344_, new_n44338_ );
and  ( new_n44350_, new_n44349_, new_n44348_ );
or   ( new_n44351_, new_n44350_, new_n44345_ );
xor  ( new_n44352_, new_n44333_, new_n44317_ );
and  ( new_n44353_, new_n44352_, new_n44351_ );
or   ( new_n44354_, new_n44353_, new_n44334_ );
xor  ( new_n44355_, new_n44197_, new_n44190_ );
nand ( new_n44356_, new_n44355_, new_n44354_ );
or   ( new_n44357_, new_n44355_, new_n44354_ );
xor  ( new_n44358_, new_n44252_, new_n44251_ );
nand ( new_n44359_, new_n44358_, new_n44357_ );
and  ( new_n44360_, new_n44359_, new_n44356_ );
nor  ( new_n44361_, new_n44360_, new_n44304_ );
xor  ( new_n44362_, new_n44248_, new_n44247_ );
xor  ( new_n44363_, new_n44281_, new_n44280_ );
and  ( new_n44364_, new_n44363_, new_n44362_ );
xor  ( new_n44365_, new_n44363_, new_n44362_ );
xor  ( new_n44366_, new_n44231_, new_n44225_ );
and  ( new_n44367_, new_n44366_, new_n44365_ );
or   ( new_n44368_, new_n44367_, new_n44364_ );
xor  ( new_n44369_, new_n44287_, new_n44286_ );
and  ( new_n44370_, new_n44369_, new_n44368_ );
or   ( new_n44371_, new_n44277_, new_n286_ );
xor  ( new_n44372_, new_n43985_, new_n275_ );
or   ( new_n44373_, new_n44372_, new_n283_ );
and  ( new_n44374_, new_n44373_, new_n44371_ );
nor  ( new_n44375_, RIbb2eda0_19, RIbb2ee18_18 );
not  ( new_n44376_, new_n44375_ );
and  ( new_n44377_, new_n44376_, new_n747_ );
xor  ( new_n44378_, new_n43793_, new_n745_ );
and  ( new_n44379_, new_n44378_, new_n822_ );
nor  ( new_n44380_, new_n44379_, new_n44377_ );
or   ( new_n44381_, new_n44380_, new_n44374_ );
xor  ( new_n44382_, new_n43884_, new_n325_ );
or   ( new_n44383_, new_n44382_, new_n409_ );
nand ( new_n44384_, new_n44310_, new_n371_ );
and  ( new_n44385_, new_n44384_, new_n44383_ );
xor  ( new_n44386_, new_n44319_, new_n43950_ );
or   ( new_n44387_, new_n44386_, new_n43983_ );
nor  ( new_n44388_, new_n44218_, new_n43880_ );
or   ( new_n44389_, new_n44219_, new_n43977_ );
or   ( new_n44390_, new_n44389_, new_n44388_ );
and  ( new_n44391_, new_n44390_, new_n44387_ );
nor  ( new_n44392_, new_n44391_, new_n44385_ );
and  ( new_n44393_, new_n44226_, new_n43949_ );
and  ( new_n44394_, new_n44192_, new_n295_ );
or   ( new_n44395_, new_n44394_, new_n44393_ );
xor  ( new_n44396_, new_n44391_, new_n44385_ );
and  ( new_n44397_, new_n44396_, new_n44395_ );
or   ( new_n44398_, new_n44397_, new_n44392_ );
xor  ( new_n44399_, new_n44380_, new_n44374_ );
nand ( new_n44400_, new_n44399_, new_n44398_ );
and  ( new_n44401_, new_n44400_, new_n44381_ );
xor  ( new_n44402_, RIbb31d70_145, RIbb2d090_81 );
nor  ( new_n44403_, new_n43740_, new_n43727_ );
not  ( new_n44404_, new_n44403_ );
nand ( new_n44405_, new_n44404_, new_n43483_ );
and  ( new_n44406_, new_n44405_, new_n43750_ );
xnor ( new_n44407_, new_n44406_, new_n44402_ );
and  ( new_n44408_, new_n44407_, new_n43880_ );
not  ( new_n44409_, new_n44408_ );
xor  ( new_n44410_, new_n43937_, new_n329_ );
or   ( new_n44411_, new_n44410_, new_n337_ );
or   ( new_n44412_, new_n44336_, new_n340_ );
and  ( new_n44413_, new_n44412_, new_n44411_ );
or   ( new_n44414_, new_n44413_, new_n44409_ );
xor  ( new_n44415_, new_n43898_, new_n520_ );
nor  ( new_n44416_, new_n44415_, new_n755_ );
and  ( new_n44417_, new_n44305_, new_n660_ );
or   ( new_n44418_, new_n44417_, new_n44416_ );
xor  ( new_n44419_, new_n44413_, new_n44409_ );
nand ( new_n44420_, new_n44419_, new_n44418_ );
and  ( new_n44421_, new_n44420_, new_n44414_ );
xor  ( new_n44422_, new_n43812_, new_n275_ );
or   ( new_n44423_, new_n44422_, new_n283_ );
or   ( new_n44424_, new_n44372_, new_n286_ );
and  ( new_n44425_, new_n44424_, new_n44423_ );
xor  ( new_n44426_, new_n43799_, new_n400_ );
or   ( new_n44427_, new_n44426_, new_n524_ );
or   ( new_n44428_, new_n44322_, new_n526_ );
and  ( new_n44429_, new_n44428_, new_n44427_ );
or   ( new_n44430_, new_n44429_, new_n44425_ );
xor  ( new_n44431_, new_n43952_, new_n309_ );
nor  ( new_n44432_, new_n44431_, new_n317_ );
nor  ( new_n44433_, new_n44327_, new_n320_ );
or   ( new_n44434_, new_n44433_, new_n44432_ );
xor  ( new_n44435_, new_n44429_, new_n44425_ );
nand ( new_n44436_, new_n44435_, new_n44434_ );
and  ( new_n44437_, new_n44436_, new_n44430_ );
or   ( new_n44438_, new_n44437_, new_n44421_ );
xor  ( new_n44439_, new_n44437_, new_n44421_ );
xor  ( new_n44440_, new_n44331_, new_n44330_ );
nand ( new_n44441_, new_n44440_, new_n44439_ );
and  ( new_n44442_, new_n44441_, new_n44438_ );
nor  ( new_n44443_, new_n44442_, new_n44401_ );
xor  ( new_n44444_, new_n44352_, new_n44351_ );
xor  ( new_n44445_, new_n44442_, new_n44401_ );
and  ( new_n44446_, new_n44445_, new_n44444_ );
or   ( new_n44447_, new_n44446_, new_n44443_ );
xor  ( new_n44448_, new_n44369_, new_n44368_ );
and  ( new_n44449_, new_n44448_, new_n44447_ );
nor  ( new_n44450_, new_n44449_, new_n44370_ );
not  ( new_n44451_, new_n44450_ );
xor  ( new_n44452_, new_n44360_, new_n44304_ );
and  ( new_n44453_, new_n44452_, new_n44451_ );
or   ( new_n44454_, new_n44453_, new_n44361_ );
xor  ( new_n44455_, new_n44297_, new_n44296_ );
nor  ( new_n44456_, new_n44455_, new_n44454_ );
xor  ( new_n44457_, new_n44355_, new_n44354_ );
xor  ( new_n44458_, new_n44457_, new_n44358_ );
not  ( new_n44459_, new_n44458_ );
xor  ( new_n44460_, new_n44315_, new_n44314_ );
xor  ( new_n44461_, new_n44349_, new_n44348_ );
and  ( new_n44462_, new_n44461_, new_n44460_ );
xor  ( new_n44463_, new_n44461_, new_n44460_ );
xor  ( new_n44464_, new_n44399_, new_n44398_ );
and  ( new_n44465_, new_n44464_, new_n44463_ );
or   ( new_n44466_, new_n44465_, new_n44462_ );
xor  ( new_n44467_, new_n44366_, new_n44365_ );
nand ( new_n44468_, new_n44467_, new_n44466_ );
nor  ( new_n44469_, new_n44467_, new_n44466_ );
xor  ( new_n44470_, new_n43787_, RIbb2ee90_17 );
nand ( new_n44471_, new_n44470_, new_n822_ );
nand ( new_n44472_, new_n44378_, new_n820_ );
and  ( new_n44473_, new_n44472_, new_n44471_ );
or   ( new_n44474_, new_n44473_, new_n895_ );
xor  ( new_n44475_, new_n43803_, RIbb2f070_13 );
and  ( new_n44476_, new_n44475_, new_n456_ );
nor  ( new_n44477_, new_n44426_, new_n526_ );
or   ( new_n44478_, new_n44477_, new_n44476_ );
xor  ( new_n44479_, new_n44473_, new_n895_ );
nand ( new_n44480_, new_n44479_, new_n44478_ );
nand ( new_n44481_, new_n44480_, new_n44474_ );
nand ( new_n44482_, new_n44481_, new_n44380_ );
xor  ( new_n44483_, new_n43888_, new_n325_ );
or   ( new_n44484_, new_n44483_, new_n409_ );
or   ( new_n44485_, new_n44382_, new_n411_ );
and  ( new_n44486_, new_n44485_, new_n44484_ );
xor  ( new_n44487_, new_n43914_, new_n275_ );
or   ( new_n44488_, new_n44487_, new_n283_ );
or   ( new_n44489_, new_n44422_, new_n286_ );
and  ( new_n44490_, new_n44489_, new_n44488_ );
nor  ( new_n44491_, new_n44490_, new_n44486_ );
and  ( new_n44492_, new_n44339_, new_n43949_ );
and  ( new_n44493_, new_n44226_, new_n295_ );
or   ( new_n44494_, new_n44493_, new_n44492_ );
xor  ( new_n44495_, new_n44490_, new_n44486_ );
and  ( new_n44496_, new_n44495_, new_n44494_ );
or   ( new_n44497_, new_n44496_, new_n44491_ );
xor  ( new_n44498_, new_n44481_, new_n44380_ );
nand ( new_n44499_, new_n44498_, new_n44497_ );
and  ( new_n44500_, new_n44499_, new_n44482_ );
xor  ( new_n44501_, RIbb31de8_146, RIbb2d018_82 );
and  ( new_n44502_, new_n44404_, new_n43479_ );
nor  ( new_n44503_, new_n44502_, new_n43746_ );
nor  ( new_n44504_, new_n44503_, new_n43481_ );
nor  ( new_n44505_, new_n44504_, new_n43745_ );
xnor ( new_n44506_, new_n44505_, new_n44501_ );
and  ( new_n44507_, new_n44506_, new_n43880_ );
not  ( new_n44508_, new_n44507_ );
xor  ( new_n44509_, new_n44407_, new_n43950_ );
or   ( new_n44510_, new_n44509_, new_n43983_ );
nor  ( new_n44511_, new_n44319_, new_n43880_ );
or   ( new_n44512_, new_n44320_, new_n43977_ );
or   ( new_n44513_, new_n44512_, new_n44511_ );
and  ( new_n44514_, new_n44513_, new_n44510_ );
nor  ( new_n44515_, new_n44514_, new_n44508_ );
xor  ( new_n44516_, new_n43894_, RIbb2ef80_15 );
and  ( new_n44517_, new_n44516_, new_n662_ );
nor  ( new_n44518_, new_n44415_, new_n757_ );
or   ( new_n44519_, new_n44518_, new_n44517_ );
xor  ( new_n44520_, new_n44514_, new_n44508_ );
and  ( new_n44521_, new_n44520_, new_n44519_ );
or   ( new_n44522_, new_n44521_, new_n44515_ );
xor  ( new_n44523_, new_n44419_, new_n44418_ );
nand ( new_n44524_, new_n44523_, new_n44522_ );
xor  ( new_n44525_, new_n44523_, new_n44522_ );
xor  ( new_n44526_, new_n44396_, new_n44395_ );
nand ( new_n44527_, new_n44526_, new_n44525_ );
and  ( new_n44528_, new_n44527_, new_n44524_ );
nor  ( new_n44529_, new_n44528_, new_n44500_ );
xor  ( new_n44530_, new_n44440_, new_n44439_ );
xor  ( new_n44531_, new_n44528_, new_n44500_ );
and  ( new_n44532_, new_n44531_, new_n44530_ );
nor  ( new_n44533_, new_n44532_, new_n44529_ );
or   ( new_n44534_, new_n44533_, new_n44469_ );
and  ( new_n44535_, new_n44534_, new_n44468_ );
nor  ( new_n44536_, new_n44535_, new_n44459_ );
xor  ( new_n44537_, new_n44535_, new_n44459_ );
xor  ( new_n44538_, new_n44448_, new_n44447_ );
and  ( new_n44539_, new_n44538_, new_n44537_ );
nor  ( new_n44540_, new_n44539_, new_n44536_ );
not  ( new_n44541_, new_n44540_ );
xor  ( new_n44542_, new_n44452_, new_n44451_ );
and  ( new_n44543_, new_n44542_, new_n44541_ );
nor  ( new_n44544_, new_n44542_, new_n44541_ );
xor  ( new_n44545_, new_n44479_, new_n44478_ );
xor  ( new_n44546_, new_n44520_, new_n44519_ );
and  ( new_n44547_, new_n44546_, new_n44545_ );
xor  ( new_n44548_, new_n44495_, new_n44494_ );
xor  ( new_n44549_, new_n44546_, new_n44545_ );
and  ( new_n44550_, new_n44549_, new_n44548_ );
or   ( new_n44551_, new_n44550_, new_n44547_ );
xor  ( new_n44552_, new_n44498_, new_n44497_ );
and  ( new_n44553_, new_n44552_, new_n44551_ );
xor  ( new_n44554_, new_n44552_, new_n44551_ );
xor  ( new_n44555_, new_n44526_, new_n44525_ );
and  ( new_n44556_, new_n44555_, new_n44554_ );
or   ( new_n44557_, new_n44556_, new_n44553_ );
xnor ( new_n44558_, new_n44464_, new_n44463_ );
or   ( new_n44559_, new_n44410_, new_n340_ );
xor  ( new_n44560_, new_n43956_, new_n329_ );
or   ( new_n44561_, new_n44560_, new_n337_ );
and  ( new_n44562_, new_n44561_, new_n44559_ );
not  ( new_n44563_, RIbb2ed28_20 );
and  ( new_n44564_, new_n1126_, new_n44563_ );
not  ( new_n44565_, new_n44564_ );
and  ( new_n44566_, new_n44565_, new_n895_ );
xor  ( new_n44567_, new_n43793_, new_n893_ );
and  ( new_n44568_, new_n44567_, new_n1042_ );
nor  ( new_n44569_, new_n44568_, new_n44566_ );
nor  ( new_n44570_, new_n44569_, new_n44562_ );
xor  ( new_n44571_, new_n43985_, RIbb2f340_7 );
and  ( new_n44572_, new_n44571_, new_n316_ );
nor  ( new_n44573_, new_n44431_, new_n320_ );
or   ( new_n44574_, new_n44573_, new_n44572_ );
xor  ( new_n44575_, new_n44569_, new_n44562_ );
and  ( new_n44576_, new_n44575_, new_n44574_ );
or   ( new_n44577_, new_n44576_, new_n44570_ );
xor  ( new_n44578_, new_n44435_, new_n44434_ );
nand ( new_n44579_, new_n44578_, new_n44577_ );
nor  ( new_n44580_, new_n44578_, new_n44577_ );
or   ( new_n44581_, new_n44483_, new_n411_ );
xor  ( new_n44582_, new_n43937_, new_n325_ );
or   ( new_n44583_, new_n44582_, new_n409_ );
and  ( new_n44584_, new_n44583_, new_n44581_ );
xor  ( new_n44585_, new_n44506_, new_n43950_ );
or   ( new_n44586_, new_n44585_, new_n43983_ );
not  ( new_n44587_, new_n44407_ );
and  ( new_n44588_, new_n44587_, new_n43879_ );
or   ( new_n44589_, new_n44408_, new_n43977_ );
or   ( new_n44590_, new_n44589_, new_n44588_ );
and  ( new_n44591_, new_n44590_, new_n44586_ );
or   ( new_n44592_, new_n44591_, new_n44584_ );
and  ( new_n44593_, new_n44386_, new_n43949_ );
and  ( new_n44594_, new_n44339_, new_n295_ );
or   ( new_n44595_, new_n44594_, new_n44593_ );
xor  ( new_n44596_, new_n44591_, new_n44584_ );
nand ( new_n44597_, new_n44596_, new_n44595_ );
and  ( new_n44598_, new_n44597_, new_n44592_ );
xor  ( new_n44599_, RIbb31e60_147, RIbb2cfa0_83 );
xnor ( new_n44600_, new_n44599_, new_n44503_ );
and  ( new_n44601_, new_n44600_, new_n43880_ );
not  ( new_n44602_, new_n44601_ );
or   ( new_n44603_, new_n44560_, new_n340_ );
xor  ( new_n44604_, new_n43952_, new_n329_ );
or   ( new_n44605_, new_n44604_, new_n337_ );
and  ( new_n44606_, new_n44605_, new_n44603_ );
or   ( new_n44607_, new_n44606_, new_n44602_ );
and  ( new_n44608_, new_n44516_, new_n660_ );
xor  ( new_n44609_, new_n43799_, new_n520_ );
nor  ( new_n44610_, new_n44609_, new_n755_ );
or   ( new_n44611_, new_n44610_, new_n44608_ );
xor  ( new_n44612_, new_n44606_, new_n44602_ );
nand ( new_n44613_, new_n44612_, new_n44611_ );
and  ( new_n44614_, new_n44613_, new_n44607_ );
nor  ( new_n44615_, new_n44614_, new_n44598_ );
nand ( new_n44616_, new_n44475_, new_n454_ );
xor  ( new_n44617_, new_n43884_, new_n400_ );
or   ( new_n44618_, new_n44617_, new_n524_ );
and  ( new_n44619_, new_n44618_, new_n44616_ );
or   ( new_n44620_, new_n44487_, new_n286_ );
xor  ( new_n44621_, new_n44183_, RIbb2f430_5 );
nand ( new_n44622_, new_n44621_, new_n282_ );
and  ( new_n44623_, new_n44622_, new_n44620_ );
nor  ( new_n44624_, new_n44623_, new_n44619_ );
and  ( new_n44625_, new_n44470_, new_n820_ );
xor  ( new_n44626_, new_n43898_, new_n745_ );
nor  ( new_n44627_, new_n44626_, new_n897_ );
or   ( new_n44628_, new_n44627_, new_n44625_ );
xor  ( new_n44629_, new_n44623_, new_n44619_ );
and  ( new_n44630_, new_n44629_, new_n44628_ );
or   ( new_n44631_, new_n44630_, new_n44624_ );
xor  ( new_n44632_, new_n44614_, new_n44598_ );
and  ( new_n44633_, new_n44632_, new_n44631_ );
nor  ( new_n44634_, new_n44633_, new_n44615_ );
or   ( new_n44635_, new_n44634_, new_n44580_ );
and  ( new_n44636_, new_n44635_, new_n44579_ );
xor  ( new_n44637_, new_n44636_, new_n44558_ );
xor  ( new_n44638_, new_n44637_, new_n44557_ );
xor  ( new_n44639_, new_n44531_, new_n44530_ );
and  ( new_n44640_, new_n44639_, new_n44638_ );
nand ( new_n44641_, new_n44571_, new_n314_ );
xor  ( new_n44642_, new_n43812_, new_n309_ );
or   ( new_n44643_, new_n44642_, new_n317_ );
nand ( new_n44644_, new_n44643_, new_n44641_ );
and  ( new_n44645_, new_n44644_, new_n44569_ );
xor  ( new_n44646_, new_n43894_, RIbb2ee90_17 );
nand ( new_n44647_, new_n44646_, new_n822_ );
or   ( new_n44648_, new_n44626_, new_n899_ );
and  ( new_n44649_, new_n44648_, new_n44647_ );
xor  ( new_n44650_, new_n44600_, new_n43950_ );
or   ( new_n44651_, new_n44650_, new_n43983_ );
nor  ( new_n44652_, new_n44506_, new_n43880_ );
or   ( new_n44653_, new_n44507_, new_n43977_ );
or   ( new_n44654_, new_n44653_, new_n44652_ );
and  ( new_n44655_, new_n44654_, new_n44651_ );
nor  ( new_n44656_, new_n44655_, new_n44649_ );
and  ( new_n44657_, new_n44386_, new_n295_ );
and  ( new_n44658_, new_n44509_, new_n43949_ );
or   ( new_n44659_, new_n44658_, new_n44657_ );
xor  ( new_n44660_, new_n44655_, new_n44649_ );
and  ( new_n44661_, new_n44660_, new_n44659_ );
or   ( new_n44662_, new_n44661_, new_n44656_ );
xor  ( new_n44663_, new_n44644_, new_n44569_ );
and  ( new_n44664_, new_n44663_, new_n44662_ );
or   ( new_n44665_, new_n44664_, new_n44645_ );
xor  ( new_n44666_, new_n44575_, new_n44574_ );
and  ( new_n44667_, new_n44666_, new_n44665_ );
xor  ( new_n44668_, new_n43787_, new_n893_ );
or   ( new_n44669_, new_n44668_, new_n1135_ );
nand ( new_n44670_, new_n44567_, new_n1040_ );
and  ( new_n44671_, new_n44670_, new_n44669_ );
or   ( new_n44672_, new_n44671_, new_n1128_ );
xor  ( new_n44673_, new_n43803_, RIbb2ef80_15 );
and  ( new_n44674_, new_n44673_, new_n662_ );
nor  ( new_n44675_, new_n44609_, new_n757_ );
or   ( new_n44676_, new_n44675_, new_n44674_ );
xor  ( new_n44677_, new_n44671_, new_n1128_ );
nand ( new_n44678_, new_n44677_, new_n44676_ );
and  ( new_n44679_, new_n44678_, new_n44672_ );
xor  ( new_n44680_, RIbb31ed8_148, RIbb2cf28_84 );
xor  ( new_n44681_, new_n44680_, new_n44404_ );
and  ( new_n44682_, new_n44681_, new_n43880_ );
not  ( new_n44683_, new_n44682_ );
xor  ( new_n44684_, new_n43956_, new_n325_ );
or   ( new_n44685_, new_n44684_, new_n409_ );
or   ( new_n44686_, new_n44582_, new_n411_ );
and  ( new_n44687_, new_n44686_, new_n44685_ );
or   ( new_n44688_, new_n44687_, new_n44683_ );
xor  ( new_n44689_, new_n43985_, RIbb2f250_9 );
and  ( new_n44690_, new_n44689_, new_n336_ );
nor  ( new_n44691_, new_n44604_, new_n340_ );
or   ( new_n44692_, new_n44691_, new_n44690_ );
xor  ( new_n44693_, new_n44687_, new_n44683_ );
nand ( new_n44694_, new_n44693_, new_n44692_ );
and  ( new_n44695_, new_n44694_, new_n44688_ );
nor  ( new_n44696_, new_n44695_, new_n44679_ );
xor  ( new_n44697_, new_n43914_, RIbb2f340_7 );
nand ( new_n44698_, new_n44697_, new_n316_ );
or   ( new_n44699_, new_n44642_, new_n320_ );
and  ( new_n44700_, new_n44699_, new_n44698_ );
xor  ( new_n44701_, new_n43888_, new_n400_ );
or   ( new_n44702_, new_n44701_, new_n524_ );
or   ( new_n44703_, new_n44617_, new_n526_ );
and  ( new_n44704_, new_n44703_, new_n44702_ );
nor  ( new_n44705_, new_n44704_, new_n44700_ );
xor  ( new_n44706_, new_n44218_, RIbb2f430_5 );
and  ( new_n44707_, new_n44706_, new_n282_ );
and  ( new_n44708_, new_n44621_, new_n280_ );
or   ( new_n44709_, new_n44708_, new_n44707_ );
xor  ( new_n44710_, new_n44704_, new_n44700_ );
and  ( new_n44711_, new_n44710_, new_n44709_ );
or   ( new_n44712_, new_n44711_, new_n44705_ );
xor  ( new_n44713_, new_n44695_, new_n44679_ );
and  ( new_n44714_, new_n44713_, new_n44712_ );
or   ( new_n44715_, new_n44714_, new_n44696_ );
xor  ( new_n44716_, new_n44666_, new_n44665_ );
and  ( new_n44717_, new_n44716_, new_n44715_ );
or   ( new_n44718_, new_n44717_, new_n44667_ );
xnor ( new_n44719_, new_n44578_, new_n44577_ );
xor  ( new_n44720_, new_n44719_, new_n44634_ );
and  ( new_n44721_, new_n44720_, new_n44718_ );
xor  ( new_n44722_, new_n44596_, new_n44595_ );
xor  ( new_n44723_, new_n44612_, new_n44611_ );
and  ( new_n44724_, new_n44723_, new_n44722_ );
xor  ( new_n44725_, new_n44629_, new_n44628_ );
xor  ( new_n44726_, new_n44723_, new_n44722_ );
and  ( new_n44727_, new_n44726_, new_n44725_ );
or   ( new_n44728_, new_n44727_, new_n44724_ );
xor  ( new_n44729_, new_n44632_, new_n44631_ );
and  ( new_n44730_, new_n44729_, new_n44728_ );
xor  ( new_n44731_, new_n44729_, new_n44728_ );
xor  ( new_n44732_, new_n44549_, new_n44548_ );
and  ( new_n44733_, new_n44732_, new_n44731_ );
or   ( new_n44734_, new_n44733_, new_n44730_ );
xor  ( new_n44735_, new_n44720_, new_n44718_ );
and  ( new_n44736_, new_n44735_, new_n44734_ );
nor  ( new_n44737_, new_n44736_, new_n44721_ );
not  ( new_n44738_, new_n44737_ );
xor  ( new_n44739_, new_n44639_, new_n44638_ );
and  ( new_n44740_, new_n44739_, new_n44738_ );
or   ( new_n44741_, new_n44740_, new_n44640_ );
nor  ( new_n44742_, new_n44636_, new_n44558_ );
and  ( new_n44743_, new_n44637_, new_n44557_ );
or   ( new_n44744_, new_n44743_, new_n44742_ );
xor  ( new_n44745_, new_n44445_, new_n44444_ );
xor  ( new_n44746_, new_n44745_, new_n44744_ );
xnor ( new_n44747_, new_n44467_, new_n44466_ );
xor  ( new_n44748_, new_n44747_, new_n44533_ );
xor  ( new_n44749_, new_n44748_, new_n44746_ );
nor  ( new_n44750_, new_n44749_, new_n44741_ );
and  ( new_n44751_, new_n44745_, new_n44744_ );
and  ( new_n44752_, new_n44748_, new_n44746_ );
nor  ( new_n44753_, new_n44752_, new_n44751_ );
xor  ( new_n44754_, new_n44538_, new_n44537_ );
not  ( new_n44755_, new_n44754_ );
and  ( new_n44756_, new_n44755_, new_n44753_ );
nor  ( new_n44757_, new_n44756_, new_n44750_ );
xor  ( new_n44758_, new_n43812_, RIbb2f250_9 );
nand ( new_n44759_, new_n44758_, new_n334_ );
xor  ( new_n44760_, new_n43914_, new_n329_ );
or   ( new_n44761_, new_n44760_, new_n337_ );
and  ( new_n44762_, new_n44761_, new_n44759_ );
xor  ( new_n44763_, new_n43888_, RIbb2ef80_15 );
nand ( new_n44764_, new_n44763_, new_n662_ );
xor  ( new_n44765_, new_n43884_, new_n520_ );
or   ( new_n44766_, new_n44765_, new_n757_ );
and  ( new_n44767_, new_n44766_, new_n44764_ );
nor  ( new_n44768_, new_n44767_, new_n44762_ );
xor  ( new_n44769_, new_n44183_, RIbb2f340_7 );
and  ( new_n44770_, new_n44769_, new_n314_ );
xor  ( new_n44771_, new_n44218_, RIbb2f340_7 );
and  ( new_n44772_, new_n44771_, new_n316_ );
or   ( new_n44773_, new_n44772_, new_n44770_ );
xor  ( new_n44774_, new_n44767_, new_n44762_ );
and  ( new_n44775_, new_n44774_, new_n44773_ );
or   ( new_n44776_, new_n44775_, new_n44768_ );
and  ( new_n44777_, new_n44646_, new_n820_ );
xor  ( new_n44778_, new_n43799_, new_n745_ );
nor  ( new_n44779_, new_n44778_, new_n897_ );
or   ( new_n44780_, new_n44779_, new_n44777_ );
xor  ( new_n44781_, RIbb31f50_149, RIbb2ceb0_85 );
nor  ( new_n44782_, new_n43735_, new_n43723_ );
nor  ( new_n44783_, new_n44782_, new_n43724_ );
nor  ( new_n44784_, new_n44783_, new_n43731_ );
xnor ( new_n44785_, new_n44784_, new_n44781_ );
and  ( new_n44786_, new_n44785_, new_n43880_ );
not  ( new_n44787_, new_n44786_ );
xor  ( new_n44788_, new_n44681_, new_n43945_ );
not  ( new_n44789_, new_n44788_ );
or   ( new_n44790_, new_n44789_, new_n43983_ );
nor  ( new_n44791_, new_n44600_, new_n43880_ );
or   ( new_n44792_, new_n44601_, new_n43977_ );
or   ( new_n44793_, new_n44792_, new_n44791_ );
and  ( new_n44794_, new_n44793_, new_n44790_ );
xor  ( new_n44795_, new_n44794_, new_n44787_ );
xor  ( new_n44796_, new_n44795_, new_n44780_ );
xor  ( new_n44797_, new_n44796_, new_n44776_ );
and  ( new_n44798_, new_n44758_, new_n336_ );
and  ( new_n44799_, new_n44689_, new_n334_ );
or   ( new_n44800_, new_n44799_, new_n44798_ );
nor  ( new_n44801_, RIbb2ebc0_23, RIbb2ec38_22 );
not  ( new_n44802_, new_n44801_ );
and  ( new_n44803_, new_n44802_, new_n1128_ );
xor  ( new_n44804_, new_n43793_, new_n1126_ );
and  ( new_n44805_, new_n44804_, new_n1253_ );
nor  ( new_n44806_, new_n44805_, new_n44803_ );
not  ( new_n44807_, new_n44806_ );
xor  ( new_n44808_, new_n43952_, new_n325_ );
or   ( new_n44809_, new_n44808_, new_n409_ );
or   ( new_n44810_, new_n44684_, new_n411_ );
and  ( new_n44811_, new_n44810_, new_n44809_ );
xor  ( new_n44812_, new_n44811_, new_n44807_ );
xor  ( new_n44813_, new_n44812_, new_n44800_ );
xor  ( new_n44814_, new_n44813_, new_n44797_ );
and  ( new_n44815_, new_n44769_, new_n316_ );
and  ( new_n44816_, new_n44697_, new_n314_ );
or   ( new_n44817_, new_n44816_, new_n44815_ );
or   ( new_n44818_, new_n44765_, new_n755_ );
nand ( new_n44819_, new_n44673_, new_n660_ );
and  ( new_n44820_, new_n44819_, new_n44818_ );
xor  ( new_n44821_, new_n43898_, new_n893_ );
or   ( new_n44822_, new_n44821_, new_n1135_ );
or   ( new_n44823_, new_n44668_, new_n1137_ );
and  ( new_n44824_, new_n44823_, new_n44822_ );
xor  ( new_n44825_, new_n44824_, new_n44820_ );
xor  ( new_n44826_, new_n44825_, new_n44817_ );
xor  ( new_n44827_, new_n43985_, new_n325_ );
or   ( new_n44828_, new_n44827_, new_n409_ );
or   ( new_n44829_, new_n44808_, new_n411_ );
and  ( new_n44830_, new_n44829_, new_n44828_ );
not  ( new_n44831_, RIbb2eb48_24 );
and  ( new_n44832_, new_n1583_, new_n44831_ );
not  ( new_n44833_, new_n44832_ );
and  ( new_n44834_, new_n44833_, new_n1357_ );
xor  ( new_n44835_, new_n43793_, RIbb2ebc0_23 );
nor  ( new_n44836_, new_n44835_, new_n1593_ );
nor  ( new_n44837_, new_n44836_, new_n44834_ );
nor  ( new_n44838_, new_n44837_, new_n44830_ );
xor  ( new_n44839_, new_n44506_, new_n275_ );
or   ( new_n44840_, new_n44839_, new_n283_ );
xor  ( new_n44841_, new_n44407_, new_n275_ );
or   ( new_n44842_, new_n44841_, new_n286_ );
and  ( new_n44843_, new_n44842_, new_n44840_ );
xor  ( new_n44844_, new_n44319_, new_n309_ );
or   ( new_n44845_, new_n44844_, new_n317_ );
nand ( new_n44846_, new_n44771_, new_n314_ );
and  ( new_n44847_, new_n44846_, new_n44845_ );
nor  ( new_n44848_, new_n44847_, new_n44843_ );
xor  ( new_n44849_, new_n43937_, RIbb2ef80_15 );
and  ( new_n44850_, new_n44849_, new_n662_ );
and  ( new_n44851_, new_n44763_, new_n660_ );
or   ( new_n44852_, new_n44851_, new_n44850_ );
xor  ( new_n44853_, new_n44847_, new_n44843_ );
and  ( new_n44854_, new_n44853_, new_n44852_ );
or   ( new_n44855_, new_n44854_, new_n44848_ );
xor  ( new_n44856_, new_n44837_, new_n44830_ );
and  ( new_n44857_, new_n44856_, new_n44855_ );
or   ( new_n44858_, new_n44857_, new_n44838_ );
and  ( new_n44859_, new_n44585_, new_n43949_ );
and  ( new_n44860_, new_n44509_, new_n295_ );
or   ( new_n44861_, new_n44860_, new_n44859_ );
xor  ( new_n44862_, new_n43937_, new_n400_ );
or   ( new_n44863_, new_n44862_, new_n524_ );
or   ( new_n44864_, new_n44701_, new_n526_ );
and  ( new_n44865_, new_n44864_, new_n44863_ );
xor  ( new_n44866_, new_n44319_, new_n275_ );
or   ( new_n44867_, new_n44866_, new_n283_ );
nand ( new_n44868_, new_n44706_, new_n280_ );
and  ( new_n44869_, new_n44868_, new_n44867_ );
xor  ( new_n44870_, new_n44869_, new_n44865_ );
xor  ( new_n44871_, new_n44870_, new_n44861_ );
xor  ( new_n44872_, new_n44871_, new_n44858_ );
xor  ( new_n44873_, new_n44872_, new_n44826_ );
and  ( new_n44874_, new_n44873_, new_n44814_ );
xor  ( new_n44875_, new_n44856_, new_n44855_ );
xor  ( new_n44876_, RIbb31fc8_150, RIbb2ce38_86 );
xnor ( new_n44877_, new_n44876_, new_n44782_ );
and  ( new_n44878_, new_n44877_, new_n43880_ );
or   ( new_n44879_, new_n44862_, new_n526_ );
xor  ( new_n44880_, new_n43956_, new_n400_ );
or   ( new_n44881_, new_n44880_, new_n524_ );
nand ( new_n44882_, new_n44881_, new_n44879_ );
xnor ( new_n44883_, new_n44882_, new_n44878_ );
xor  ( new_n44884_, new_n44785_, new_n43945_ );
nand ( new_n44885_, new_n44884_, new_n43982_ );
nor  ( new_n44886_, new_n44681_, new_n43880_ );
or   ( new_n44887_, new_n44682_, new_n43977_ );
or   ( new_n44888_, new_n44887_, new_n44886_ );
and  ( new_n44889_, new_n44888_, new_n44885_ );
xor  ( new_n44890_, new_n44889_, new_n44883_ );
and  ( new_n44891_, new_n44890_, new_n44875_ );
xor  ( new_n44892_, new_n44183_, new_n329_ );
or   ( new_n44893_, new_n44892_, new_n340_ );
xor  ( new_n44894_, new_n44218_, RIbb2f250_9 );
nand ( new_n44895_, new_n44894_, new_n336_ );
and  ( new_n44896_, new_n44895_, new_n44893_ );
xor  ( new_n44897_, new_n43884_, new_n745_ );
or   ( new_n44898_, new_n44897_, new_n899_ );
xor  ( new_n44899_, new_n43888_, new_n745_ );
or   ( new_n44900_, new_n44899_, new_n897_ );
and  ( new_n44901_, new_n44900_, new_n44898_ );
or   ( new_n44902_, new_n44901_, new_n44896_ );
xor  ( new_n44903_, new_n43914_, RIbb2f160_11 );
and  ( new_n44904_, new_n44903_, new_n373_ );
xor  ( new_n44905_, new_n43812_, RIbb2f160_11 );
and  ( new_n44906_, new_n44905_, new_n371_ );
or   ( new_n44907_, new_n44906_, new_n44904_ );
xor  ( new_n44908_, new_n44901_, new_n44896_ );
nand ( new_n44909_, new_n44908_, new_n44907_ );
nand ( new_n44910_, new_n44909_, new_n44902_ );
and  ( new_n44911_, new_n44910_, new_n44837_ );
or   ( new_n44912_, new_n44844_, new_n320_ );
xor  ( new_n44913_, new_n44407_, new_n309_ );
or   ( new_n44914_, new_n44913_, new_n317_ );
and  ( new_n44915_, new_n44914_, new_n44912_ );
or   ( new_n44916_, new_n44839_, new_n286_ );
xor  ( new_n44917_, new_n44600_, new_n275_ );
or   ( new_n44918_, new_n44917_, new_n283_ );
and  ( new_n44919_, new_n44918_, new_n44916_ );
nor  ( new_n44920_, new_n44919_, new_n44915_ );
xor  ( new_n44921_, new_n43894_, RIbb2ecb0_21 );
and  ( new_n44922_, new_n44921_, new_n1253_ );
xor  ( new_n44923_, new_n43898_, new_n1126_ );
nor  ( new_n44924_, new_n44923_, new_n1366_ );
or   ( new_n44925_, new_n44924_, new_n44922_ );
xor  ( new_n44926_, new_n44919_, new_n44915_ );
and  ( new_n44927_, new_n44926_, new_n44925_ );
or   ( new_n44928_, new_n44927_, new_n44920_ );
xor  ( new_n44929_, new_n44910_, new_n44837_ );
and  ( new_n44930_, new_n44929_, new_n44928_ );
or   ( new_n44931_, new_n44930_, new_n44911_ );
xor  ( new_n44932_, new_n44890_, new_n44875_ );
and  ( new_n44933_, new_n44932_, new_n44931_ );
or   ( new_n44934_, new_n44933_, new_n44891_ );
xor  ( new_n44935_, new_n44873_, new_n44814_ );
and  ( new_n44936_, new_n44935_, new_n44934_ );
or   ( new_n44937_, new_n44936_, new_n44874_ );
xor  ( new_n44938_, new_n43952_, new_n400_ );
or   ( new_n44939_, new_n44938_, new_n524_ );
or   ( new_n44940_, new_n44880_, new_n526_ );
and  ( new_n44941_, new_n44940_, new_n44939_ );
xor  ( new_n44942_, new_n44877_, new_n43945_ );
nand ( new_n44943_, new_n44942_, new_n43982_ );
not  ( new_n44944_, new_n44785_ );
and  ( new_n44945_, new_n44944_, new_n43879_ );
or   ( new_n44946_, new_n44786_, new_n43977_ );
or   ( new_n44947_, new_n44946_, new_n44945_ );
and  ( new_n44948_, new_n44947_, new_n44943_ );
or   ( new_n44949_, new_n44948_, new_n44941_ );
and  ( new_n44950_, new_n44789_, new_n43949_ );
and  ( new_n44951_, new_n44650_, new_n295_ );
or   ( new_n44952_, new_n44951_, new_n44950_ );
xor  ( new_n44953_, new_n44948_, new_n44941_ );
nand ( new_n44954_, new_n44953_, new_n44952_ );
and  ( new_n44955_, new_n44954_, new_n44949_ );
xor  ( new_n44956_, new_n43803_, RIbb2ee90_17 );
nand ( new_n44957_, new_n44956_, new_n820_ );
or   ( new_n44958_, new_n44897_, new_n897_ );
and  ( new_n44959_, new_n44958_, new_n44957_ );
or   ( new_n44960_, new_n44892_, new_n337_ );
or   ( new_n44961_, new_n44760_, new_n340_ );
and  ( new_n44962_, new_n44961_, new_n44960_ );
or   ( new_n44963_, new_n44962_, new_n44959_ );
nor  ( new_n44964_, new_n44923_, new_n1364_ );
xor  ( new_n44965_, new_n43787_, RIbb2ecb0_21 );
and  ( new_n44966_, new_n44965_, new_n1251_ );
or   ( new_n44967_, new_n44966_, new_n44964_ );
xor  ( new_n44968_, new_n44962_, new_n44959_ );
nand ( new_n44969_, new_n44968_, new_n44967_ );
and  ( new_n44970_, new_n44969_, new_n44963_ );
or   ( new_n44971_, new_n44970_, new_n44955_ );
xor  ( new_n44972_, RIbb32040_151, RIbb2cdc0_87 );
nor  ( new_n44973_, new_n43733_, new_n43722_ );
xnor ( new_n44974_, new_n44973_, new_n44972_ );
and  ( new_n44975_, new_n44974_, new_n43880_ );
not  ( new_n44976_, new_n44975_ );
nand ( new_n44977_, new_n44905_, new_n373_ );
or   ( new_n44978_, new_n44827_, new_n411_ );
and  ( new_n44979_, new_n44978_, new_n44977_ );
nor  ( new_n44980_, new_n44979_, new_n44976_ );
xor  ( new_n44981_, new_n43799_, new_n893_ );
nor  ( new_n44982_, new_n44981_, new_n1135_ );
xor  ( new_n44983_, new_n43894_, RIbb2eda0_19 );
and  ( new_n44984_, new_n44983_, new_n1040_ );
or   ( new_n44985_, new_n44984_, new_n44982_ );
xor  ( new_n44986_, new_n44979_, new_n44976_ );
and  ( new_n44987_, new_n44986_, new_n44985_ );
or   ( new_n44988_, new_n44987_, new_n44980_ );
xor  ( new_n44989_, new_n44970_, new_n44955_ );
nand ( new_n44990_, new_n44989_, new_n44988_ );
and  ( new_n44991_, new_n44990_, new_n44971_ );
and  ( new_n44992_, new_n44956_, new_n822_ );
nor  ( new_n44993_, new_n44778_, new_n899_ );
or   ( new_n44994_, new_n44993_, new_n44992_ );
nand ( new_n44995_, new_n44965_, new_n1253_ );
nand ( new_n44996_, new_n44804_, new_n1251_ );
and  ( new_n44997_, new_n44996_, new_n44995_ );
xor  ( new_n44998_, new_n44997_, new_n1357_ );
xor  ( new_n44999_, new_n44998_, new_n44994_ );
and  ( new_n45000_, new_n44650_, new_n43949_ );
and  ( new_n45001_, new_n44585_, new_n295_ );
or   ( new_n45002_, new_n45001_, new_n45000_ );
or   ( new_n45003_, new_n44821_, new_n1137_ );
nand ( new_n45004_, new_n44983_, new_n1042_ );
and  ( new_n45005_, new_n45004_, new_n45003_ );
or   ( new_n45006_, new_n44866_, new_n286_ );
or   ( new_n45007_, new_n44841_, new_n283_ );
and  ( new_n45008_, new_n45007_, new_n45006_ );
xor  ( new_n45009_, new_n45008_, new_n45005_ );
xor  ( new_n45010_, new_n45009_, new_n45002_ );
nand ( new_n45011_, new_n45010_, new_n44999_ );
xor  ( new_n45012_, new_n45010_, new_n44999_ );
xor  ( new_n45013_, new_n44774_, new_n44773_ );
nand ( new_n45014_, new_n45013_, new_n45012_ );
and  ( new_n45015_, new_n45014_, new_n45011_ );
nor  ( new_n45016_, new_n45015_, new_n44991_ );
nor  ( new_n45017_, new_n45008_, new_n45005_ );
and  ( new_n45018_, new_n45009_, new_n45002_ );
or   ( new_n45019_, new_n45018_, new_n45017_ );
nand ( new_n45020_, new_n44882_, new_n44878_ );
or   ( new_n45021_, new_n44889_, new_n44883_ );
and  ( new_n45022_, new_n45021_, new_n45020_ );
or   ( new_n45023_, new_n44997_, new_n1357_ );
nand ( new_n45024_, new_n44998_, new_n44994_ );
and  ( new_n45025_, new_n45024_, new_n45023_ );
xor  ( new_n45026_, new_n45025_, new_n45022_ );
xor  ( new_n45027_, new_n45026_, new_n45019_ );
xor  ( new_n45028_, new_n45015_, new_n44991_ );
and  ( new_n45029_, new_n45028_, new_n45027_ );
or   ( new_n45030_, new_n45029_, new_n45016_ );
nor  ( new_n45031_, new_n44824_, new_n44820_ );
and  ( new_n45032_, new_n44825_, new_n44817_ );
or   ( new_n45033_, new_n45032_, new_n45031_ );
or   ( new_n45034_, new_n44794_, new_n44787_ );
nand ( new_n45035_, new_n44795_, new_n44780_ );
and  ( new_n45036_, new_n45035_, new_n45034_ );
xor  ( new_n45037_, new_n45036_, new_n44806_ );
xor  ( new_n45038_, new_n45037_, new_n45033_ );
or   ( new_n45039_, new_n45025_, new_n45022_ );
nand ( new_n45040_, new_n45026_, new_n45019_ );
and  ( new_n45041_, new_n45040_, new_n45039_ );
nand ( new_n45042_, new_n44796_, new_n44776_ );
nand ( new_n45043_, new_n44813_, new_n44797_ );
and  ( new_n45044_, new_n45043_, new_n45042_ );
xor  ( new_n45045_, new_n45044_, new_n45041_ );
xor  ( new_n45046_, new_n45045_, new_n45038_ );
xor  ( new_n45047_, new_n45046_, new_n45030_ );
nor  ( new_n45048_, new_n44811_, new_n44807_ );
and  ( new_n45049_, new_n44812_, new_n44800_ );
or   ( new_n45050_, new_n45049_, new_n45048_ );
nor  ( new_n45051_, new_n44869_, new_n44865_ );
and  ( new_n45052_, new_n44870_, new_n44861_ );
or   ( new_n45053_, new_n45052_, new_n45051_ );
xor  ( new_n45054_, new_n44693_, new_n44692_ );
xor  ( new_n45055_, new_n45054_, new_n45053_ );
xor  ( new_n45056_, new_n45055_, new_n45050_ );
or   ( new_n45057_, new_n44871_, new_n44858_ );
and  ( new_n45058_, new_n44871_, new_n44858_ );
or   ( new_n45059_, new_n45058_, new_n44826_ );
and  ( new_n45060_, new_n45059_, new_n45057_ );
xor  ( new_n45061_, new_n45060_, new_n45056_ );
xor  ( new_n45062_, new_n44677_, new_n44676_ );
xor  ( new_n45063_, new_n44710_, new_n44709_ );
xor  ( new_n45064_, new_n45063_, new_n45062_ );
xor  ( new_n45065_, new_n44660_, new_n44659_ );
xor  ( new_n45066_, new_n45065_, new_n45064_ );
xor  ( new_n45067_, new_n45066_, new_n45061_ );
xor  ( new_n45068_, new_n45067_, new_n45047_ );
nand ( new_n45069_, new_n45068_, new_n44937_ );
xor  ( new_n45070_, new_n43787_, new_n1355_ );
or   ( new_n45071_, new_n45070_, new_n1593_ );
or   ( new_n45072_, new_n44835_, new_n1595_ );
and  ( new_n45073_, new_n45072_, new_n45071_ );
or   ( new_n45074_, new_n45073_, new_n1585_ );
nor  ( new_n45075_, new_n44981_, new_n1137_ );
xor  ( new_n45076_, new_n43803_, RIbb2eda0_19 );
and  ( new_n45077_, new_n45076_, new_n1042_ );
or   ( new_n45078_, new_n45077_, new_n45075_ );
xor  ( new_n45079_, new_n45073_, new_n1585_ );
nand ( new_n45080_, new_n45079_, new_n45078_ );
and  ( new_n45081_, new_n45080_, new_n45074_ );
or   ( new_n45082_, new_n44788_, new_n302_ );
or   ( new_n45083_, new_n44884_, new_n44007_ );
and  ( new_n45084_, new_n45083_, new_n45082_ );
xor  ( new_n45085_, new_n44974_, new_n43945_ );
nand ( new_n45086_, new_n45085_, new_n43982_ );
nor  ( new_n45087_, new_n44877_, new_n43880_ );
or   ( new_n45088_, new_n44878_, new_n43977_ );
or   ( new_n45089_, new_n45088_, new_n45087_ );
and  ( new_n45090_, new_n45089_, new_n45086_ );
or   ( new_n45091_, new_n45090_, new_n45084_ );
and  ( new_n45092_, new_n44849_, new_n660_ );
xor  ( new_n45093_, new_n43956_, new_n520_ );
nor  ( new_n45094_, new_n45093_, new_n755_ );
or   ( new_n45095_, new_n45094_, new_n45092_ );
xor  ( new_n45096_, new_n45090_, new_n45084_ );
nand ( new_n45097_, new_n45096_, new_n45095_ );
and  ( new_n45098_, new_n45097_, new_n45091_ );
or   ( new_n45099_, new_n45098_, new_n45081_ );
xor  ( new_n45100_, new_n45098_, new_n45081_ );
xor  ( new_n45101_, new_n44986_, new_n44985_ );
nand ( new_n45102_, new_n45101_, new_n45100_ );
and  ( new_n45103_, new_n45102_, new_n45099_ );
xor  ( new_n45104_, new_n44953_, new_n44952_ );
xor  ( new_n45105_, new_n44853_, new_n44852_ );
nand ( new_n45106_, new_n45105_, new_n45104_ );
xor  ( new_n45107_, new_n45105_, new_n45104_ );
xor  ( new_n45108_, new_n44968_, new_n44967_ );
nand ( new_n45109_, new_n45108_, new_n45107_ );
and  ( new_n45110_, new_n45109_, new_n45106_ );
nor  ( new_n45111_, new_n45110_, new_n45103_ );
xor  ( new_n45112_, new_n44989_, new_n44988_ );
xor  ( new_n45113_, new_n45110_, new_n45103_ );
and  ( new_n45114_, new_n45113_, new_n45112_ );
or   ( new_n45115_, new_n45114_, new_n45111_ );
xor  ( new_n45116_, new_n45028_, new_n45027_ );
and  ( new_n45117_, new_n45116_, new_n45115_ );
xor  ( new_n45118_, RIbb320b8_152, RIbb2cd48_88 );
xnor ( new_n45119_, new_n45118_, new_n43721_ );
and  ( new_n45120_, new_n45119_, new_n43880_ );
not  ( new_n45121_, new_n45120_ );
nor  ( new_n45122_, RIbb2e9e0_27, RIbb2ea58_26 );
not  ( new_n45123_, new_n45122_ );
and  ( new_n45124_, new_n45123_, new_n1585_ );
xor  ( new_n45125_, new_n43793_, new_n1583_ );
and  ( new_n45126_, new_n45125_, new_n1741_ );
nor  ( new_n45127_, new_n45126_, new_n45124_ );
or   ( new_n45128_, new_n45127_, new_n45121_ );
nor  ( new_n45129_, new_n44938_, new_n526_ );
xor  ( new_n45130_, new_n43985_, RIbb2f070_13 );
and  ( new_n45131_, new_n45130_, new_n456_ );
or   ( new_n45132_, new_n45131_, new_n45129_ );
xor  ( new_n45133_, new_n45127_, new_n45121_ );
nand ( new_n45134_, new_n45133_, new_n45132_ );
and  ( new_n45135_, new_n45134_, new_n45128_ );
or   ( new_n45136_, new_n44884_, new_n302_ );
or   ( new_n45137_, new_n44942_, new_n44007_ );
and  ( new_n45138_, new_n45137_, new_n45136_ );
xor  ( new_n45139_, new_n44681_, new_n275_ );
or   ( new_n45140_, new_n45139_, new_n283_ );
or   ( new_n45141_, new_n44917_, new_n286_ );
and  ( new_n45142_, new_n45141_, new_n45140_ );
nor  ( new_n45143_, new_n45142_, new_n45138_ );
xor  ( new_n45144_, new_n43952_, new_n520_ );
nor  ( new_n45145_, new_n45144_, new_n755_ );
nor  ( new_n45146_, new_n45093_, new_n757_ );
nor  ( new_n45147_, new_n45146_, new_n45145_ );
and  ( new_n45148_, new_n45142_, new_n45138_ );
nor  ( new_n45149_, new_n45148_, new_n45147_ );
nor  ( new_n45150_, new_n45149_, new_n45143_ );
or   ( new_n45151_, new_n44899_, new_n899_ );
xor  ( new_n45152_, new_n43937_, RIbb2ee90_17 );
nand ( new_n45153_, new_n45152_, new_n822_ );
and  ( new_n45154_, new_n45153_, new_n45151_ );
xor  ( new_n45155_, new_n44506_, new_n309_ );
or   ( new_n45156_, new_n45155_, new_n317_ );
or   ( new_n45157_, new_n44913_, new_n320_ );
and  ( new_n45158_, new_n45157_, new_n45156_ );
or   ( new_n45159_, new_n45158_, new_n45154_ );
xor  ( new_n45160_, new_n44319_, RIbb2f250_9 );
and  ( new_n45161_, new_n45160_, new_n336_ );
and  ( new_n45162_, new_n44894_, new_n334_ );
or   ( new_n45163_, new_n45162_, new_n45161_ );
xor  ( new_n45164_, new_n45158_, new_n45154_ );
nand ( new_n45165_, new_n45164_, new_n45163_ );
and  ( new_n45166_, new_n45165_, new_n45159_ );
or   ( new_n45167_, new_n45166_, new_n45150_ );
nand ( new_n45168_, new_n45076_, new_n1040_ );
xor  ( new_n45169_, new_n43884_, RIbb2eda0_19 );
nand ( new_n45170_, new_n45169_, new_n1042_ );
and  ( new_n45171_, new_n45170_, new_n45168_ );
or   ( new_n45172_, new_n45070_, new_n1595_ );
xor  ( new_n45173_, new_n43898_, new_n1355_ );
or   ( new_n45174_, new_n45173_, new_n1593_ );
and  ( new_n45175_, new_n45174_, new_n45172_ );
nor  ( new_n45176_, new_n45175_, new_n45171_ );
and  ( new_n45177_, new_n44903_, new_n371_ );
xor  ( new_n45178_, new_n44183_, RIbb2f160_11 );
and  ( new_n45179_, new_n45178_, new_n373_ );
or   ( new_n45180_, new_n45179_, new_n45177_ );
xor  ( new_n45181_, new_n45175_, new_n45171_ );
and  ( new_n45182_, new_n45181_, new_n45180_ );
or   ( new_n45183_, new_n45182_, new_n45176_ );
xor  ( new_n45184_, new_n45166_, new_n45150_ );
nand ( new_n45185_, new_n45184_, new_n45183_ );
and  ( new_n45186_, new_n45185_, new_n45167_ );
nor  ( new_n45187_, new_n45186_, new_n45135_ );
xor  ( new_n45188_, new_n45186_, new_n45135_ );
xor  ( new_n45189_, new_n44929_, new_n44928_ );
and  ( new_n45190_, new_n45189_, new_n45188_ );
or   ( new_n45191_, new_n45190_, new_n45187_ );
xor  ( new_n45192_, new_n45013_, new_n45012_ );
and  ( new_n45193_, new_n45192_, new_n45191_ );
xor  ( new_n45194_, RIbb32130_153, RIbb2ccd0_89 );
nor  ( new_n45195_, new_n43707_, new_n43685_ );
not  ( new_n45196_, new_n45195_ );
and  ( new_n45197_, new_n45196_, new_n43692_ );
nor  ( new_n45198_, new_n45197_, new_n43712_ );
not  ( new_n45199_, new_n45198_ );
and  ( new_n45200_, new_n45199_, new_n43690_ );
nor  ( new_n45201_, new_n45200_, new_n43711_ );
nor  ( new_n45202_, new_n45201_, new_n43686_ );
nor  ( new_n45203_, new_n45202_, new_n43710_ );
xnor ( new_n45204_, new_n45203_, new_n45194_ );
and  ( new_n45205_, new_n45204_, new_n43880_ );
not  ( new_n45206_, new_n45205_ );
xor  ( new_n45207_, new_n45119_, new_n43945_ );
nand ( new_n45208_, new_n45207_, new_n43982_ );
not  ( new_n45209_, new_n44974_ );
and  ( new_n45210_, new_n45209_, new_n43879_ );
or   ( new_n45211_, new_n44975_, new_n43977_ );
or   ( new_n45212_, new_n45211_, new_n45210_ );
and  ( new_n45213_, new_n45212_, new_n45208_ );
nor  ( new_n45214_, new_n45213_, new_n45206_ );
xor  ( new_n45215_, new_n43799_, new_n1126_ );
nor  ( new_n45216_, new_n45215_, new_n1364_ );
and  ( new_n45217_, new_n44921_, new_n1251_ );
or   ( new_n45218_, new_n45217_, new_n45216_ );
xor  ( new_n45219_, new_n45213_, new_n45206_ );
and  ( new_n45220_, new_n45219_, new_n45218_ );
or   ( new_n45221_, new_n45220_, new_n45214_ );
xor  ( new_n45222_, new_n45133_, new_n45132_ );
and  ( new_n45223_, new_n45222_, new_n45221_ );
xor  ( new_n45224_, new_n45222_, new_n45221_ );
xor  ( new_n45225_, new_n44908_, new_n44907_ );
and  ( new_n45226_, new_n45225_, new_n45224_ );
or   ( new_n45227_, new_n45226_, new_n45223_ );
xor  ( new_n45228_, new_n45101_, new_n45100_ );
and  ( new_n45229_, new_n45228_, new_n45227_ );
xor  ( new_n45230_, new_n45079_, new_n45078_ );
xor  ( new_n45231_, new_n45096_, new_n45095_ );
and  ( new_n45232_, new_n45231_, new_n45230_ );
xor  ( new_n45233_, new_n45231_, new_n45230_ );
xor  ( new_n45234_, new_n44926_, new_n44925_ );
and  ( new_n45235_, new_n45234_, new_n45233_ );
or   ( new_n45236_, new_n45235_, new_n45232_ );
xor  ( new_n45237_, new_n45228_, new_n45227_ );
and  ( new_n45238_, new_n45237_, new_n45236_ );
or   ( new_n45239_, new_n45238_, new_n45229_ );
xor  ( new_n45240_, new_n45192_, new_n45191_ );
and  ( new_n45241_, new_n45240_, new_n45239_ );
or   ( new_n45242_, new_n45241_, new_n45193_ );
xor  ( new_n45243_, new_n45116_, new_n45115_ );
and  ( new_n45244_, new_n45243_, new_n45242_ );
nor  ( new_n45245_, new_n45244_, new_n45117_ );
xnor ( new_n45246_, new_n45068_, new_n44937_ );
or   ( new_n45247_, new_n45246_, new_n45245_ );
and  ( new_n45248_, new_n45247_, new_n45069_ );
and  ( new_n45249_, new_n45046_, new_n45030_ );
and  ( new_n45250_, new_n45067_, new_n45047_ );
nor  ( new_n45251_, new_n45250_, new_n45249_ );
and  ( new_n45252_, new_n45060_, new_n45056_ );
and  ( new_n45253_, new_n45066_, new_n45061_ );
or   ( new_n45254_, new_n45253_, new_n45252_ );
nor  ( new_n45255_, new_n45044_, new_n45041_ );
and  ( new_n45256_, new_n45045_, new_n45038_ );
or   ( new_n45257_, new_n45256_, new_n45255_ );
and  ( new_n45258_, new_n45063_, new_n45062_ );
and  ( new_n45259_, new_n45065_, new_n45064_ );
or   ( new_n45260_, new_n45259_, new_n45258_ );
nor  ( new_n45261_, new_n45036_, new_n44806_ );
and  ( new_n45262_, new_n45037_, new_n45033_ );
or   ( new_n45263_, new_n45262_, new_n45261_ );
xor  ( new_n45264_, new_n44663_, new_n44662_ );
xor  ( new_n45265_, new_n45264_, new_n45263_ );
xor  ( new_n45266_, new_n45265_, new_n45260_ );
xor  ( new_n45267_, new_n45266_, new_n45257_ );
and  ( new_n45268_, new_n45054_, new_n45053_ );
and  ( new_n45269_, new_n45055_, new_n45050_ );
or   ( new_n45270_, new_n45269_, new_n45268_ );
xor  ( new_n45271_, new_n44713_, new_n44712_ );
xor  ( new_n45272_, new_n45271_, new_n45270_ );
xor  ( new_n45273_, new_n44726_, new_n44725_ );
xor  ( new_n45274_, new_n45273_, new_n45272_ );
xor  ( new_n45275_, new_n45274_, new_n45267_ );
xnor ( new_n45276_, new_n45275_, new_n45254_ );
xnor ( new_n45277_, new_n45276_, new_n45251_ );
and  ( new_n45278_, new_n45277_, new_n45248_ );
nand ( new_n45279_, new_n45275_, new_n45254_ );
or   ( new_n45280_, new_n45276_, new_n45251_ );
and  ( new_n45281_, new_n45280_, new_n45279_ );
and  ( new_n45282_, new_n45266_, new_n45257_ );
and  ( new_n45283_, new_n45274_, new_n45267_ );
nor  ( new_n45284_, new_n45283_, new_n45282_ );
and  ( new_n45285_, new_n45271_, new_n45270_ );
and  ( new_n45286_, new_n45273_, new_n45272_ );
or   ( new_n45287_, new_n45286_, new_n45285_ );
and  ( new_n45288_, new_n45264_, new_n45263_ );
and  ( new_n45289_, new_n45265_, new_n45260_ );
or   ( new_n45290_, new_n45289_, new_n45288_ );
xor  ( new_n45291_, new_n44716_, new_n44715_ );
xor  ( new_n45292_, new_n45291_, new_n45290_ );
xor  ( new_n45293_, new_n44732_, new_n44731_ );
xor  ( new_n45294_, new_n45293_, new_n45292_ );
xnor ( new_n45295_, new_n45294_, new_n45287_ );
xnor ( new_n45296_, new_n45295_, new_n45284_ );
and  ( new_n45297_, new_n45296_, new_n45281_ );
or   ( new_n45298_, new_n45297_, new_n45278_ );
xor  ( new_n45299_, new_n44932_, new_n44931_ );
xor  ( new_n45300_, new_n45113_, new_n45112_ );
and  ( new_n45301_, new_n45300_, new_n45299_ );
nand ( new_n45302_, new_n45130_, new_n454_ );
xor  ( new_n45303_, new_n43812_, new_n400_ );
or   ( new_n45304_, new_n45303_, new_n524_ );
nand ( new_n45305_, new_n45304_, new_n45302_ );
nand ( new_n45306_, new_n45305_, new_n45127_ );
xor  ( new_n45307_, new_n44785_, new_n275_ );
or   ( new_n45308_, new_n45307_, new_n283_ );
or   ( new_n45309_, new_n45139_, new_n286_ );
and  ( new_n45310_, new_n45309_, new_n45308_ );
or   ( new_n45311_, new_n45085_, new_n44007_ );
or   ( new_n45312_, new_n44942_, new_n302_ );
and  ( new_n45313_, new_n45312_, new_n45311_ );
nor  ( new_n45314_, new_n45313_, new_n45310_ );
xor  ( new_n45315_, new_n43956_, new_n745_ );
nor  ( new_n45316_, new_n45315_, new_n897_ );
and  ( new_n45317_, new_n45152_, new_n820_ );
nor  ( new_n45318_, new_n45317_, new_n45316_ );
and  ( new_n45319_, new_n45313_, new_n45310_ );
nor  ( new_n45320_, new_n45319_, new_n45318_ );
or   ( new_n45321_, new_n45320_, new_n45314_ );
xor  ( new_n45322_, new_n45305_, new_n45127_ );
nand ( new_n45323_, new_n45322_, new_n45321_ );
and  ( new_n45324_, new_n45323_, new_n45306_ );
xor  ( new_n45325_, new_n43787_, new_n1583_ );
or   ( new_n45326_, new_n45325_, new_n1844_ );
nand ( new_n45327_, new_n45125_, new_n1739_ );
and  ( new_n45328_, new_n45327_, new_n45326_ );
or   ( new_n45329_, new_n45328_, new_n1842_ );
nor  ( new_n45330_, new_n45215_, new_n1366_ );
xor  ( new_n45331_, new_n43803_, RIbb2ecb0_21 );
and  ( new_n45332_, new_n45331_, new_n1253_ );
or   ( new_n45333_, new_n45332_, new_n45330_ );
xor  ( new_n45334_, new_n45328_, new_n1842_ );
nand ( new_n45335_, new_n45334_, new_n45333_ );
and  ( new_n45336_, new_n45335_, new_n45329_ );
nand ( new_n45337_, new_n45178_, new_n371_ );
xor  ( new_n45338_, new_n44218_, new_n325_ );
or   ( new_n45339_, new_n45338_, new_n409_ );
and  ( new_n45340_, new_n45339_, new_n45337_ );
or   ( new_n45341_, new_n45303_, new_n526_ );
xor  ( new_n45342_, new_n43914_, RIbb2f070_13 );
nand ( new_n45343_, new_n45342_, new_n456_ );
and  ( new_n45344_, new_n45343_, new_n45341_ );
or   ( new_n45345_, new_n45344_, new_n45340_ );
and  ( new_n45346_, new_n45344_, new_n45340_ );
and  ( new_n45347_, new_n45169_, new_n1040_ );
xor  ( new_n45348_, new_n43888_, RIbb2eda0_19 );
and  ( new_n45349_, new_n45348_, new_n1042_ );
nor  ( new_n45350_, new_n45349_, new_n45347_ );
or   ( new_n45351_, new_n45350_, new_n45346_ );
and  ( new_n45352_, new_n45351_, new_n45345_ );
or   ( new_n45353_, new_n45352_, new_n45336_ );
and  ( new_n45354_, new_n45352_, new_n45336_ );
or   ( new_n45355_, new_n45155_, new_n320_ );
xor  ( new_n45356_, new_n44600_, new_n309_ );
or   ( new_n45357_, new_n45356_, new_n317_ );
and  ( new_n45358_, new_n45357_, new_n45355_ );
nand ( new_n45359_, new_n45160_, new_n334_ );
xor  ( new_n45360_, new_n44407_, RIbb2f250_9 );
nand ( new_n45361_, new_n45360_, new_n336_ );
and  ( new_n45362_, new_n45361_, new_n45359_ );
nor  ( new_n45363_, new_n45362_, new_n45358_ );
xor  ( new_n45364_, new_n43894_, RIbb2ebc0_23 );
and  ( new_n45365_, new_n45364_, new_n1476_ );
nor  ( new_n45366_, new_n45173_, new_n1595_ );
nor  ( new_n45367_, new_n45366_, new_n45365_ );
and  ( new_n45368_, new_n45362_, new_n45358_ );
nor  ( new_n45369_, new_n45368_, new_n45367_ );
nor  ( new_n45370_, new_n45369_, new_n45363_ );
or   ( new_n45371_, new_n45370_, new_n45354_ );
and  ( new_n45372_, new_n45371_, new_n45353_ );
nor  ( new_n45373_, new_n45372_, new_n45324_ );
xor  ( new_n45374_, new_n45184_, new_n45183_ );
xor  ( new_n45375_, new_n45372_, new_n45324_ );
and  ( new_n45376_, new_n45375_, new_n45374_ );
or   ( new_n45377_, new_n45376_, new_n45373_ );
xor  ( new_n45378_, new_n45108_, new_n45107_ );
and  ( new_n45379_, new_n45378_, new_n45377_ );
xor  ( new_n45380_, new_n45189_, new_n45188_ );
xor  ( new_n45381_, new_n45378_, new_n45377_ );
and  ( new_n45382_, new_n45381_, new_n45380_ );
or   ( new_n45383_, new_n45382_, new_n45379_ );
xor  ( new_n45384_, new_n45300_, new_n45299_ );
and  ( new_n45385_, new_n45384_, new_n45383_ );
nor  ( new_n45386_, new_n45385_, new_n45301_ );
not  ( new_n45387_, new_n45386_ );
xor  ( new_n45388_, new_n44935_, new_n44934_ );
nand ( new_n45389_, new_n45388_, new_n45387_ );
xor  ( new_n45390_, new_n45388_, new_n45387_ );
xor  ( new_n45391_, new_n45243_, new_n45242_ );
nand ( new_n45392_, new_n45391_, new_n45390_ );
and  ( new_n45393_, new_n45392_, new_n45389_ );
xnor ( new_n45394_, new_n45246_, new_n45245_ );
and  ( new_n45395_, new_n45394_, new_n45393_ );
or   ( new_n45396_, new_n45395_, new_n45298_ );
xnor ( new_n45397_, new_n45391_, new_n45390_ );
xor  ( new_n45398_, new_n45240_, new_n45239_ );
xor  ( new_n45399_, new_n45384_, new_n45383_ );
nand ( new_n45400_, new_n45399_, new_n45398_ );
nor  ( new_n45401_, new_n45399_, new_n45398_ );
xor  ( new_n45402_, RIbb321a8_154, RIbb2cc58_90 );
xnor ( new_n45403_, new_n45402_, new_n45201_ );
and  ( new_n45404_, new_n45403_, new_n43880_ );
not  ( new_n45405_, new_n45404_ );
xor  ( new_n45406_, new_n45204_, new_n43945_ );
nand ( new_n45407_, new_n45406_, new_n43982_ );
nor  ( new_n45408_, new_n45119_, new_n43880_ );
or   ( new_n45409_, new_n45120_, new_n43977_ );
or   ( new_n45410_, new_n45409_, new_n45408_ );
and  ( new_n45411_, new_n45410_, new_n45407_ );
nor  ( new_n45412_, new_n45411_, new_n45405_ );
nor  ( new_n45413_, new_n45144_, new_n757_ );
xor  ( new_n45414_, new_n43985_, RIbb2ef80_15 );
and  ( new_n45415_, new_n45414_, new_n662_ );
or   ( new_n45416_, new_n45415_, new_n45413_ );
xor  ( new_n45417_, new_n45411_, new_n45405_ );
and  ( new_n45418_, new_n45417_, new_n45416_ );
or   ( new_n45419_, new_n45418_, new_n45412_ );
xor  ( new_n45420_, new_n45219_, new_n45218_ );
and  ( new_n45421_, new_n45420_, new_n45419_ );
xor  ( new_n45422_, new_n45420_, new_n45419_ );
xor  ( new_n45423_, new_n45181_, new_n45180_ );
and  ( new_n45424_, new_n45423_, new_n45422_ );
or   ( new_n45425_, new_n45424_, new_n45421_ );
xor  ( new_n45426_, new_n45225_, new_n45224_ );
and  ( new_n45427_, new_n45426_, new_n45425_ );
xor  ( new_n45428_, new_n45426_, new_n45425_ );
xor  ( new_n45429_, new_n45234_, new_n45233_ );
and  ( new_n45430_, new_n45429_, new_n45428_ );
or   ( new_n45431_, new_n45430_, new_n45427_ );
xor  ( new_n45432_, new_n45237_, new_n45236_ );
nand ( new_n45433_, new_n45432_, new_n45431_ );
xor  ( new_n45434_, new_n45164_, new_n45163_ );
xnor ( new_n45435_, new_n45142_, new_n45138_ );
nand ( new_n45436_, new_n45435_, new_n45147_ );
not  ( new_n45437_, new_n45149_ );
or   ( new_n45438_, new_n45437_, new_n45143_ );
and  ( new_n45439_, new_n45438_, new_n45436_ );
nand ( new_n45440_, new_n45439_, new_n45434_ );
not  ( new_n45441_, RIbb2e968_28 );
and  ( new_n45442_, new_n2118_, new_n45441_ );
not  ( new_n45443_, new_n45442_ );
and  ( new_n45444_, new_n45443_, new_n1842_ );
xor  ( new_n45445_, new_n43793_, new_n1840_ );
and  ( new_n45446_, new_n45445_, new_n2002_ );
nor  ( new_n45447_, new_n45446_, new_n45444_ );
nand ( new_n45448_, new_n45348_, new_n1040_ );
xor  ( new_n45449_, new_n43937_, RIbb2eda0_19 );
nand ( new_n45450_, new_n45449_, new_n1042_ );
and  ( new_n45451_, new_n45450_, new_n45448_ );
xor  ( new_n45452_, new_n44319_, new_n325_ );
or   ( new_n45453_, new_n45452_, new_n409_ );
or   ( new_n45454_, new_n45338_, new_n411_ );
and  ( new_n45455_, new_n45454_, new_n45453_ );
or   ( new_n45456_, new_n45455_, new_n45451_ );
and  ( new_n45457_, new_n45360_, new_n334_ );
xor  ( new_n45458_, new_n44506_, RIbb2f250_9 );
and  ( new_n45459_, new_n45458_, new_n336_ );
nor  ( new_n45460_, new_n45459_, new_n45457_ );
and  ( new_n45461_, new_n45455_, new_n45451_ );
or   ( new_n45462_, new_n45461_, new_n45460_ );
and  ( new_n45463_, new_n45462_, new_n45456_ );
nor  ( new_n45464_, new_n45463_, new_n45447_ );
or   ( new_n45465_, new_n45325_, new_n1846_ );
xor  ( new_n45466_, new_n43898_, new_n1583_ );
or   ( new_n45467_, new_n45466_, new_n1844_ );
and  ( new_n45468_, new_n45467_, new_n45465_ );
nand ( new_n45469_, new_n45331_, new_n1251_ );
xor  ( new_n45470_, new_n43884_, RIbb2ecb0_21 );
nand ( new_n45471_, new_n45470_, new_n1253_ );
and  ( new_n45472_, new_n45471_, new_n45469_ );
nor  ( new_n45473_, new_n45472_, new_n45468_ );
and  ( new_n45474_, new_n45342_, new_n454_ );
xor  ( new_n45475_, new_n44183_, RIbb2f070_13 );
and  ( new_n45476_, new_n45475_, new_n456_ );
or   ( new_n45477_, new_n45476_, new_n45474_ );
xor  ( new_n45478_, new_n45472_, new_n45468_ );
and  ( new_n45479_, new_n45478_, new_n45477_ );
or   ( new_n45480_, new_n45479_, new_n45473_ );
xor  ( new_n45481_, new_n45463_, new_n45447_ );
and  ( new_n45482_, new_n45481_, new_n45480_ );
or   ( new_n45483_, new_n45482_, new_n45464_ );
xor  ( new_n45484_, new_n45439_, new_n45434_ );
nand ( new_n45485_, new_n45484_, new_n45483_ );
and  ( new_n45486_, new_n45485_, new_n45440_ );
xor  ( new_n45487_, new_n45322_, new_n45321_ );
xnor ( new_n45488_, new_n45352_, new_n45336_ );
xor  ( new_n45489_, new_n45488_, new_n45370_ );
nand ( new_n45490_, new_n45489_, new_n45487_ );
xor  ( new_n45491_, new_n45334_, new_n45333_ );
xnor ( new_n45492_, new_n45313_, new_n45310_ );
nand ( new_n45493_, new_n45492_, new_n45318_ );
not  ( new_n45494_, new_n45314_ );
nand ( new_n45495_, new_n45320_, new_n45494_ );
and  ( new_n45496_, new_n45495_, new_n45493_ );
and  ( new_n45497_, new_n45496_, new_n45491_ );
xor  ( new_n45498_, new_n45496_, new_n45491_ );
xor  ( new_n45499_, new_n45417_, new_n45416_ );
and  ( new_n45500_, new_n45499_, new_n45498_ );
or   ( new_n45501_, new_n45500_, new_n45497_ );
xor  ( new_n45502_, new_n45489_, new_n45487_ );
nand ( new_n45503_, new_n45502_, new_n45501_ );
and  ( new_n45504_, new_n45503_, new_n45490_ );
nor  ( new_n45505_, new_n45504_, new_n45486_ );
xor  ( new_n45506_, new_n45504_, new_n45486_ );
xor  ( new_n45507_, new_n45375_, new_n45374_ );
and  ( new_n45508_, new_n45507_, new_n45506_ );
nor  ( new_n45509_, new_n45508_, new_n45505_ );
not  ( new_n45510_, new_n45509_ );
xor  ( new_n45511_, new_n45432_, new_n45431_ );
nand ( new_n45512_, new_n45511_, new_n45510_ );
and  ( new_n45513_, new_n45512_, new_n45433_ );
or   ( new_n45514_, new_n45513_, new_n45401_ );
and  ( new_n45515_, new_n45514_, new_n45400_ );
and  ( new_n45516_, new_n45515_, new_n45397_ );
xor  ( new_n45517_, new_n44681_, new_n309_ );
or   ( new_n45518_, new_n45517_, new_n317_ );
or   ( new_n45519_, new_n45356_, new_n320_ );
and  ( new_n45520_, new_n45519_, new_n45518_ );
xor  ( new_n45521_, new_n43952_, new_n745_ );
or   ( new_n45522_, new_n45521_, new_n897_ );
or   ( new_n45523_, new_n45315_, new_n899_ );
and  ( new_n45524_, new_n45523_, new_n45522_ );
nor  ( new_n45525_, new_n45524_, new_n45520_ );
and  ( new_n45526_, new_n45364_, new_n1474_ );
xor  ( new_n45527_, new_n43799_, new_n1355_ );
nor  ( new_n45528_, new_n45527_, new_n1593_ );
nor  ( new_n45529_, new_n45528_, new_n45526_ );
and  ( new_n45530_, new_n45524_, new_n45520_ );
nor  ( new_n45531_, new_n45530_, new_n45529_ );
nor  ( new_n45532_, new_n45531_, new_n45525_ );
or   ( new_n45533_, new_n45307_, new_n286_ );
xor  ( new_n45534_, new_n44877_, new_n275_ );
or   ( new_n45535_, new_n45534_, new_n283_ );
and  ( new_n45536_, new_n45535_, new_n45533_ );
or   ( new_n45537_, new_n45207_, new_n44007_ );
or   ( new_n45538_, new_n45085_, new_n302_ );
and  ( new_n45539_, new_n45538_, new_n45537_ );
or   ( new_n45540_, new_n45539_, new_n45536_ );
and  ( new_n45541_, new_n45414_, new_n660_ );
xor  ( new_n45542_, new_n43812_, RIbb2ef80_15 );
and  ( new_n45543_, new_n45542_, new_n662_ );
or   ( new_n45544_, new_n45543_, new_n45541_ );
xor  ( new_n45545_, new_n45539_, new_n45536_ );
nand ( new_n45546_, new_n45545_, new_n45544_ );
and  ( new_n45547_, new_n45546_, new_n45540_ );
nor  ( new_n45548_, new_n45547_, new_n45532_ );
xor  ( new_n45549_, new_n45547_, new_n45532_ );
xnor ( new_n45550_, new_n45344_, new_n45340_ );
xor  ( new_n45551_, new_n45550_, new_n45350_ );
and  ( new_n45552_, new_n45551_, new_n45549_ );
or   ( new_n45553_, new_n45552_, new_n45548_ );
xor  ( new_n45554_, new_n45423_, new_n45422_ );
and  ( new_n45555_, new_n45554_, new_n45553_ );
xor  ( new_n45556_, new_n45554_, new_n45553_ );
xor  ( new_n45557_, new_n45484_, new_n45483_ );
and  ( new_n45558_, new_n45557_, new_n45556_ );
nor  ( new_n45559_, new_n45558_, new_n45555_ );
not  ( new_n45560_, new_n45559_ );
xor  ( new_n45561_, new_n45429_, new_n45428_ );
and  ( new_n45562_, new_n45561_, new_n45560_ );
xor  ( new_n45563_, new_n45561_, new_n45560_ );
xor  ( new_n45564_, new_n45507_, new_n45506_ );
and  ( new_n45565_, new_n45564_, new_n45563_ );
or   ( new_n45566_, new_n45565_, new_n45562_ );
xor  ( new_n45567_, new_n45381_, new_n45380_ );
nand ( new_n45568_, new_n45567_, new_n45566_ );
xor  ( new_n45569_, new_n45511_, new_n45510_ );
xor  ( new_n45570_, new_n45567_, new_n45566_ );
nand ( new_n45571_, new_n45570_, new_n45569_ );
and  ( new_n45572_, new_n45571_, new_n45568_ );
xor  ( new_n45573_, new_n45399_, new_n45398_ );
xor  ( new_n45574_, new_n45573_, new_n45513_ );
and  ( new_n45575_, new_n45574_, new_n45572_ );
or   ( new_n45576_, new_n45575_, new_n45516_ );
nor  ( new_n45577_, RIbb2e800_31, RIbb2e878_30 );
not  ( new_n45578_, new_n45577_ );
and  ( new_n45579_, new_n45578_, new_n2120_ );
xor  ( new_n45580_, new_n43793_, new_n2118_ );
and  ( new_n45581_, new_n45580_, new_n2244_ );
nor  ( new_n45582_, new_n45581_, new_n45579_ );
xor  ( new_n45583_, RIbb32220_155, RIbb2cbe0_91 );
xor  ( new_n45584_, new_n45583_, new_n45199_ );
xor  ( new_n45585_, new_n45584_, new_n43945_ );
not  ( new_n45586_, new_n45585_ );
or   ( new_n45587_, new_n45586_, new_n43983_ );
nor  ( new_n45588_, new_n45403_, new_n43880_ );
or   ( new_n45589_, new_n45404_, new_n43977_ );
or   ( new_n45590_, new_n45589_, new_n45588_ );
and  ( new_n45591_, new_n45590_, new_n45587_ );
nor  ( new_n45592_, new_n45591_, new_n45582_ );
xor  ( new_n45593_, RIbb32310_157, RIbb2caf0_93 );
nor  ( new_n45594_, new_n43702_, new_n43684_ );
nor  ( new_n45595_, new_n45594_, new_n43488_ );
nor  ( new_n45596_, new_n45595_, new_n43698_ );
xnor ( new_n45597_, new_n45596_, new_n45593_ );
and  ( new_n45598_, new_n45597_, new_n43880_ );
not  ( new_n45599_, new_n45598_ );
xor  ( new_n45600_, new_n43787_, new_n1840_ );
or   ( new_n45601_, new_n45600_, new_n2124_ );
xor  ( new_n45602_, new_n43898_, new_n1840_ );
or   ( new_n45603_, new_n45602_, new_n2122_ );
and  ( new_n45604_, new_n45603_, new_n45601_ );
nor  ( new_n45605_, new_n45604_, new_n45599_ );
xor  ( new_n45606_, new_n43803_, RIbb2ebc0_23 );
and  ( new_n45607_, new_n45606_, new_n1474_ );
xor  ( new_n45608_, new_n43884_, RIbb2ebc0_23 );
and  ( new_n45609_, new_n45608_, new_n1476_ );
or   ( new_n45610_, new_n45609_, new_n45607_ );
xor  ( new_n45611_, new_n45604_, new_n45599_ );
and  ( new_n45612_, new_n45611_, new_n45610_ );
or   ( new_n45613_, new_n45612_, new_n45605_ );
xor  ( new_n45614_, new_n45591_, new_n45582_ );
and  ( new_n45615_, new_n45614_, new_n45613_ );
or   ( new_n45616_, new_n45615_, new_n45592_ );
xnor ( new_n45617_, new_n45524_, new_n45520_ );
nand ( new_n45618_, new_n45617_, new_n45529_ );
not  ( new_n45619_, new_n45531_ );
or   ( new_n45620_, new_n45619_, new_n45525_ );
and  ( new_n45621_, new_n45620_, new_n45618_ );
and  ( new_n45622_, new_n45621_, new_n45616_ );
xor  ( new_n45623_, new_n43888_, RIbb2ecb0_21 );
nand ( new_n45624_, new_n45623_, new_n1251_ );
xor  ( new_n45625_, new_n43937_, new_n1126_ );
or   ( new_n45626_, new_n45625_, new_n1364_ );
and  ( new_n45627_, new_n45626_, new_n45624_ );
xor  ( new_n45628_, new_n44319_, RIbb2f070_13 );
nand ( new_n45629_, new_n45628_, new_n456_ );
xor  ( new_n45630_, new_n44218_, new_n400_ );
or   ( new_n45631_, new_n45630_, new_n526_ );
and  ( new_n45632_, new_n45631_, new_n45629_ );
or   ( new_n45633_, new_n45632_, new_n45627_ );
xor  ( new_n45634_, new_n44183_, RIbb2ef80_15 );
and  ( new_n45635_, new_n45634_, new_n662_ );
xor  ( new_n45636_, new_n43914_, RIbb2ef80_15 );
and  ( new_n45637_, new_n45636_, new_n660_ );
or   ( new_n45638_, new_n45637_, new_n45635_ );
xor  ( new_n45639_, new_n45632_, new_n45627_ );
nand ( new_n45640_, new_n45639_, new_n45638_ );
and  ( new_n45641_, new_n45640_, new_n45633_ );
xor  ( new_n45642_, new_n44407_, new_n325_ );
or   ( new_n45643_, new_n45642_, new_n411_ );
xor  ( new_n45644_, new_n44506_, RIbb2f160_11 );
nand ( new_n45645_, new_n45644_, new_n373_ );
and  ( new_n45646_, new_n45645_, new_n45643_ );
xor  ( new_n45647_, new_n43894_, new_n1583_ );
or   ( new_n45648_, new_n45647_, new_n1846_ );
xor  ( new_n45649_, new_n43799_, new_n1583_ );
or   ( new_n45650_, new_n45649_, new_n1844_ );
and  ( new_n45651_, new_n45650_, new_n45648_ );
or   ( new_n45652_, new_n45651_, new_n45646_ );
xor  ( new_n45653_, new_n44681_, RIbb2f250_9 );
and  ( new_n45654_, new_n45653_, new_n336_ );
xor  ( new_n45655_, new_n44600_, RIbb2f250_9 );
and  ( new_n45656_, new_n45655_, new_n334_ );
or   ( new_n45657_, new_n45656_, new_n45654_ );
xor  ( new_n45658_, new_n45651_, new_n45646_ );
nand ( new_n45659_, new_n45658_, new_n45657_ );
and  ( new_n45660_, new_n45659_, new_n45652_ );
nor  ( new_n45661_, new_n45660_, new_n45641_ );
xor  ( new_n45662_, new_n43952_, new_n893_ );
or   ( new_n45663_, new_n45662_, new_n1135_ );
xor  ( new_n45664_, new_n43956_, new_n893_ );
or   ( new_n45665_, new_n45664_, new_n1137_ );
and  ( new_n45666_, new_n45665_, new_n45663_ );
xor  ( new_n45667_, new_n44877_, new_n309_ );
or   ( new_n45668_, new_n45667_, new_n317_ );
xor  ( new_n45669_, new_n44785_, new_n309_ );
or   ( new_n45670_, new_n45669_, new_n320_ );
and  ( new_n45671_, new_n45670_, new_n45668_ );
nor  ( new_n45672_, new_n45671_, new_n45666_ );
xor  ( new_n45673_, new_n45119_, new_n275_ );
nor  ( new_n45674_, new_n45673_, new_n283_ );
xor  ( new_n45675_, new_n44974_, RIbb2f430_5 );
and  ( new_n45676_, new_n45675_, new_n280_ );
or   ( new_n45677_, new_n45676_, new_n45674_ );
xor  ( new_n45678_, new_n45671_, new_n45666_ );
and  ( new_n45679_, new_n45678_, new_n45677_ );
or   ( new_n45680_, new_n45679_, new_n45672_ );
xor  ( new_n45681_, new_n45660_, new_n45641_ );
and  ( new_n45682_, new_n45681_, new_n45680_ );
nor  ( new_n45683_, new_n45682_, new_n45661_ );
xnor ( new_n45684_, new_n45621_, new_n45616_ );
nor  ( new_n45685_, new_n45684_, new_n45683_ );
nor  ( new_n45686_, new_n45685_, new_n45622_ );
not  ( new_n45687_, new_n45686_ );
xor  ( new_n45688_, new_n45551_, new_n45549_ );
nand ( new_n45689_, new_n45675_, new_n282_ );
or   ( new_n45690_, new_n45534_, new_n286_ );
and  ( new_n45691_, new_n45690_, new_n45689_ );
or   ( new_n45692_, new_n45207_, new_n302_ );
or   ( new_n45693_, new_n45406_, new_n44007_ );
and  ( new_n45694_, new_n45693_, new_n45692_ );
or   ( new_n45695_, new_n45694_, new_n45691_ );
nor  ( new_n45696_, new_n45521_, new_n899_ );
xor  ( new_n45697_, new_n43985_, RIbb2ee90_17 );
and  ( new_n45698_, new_n45697_, new_n822_ );
or   ( new_n45699_, new_n45698_, new_n45696_ );
xor  ( new_n45700_, new_n45694_, new_n45691_ );
nand ( new_n45701_, new_n45700_, new_n45699_ );
and  ( new_n45702_, new_n45701_, new_n45695_ );
or   ( new_n45703_, new_n45517_, new_n320_ );
or   ( new_n45704_, new_n45669_, new_n317_ );
and  ( new_n45705_, new_n45704_, new_n45703_ );
or   ( new_n45706_, new_n45647_, new_n1844_ );
or   ( new_n45707_, new_n45466_, new_n1846_ );
and  ( new_n45708_, new_n45707_, new_n45706_ );
nor  ( new_n45709_, new_n45708_, new_n45705_ );
nor  ( new_n45710_, new_n45664_, new_n1135_ );
and  ( new_n45711_, new_n45449_, new_n1040_ );
nor  ( new_n45712_, new_n45711_, new_n45710_ );
and  ( new_n45713_, new_n45708_, new_n45705_ );
nor  ( new_n45714_, new_n45713_, new_n45712_ );
nor  ( new_n45715_, new_n45714_, new_n45709_ );
nor  ( new_n45716_, new_n45715_, new_n45702_ );
and  ( new_n45717_, new_n45584_, new_n43880_ );
xnor ( new_n45718_, new_n45717_, new_n45447_ );
xor  ( new_n45719_, new_n45403_, new_n43945_ );
not  ( new_n45720_, new_n45719_ );
or   ( new_n45721_, new_n45720_, new_n43983_ );
not  ( new_n45722_, new_n45204_ );
and  ( new_n45723_, new_n45722_, new_n43879_ );
or   ( new_n45724_, new_n45205_, new_n43977_ );
or   ( new_n45725_, new_n45724_, new_n45723_ );
and  ( new_n45726_, new_n45725_, new_n45721_ );
xor  ( new_n45727_, new_n45726_, new_n45718_ );
xor  ( new_n45728_, new_n45715_, new_n45702_ );
and  ( new_n45729_, new_n45728_, new_n45727_ );
or   ( new_n45730_, new_n45729_, new_n45716_ );
xor  ( new_n45731_, new_n45481_, new_n45480_ );
xor  ( new_n45732_, new_n45731_, new_n45730_ );
xor  ( new_n45733_, new_n45732_, new_n45688_ );
and  ( new_n45734_, new_n45733_, new_n45687_ );
xor  ( new_n45735_, new_n45733_, new_n45687_ );
xor  ( new_n45736_, new_n45728_, new_n45727_ );
xor  ( new_n45737_, RIbb32298_156, RIbb2cb68_92 );
xor  ( new_n45738_, new_n45737_, new_n45196_ );
and  ( new_n45739_, new_n45738_, new_n43880_ );
not  ( new_n45740_, new_n45739_ );
nand ( new_n45741_, new_n45475_, new_n454_ );
or   ( new_n45742_, new_n45630_, new_n524_ );
and  ( new_n45743_, new_n45742_, new_n45741_ );
nor  ( new_n45744_, new_n45743_, new_n45740_ );
and  ( new_n45745_, new_n45636_, new_n662_ );
and  ( new_n45746_, new_n45542_, new_n660_ );
or   ( new_n45747_, new_n45746_, new_n45745_ );
xor  ( new_n45748_, new_n45743_, new_n45740_ );
and  ( new_n45749_, new_n45748_, new_n45747_ );
nor  ( new_n45750_, new_n45749_, new_n45744_ );
or   ( new_n45751_, new_n45600_, new_n2122_ );
nand ( new_n45752_, new_n45445_, new_n2000_ );
and  ( new_n45753_, new_n45752_, new_n45751_ );
or   ( new_n45754_, new_n45753_, new_n2120_ );
nor  ( new_n45755_, new_n45527_, new_n1595_ );
and  ( new_n45756_, new_n45606_, new_n1476_ );
or   ( new_n45757_, new_n45756_, new_n45755_ );
xor  ( new_n45758_, new_n45753_, new_n2120_ );
nand ( new_n45759_, new_n45758_, new_n45757_ );
and  ( new_n45760_, new_n45759_, new_n45754_ );
xnor ( new_n45761_, new_n45760_, new_n45750_ );
and  ( new_n45762_, new_n45470_, new_n1251_ );
and  ( new_n45763_, new_n45623_, new_n1253_ );
nor  ( new_n45764_, new_n45763_, new_n45762_ );
or   ( new_n45765_, new_n45452_, new_n411_ );
or   ( new_n45766_, new_n45642_, new_n409_ );
and  ( new_n45767_, new_n45766_, new_n45765_ );
nor  ( new_n45768_, new_n45767_, new_n45764_ );
and  ( new_n45769_, new_n45767_, new_n45764_ );
and  ( new_n45770_, new_n45655_, new_n336_ );
and  ( new_n45771_, new_n45458_, new_n334_ );
nor  ( new_n45772_, new_n45771_, new_n45770_ );
nor  ( new_n45773_, new_n45772_, new_n45769_ );
nor  ( new_n45774_, new_n45773_, new_n45768_ );
xor  ( new_n45775_, new_n45774_, new_n45761_ );
or   ( new_n45776_, new_n45775_, new_n45736_ );
and  ( new_n45777_, new_n45775_, new_n45736_ );
xor  ( new_n45778_, new_n45700_, new_n45699_ );
xnor ( new_n45779_, new_n45708_, new_n45705_ );
nand ( new_n45780_, new_n45779_, new_n45712_ );
not  ( new_n45781_, new_n45714_ );
or   ( new_n45782_, new_n45781_, new_n45709_ );
and  ( new_n45783_, new_n45782_, new_n45780_ );
nor  ( new_n45784_, new_n45783_, new_n45778_ );
and  ( new_n45785_, new_n45783_, new_n45778_ );
xor  ( new_n45786_, new_n45767_, new_n45764_ );
not  ( new_n45787_, new_n45786_ );
and  ( new_n45788_, new_n45787_, new_n45772_ );
not  ( new_n45789_, new_n45768_ );
and  ( new_n45790_, new_n45773_, new_n45789_ );
nor  ( new_n45791_, new_n45790_, new_n45788_ );
nor  ( new_n45792_, new_n45791_, new_n45785_ );
nor  ( new_n45793_, new_n45792_, new_n45784_ );
or   ( new_n45794_, new_n45793_, new_n45777_ );
and  ( new_n45795_, new_n45794_, new_n45776_ );
and  ( new_n45796_, new_n45795_, new_n45735_ );
nor  ( new_n45797_, new_n45796_, new_n45734_ );
not  ( new_n45798_, new_n45797_ );
xor  ( new_n45799_, new_n45499_, new_n45498_ );
xor  ( new_n45800_, new_n45545_, new_n45544_ );
xnor ( new_n45801_, new_n45455_, new_n45451_ );
xor  ( new_n45802_, new_n45801_, new_n45460_ );
or   ( new_n45803_, new_n45802_, new_n45800_ );
and  ( new_n45804_, new_n45802_, new_n45800_ );
xor  ( new_n45805_, new_n45478_, new_n45477_ );
or   ( new_n45806_, new_n45805_, new_n45804_ );
and  ( new_n45807_, new_n45806_, new_n45803_ );
and  ( new_n45808_, new_n45807_, new_n45799_ );
xor  ( new_n45809_, new_n45807_, new_n45799_ );
and  ( new_n45810_, new_n45717_, new_n45447_ );
nor  ( new_n45811_, new_n45726_, new_n45718_ );
nor  ( new_n45812_, new_n45811_, new_n45810_ );
xnor ( new_n45813_, new_n45362_, new_n45358_ );
xnor ( new_n45814_, new_n45813_, new_n45367_ );
xnor ( new_n45815_, new_n45814_, new_n45812_ );
or   ( new_n45816_, new_n45760_, new_n45750_ );
and  ( new_n45817_, new_n45760_, new_n45750_ );
or   ( new_n45818_, new_n45774_, new_n45817_ );
and  ( new_n45819_, new_n45818_, new_n45816_ );
xor  ( new_n45820_, new_n45819_, new_n45815_ );
and  ( new_n45821_, new_n45820_, new_n45809_ );
or   ( new_n45822_, new_n45821_, new_n45808_ );
xor  ( new_n45823_, new_n45557_, new_n45556_ );
xor  ( new_n45824_, new_n45823_, new_n45822_ );
and  ( new_n45825_, new_n45731_, new_n45730_ );
and  ( new_n45826_, new_n45732_, new_n45688_ );
or   ( new_n45827_, new_n45826_, new_n45825_ );
nor  ( new_n45828_, new_n45814_, new_n45812_ );
nor  ( new_n45829_, new_n45819_, new_n45815_ );
or   ( new_n45830_, new_n45829_, new_n45828_ );
xor  ( new_n45831_, new_n45502_, new_n45501_ );
xor  ( new_n45832_, new_n45831_, new_n45830_ );
xor  ( new_n45833_, new_n45832_, new_n45827_ );
xor  ( new_n45834_, new_n45833_, new_n45824_ );
nand ( new_n45835_, new_n45834_, new_n45798_ );
xor  ( new_n45836_, new_n45834_, new_n45798_ );
xor  ( new_n45837_, new_n45820_, new_n45809_ );
xnor ( new_n45838_, new_n45684_, new_n45683_ );
or   ( new_n45839_, new_n45673_, new_n286_ );
xor  ( new_n45840_, new_n45204_, new_n275_ );
or   ( new_n45841_, new_n45840_, new_n283_ );
and  ( new_n45842_, new_n45841_, new_n45839_ );
not  ( new_n45843_, RIbb2e788_32 );
and  ( new_n45844_, new_n2797_, new_n45843_ );
not  ( new_n45845_, new_n45844_ );
and  ( new_n45846_, new_n45845_, new_n2423_ );
xor  ( new_n45847_, new_n43793_, new_n2421_ );
and  ( new_n45848_, new_n45847_, new_n2615_ );
nor  ( new_n45849_, new_n45848_, new_n45846_ );
nor  ( new_n45850_, new_n45849_, new_n45842_ );
and  ( new_n45851_, new_n45720_, new_n295_ );
and  ( new_n45852_, new_n45586_, new_n43949_ );
or   ( new_n45853_, new_n45852_, new_n45851_ );
xor  ( new_n45854_, new_n45849_, new_n45842_ );
and  ( new_n45855_, new_n45854_, new_n45853_ );
nor  ( new_n45856_, new_n45855_, new_n45850_ );
not  ( new_n45857_, new_n45856_ );
xor  ( new_n45858_, new_n45678_, new_n45677_ );
and  ( new_n45859_, new_n45858_, new_n45857_ );
xor  ( new_n45860_, new_n45858_, new_n45857_ );
xor  ( new_n45861_, new_n45658_, new_n45657_ );
and  ( new_n45862_, new_n45861_, new_n45860_ );
or   ( new_n45863_, new_n45862_, new_n45859_ );
xor  ( new_n45864_, new_n45681_, new_n45680_ );
nand ( new_n45865_, new_n45864_, new_n45863_ );
xor  ( new_n45866_, new_n43812_, RIbb2ee90_17 );
and  ( new_n45867_, new_n45866_, new_n822_ );
and  ( new_n45868_, new_n45697_, new_n820_ );
nor  ( new_n45869_, new_n45868_, new_n45867_ );
or   ( new_n45870_, new_n45406_, new_n302_ );
or   ( new_n45871_, new_n45719_, new_n44007_ );
and  ( new_n45872_, new_n45871_, new_n45870_ );
xnor ( new_n45873_, new_n45872_, new_n45869_ );
xor  ( new_n45874_, new_n45738_, new_n43945_ );
nand ( new_n45875_, new_n45874_, new_n43982_ );
nor  ( new_n45876_, new_n45584_, new_n43880_ );
or   ( new_n45877_, new_n45717_, new_n43977_ );
or   ( new_n45878_, new_n45877_, new_n45876_ );
and  ( new_n45879_, new_n45878_, new_n45875_ );
xor  ( new_n45880_, new_n45879_, new_n45873_ );
xor  ( new_n45881_, new_n45611_, new_n45610_ );
and  ( new_n45882_, new_n45881_, new_n45880_ );
xor  ( new_n45883_, new_n45639_, new_n45638_ );
xor  ( new_n45884_, new_n45881_, new_n45880_ );
and  ( new_n45885_, new_n45884_, new_n45883_ );
or   ( new_n45886_, new_n45885_, new_n45882_ );
xor  ( new_n45887_, new_n45864_, new_n45863_ );
nand ( new_n45888_, new_n45887_, new_n45886_ );
and  ( new_n45889_, new_n45888_, new_n45865_ );
nand ( new_n45890_, new_n45889_, new_n45838_ );
or   ( new_n45891_, new_n45889_, new_n45838_ );
xor  ( new_n45892_, new_n45775_, new_n45736_ );
xnor ( new_n45893_, new_n45892_, new_n45793_ );
nand ( new_n45894_, new_n45893_, new_n45891_ );
and  ( new_n45895_, new_n45894_, new_n45890_ );
or   ( new_n45896_, new_n45895_, new_n45837_ );
and  ( new_n45897_, new_n45895_, new_n45837_ );
nor  ( new_n45898_, new_n45872_, new_n45869_ );
nor  ( new_n45899_, new_n45879_, new_n45873_ );
nor  ( new_n45900_, new_n45899_, new_n45898_ );
not  ( new_n45901_, new_n45900_ );
xor  ( new_n45902_, new_n45758_, new_n45757_ );
and  ( new_n45903_, new_n45902_, new_n45901_ );
xor  ( new_n45904_, new_n45902_, new_n45901_ );
xor  ( new_n45905_, new_n45748_, new_n45747_ );
and  ( new_n45906_, new_n45905_, new_n45904_ );
or   ( new_n45907_, new_n45906_, new_n45903_ );
xor  ( new_n45908_, new_n45802_, new_n45800_ );
xor  ( new_n45909_, new_n45908_, new_n45805_ );
nor  ( new_n45910_, new_n45909_, new_n45907_ );
and  ( new_n45911_, new_n45909_, new_n45907_ );
not  ( new_n45912_, new_n45911_ );
not  ( new_n45913_, new_n45582_ );
xor  ( new_n45914_, new_n43787_, new_n2118_ );
or   ( new_n45915_, new_n45914_, new_n2425_ );
nand ( new_n45916_, new_n45580_, new_n2242_ );
and  ( new_n45917_, new_n45916_, new_n45915_ );
or   ( new_n45918_, new_n45917_, new_n2423_ );
nor  ( new_n45919_, new_n45649_, new_n1846_ );
xor  ( new_n45920_, new_n43803_, RIbb2ead0_25 );
and  ( new_n45921_, new_n45920_, new_n1741_ );
or   ( new_n45922_, new_n45921_, new_n45919_ );
xor  ( new_n45923_, new_n45917_, new_n2423_ );
nand ( new_n45924_, new_n45923_, new_n45922_ );
and  ( new_n45925_, new_n45924_, new_n45918_ );
nor  ( new_n45926_, new_n45925_, new_n45913_ );
xor  ( new_n45927_, RIbb32388_158, RIbb2ca78_94 );
xnor ( new_n45928_, new_n45927_, new_n45594_ );
and  ( new_n45929_, new_n45928_, new_n43880_ );
not  ( new_n45930_, new_n45929_ );
xor  ( new_n45931_, new_n45597_, new_n43945_ );
not  ( new_n45932_, new_n45931_ );
or   ( new_n45933_, new_n45932_, new_n43983_ );
nor  ( new_n45934_, new_n45738_, new_n43880_ );
or   ( new_n45935_, new_n45739_, new_n43977_ );
or   ( new_n45936_, new_n45935_, new_n45934_ );
and  ( new_n45937_, new_n45936_, new_n45933_ );
nor  ( new_n45938_, new_n45937_, new_n45930_ );
and  ( new_n45939_, new_n45866_, new_n820_ );
xor  ( new_n45940_, new_n43914_, RIbb2ee90_17 );
and  ( new_n45941_, new_n45940_, new_n822_ );
or   ( new_n45942_, new_n45941_, new_n45939_ );
xor  ( new_n45943_, new_n45937_, new_n45930_ );
and  ( new_n45944_, new_n45943_, new_n45942_ );
or   ( new_n45945_, new_n45944_, new_n45938_ );
xor  ( new_n45946_, new_n45925_, new_n45913_ );
and  ( new_n45947_, new_n45946_, new_n45945_ );
or   ( new_n45948_, new_n45947_, new_n45926_ );
xor  ( new_n45949_, new_n45614_, new_n45613_ );
and  ( new_n45950_, new_n45949_, new_n45948_ );
nand ( new_n45951_, new_n45608_, new_n1474_ );
xor  ( new_n45952_, new_n43888_, RIbb2ebc0_23 );
nand ( new_n45953_, new_n45952_, new_n1476_ );
and  ( new_n45954_, new_n45953_, new_n45951_ );
xor  ( new_n45955_, new_n44218_, RIbb2ef80_15 );
nand ( new_n45956_, new_n45955_, new_n662_ );
nand ( new_n45957_, new_n45634_, new_n660_ );
and  ( new_n45958_, new_n45957_, new_n45956_ );
or   ( new_n45959_, new_n45958_, new_n45954_ );
and  ( new_n45960_, new_n45628_, new_n454_ );
xor  ( new_n45961_, new_n44407_, RIbb2f070_13 );
and  ( new_n45962_, new_n45961_, new_n456_ );
or   ( new_n45963_, new_n45962_, new_n45960_ );
xor  ( new_n45964_, new_n45958_, new_n45954_ );
nand ( new_n45965_, new_n45964_, new_n45963_ );
and  ( new_n45966_, new_n45965_, new_n45959_ );
or   ( new_n45967_, new_n45667_, new_n320_ );
xor  ( new_n45968_, new_n44974_, new_n309_ );
or   ( new_n45969_, new_n45968_, new_n317_ );
and  ( new_n45970_, new_n45969_, new_n45967_ );
nand ( new_n45971_, new_n45653_, new_n334_ );
xor  ( new_n45972_, new_n44785_, new_n329_ );
or   ( new_n45973_, new_n45972_, new_n337_ );
and  ( new_n45974_, new_n45973_, new_n45971_ );
or   ( new_n45975_, new_n45974_, new_n45970_ );
nor  ( new_n45976_, new_n45662_, new_n1137_ );
xor  ( new_n45977_, new_n43985_, RIbb2eda0_19 );
and  ( new_n45978_, new_n45977_, new_n1042_ );
nor  ( new_n45979_, new_n45978_, new_n45976_ );
and  ( new_n45980_, new_n45974_, new_n45970_ );
or   ( new_n45981_, new_n45980_, new_n45979_ );
and  ( new_n45982_, new_n45981_, new_n45975_ );
nor  ( new_n45983_, new_n45982_, new_n45966_ );
xor  ( new_n45984_, new_n43894_, RIbb2e9e0_27 );
nand ( new_n45985_, new_n45984_, new_n2002_ );
or   ( new_n45986_, new_n45602_, new_n2124_ );
and  ( new_n45987_, new_n45986_, new_n45985_ );
or   ( new_n45988_, new_n45625_, new_n1366_ );
xor  ( new_n45989_, new_n43956_, new_n1126_ );
or   ( new_n45990_, new_n45989_, new_n1364_ );
and  ( new_n45991_, new_n45990_, new_n45988_ );
nor  ( new_n45992_, new_n45991_, new_n45987_ );
and  ( new_n45993_, new_n45644_, new_n371_ );
xor  ( new_n45994_, new_n44600_, RIbb2f160_11 );
and  ( new_n45995_, new_n45994_, new_n373_ );
or   ( new_n45996_, new_n45995_, new_n45993_ );
xor  ( new_n45997_, new_n45991_, new_n45987_ );
and  ( new_n45998_, new_n45997_, new_n45996_ );
nor  ( new_n45999_, new_n45998_, new_n45992_ );
not  ( new_n46000_, new_n45999_ );
xor  ( new_n46001_, new_n45982_, new_n45966_ );
and  ( new_n46002_, new_n46001_, new_n46000_ );
or   ( new_n46003_, new_n46002_, new_n45983_ );
xor  ( new_n46004_, new_n45949_, new_n45948_ );
and  ( new_n46005_, new_n46004_, new_n46003_ );
nor  ( new_n46006_, new_n46005_, new_n45950_ );
and  ( new_n46007_, new_n46006_, new_n45912_ );
nor  ( new_n46008_, new_n46007_, new_n45910_ );
or   ( new_n46009_, new_n46008_, new_n45897_ );
and  ( new_n46010_, new_n46009_, new_n45896_ );
nand ( new_n46011_, new_n46010_, new_n45836_ );
and  ( new_n46012_, new_n46011_, new_n45835_ );
xor  ( new_n46013_, new_n45564_, new_n45563_ );
nand ( new_n46014_, new_n45831_, new_n45830_ );
nand ( new_n46015_, new_n45832_, new_n45827_ );
and  ( new_n46016_, new_n46015_, new_n46014_ );
nand ( new_n46017_, new_n45823_, new_n45822_ );
nand ( new_n46018_, new_n45833_, new_n45824_ );
and  ( new_n46019_, new_n46018_, new_n46017_ );
xor  ( new_n46020_, new_n46019_, new_n46016_ );
xnor ( new_n46021_, new_n46020_, new_n46013_ );
and  ( new_n46022_, new_n46021_, new_n46012_ );
or   ( new_n46023_, new_n46019_, new_n46016_ );
nand ( new_n46024_, new_n46020_, new_n46013_ );
and  ( new_n46025_, new_n46024_, new_n46023_ );
xnor ( new_n46026_, new_n45570_, new_n45569_ );
and  ( new_n46027_, new_n46026_, new_n46025_ );
or   ( new_n46028_, new_n46027_, new_n46022_ );
or   ( new_n46029_, new_n46028_, new_n45576_ );
or   ( new_n46030_, new_n46029_, new_n45396_ );
xor  ( new_n46031_, new_n45905_, new_n45904_ );
xor  ( new_n46032_, new_n45783_, new_n45778_ );
xor  ( new_n46033_, new_n46032_, new_n45791_ );
xor  ( new_n46034_, new_n46033_, new_n46031_ );
nor  ( new_n46035_, new_n43700_, new_n43683_ );
xor  ( new_n46036_, RIbb32400_159, RIbb2ca00_95 );
xnor ( new_n46037_, new_n46036_, new_n46035_ );
and  ( new_n46038_, new_n46037_, new_n43880_ );
not  ( new_n46039_, new_n46038_ );
nand ( new_n46040_, new_n45920_, new_n1739_ );
xor  ( new_n46041_, new_n43884_, new_n1583_ );
or   ( new_n46042_, new_n46041_, new_n1844_ );
and  ( new_n46043_, new_n46042_, new_n46040_ );
or   ( new_n46044_, new_n46043_, new_n46039_ );
and  ( new_n46045_, new_n45955_, new_n660_ );
xor  ( new_n46046_, new_n44319_, RIbb2ef80_15 );
and  ( new_n46047_, new_n46046_, new_n662_ );
or   ( new_n46048_, new_n46047_, new_n46045_ );
xor  ( new_n46049_, new_n46043_, new_n46039_ );
nand ( new_n46050_, new_n46049_, new_n46048_ );
and  ( new_n46051_, new_n46050_, new_n46044_ );
or   ( new_n46052_, new_n45840_, new_n286_ );
xor  ( new_n46053_, new_n45403_, new_n275_ );
or   ( new_n46054_, new_n46053_, new_n283_ );
and  ( new_n46055_, new_n46054_, new_n46052_ );
xor  ( new_n46056_, new_n45119_, new_n309_ );
or   ( new_n46057_, new_n46056_, new_n317_ );
or   ( new_n46058_, new_n45968_, new_n320_ );
and  ( new_n46059_, new_n46058_, new_n46057_ );
or   ( new_n46060_, new_n46059_, new_n46055_ );
and  ( new_n46061_, new_n45977_, new_n1040_ );
xor  ( new_n46062_, new_n43812_, RIbb2eda0_19 );
and  ( new_n46063_, new_n46062_, new_n1042_ );
nor  ( new_n46064_, new_n46063_, new_n46061_ );
and  ( new_n46065_, new_n46059_, new_n46055_ );
or   ( new_n46066_, new_n46065_, new_n46064_ );
and  ( new_n46067_, new_n46066_, new_n46060_ );
nor  ( new_n46068_, new_n46067_, new_n46051_ );
xor  ( new_n46069_, new_n43898_, new_n2118_ );
or   ( new_n46070_, new_n46069_, new_n2425_ );
or   ( new_n46071_, new_n45914_, new_n2427_ );
and  ( new_n46072_, new_n46071_, new_n46070_ );
xor  ( new_n46073_, new_n45928_, new_n43945_ );
not  ( new_n46074_, new_n46073_ );
or   ( new_n46075_, new_n46074_, new_n43983_ );
not  ( new_n46076_, new_n45597_ );
and  ( new_n46077_, new_n46076_, new_n43879_ );
or   ( new_n46078_, new_n45598_, new_n43977_ );
or   ( new_n46079_, new_n46078_, new_n46077_ );
and  ( new_n46080_, new_n46079_, new_n46075_ );
nor  ( new_n46081_, new_n46080_, new_n46072_ );
xor  ( new_n46082_, new_n44183_, RIbb2ee90_17 );
and  ( new_n46083_, new_n46082_, new_n822_ );
and  ( new_n46084_, new_n45940_, new_n820_ );
or   ( new_n46085_, new_n46084_, new_n46083_ );
xor  ( new_n46086_, new_n46080_, new_n46072_ );
and  ( new_n46087_, new_n46086_, new_n46085_ );
or   ( new_n46088_, new_n46087_, new_n46081_ );
xor  ( new_n46089_, new_n46067_, new_n46051_ );
and  ( new_n46090_, new_n46089_, new_n46088_ );
or   ( new_n46091_, new_n46090_, new_n46068_ );
xor  ( new_n46092_, new_n45946_, new_n45945_ );
nand ( new_n46093_, new_n46092_, new_n46091_ );
or   ( new_n46094_, new_n46092_, new_n46091_ );
xor  ( new_n46095_, new_n46001_, new_n46000_ );
nand ( new_n46096_, new_n46095_, new_n46094_ );
nand ( new_n46097_, new_n46096_, new_n46093_ );
xnor ( new_n46098_, new_n46097_, new_n46034_ );
xnor ( new_n46099_, new_n45861_, new_n45860_ );
xor  ( new_n46100_, new_n45997_, new_n45996_ );
xnor ( new_n46101_, new_n45974_, new_n45970_ );
xor  ( new_n46102_, new_n46101_, new_n45979_ );
nand ( new_n46103_, new_n46102_, new_n46100_ );
nor  ( new_n46104_, new_n46102_, new_n46100_ );
not  ( new_n46105_, new_n45849_ );
or   ( new_n46106_, new_n45585_, new_n302_ );
or   ( new_n46107_, new_n45874_, new_n44007_ );
and  ( new_n46108_, new_n46107_, new_n46106_ );
nor  ( new_n46109_, new_n46108_, new_n46105_ );
and  ( new_n46110_, new_n46108_, new_n46105_ );
xor  ( new_n46111_, new_n44681_, RIbb2f160_11 );
and  ( new_n46112_, new_n46111_, new_n371_ );
xor  ( new_n46113_, new_n44785_, RIbb2f160_11 );
and  ( new_n46114_, new_n46113_, new_n373_ );
nor  ( new_n46115_, new_n46114_, new_n46112_ );
xor  ( new_n46116_, new_n44877_, new_n329_ );
or   ( new_n46117_, new_n46116_, new_n340_ );
xor  ( new_n46118_, new_n44974_, RIbb2f250_9 );
nand ( new_n46119_, new_n46118_, new_n336_ );
and  ( new_n46120_, new_n46119_, new_n46117_ );
nor  ( new_n46121_, new_n46120_, new_n46115_ );
xor  ( new_n46122_, new_n43937_, RIbb2ebc0_23 );
and  ( new_n46123_, new_n46122_, new_n1474_ );
xor  ( new_n46124_, new_n43956_, new_n1355_ );
nor  ( new_n46125_, new_n46124_, new_n1593_ );
nor  ( new_n46126_, new_n46125_, new_n46123_ );
and  ( new_n46127_, new_n46120_, new_n46115_ );
nor  ( new_n46128_, new_n46127_, new_n46126_ );
nor  ( new_n46129_, new_n46128_, new_n46121_ );
nor  ( new_n46130_, new_n46129_, new_n46110_ );
nor  ( new_n46131_, new_n46130_, new_n46109_ );
or   ( new_n46132_, new_n46131_, new_n46104_ );
and  ( new_n46133_, new_n46132_, new_n46103_ );
or   ( new_n46134_, new_n46133_, new_n46099_ );
and  ( new_n46135_, new_n46133_, new_n46099_ );
xor  ( new_n46136_, RIbb32478_160, RIbb2c988_96 );
xnor ( new_n46137_, new_n46136_, new_n43682_ );
and  ( new_n46138_, new_n46137_, new_n43880_ );
nand ( new_n46139_, new_n46138_, new_n2800_ );
xor  ( new_n46140_, new_n43787_, RIbb2e800_31 );
and  ( new_n46141_, new_n46140_, new_n2615_ );
and  ( new_n46142_, new_n45847_, new_n2613_ );
nor  ( new_n46143_, new_n46142_, new_n46141_ );
not  ( new_n46144_, new_n46143_ );
xor  ( new_n46145_, new_n46138_, new_n2800_ );
nand ( new_n46146_, new_n46145_, new_n46144_ );
and  ( new_n46147_, new_n46146_, new_n46139_ );
xor  ( new_n46148_, new_n43888_, new_n1583_ );
or   ( new_n46149_, new_n46148_, new_n1844_ );
or   ( new_n46150_, new_n46041_, new_n1846_ );
and  ( new_n46151_, new_n46150_, new_n46149_ );
xor  ( new_n46152_, new_n43799_, new_n1840_ );
or   ( new_n46153_, new_n46152_, new_n2124_ );
xor  ( new_n46154_, new_n43803_, RIbb2e9e0_27 );
nand ( new_n46155_, new_n46154_, new_n2002_ );
and  ( new_n46156_, new_n46155_, new_n46153_ );
or   ( new_n46157_, new_n46156_, new_n46151_ );
xor  ( new_n46158_, new_n44218_, RIbb2ee90_17 );
and  ( new_n46159_, new_n46158_, new_n822_ );
and  ( new_n46160_, new_n46082_, new_n820_ );
or   ( new_n46161_, new_n46160_, new_n46159_ );
xor  ( new_n46162_, new_n46156_, new_n46151_ );
nand ( new_n46163_, new_n46162_, new_n46161_ );
and  ( new_n46164_, new_n46163_, new_n46157_ );
nor  ( new_n46165_, new_n46164_, new_n46147_ );
xor  ( new_n46166_, new_n43914_, RIbb2eda0_19 );
and  ( new_n46167_, new_n46166_, new_n1042_ );
and  ( new_n46168_, new_n46062_, new_n1040_ );
nor  ( new_n46169_, new_n46168_, new_n46167_ );
or   ( new_n46170_, new_n45874_, new_n302_ );
or   ( new_n46171_, new_n45931_, new_n44007_ );
and  ( new_n46172_, new_n46171_, new_n46170_ );
nor  ( new_n46173_, new_n46172_, new_n46169_ );
xnor ( new_n46174_, new_n46172_, new_n46169_ );
xor  ( new_n46175_, new_n46037_, new_n43945_ );
nand ( new_n46176_, new_n46175_, new_n43982_ );
nor  ( new_n46177_, new_n45928_, new_n43880_ );
or   ( new_n46178_, new_n45929_, new_n43977_ );
or   ( new_n46179_, new_n46178_, new_n46177_ );
and  ( new_n46180_, new_n46179_, new_n46176_ );
nor  ( new_n46181_, new_n46180_, new_n46174_ );
nor  ( new_n46182_, new_n46181_, new_n46173_ );
xnor ( new_n46183_, new_n46164_, new_n46147_ );
nor  ( new_n46184_, new_n46183_, new_n46182_ );
or   ( new_n46185_, new_n46184_, new_n46165_ );
xor  ( new_n46186_, new_n46089_, new_n46088_ );
nor  ( new_n46187_, new_n46186_, new_n46185_ );
nand ( new_n46188_, new_n46111_, new_n373_ );
nand ( new_n46189_, new_n45994_, new_n371_ );
and  ( new_n46190_, new_n46189_, new_n46188_ );
nand ( new_n46191_, new_n45961_, new_n454_ );
xor  ( new_n46192_, new_n44506_, new_n400_ );
or   ( new_n46193_, new_n46192_, new_n524_ );
and  ( new_n46194_, new_n46193_, new_n46191_ );
nor  ( new_n46195_, new_n46194_, new_n46190_ );
and  ( new_n46196_, new_n46122_, new_n1476_ );
and  ( new_n46197_, new_n45952_, new_n1474_ );
or   ( new_n46198_, new_n46197_, new_n46196_ );
xor  ( new_n46199_, new_n46194_, new_n46190_ );
and  ( new_n46200_, new_n46199_, new_n46198_ );
nor  ( new_n46201_, new_n46200_, new_n46195_ );
or   ( new_n46202_, new_n46116_, new_n337_ );
or   ( new_n46203_, new_n45972_, new_n340_ );
and  ( new_n46204_, new_n46203_, new_n46202_ );
or   ( new_n46205_, new_n45989_, new_n1366_ );
xor  ( new_n46206_, new_n43952_, new_n1126_ );
or   ( new_n46207_, new_n46206_, new_n1364_ );
and  ( new_n46208_, new_n46207_, new_n46205_ );
or   ( new_n46209_, new_n46208_, new_n46204_ );
and  ( new_n46210_, new_n45984_, new_n2000_ );
nor  ( new_n46211_, new_n46152_, new_n2122_ );
nor  ( new_n46212_, new_n46211_, new_n46210_ );
and  ( new_n46213_, new_n46208_, new_n46204_ );
or   ( new_n46214_, new_n46213_, new_n46212_ );
and  ( new_n46215_, new_n46214_, new_n46209_ );
xor  ( new_n46216_, new_n46215_, new_n46201_ );
xor  ( new_n46217_, new_n45943_, new_n45942_ );
xor  ( new_n46218_, new_n46217_, new_n46216_ );
not  ( new_n46219_, new_n46218_ );
nand ( new_n46220_, new_n46186_, new_n46185_ );
and  ( new_n46221_, new_n46220_, new_n46219_ );
or   ( new_n46222_, new_n46221_, new_n46187_ );
or   ( new_n46223_, new_n46222_, new_n46135_ );
and  ( new_n46224_, new_n46223_, new_n46134_ );
nor  ( new_n46225_, new_n46224_, new_n46098_ );
xor  ( new_n46226_, new_n46224_, new_n46098_ );
nor  ( new_n46227_, new_n46215_, new_n46201_ );
and  ( new_n46228_, new_n46217_, new_n46216_ );
nor  ( new_n46229_, new_n46228_, new_n46227_ );
xor  ( new_n46230_, new_n45923_, new_n45922_ );
xor  ( new_n46231_, new_n45854_, new_n45853_ );
nand ( new_n46232_, new_n46231_, new_n46230_ );
xor  ( new_n46233_, new_n46231_, new_n46230_ );
xor  ( new_n46234_, new_n45964_, new_n45963_ );
nand ( new_n46235_, new_n46234_, new_n46233_ );
and  ( new_n46236_, new_n46235_, new_n46232_ );
xor  ( new_n46237_, new_n46236_, new_n46229_ );
xor  ( new_n46238_, new_n45884_, new_n45883_ );
xnor ( new_n46239_, new_n46238_, new_n46237_ );
xor  ( new_n46240_, new_n45584_, new_n275_ );
or   ( new_n46241_, new_n46240_, new_n283_ );
or   ( new_n46242_, new_n46053_, new_n286_ );
and  ( new_n46243_, new_n46242_, new_n46241_ );
or   ( new_n46244_, new_n46206_, new_n1366_ );
xor  ( new_n46245_, new_n43985_, new_n1126_ );
or   ( new_n46246_, new_n46245_, new_n1364_ );
and  ( new_n46247_, new_n46246_, new_n46244_ );
or   ( new_n46248_, new_n46247_, new_n46243_ );
nor  ( new_n46249_, new_n46056_, new_n320_ );
xor  ( new_n46250_, new_n45204_, RIbb2f340_7 );
and  ( new_n46251_, new_n46250_, new_n316_ );
or   ( new_n46252_, new_n46251_, new_n46249_ );
xor  ( new_n46253_, new_n46247_, new_n46243_ );
nand ( new_n46254_, new_n46253_, new_n46252_ );
and  ( new_n46255_, new_n46254_, new_n46248_ );
or   ( new_n46256_, new_n46069_, new_n2427_ );
xor  ( new_n46257_, new_n43894_, RIbb2e8f0_29 );
nand ( new_n46258_, new_n46257_, new_n2244_ );
and  ( new_n46259_, new_n46258_, new_n46256_ );
xor  ( new_n46260_, new_n44600_, new_n400_ );
or   ( new_n46261_, new_n46260_, new_n524_ );
or   ( new_n46262_, new_n46192_, new_n526_ );
and  ( new_n46263_, new_n46262_, new_n46261_ );
or   ( new_n46264_, new_n46263_, new_n46259_ );
and  ( new_n46265_, new_n46046_, new_n660_ );
xor  ( new_n46266_, new_n44407_, RIbb2ef80_15 );
and  ( new_n46267_, new_n46266_, new_n662_ );
or   ( new_n46268_, new_n46267_, new_n46265_ );
xor  ( new_n46269_, new_n46263_, new_n46259_ );
nand ( new_n46270_, new_n46269_, new_n46268_ );
and  ( new_n46271_, new_n46270_, new_n46264_ );
nor  ( new_n46272_, new_n46271_, new_n46255_ );
xor  ( new_n46273_, new_n46086_, new_n46085_ );
xor  ( new_n46274_, new_n46271_, new_n46255_ );
and  ( new_n46275_, new_n46274_, new_n46273_ );
or   ( new_n46276_, new_n46275_, new_n46272_ );
xor  ( new_n46277_, new_n46234_, new_n46233_ );
nand ( new_n46278_, new_n46277_, new_n46276_ );
nor  ( new_n46279_, new_n46277_, new_n46276_ );
xor  ( new_n46280_, new_n46199_, new_n46198_ );
xor  ( new_n46281_, new_n46049_, new_n46048_ );
nand ( new_n46282_, new_n46281_, new_n46280_ );
xor  ( new_n46283_, new_n46281_, new_n46280_ );
xnor ( new_n46284_, new_n46059_, new_n46055_ );
xor  ( new_n46285_, new_n46284_, new_n46064_ );
nand ( new_n46286_, new_n46285_, new_n46283_ );
and  ( new_n46287_, new_n46286_, new_n46282_ );
or   ( new_n46288_, new_n46287_, new_n46279_ );
and  ( new_n46289_, new_n46288_, new_n46278_ );
nand ( new_n46290_, new_n46289_, new_n46239_ );
nor  ( new_n46291_, new_n46289_, new_n46239_ );
xor  ( new_n46292_, new_n46092_, new_n46091_ );
xor  ( new_n46293_, new_n46292_, new_n46095_ );
or   ( new_n46294_, new_n46293_, new_n46291_ );
and  ( new_n46295_, new_n46294_, new_n46290_ );
and  ( new_n46296_, new_n46295_, new_n46226_ );
nor  ( new_n46297_, new_n46296_, new_n46225_ );
xor  ( new_n46298_, new_n45889_, new_n45838_ );
xor  ( new_n46299_, new_n46298_, new_n45893_ );
nand ( new_n46300_, new_n46299_, new_n46297_ );
xor  ( new_n46301_, new_n46299_, new_n46297_ );
nor  ( new_n46302_, new_n46236_, new_n46229_ );
and  ( new_n46303_, new_n46238_, new_n46237_ );
nor  ( new_n46304_, new_n46303_, new_n46302_ );
not  ( new_n46305_, new_n46304_ );
xor  ( new_n46306_, new_n46004_, new_n46003_ );
and  ( new_n46307_, new_n46306_, new_n46305_ );
xor  ( new_n46308_, new_n46306_, new_n46305_ );
xor  ( new_n46309_, new_n45887_, new_n45886_ );
and  ( new_n46310_, new_n46309_, new_n46308_ );
nor  ( new_n46311_, new_n46310_, new_n46307_ );
nand ( new_n46312_, new_n46033_, new_n46031_ );
nand ( new_n46313_, new_n46097_, new_n46034_ );
and  ( new_n46314_, new_n46313_, new_n46312_ );
xor  ( new_n46315_, new_n45909_, new_n45907_ );
xor  ( new_n46316_, new_n46315_, new_n46006_ );
xnor ( new_n46317_, new_n46316_, new_n46314_ );
xnor ( new_n46318_, new_n46317_, new_n46311_ );
nand ( new_n46319_, new_n46318_, new_n46301_ );
and  ( new_n46320_, new_n46319_, new_n46300_ );
xor  ( new_n46321_, new_n45795_, new_n45735_ );
xnor ( new_n46322_, new_n45895_, new_n45837_ );
xor  ( new_n46323_, new_n46322_, new_n46008_ );
xor  ( new_n46324_, new_n46323_, new_n46321_ );
or   ( new_n46325_, new_n46316_, new_n46314_ );
and  ( new_n46326_, new_n46316_, new_n46314_ );
or   ( new_n46327_, new_n46326_, new_n46311_ );
and  ( new_n46328_, new_n46327_, new_n46325_ );
xor  ( new_n46329_, new_n46328_, new_n46324_ );
or   ( new_n46330_, new_n46329_, new_n46320_ );
xnor ( new_n46331_, new_n46010_, new_n45836_ );
not  ( new_n46332_, new_n46321_ );
or   ( new_n46333_, new_n46323_, new_n46332_ );
and  ( new_n46334_, new_n46323_, new_n46332_ );
or   ( new_n46335_, new_n46328_, new_n46334_ );
and  ( new_n46336_, new_n46335_, new_n46333_ );
nand ( new_n46337_, new_n46336_, new_n46331_ );
and  ( new_n46338_, new_n46337_, new_n46330_ );
xor  ( new_n46339_, new_n46309_, new_n46308_ );
xor  ( new_n46340_, new_n46295_, new_n46226_ );
and  ( new_n46341_, new_n46340_, new_n46339_ );
xnor ( new_n46342_, new_n46340_, new_n46339_ );
xor  ( new_n46343_, new_n46133_, new_n46099_ );
xor  ( new_n46344_, new_n46343_, new_n46222_ );
xnor ( new_n46345_, new_n46208_, new_n46204_ );
xor  ( new_n46346_, new_n46345_, new_n46212_ );
xor  ( new_n46347_, new_n46108_, new_n45849_ );
xor  ( new_n46348_, new_n46347_, new_n46129_ );
and  ( new_n46349_, new_n46348_, new_n46346_ );
nor  ( new_n46350_, new_n46348_, new_n46346_ );
xor  ( new_n46351_, new_n46145_, new_n46144_ );
not  ( new_n46352_, new_n46351_ );
not  ( new_n46353_, RIbb2e698_34 );
and  ( new_n46354_, new_n3113_, new_n46353_ );
not  ( new_n46355_, new_n46354_ );
and  ( new_n46356_, new_n46355_, new_n2799_ );
xor  ( new_n46357_, new_n43793_, new_n2797_ );
and  ( new_n46358_, new_n46357_, new_n2930_ );
nor  ( new_n46359_, new_n46358_, new_n46356_ );
nor  ( new_n46360_, new_n46359_, new_n46352_ );
xor  ( new_n46361_, new_n46359_, new_n46351_ );
xor  ( new_n46362_, new_n44681_, new_n400_ );
or   ( new_n46363_, new_n46362_, new_n524_ );
or   ( new_n46364_, new_n46260_, new_n526_ );
and  ( new_n46365_, new_n46364_, new_n46363_ );
xor  ( new_n46366_, new_n43952_, new_n1355_ );
or   ( new_n46367_, new_n46366_, new_n1593_ );
or   ( new_n46368_, new_n46124_, new_n1595_ );
and  ( new_n46369_, new_n46368_, new_n46367_ );
nor  ( new_n46370_, new_n46369_, new_n46365_ );
and  ( new_n46371_, new_n46257_, new_n2242_ );
xor  ( new_n46372_, new_n43799_, new_n2118_ );
nor  ( new_n46373_, new_n46372_, new_n2425_ );
nor  ( new_n46374_, new_n46373_, new_n46371_ );
and  ( new_n46375_, new_n46369_, new_n46365_ );
nor  ( new_n46376_, new_n46375_, new_n46374_ );
nor  ( new_n46377_, new_n46376_, new_n46370_ );
nor  ( new_n46378_, new_n46377_, new_n46361_ );
nor  ( new_n46379_, new_n46378_, new_n46360_ );
nor  ( new_n46380_, new_n46379_, new_n46350_ );
or   ( new_n46381_, new_n46380_, new_n46349_ );
xnor ( new_n46382_, new_n46102_, new_n46100_ );
xor  ( new_n46383_, new_n46382_, new_n46131_ );
nand ( new_n46384_, new_n46383_, new_n46381_ );
nor  ( new_n46385_, new_n46383_, new_n46381_ );
xnor ( new_n46386_, new_n46183_, new_n46182_ );
nand ( new_n46387_, new_n46140_, new_n2613_ );
xor  ( new_n46388_, new_n43898_, new_n2421_ );
or   ( new_n46389_, new_n46388_, new_n2807_ );
and  ( new_n46390_, new_n46389_, new_n46387_ );
xor  ( new_n46391_, new_n46137_, new_n43945_ );
not  ( new_n46392_, new_n46391_ );
or   ( new_n46393_, new_n46392_, new_n43983_ );
nor  ( new_n46394_, new_n46037_, new_n43880_ );
or   ( new_n46395_, new_n46038_, new_n43977_ );
or   ( new_n46396_, new_n46395_, new_n46394_ );
and  ( new_n46397_, new_n46396_, new_n46393_ );
nor  ( new_n46398_, new_n46397_, new_n46390_ );
and  ( new_n46399_, new_n46158_, new_n820_ );
xor  ( new_n46400_, new_n44319_, RIbb2ee90_17 );
and  ( new_n46401_, new_n46400_, new_n822_ );
or   ( new_n46402_, new_n46401_, new_n46399_ );
xor  ( new_n46403_, new_n46397_, new_n46390_ );
and  ( new_n46404_, new_n46403_, new_n46402_ );
nor  ( new_n46405_, new_n46404_, new_n46398_ );
not  ( new_n46406_, new_n46405_ );
xor  ( new_n46407_, RIbb324f0_161, RIbb2c910_97 );
nor  ( new_n46408_, new_n43634_, new_n43548_ );
not  ( new_n46409_, new_n46408_ );
and  ( new_n46410_, new_n46409_, new_n43557_ );
nor  ( new_n46411_, new_n46410_, new_n43607_ );
not  ( new_n46412_, new_n46411_ );
and  ( new_n46413_, new_n46412_, new_n43568_ );
nor  ( new_n46414_, new_n46413_, new_n43651_ );
not  ( new_n46415_, new_n46414_ );
and  ( new_n46416_, new_n46415_, new_n43590_ );
nor  ( new_n46417_, new_n46416_, new_n43664_ );
not  ( new_n46418_, new_n46417_ );
and  ( new_n46419_, new_n46418_, new_n43572_ );
nor  ( new_n46420_, new_n46419_, new_n43671_ );
not  ( new_n46421_, new_n46420_ );
and  ( new_n46422_, new_n46421_, new_n43575_ );
nor  ( new_n46423_, new_n46422_, new_n43670_ );
not  ( new_n46424_, new_n46423_ );
and  ( new_n46425_, new_n46424_, new_n43570_ );
nor  ( new_n46426_, new_n46425_, new_n43669_ );
xnor ( new_n46427_, new_n46426_, new_n46407_ );
and  ( new_n46428_, new_n46427_, new_n43880_ );
not  ( new_n46429_, new_n46428_ );
xor  ( new_n46430_, new_n44183_, RIbb2eda0_19 );
nand ( new_n46431_, new_n46430_, new_n1042_ );
nand ( new_n46432_, new_n46166_, new_n1040_ );
and  ( new_n46433_, new_n46432_, new_n46431_ );
nor  ( new_n46434_, new_n46433_, new_n46429_ );
and  ( new_n46435_, new_n45932_, new_n295_ );
and  ( new_n46436_, new_n46074_, new_n43949_ );
or   ( new_n46437_, new_n46436_, new_n46435_ );
xor  ( new_n46438_, new_n46433_, new_n46429_ );
and  ( new_n46439_, new_n46438_, new_n46437_ );
nor  ( new_n46440_, new_n46439_, new_n46434_ );
not  ( new_n46441_, new_n46440_ );
and  ( new_n46442_, new_n46441_, new_n46406_ );
and  ( new_n46443_, new_n46440_, new_n46405_ );
nand ( new_n46444_, new_n46266_, new_n660_ );
xor  ( new_n46445_, new_n44506_, new_n520_ );
or   ( new_n46446_, new_n46445_, new_n755_ );
and  ( new_n46447_, new_n46446_, new_n46444_ );
or   ( new_n46448_, new_n46148_, new_n1846_ );
xor  ( new_n46449_, new_n43937_, RIbb2ead0_25 );
nand ( new_n46450_, new_n46449_, new_n1741_ );
and  ( new_n46451_, new_n46450_, new_n46448_ );
nor  ( new_n46452_, new_n46451_, new_n46447_ );
xor  ( new_n46453_, new_n43884_, RIbb2e9e0_27 );
and  ( new_n46454_, new_n46453_, new_n2002_ );
and  ( new_n46455_, new_n46154_, new_n2000_ );
nor  ( new_n46456_, new_n46455_, new_n46454_ );
and  ( new_n46457_, new_n46451_, new_n46447_ );
nor  ( new_n46458_, new_n46457_, new_n46456_ );
nor  ( new_n46459_, new_n46458_, new_n46452_ );
nor  ( new_n46460_, new_n46459_, new_n46443_ );
nor  ( new_n46461_, new_n46460_, new_n46442_ );
nor  ( new_n46462_, new_n46461_, new_n46386_ );
xor  ( new_n46463_, new_n46461_, new_n46386_ );
xor  ( new_n46464_, new_n46274_, new_n46273_ );
and  ( new_n46465_, new_n46464_, new_n46463_ );
nor  ( new_n46466_, new_n46465_, new_n46462_ );
or   ( new_n46467_, new_n46466_, new_n46385_ );
and  ( new_n46468_, new_n46467_, new_n46384_ );
or   ( new_n46469_, new_n46468_, new_n46344_ );
and  ( new_n46470_, new_n46468_, new_n46344_ );
or   ( new_n46471_, new_n46240_, new_n286_ );
xor  ( new_n46472_, new_n45738_, new_n275_ );
or   ( new_n46473_, new_n46472_, new_n283_ );
nand ( new_n46474_, new_n46473_, new_n46471_ );
and  ( new_n46475_, new_n46474_, new_n46359_ );
and  ( new_n46476_, new_n46250_, new_n314_ );
xor  ( new_n46477_, new_n45403_, new_n309_ );
nor  ( new_n46478_, new_n46477_, new_n317_ );
nor  ( new_n46479_, new_n46478_, new_n46476_ );
not  ( new_n46480_, new_n46479_ );
xor  ( new_n46481_, new_n46474_, new_n46359_ );
and  ( new_n46482_, new_n46481_, new_n46480_ );
or   ( new_n46483_, new_n46482_, new_n46475_ );
xor  ( new_n46484_, new_n46269_, new_n46268_ );
nand ( new_n46485_, new_n46484_, new_n46483_ );
xor  ( new_n46486_, new_n46253_, new_n46252_ );
xor  ( new_n46487_, new_n46484_, new_n46483_ );
nand ( new_n46488_, new_n46487_, new_n46486_ );
and  ( new_n46489_, new_n46488_, new_n46485_ );
nand ( new_n46490_, new_n46113_, new_n371_ );
xor  ( new_n46491_, new_n44877_, new_n325_ );
or   ( new_n46492_, new_n46491_, new_n409_ );
and  ( new_n46493_, new_n46492_, new_n46490_ );
xor  ( new_n46494_, new_n43812_, RIbb2ecb0_21 );
nand ( new_n46495_, new_n46494_, new_n1253_ );
or   ( new_n46496_, new_n46245_, new_n1366_ );
and  ( new_n46497_, new_n46496_, new_n46495_ );
nor  ( new_n46498_, new_n46497_, new_n46493_ );
and  ( new_n46499_, new_n46118_, new_n334_ );
xor  ( new_n46500_, new_n45119_, new_n329_ );
nor  ( new_n46501_, new_n46500_, new_n337_ );
or   ( new_n46502_, new_n46501_, new_n46499_ );
xor  ( new_n46503_, new_n46497_, new_n46493_ );
and  ( new_n46504_, new_n46503_, new_n46502_ );
or   ( new_n46505_, new_n46504_, new_n46498_ );
xor  ( new_n46506_, new_n46162_, new_n46161_ );
nand ( new_n46507_, new_n46506_, new_n46505_ );
xor  ( new_n46508_, new_n46506_, new_n46505_ );
xor  ( new_n46509_, new_n46180_, new_n46174_ );
nand ( new_n46510_, new_n46509_, new_n46508_ );
and  ( new_n46511_, new_n46510_, new_n46507_ );
or   ( new_n46512_, new_n46511_, new_n46489_ );
xor  ( new_n46513_, new_n46285_, new_n46283_ );
xor  ( new_n46514_, new_n46511_, new_n46489_ );
nand ( new_n46515_, new_n46514_, new_n46513_ );
and  ( new_n46516_, new_n46515_, new_n46512_ );
xor  ( new_n46517_, new_n46277_, new_n46276_ );
xor  ( new_n46518_, new_n46517_, new_n46287_ );
nor  ( new_n46519_, new_n46518_, new_n46516_ );
and  ( new_n46520_, new_n46518_, new_n46516_ );
xor  ( new_n46521_, new_n46186_, new_n46185_ );
xor  ( new_n46522_, new_n46521_, new_n46219_ );
nor  ( new_n46523_, new_n46522_, new_n46520_ );
nor  ( new_n46524_, new_n46523_, new_n46519_ );
or   ( new_n46525_, new_n46524_, new_n46470_ );
and  ( new_n46526_, new_n46525_, new_n46469_ );
nor  ( new_n46527_, new_n46526_, new_n46342_ );
or   ( new_n46528_, new_n46527_, new_n46341_ );
xnor ( new_n46529_, new_n46318_, new_n46301_ );
or   ( new_n46530_, new_n46529_, new_n46528_ );
xor  ( new_n46531_, new_n46289_, new_n46239_ );
xor  ( new_n46532_, new_n46531_, new_n46293_ );
xnor ( new_n46533_, new_n46468_, new_n46344_ );
xor  ( new_n46534_, new_n46533_, new_n46524_ );
and  ( new_n46535_, new_n46534_, new_n46532_ );
xor  ( new_n46536_, new_n46534_, new_n46532_ );
xor  ( new_n46537_, new_n46464_, new_n46463_ );
xor  ( new_n46538_, new_n46481_, new_n46480_ );
xor  ( new_n46539_, new_n46438_, new_n46437_ );
and  ( new_n46540_, new_n46539_, new_n46538_ );
xor  ( new_n46541_, new_n46539_, new_n46538_ );
xor  ( new_n46542_, new_n46403_, new_n46402_ );
and  ( new_n46543_, new_n46542_, new_n46541_ );
or   ( new_n46544_, new_n46543_, new_n46540_ );
xor  ( new_n46545_, new_n46487_, new_n46486_ );
or   ( new_n46546_, new_n46545_, new_n46544_ );
xor  ( new_n46547_, new_n46509_, new_n46508_ );
and  ( new_n46548_, new_n46545_, new_n46544_ );
or   ( new_n46549_, new_n46548_, new_n46547_ );
and  ( new_n46550_, new_n46549_, new_n46546_ );
and  ( new_n46551_, new_n46550_, new_n46537_ );
xor  ( new_n46552_, new_n46550_, new_n46537_ );
xor  ( new_n46553_, new_n46514_, new_n46513_ );
and  ( new_n46554_, new_n46553_, new_n46552_ );
or   ( new_n46555_, new_n46554_, new_n46551_ );
xnor ( new_n46556_, new_n46383_, new_n46381_ );
xor  ( new_n46557_, new_n46556_, new_n46466_ );
or   ( new_n46558_, new_n46557_, new_n46555_ );
nand ( new_n46559_, new_n46557_, new_n46555_ );
xnor ( new_n46560_, new_n46120_, new_n46115_ );
and  ( new_n46561_, new_n46560_, new_n46126_ );
not  ( new_n46562_, new_n46121_ );
and  ( new_n46563_, new_n46128_, new_n46562_ );
or   ( new_n46564_, new_n46563_, new_n46561_ );
nand ( new_n46565_, new_n46453_, new_n2000_ );
xor  ( new_n46566_, new_n43888_, RIbb2e9e0_27 );
nand ( new_n46567_, new_n46566_, new_n2002_ );
and  ( new_n46568_, new_n46567_, new_n46565_ );
or   ( new_n46569_, new_n46445_, new_n757_ );
xor  ( new_n46570_, new_n44600_, RIbb2ef80_15 );
nand ( new_n46571_, new_n46570_, new_n662_ );
and  ( new_n46572_, new_n46571_, new_n46569_ );
nor  ( new_n46573_, new_n46572_, new_n46568_ );
and  ( new_n46574_, new_n46400_, new_n820_ );
xor  ( new_n46575_, new_n44407_, RIbb2ee90_17 );
and  ( new_n46576_, new_n46575_, new_n822_ );
nor  ( new_n46577_, new_n46576_, new_n46574_ );
and  ( new_n46578_, new_n46572_, new_n46568_ );
nor  ( new_n46579_, new_n46578_, new_n46577_ );
nor  ( new_n46580_, new_n46579_, new_n46573_ );
xor  ( new_n46581_, new_n43894_, new_n2421_ );
or   ( new_n46582_, new_n46581_, new_n2807_ );
or   ( new_n46583_, new_n46388_, new_n2809_ );
and  ( new_n46584_, new_n46583_, new_n46582_ );
or   ( new_n46585_, new_n46362_, new_n526_ );
xor  ( new_n46586_, new_n44785_, new_n400_ );
or   ( new_n46587_, new_n46586_, new_n524_ );
and  ( new_n46588_, new_n46587_, new_n46585_ );
nor  ( new_n46589_, new_n46588_, new_n46584_ );
xor  ( new_n46590_, new_n43956_, new_n1583_ );
nor  ( new_n46591_, new_n46590_, new_n1844_ );
and  ( new_n46592_, new_n46449_, new_n1739_ );
nor  ( new_n46593_, new_n46592_, new_n46591_ );
and  ( new_n46594_, new_n46588_, new_n46584_ );
nor  ( new_n46595_, new_n46594_, new_n46593_ );
nor  ( new_n46596_, new_n46595_, new_n46589_ );
or   ( new_n46597_, new_n46596_, new_n46580_ );
and  ( new_n46598_, new_n46596_, new_n46580_ );
or   ( new_n46599_, new_n46500_, new_n340_ );
xor  ( new_n46600_, new_n45204_, new_n329_ );
or   ( new_n46601_, new_n46600_, new_n337_ );
and  ( new_n46602_, new_n46601_, new_n46599_ );
or   ( new_n46603_, new_n46491_, new_n411_ );
xor  ( new_n46604_, new_n44974_, new_n325_ );
or   ( new_n46605_, new_n46604_, new_n409_ );
and  ( new_n46606_, new_n46605_, new_n46603_ );
nor  ( new_n46607_, new_n46606_, new_n46602_ );
nor  ( new_n46608_, new_n46366_, new_n1595_ );
xor  ( new_n46609_, new_n43985_, RIbb2ebc0_23 );
and  ( new_n46610_, new_n46609_, new_n1476_ );
nor  ( new_n46611_, new_n46610_, new_n46608_ );
and  ( new_n46612_, new_n46606_, new_n46602_ );
nor  ( new_n46613_, new_n46612_, new_n46611_ );
nor  ( new_n46614_, new_n46613_, new_n46607_ );
or   ( new_n46615_, new_n46614_, new_n46598_ );
and  ( new_n46616_, new_n46615_, new_n46597_ );
or   ( new_n46617_, new_n46616_, new_n46564_ );
xor  ( new_n46618_, RIbb32568_162, RIbb2c898_98 );
xor  ( new_n46619_, new_n46618_, new_n46424_ );
and  ( new_n46620_, new_n46619_, new_n43880_ );
nor  ( new_n46621_, new_n46620_, new_n3116_ );
nand ( new_n46622_, new_n46620_, new_n3116_ );
xor  ( new_n46623_, new_n46427_, new_n43945_ );
and  ( new_n46624_, new_n46623_, new_n43982_ );
nor  ( new_n46625_, new_n46137_, new_n43880_ );
not  ( new_n46626_, new_n46625_ );
nor  ( new_n46627_, new_n46138_, new_n43977_ );
and  ( new_n46628_, new_n46627_, new_n46626_ );
nor  ( new_n46629_, new_n46628_, new_n46624_ );
and  ( new_n46630_, new_n46629_, new_n46622_ );
or   ( new_n46631_, new_n46630_, new_n46621_ );
or   ( new_n46632_, new_n46472_, new_n286_ );
xor  ( new_n46633_, new_n45597_, new_n275_ );
or   ( new_n46634_, new_n46633_, new_n283_ );
and  ( new_n46635_, new_n46634_, new_n46632_ );
or   ( new_n46636_, new_n46175_, new_n44007_ );
or   ( new_n46637_, new_n46073_, new_n302_ );
and  ( new_n46638_, new_n46637_, new_n46636_ );
or   ( new_n46639_, new_n46638_, new_n46635_ );
xor  ( new_n46640_, new_n43914_, RIbb2ecb0_21 );
and  ( new_n46641_, new_n46640_, new_n1253_ );
and  ( new_n46642_, new_n46494_, new_n1251_ );
nor  ( new_n46643_, new_n46642_, new_n46641_ );
and  ( new_n46644_, new_n46638_, new_n46635_ );
or   ( new_n46645_, new_n46644_, new_n46643_ );
and  ( new_n46646_, new_n46645_, new_n46639_ );
nor  ( new_n46647_, new_n46646_, new_n46631_ );
xor  ( new_n46648_, new_n43787_, RIbb2e710_33 );
nand ( new_n46649_, new_n46648_, new_n2930_ );
nand ( new_n46650_, new_n46357_, new_n2928_ );
and  ( new_n46651_, new_n46650_, new_n46649_ );
or   ( new_n46652_, new_n46372_, new_n2427_ );
xor  ( new_n46653_, new_n43803_, new_n2118_ );
or   ( new_n46654_, new_n46653_, new_n2425_ );
and  ( new_n46655_, new_n46654_, new_n46652_ );
nor  ( new_n46656_, new_n46655_, new_n46651_ );
and  ( new_n46657_, new_n46430_, new_n1040_ );
xor  ( new_n46658_, new_n44218_, RIbb2eda0_19 );
and  ( new_n46659_, new_n46658_, new_n1042_ );
nor  ( new_n46660_, new_n46659_, new_n46657_ );
not  ( new_n46661_, new_n46660_ );
xor  ( new_n46662_, new_n46655_, new_n46651_ );
and  ( new_n46663_, new_n46662_, new_n46661_ );
or   ( new_n46664_, new_n46663_, new_n46656_ );
xor  ( new_n46665_, new_n46646_, new_n46631_ );
and  ( new_n46666_, new_n46665_, new_n46664_ );
or   ( new_n46667_, new_n46666_, new_n46647_ );
xor  ( new_n46668_, new_n46616_, new_n46564_ );
nand ( new_n46669_, new_n46668_, new_n46667_ );
and  ( new_n46670_, new_n46669_, new_n46617_ );
xor  ( new_n46671_, new_n46348_, new_n46346_ );
xor  ( new_n46672_, new_n46671_, new_n46379_ );
nor  ( new_n46673_, new_n46672_, new_n46670_ );
xor  ( new_n46674_, new_n46377_, new_n46361_ );
xnor ( new_n46675_, new_n46451_, new_n46447_ );
nand ( new_n46676_, new_n46675_, new_n46456_ );
not  ( new_n46677_, new_n46458_ );
or   ( new_n46678_, new_n46677_, new_n46452_ );
and  ( new_n46679_, new_n46678_, new_n46676_ );
xor  ( new_n46680_, new_n46503_, new_n46502_ );
or   ( new_n46681_, new_n46680_, new_n46679_ );
xnor ( new_n46682_, new_n46369_, new_n46365_ );
nand ( new_n46683_, new_n46682_, new_n46374_ );
not  ( new_n46684_, new_n46376_ );
or   ( new_n46685_, new_n46684_, new_n46370_ );
and  ( new_n46686_, new_n46685_, new_n46683_ );
and  ( new_n46687_, new_n46680_, new_n46679_ );
or   ( new_n46688_, new_n46687_, new_n46686_ );
and  ( new_n46689_, new_n46688_, new_n46681_ );
and  ( new_n46690_, new_n46689_, new_n46674_ );
xor  ( new_n46691_, new_n46689_, new_n46674_ );
xor  ( new_n46692_, new_n46440_, new_n46406_ );
nand ( new_n46693_, new_n46692_, new_n46459_ );
or   ( new_n46694_, new_n46459_, new_n46443_ );
or   ( new_n46695_, new_n46694_, new_n46442_ );
and  ( new_n46696_, new_n46695_, new_n46693_ );
and  ( new_n46697_, new_n46696_, new_n46691_ );
or   ( new_n46698_, new_n46697_, new_n46690_ );
xor  ( new_n46699_, new_n46672_, new_n46670_ );
and  ( new_n46700_, new_n46699_, new_n46698_ );
nor  ( new_n46701_, new_n46700_, new_n46673_ );
nand ( new_n46702_, new_n46701_, new_n46559_ );
and  ( new_n46703_, new_n46702_, new_n46558_ );
and  ( new_n46704_, new_n46703_, new_n46536_ );
or   ( new_n46705_, new_n46704_, new_n46535_ );
xor  ( new_n46706_, new_n46526_, new_n46342_ );
or   ( new_n46707_, new_n46706_, new_n46705_ );
and  ( new_n46708_, new_n46707_, new_n46530_ );
and  ( new_n46709_, new_n46708_, new_n46338_ );
xor  ( new_n46710_, new_n46703_, new_n46536_ );
not  ( new_n46711_, new_n46710_ );
xor  ( new_n46712_, new_n46518_, new_n46516_ );
xor  ( new_n46713_, new_n46712_, new_n46522_ );
xor  ( new_n46714_, new_n46557_, new_n46555_ );
xor  ( new_n46715_, new_n46714_, new_n46701_ );
nor  ( new_n46716_, new_n46715_, new_n46713_ );
and  ( new_n46717_, new_n46715_, new_n46713_ );
nor  ( new_n46718_, RIbb2e530_37, RIbb2e5a8_36 );
not  ( new_n46719_, new_n46718_ );
and  ( new_n46720_, new_n46719_, new_n3115_ );
xor  ( new_n46721_, new_n43793_, new_n3113_ );
and  ( new_n46722_, new_n46721_, new_n3293_ );
nor  ( new_n46723_, new_n46722_, new_n46720_ );
or   ( new_n46724_, new_n46477_, new_n320_ );
xor  ( new_n46725_, new_n45584_, new_n309_ );
or   ( new_n46726_, new_n46725_, new_n317_ );
and  ( new_n46727_, new_n46726_, new_n46724_ );
or   ( new_n46728_, new_n46727_, new_n46723_ );
xor  ( new_n46729_, new_n46727_, new_n46723_ );
xnor ( new_n46730_, new_n46620_, new_n3116_ );
xor  ( new_n46731_, new_n46730_, new_n46629_ );
nand ( new_n46732_, new_n46731_, new_n46729_ );
and  ( new_n46733_, new_n46732_, new_n46728_ );
xor  ( new_n46734_, new_n45119_, new_n325_ );
or   ( new_n46735_, new_n46734_, new_n409_ );
or   ( new_n46736_, new_n46604_, new_n411_ );
and  ( new_n46737_, new_n46736_, new_n46735_ );
xor  ( new_n46738_, new_n44877_, RIbb2f070_13 );
nand ( new_n46739_, new_n46738_, new_n456_ );
or   ( new_n46740_, new_n46586_, new_n526_ );
and  ( new_n46741_, new_n46740_, new_n46739_ );
or   ( new_n46742_, new_n46741_, new_n46737_ );
xor  ( new_n46743_, new_n43952_, new_n1583_ );
or   ( new_n46744_, new_n46743_, new_n1844_ );
or   ( new_n46745_, new_n46590_, new_n1846_ );
and  ( new_n46746_, new_n46745_, new_n46744_ );
and  ( new_n46747_, new_n46741_, new_n46737_ );
or   ( new_n46748_, new_n46747_, new_n46746_ );
and  ( new_n46749_, new_n46748_, new_n46742_ );
nand ( new_n46750_, new_n46575_, new_n820_ );
xor  ( new_n46751_, new_n44506_, new_n745_ );
or   ( new_n46752_, new_n46751_, new_n897_ );
and  ( new_n46753_, new_n46752_, new_n46750_ );
xor  ( new_n46754_, new_n43799_, new_n2421_ );
or   ( new_n46755_, new_n46754_, new_n2807_ );
or   ( new_n46756_, new_n46581_, new_n2809_ );
and  ( new_n46757_, new_n46756_, new_n46755_ );
nor  ( new_n46758_, new_n46757_, new_n46753_ );
xor  ( new_n46759_, new_n44681_, RIbb2ef80_15 );
and  ( new_n46760_, new_n46759_, new_n662_ );
and  ( new_n46761_, new_n46570_, new_n660_ );
nor  ( new_n46762_, new_n46761_, new_n46760_ );
and  ( new_n46763_, new_n46757_, new_n46753_ );
nor  ( new_n46764_, new_n46763_, new_n46762_ );
nor  ( new_n46765_, new_n46764_, new_n46758_ );
or   ( new_n46766_, new_n46765_, new_n46749_ );
xor  ( new_n46767_, new_n45738_, new_n309_ );
or   ( new_n46768_, new_n46767_, new_n317_ );
or   ( new_n46769_, new_n46725_, new_n320_ );
and  ( new_n46770_, new_n46769_, new_n46768_ );
or   ( new_n46771_, new_n46600_, new_n340_ );
xor  ( new_n46772_, new_n45403_, new_n329_ );
or   ( new_n46773_, new_n46772_, new_n337_ );
and  ( new_n46774_, new_n46773_, new_n46771_ );
nor  ( new_n46775_, new_n46774_, new_n46770_ );
xor  ( new_n46776_, new_n43812_, RIbb2ebc0_23 );
and  ( new_n46777_, new_n46776_, new_n1476_ );
and  ( new_n46778_, new_n46609_, new_n1474_ );
nor  ( new_n46779_, new_n46778_, new_n46777_ );
not  ( new_n46780_, new_n46779_ );
nand ( new_n46781_, new_n46774_, new_n46770_ );
and  ( new_n46782_, new_n46781_, new_n46780_ );
or   ( new_n46783_, new_n46782_, new_n46775_ );
xor  ( new_n46784_, new_n46765_, new_n46749_ );
nand ( new_n46785_, new_n46784_, new_n46783_ );
and  ( new_n46786_, new_n46785_, new_n46766_ );
nor  ( new_n46787_, new_n46786_, new_n46733_ );
xor  ( new_n46788_, RIbb325e0_163, RIbb2c820_99 );
xor  ( new_n46789_, new_n46788_, new_n46421_ );
and  ( new_n46790_, new_n46789_, new_n43880_ );
not  ( new_n46791_, new_n46790_ );
xor  ( new_n46792_, new_n46619_, new_n43945_ );
not  ( new_n46793_, new_n46792_ );
or   ( new_n46794_, new_n46793_, new_n43983_ );
nor  ( new_n46795_, new_n46427_, new_n43880_ );
or   ( new_n46796_, new_n46428_, new_n43977_ );
or   ( new_n46797_, new_n46796_, new_n46795_ );
and  ( new_n46798_, new_n46797_, new_n46794_ );
nor  ( new_n46799_, new_n46798_, new_n46791_ );
xor  ( new_n46800_, new_n44183_, RIbb2ecb0_21 );
and  ( new_n46801_, new_n46800_, new_n1253_ );
and  ( new_n46802_, new_n46640_, new_n1251_ );
or   ( new_n46803_, new_n46802_, new_n46801_ );
xor  ( new_n46804_, new_n46798_, new_n46791_ );
and  ( new_n46805_, new_n46804_, new_n46803_ );
nor  ( new_n46806_, new_n46805_, new_n46799_ );
nand ( new_n46807_, new_n46658_, new_n1040_ );
xor  ( new_n46808_, new_n44319_, RIbb2eda0_19 );
nand ( new_n46809_, new_n46808_, new_n1042_ );
and  ( new_n46810_, new_n46809_, new_n46807_ );
xor  ( new_n46811_, new_n43884_, new_n2118_ );
or   ( new_n46812_, new_n46811_, new_n2425_ );
or   ( new_n46813_, new_n46653_, new_n2427_ );
and  ( new_n46814_, new_n46813_, new_n46812_ );
or   ( new_n46815_, new_n46814_, new_n46810_ );
xor  ( new_n46816_, new_n43937_, RIbb2e9e0_27 );
and  ( new_n46817_, new_n46816_, new_n2002_ );
and  ( new_n46818_, new_n46566_, new_n2000_ );
nor  ( new_n46819_, new_n46818_, new_n46817_ );
and  ( new_n46820_, new_n46814_, new_n46810_ );
or   ( new_n46821_, new_n46820_, new_n46819_ );
and  ( new_n46822_, new_n46821_, new_n46815_ );
nor  ( new_n46823_, new_n46822_, new_n46806_ );
xor  ( new_n46824_, new_n46822_, new_n46806_ );
not  ( new_n46825_, new_n46824_ );
or   ( new_n46826_, new_n46175_, new_n302_ );
or   ( new_n46827_, new_n46391_, new_n44007_ );
and  ( new_n46828_, new_n46827_, new_n46826_ );
or   ( new_n46829_, new_n46633_, new_n286_ );
xor  ( new_n46830_, new_n45928_, new_n275_ );
or   ( new_n46831_, new_n46830_, new_n283_ );
and  ( new_n46832_, new_n46831_, new_n46829_ );
or   ( new_n46833_, new_n46832_, new_n46828_ );
xor  ( new_n46834_, new_n43898_, new_n2797_ );
nor  ( new_n46835_, new_n46834_, new_n3117_ );
and  ( new_n46836_, new_n46648_, new_n2928_ );
nor  ( new_n46837_, new_n46836_, new_n46835_ );
and  ( new_n46838_, new_n46832_, new_n46828_ );
or   ( new_n46839_, new_n46838_, new_n46837_ );
and  ( new_n46840_, new_n46839_, new_n46833_ );
nor  ( new_n46841_, new_n46840_, new_n46825_ );
nor  ( new_n46842_, new_n46841_, new_n46823_ );
xnor ( new_n46843_, new_n46786_, new_n46733_ );
nor  ( new_n46844_, new_n46843_, new_n46842_ );
or   ( new_n46845_, new_n46844_, new_n46787_ );
xor  ( new_n46846_, new_n46668_, new_n46667_ );
and  ( new_n46847_, new_n46846_, new_n46845_ );
xor  ( new_n46848_, new_n46665_, new_n46664_ );
xnor ( new_n46849_, new_n46596_, new_n46580_ );
xor  ( new_n46850_, new_n46849_, new_n46614_ );
and  ( new_n46851_, new_n46850_, new_n46848_ );
xor  ( new_n46852_, new_n46662_, new_n46661_ );
xnor ( new_n46853_, new_n46638_, new_n46635_ );
xor  ( new_n46854_, new_n46853_, new_n46643_ );
and  ( new_n46855_, new_n46854_, new_n46852_ );
xor  ( new_n46856_, new_n46854_, new_n46852_ );
xnor ( new_n46857_, new_n46606_, new_n46602_ );
xor  ( new_n46858_, new_n46857_, new_n46611_ );
and  ( new_n46859_, new_n46858_, new_n46856_ );
nor  ( new_n46860_, new_n46859_, new_n46855_ );
not  ( new_n46861_, new_n46860_ );
xor  ( new_n46862_, new_n46850_, new_n46848_ );
and  ( new_n46863_, new_n46862_, new_n46861_ );
nor  ( new_n46864_, new_n46863_, new_n46851_ );
xnor ( new_n46865_, new_n46846_, new_n46845_ );
nor  ( new_n46866_, new_n46865_, new_n46864_ );
nor  ( new_n46867_, new_n46866_, new_n46847_ );
not  ( new_n46868_, new_n46867_ );
xor  ( new_n46869_, new_n46699_, new_n46698_ );
and  ( new_n46870_, new_n46869_, new_n46868_ );
xor  ( new_n46871_, new_n46869_, new_n46868_ );
xor  ( new_n46872_, new_n46553_, new_n46552_ );
and  ( new_n46873_, new_n46872_, new_n46871_ );
nor  ( new_n46874_, new_n46873_, new_n46870_ );
nor  ( new_n46875_, new_n46874_, new_n46717_ );
nor  ( new_n46876_, new_n46875_, new_n46716_ );
nand ( new_n46877_, new_n46876_, new_n46711_ );
xor  ( new_n46878_, new_n43894_, RIbb2e710_33 );
nand ( new_n46879_, new_n46878_, new_n2928_ );
xor  ( new_n46880_, new_n43799_, new_n2797_ );
or   ( new_n46881_, new_n46880_, new_n3117_ );
and  ( new_n46882_, new_n46881_, new_n46879_ );
xor  ( new_n46883_, new_n43952_, new_n1840_ );
or   ( new_n46884_, new_n46883_, new_n2122_ );
xor  ( new_n46885_, new_n43956_, new_n1840_ );
or   ( new_n46886_, new_n46885_, new_n2124_ );
and  ( new_n46887_, new_n46886_, new_n46884_ );
nor  ( new_n46888_, new_n46887_, new_n46882_ );
xor  ( new_n46889_, new_n44877_, RIbb2ef80_15 );
and  ( new_n46890_, new_n46889_, new_n662_ );
xor  ( new_n46891_, new_n44785_, RIbb2ef80_15 );
and  ( new_n46892_, new_n46891_, new_n660_ );
or   ( new_n46893_, new_n46892_, new_n46890_ );
xor  ( new_n46894_, new_n46887_, new_n46882_ );
and  ( new_n46895_, new_n46894_, new_n46893_ );
nor  ( new_n46896_, new_n46895_, new_n46888_ );
not  ( new_n46897_, new_n46896_ );
xor  ( new_n46898_, new_n44407_, RIbb2eda0_19 );
and  ( new_n46899_, new_n46898_, new_n1042_ );
and  ( new_n46900_, new_n46808_, new_n1040_ );
nor  ( new_n46901_, new_n46900_, new_n46899_ );
xor  ( new_n46902_, new_n43888_, new_n2118_ );
or   ( new_n46903_, new_n46902_, new_n2425_ );
or   ( new_n46904_, new_n46811_, new_n2427_ );
and  ( new_n46905_, new_n46904_, new_n46903_ );
xor  ( new_n46906_, new_n43803_, new_n2421_ );
or   ( new_n46907_, new_n46906_, new_n2807_ );
or   ( new_n46908_, new_n46754_, new_n2809_ );
and  ( new_n46909_, new_n46908_, new_n46907_ );
xnor ( new_n46910_, new_n46909_, new_n46905_ );
xor  ( new_n46911_, new_n46910_, new_n46901_ );
xor  ( new_n46912_, new_n46911_, new_n46897_ );
xor  ( new_n46913_, new_n43787_, RIbb2e620_35 );
and  ( new_n46914_, new_n46913_, new_n3293_ );
and  ( new_n46915_, new_n46721_, new_n3291_ );
nor  ( new_n46916_, new_n46915_, new_n46914_ );
xor  ( new_n46917_, new_n44218_, RIbb2ecb0_21 );
nand ( new_n46918_, new_n46917_, new_n1253_ );
nand ( new_n46919_, new_n46800_, new_n1251_ );
and  ( new_n46920_, new_n46919_, new_n46918_ );
xor  ( new_n46921_, new_n46037_, new_n275_ );
or   ( new_n46922_, new_n46921_, new_n283_ );
or   ( new_n46923_, new_n46830_, new_n286_ );
and  ( new_n46924_, new_n46923_, new_n46922_ );
xnor ( new_n46925_, new_n46924_, new_n46920_ );
xor  ( new_n46926_, new_n46925_, new_n46916_ );
xnor ( new_n46927_, new_n46926_, new_n46912_ );
xor  ( new_n46928_, new_n45204_, RIbb2f160_11 );
and  ( new_n46929_, new_n46928_, new_n371_ );
xor  ( new_n46930_, new_n45403_, new_n325_ );
nor  ( new_n46931_, new_n46930_, new_n409_ );
nor  ( new_n46932_, new_n46931_, new_n46929_ );
xor  ( new_n46933_, new_n45119_, new_n400_ );
or   ( new_n46934_, new_n46933_, new_n524_ );
xor  ( new_n46935_, new_n44974_, RIbb2f070_13 );
nand ( new_n46936_, new_n46935_, new_n454_ );
and  ( new_n46937_, new_n46936_, new_n46934_ );
nor  ( new_n46938_, new_n46937_, new_n46932_ );
not  ( new_n46939_, new_n46938_ );
xor  ( new_n46940_, new_n43812_, RIbb2ead0_25 );
and  ( new_n46941_, new_n46940_, new_n1741_ );
xor  ( new_n46942_, new_n43985_, RIbb2ead0_25 );
and  ( new_n46943_, new_n46942_, new_n1739_ );
nor  ( new_n46944_, new_n46943_, new_n46941_ );
and  ( new_n46945_, new_n46937_, new_n46932_ );
nor  ( new_n46946_, new_n46945_, new_n46944_ );
not  ( new_n46947_, new_n46946_ );
and  ( new_n46948_, new_n46947_, new_n46939_ );
xor  ( new_n46949_, RIbb326d0_165, RIbb2c730_101 );
and  ( new_n46950_, new_n46415_, new_n43583_ );
nor  ( new_n46951_, new_n46950_, new_n43656_ );
not  ( new_n46952_, new_n46951_ );
and  ( new_n46953_, new_n46952_, new_n43586_ );
nor  ( new_n46954_, new_n46953_, new_n43655_ );
not  ( new_n46955_, new_n46954_ );
and  ( new_n46956_, new_n46955_, new_n43588_ );
nor  ( new_n46957_, new_n46956_, new_n43654_ );
xnor ( new_n46958_, new_n46957_, new_n46949_ );
and  ( new_n46959_, new_n46958_, new_n43880_ );
not  ( new_n46960_, new_n46959_ );
xor  ( new_n46961_, RIbb32658_164, RIbb2c7a8_100 );
xor  ( new_n46962_, new_n46961_, new_n46418_ );
xor  ( new_n46963_, new_n46962_, new_n43879_ );
or   ( new_n46964_, new_n46963_, new_n43983_ );
nor  ( new_n46965_, new_n46789_, new_n43880_ );
or   ( new_n46966_, new_n46790_, new_n43977_ );
or   ( new_n46967_, new_n46966_, new_n46965_ );
and  ( new_n46968_, new_n46967_, new_n46964_ );
nor  ( new_n46969_, new_n46968_, new_n46960_ );
not  ( new_n46970_, new_n46623_ );
and  ( new_n46971_, new_n46970_, new_n295_ );
and  ( new_n46972_, new_n46793_, new_n43949_ );
or   ( new_n46973_, new_n46972_, new_n46971_ );
xor  ( new_n46974_, new_n46968_, new_n46960_ );
and  ( new_n46975_, new_n46974_, new_n46973_ );
or   ( new_n46976_, new_n46975_, new_n46969_ );
and  ( new_n46977_, new_n46392_, new_n295_ );
and  ( new_n46978_, new_n46970_, new_n43949_ );
nor  ( new_n46979_, new_n46978_, new_n46977_ );
xor  ( new_n46980_, new_n46789_, new_n43945_ );
nand ( new_n46981_, new_n46980_, new_n43982_ );
nor  ( new_n46982_, new_n46619_, new_n43880_ );
or   ( new_n46983_, new_n46620_, new_n43977_ );
or   ( new_n46984_, new_n46983_, new_n46982_ );
and  ( new_n46985_, new_n46984_, new_n46981_ );
xor  ( new_n46986_, new_n46985_, new_n3460_ );
xor  ( new_n46987_, new_n46986_, new_n46979_ );
xnor ( new_n46988_, new_n46987_, new_n46976_ );
xor  ( new_n46989_, new_n46988_, new_n46948_ );
or   ( new_n46990_, new_n46921_, new_n286_ );
xor  ( new_n46991_, new_n46137_, RIbb2f430_5 );
nand ( new_n46992_, new_n46991_, new_n282_ );
and  ( new_n46993_, new_n46992_, new_n46990_ );
xor  ( new_n46994_, new_n44183_, RIbb2ebc0_23 );
nand ( new_n46995_, new_n46994_, new_n1476_ );
xor  ( new_n46996_, new_n43914_, new_n1355_ );
or   ( new_n46997_, new_n46996_, new_n1595_ );
and  ( new_n46998_, new_n46997_, new_n46995_ );
nor  ( new_n46999_, new_n46998_, new_n46993_ );
xor  ( new_n47000_, new_n45928_, new_n309_ );
nor  ( new_n47001_, new_n47000_, new_n317_ );
xor  ( new_n47002_, new_n45597_, RIbb2f340_7 );
and  ( new_n47003_, new_n47002_, new_n314_ );
nor  ( new_n47004_, new_n47003_, new_n47001_ );
and  ( new_n47005_, new_n46998_, new_n46993_ );
nor  ( new_n47006_, new_n47005_, new_n47004_ );
nor  ( new_n47007_, new_n47006_, new_n46999_ );
xor  ( new_n47008_, new_n43937_, new_n2118_ );
or   ( new_n47009_, new_n47008_, new_n2425_ );
or   ( new_n47010_, new_n46902_, new_n2427_ );
and  ( new_n47011_, new_n47010_, new_n47009_ );
xor  ( new_n47012_, new_n44681_, RIbb2ee90_17 );
nand ( new_n47013_, new_n47012_, new_n822_ );
xor  ( new_n47014_, new_n44600_, new_n745_ );
or   ( new_n47015_, new_n47014_, new_n899_ );
and  ( new_n47016_, new_n47015_, new_n47013_ );
or   ( new_n47017_, new_n47016_, new_n47011_ );
and  ( new_n47018_, new_n46898_, new_n1040_ );
xor  ( new_n47019_, new_n44506_, RIbb2eda0_19 );
and  ( new_n47020_, new_n47019_, new_n1042_ );
nor  ( new_n47021_, new_n47020_, new_n47018_ );
and  ( new_n47022_, new_n47016_, new_n47011_ );
or   ( new_n47023_, new_n47022_, new_n47021_ );
and  ( new_n47024_, new_n47023_, new_n47017_ );
xnor ( new_n47025_, new_n47024_, new_n47007_ );
or   ( new_n47026_, new_n46906_, new_n2809_ );
xor  ( new_n47027_, new_n43884_, new_n2421_ );
or   ( new_n47028_, new_n47027_, new_n2807_ );
and  ( new_n47029_, new_n47028_, new_n47026_ );
nand ( new_n47030_, new_n46913_, new_n3291_ );
xor  ( new_n47031_, new_n43898_, new_n3113_ );
or   ( new_n47032_, new_n47031_, new_n3461_ );
and  ( new_n47033_, new_n47032_, new_n47030_ );
or   ( new_n47034_, new_n47033_, new_n47029_ );
and  ( new_n47035_, new_n46917_, new_n1251_ );
xor  ( new_n47036_, new_n44319_, RIbb2ecb0_21 );
and  ( new_n47037_, new_n47036_, new_n1253_ );
nor  ( new_n47038_, new_n47037_, new_n47035_ );
and  ( new_n47039_, new_n47033_, new_n47029_ );
or   ( new_n47040_, new_n47039_, new_n47038_ );
and  ( new_n47041_, new_n47040_, new_n47034_ );
xor  ( new_n47042_, new_n47041_, new_n47025_ );
xor  ( new_n47043_, new_n47042_, new_n46989_ );
xor  ( new_n47044_, new_n47043_, new_n46927_ );
xor  ( new_n47045_, RIbb327c0_167, RIbb2c640_103 );
xor  ( new_n47046_, new_n47045_, new_n46952_ );
nand ( new_n47047_, new_n47046_, new_n43880_ );
or   ( new_n47048_, new_n46980_, new_n302_ );
xor  ( new_n47049_, new_n46962_, new_n43945_ );
or   ( new_n47050_, new_n47049_, new_n44007_ );
and  ( new_n47051_, new_n47050_, new_n47048_ );
or   ( new_n47052_, new_n47051_, new_n47047_ );
xor  ( new_n47053_, new_n46427_, RIbb2f430_5 );
and  ( new_n47054_, new_n47053_, new_n280_ );
xor  ( new_n47055_, new_n46619_, new_n275_ );
nor  ( new_n47056_, new_n47055_, new_n283_ );
or   ( new_n47057_, new_n47056_, new_n47054_ );
xor  ( new_n47058_, new_n47051_, new_n47047_ );
nand ( new_n47059_, new_n47058_, new_n47057_ );
and  ( new_n47060_, new_n47059_, new_n47052_ );
nor  ( new_n47061_, RIbb2e350_41, RIbb2e3c8_40 );
not  ( new_n47062_, new_n47061_ );
and  ( new_n47063_, new_n47062_, new_n3894_ );
xor  ( new_n47064_, new_n43793_, new_n3892_ );
and  ( new_n47065_, new_n47064_, new_n4034_ );
nor  ( new_n47066_, new_n47065_, new_n47063_ );
nor  ( new_n47067_, new_n47066_, new_n47060_ );
xor  ( new_n47068_, new_n43956_, new_n2118_ );
or   ( new_n47069_, new_n47068_, new_n2427_ );
xor  ( new_n47070_, new_n43952_, new_n2118_ );
or   ( new_n47071_, new_n47070_, new_n2425_ );
and  ( new_n47072_, new_n47071_, new_n47069_ );
xor  ( new_n47073_, new_n44600_, RIbb2eda0_19 );
nand ( new_n47074_, new_n47073_, new_n1040_ );
xor  ( new_n47075_, new_n44681_, new_n893_ );
or   ( new_n47076_, new_n47075_, new_n1135_ );
and  ( new_n47077_, new_n47076_, new_n47074_ );
nor  ( new_n47078_, new_n47077_, new_n47072_ );
xor  ( new_n47079_, new_n43894_, RIbb2e620_35 );
and  ( new_n47080_, new_n47079_, new_n3291_ );
xor  ( new_n47081_, new_n43799_, new_n3113_ );
nor  ( new_n47082_, new_n47081_, new_n3461_ );
nor  ( new_n47083_, new_n47082_, new_n47080_ );
and  ( new_n47084_, new_n47077_, new_n47072_ );
nor  ( new_n47085_, new_n47084_, new_n47083_ );
or   ( new_n47086_, new_n47085_, new_n47078_ );
xor  ( new_n47087_, new_n47066_, new_n47060_ );
and  ( new_n47088_, new_n47087_, new_n47086_ );
or   ( new_n47089_, new_n47088_, new_n47067_ );
or   ( new_n47090_, new_n46980_, new_n44007_ );
or   ( new_n47091_, new_n46792_, new_n302_ );
and  ( new_n47092_, new_n47091_, new_n47090_ );
nor  ( new_n47093_, new_n47092_, new_n3894_ );
and  ( new_n47094_, new_n46991_, new_n280_ );
and  ( new_n47095_, new_n47053_, new_n282_ );
or   ( new_n47096_, new_n47095_, new_n47094_ );
xor  ( new_n47097_, new_n47092_, new_n3894_ );
and  ( new_n47098_, new_n47097_, new_n47096_ );
or   ( new_n47099_, new_n47098_, new_n47093_ );
not  ( new_n47100_, RIbb2e4b8_38 );
and  ( new_n47101_, new_n3892_, new_n47100_ );
not  ( new_n47102_, new_n47101_ );
and  ( new_n47103_, new_n47102_, new_n3459_ );
xor  ( new_n47104_, new_n43793_, new_n3457_ );
and  ( new_n47105_, new_n47104_, new_n3733_ );
nor  ( new_n47106_, new_n47105_, new_n47103_ );
xor  ( new_n47107_, new_n45584_, RIbb2f250_9 );
nand ( new_n47108_, new_n47107_, new_n334_ );
xor  ( new_n47109_, new_n45738_, new_n329_ );
or   ( new_n47110_, new_n47109_, new_n337_ );
nand ( new_n47111_, new_n47110_, new_n47108_ );
xor  ( new_n47112_, new_n47111_, new_n47106_ );
xor  ( new_n47113_, new_n47112_, new_n47099_ );
nand ( new_n47114_, new_n47113_, new_n47089_ );
xor  ( new_n47115_, new_n43888_, new_n2421_ );
or   ( new_n47116_, new_n47115_, new_n2809_ );
xor  ( new_n47117_, new_n43937_, new_n2421_ );
or   ( new_n47118_, new_n47117_, new_n2807_ );
and  ( new_n47119_, new_n47118_, new_n47116_ );
xor  ( new_n47120_, new_n43803_, new_n2797_ );
or   ( new_n47121_, new_n47120_, new_n3119_ );
xor  ( new_n47122_, new_n43884_, RIbb2e710_33 );
nand ( new_n47123_, new_n47122_, new_n2930_ );
and  ( new_n47124_, new_n47123_, new_n47121_ );
nor  ( new_n47125_, new_n47124_, new_n47119_ );
xor  ( new_n47126_, new_n44506_, RIbb2ecb0_21 );
and  ( new_n47127_, new_n47126_, new_n1253_ );
xor  ( new_n47128_, new_n44407_, RIbb2ecb0_21 );
and  ( new_n47129_, new_n47128_, new_n1251_ );
or   ( new_n47130_, new_n47129_, new_n47127_ );
xor  ( new_n47131_, new_n47124_, new_n47119_ );
and  ( new_n47132_, new_n47131_, new_n47130_ );
nor  ( new_n47133_, new_n47132_, new_n47125_ );
xor  ( new_n47134_, new_n44785_, RIbb2ee90_17 );
nand ( new_n47135_, new_n47134_, new_n820_ );
xor  ( new_n47136_, new_n44877_, RIbb2ee90_17 );
nand ( new_n47137_, new_n47136_, new_n822_ );
and  ( new_n47138_, new_n47137_, new_n47135_ );
xor  ( new_n47139_, new_n43985_, RIbb2e9e0_27 );
nand ( new_n47140_, new_n47139_, new_n2000_ );
xor  ( new_n47141_, new_n43812_, new_n1840_ );
or   ( new_n47142_, new_n47141_, new_n2122_ );
and  ( new_n47143_, new_n47142_, new_n47140_ );
or   ( new_n47144_, new_n47143_, new_n47138_ );
xor  ( new_n47145_, new_n44974_, RIbb2ef80_15 );
and  ( new_n47146_, new_n47145_, new_n660_ );
xor  ( new_n47147_, new_n45119_, new_n520_ );
nor  ( new_n47148_, new_n47147_, new_n755_ );
or   ( new_n47149_, new_n47148_, new_n47146_ );
xor  ( new_n47150_, new_n47143_, new_n47138_ );
nand ( new_n47151_, new_n47150_, new_n47149_ );
and  ( new_n47152_, new_n47151_, new_n47144_ );
nor  ( new_n47153_, new_n47152_, new_n47133_ );
xnor ( new_n47154_, new_n47152_, new_n47133_ );
xor  ( new_n47155_, new_n43787_, new_n3457_ );
or   ( new_n47156_, new_n47155_, new_n3898_ );
xor  ( new_n47157_, new_n43898_, new_n3457_ );
or   ( new_n47158_, new_n47157_, new_n3896_ );
and  ( new_n47159_, new_n47158_, new_n47156_ );
xor  ( new_n47160_, new_n46037_, new_n309_ );
or   ( new_n47161_, new_n47160_, new_n320_ );
xor  ( new_n47162_, new_n46137_, new_n309_ );
or   ( new_n47163_, new_n47162_, new_n317_ );
and  ( new_n47164_, new_n47163_, new_n47161_ );
nor  ( new_n47165_, new_n47164_, new_n47159_ );
and  ( new_n47166_, new_n47164_, new_n47159_ );
xor  ( new_n47167_, new_n44319_, RIbb2ebc0_23 );
and  ( new_n47168_, new_n47167_, new_n1476_ );
xor  ( new_n47169_, new_n44218_, RIbb2ebc0_23 );
and  ( new_n47170_, new_n47169_, new_n1474_ );
nor  ( new_n47171_, new_n47170_, new_n47168_ );
nor  ( new_n47172_, new_n47171_, new_n47166_ );
nor  ( new_n47173_, new_n47172_, new_n47165_ );
nor  ( new_n47174_, new_n47173_, new_n47154_ );
or   ( new_n47175_, new_n47174_, new_n47153_ );
xor  ( new_n47176_, new_n47113_, new_n47089_ );
nand ( new_n47177_, new_n47176_, new_n47175_ );
and  ( new_n47178_, new_n47177_, new_n47114_ );
nand ( new_n47179_, new_n47036_, new_n1251_ );
nand ( new_n47180_, new_n47128_, new_n1253_ );
and  ( new_n47181_, new_n47180_, new_n47179_ );
or   ( new_n47182_, new_n46880_, new_n3119_ );
or   ( new_n47183_, new_n47120_, new_n3117_ );
and  ( new_n47184_, new_n47183_, new_n47182_ );
nor  ( new_n47185_, new_n47184_, new_n47181_ );
and  ( new_n47186_, new_n46994_, new_n1474_ );
and  ( new_n47187_, new_n47169_, new_n1476_ );
nor  ( new_n47188_, new_n47187_, new_n47186_ );
and  ( new_n47189_, new_n47184_, new_n47181_ );
nor  ( new_n47190_, new_n47189_, new_n47188_ );
nor  ( new_n47191_, new_n47190_, new_n47185_ );
nand ( new_n47192_, new_n47079_, new_n3293_ );
or   ( new_n47193_, new_n47031_, new_n3463_ );
and  ( new_n47194_, new_n47193_, new_n47192_ );
or   ( new_n47195_, new_n47027_, new_n2809_ );
or   ( new_n47196_, new_n47115_, new_n2807_ );
and  ( new_n47197_, new_n47196_, new_n47195_ );
or   ( new_n47198_, new_n47197_, new_n47194_ );
and  ( new_n47199_, new_n47073_, new_n1042_ );
and  ( new_n47200_, new_n47019_, new_n1040_ );
nor  ( new_n47201_, new_n47200_, new_n47199_ );
and  ( new_n47202_, new_n47197_, new_n47194_ );
or   ( new_n47203_, new_n47202_, new_n47201_ );
and  ( new_n47204_, new_n47203_, new_n47198_ );
nor  ( new_n47205_, new_n47204_, new_n47191_ );
and  ( new_n47206_, new_n47204_, new_n47191_ );
or   ( new_n47207_, new_n47155_, new_n3896_ );
nand ( new_n47208_, new_n47104_, new_n3731_ );
and  ( new_n47209_, new_n47208_, new_n47207_ );
xor  ( new_n47210_, new_n45597_, new_n329_ );
or   ( new_n47211_, new_n47210_, new_n337_ );
or   ( new_n47212_, new_n47109_, new_n340_ );
and  ( new_n47213_, new_n47212_, new_n47211_ );
nor  ( new_n47214_, new_n47213_, new_n47209_ );
and  ( new_n47215_, new_n47213_, new_n47209_ );
nor  ( new_n47216_, new_n47160_, new_n317_ );
nor  ( new_n47217_, new_n47000_, new_n320_ );
nor  ( new_n47218_, new_n47217_, new_n47216_ );
nor  ( new_n47219_, new_n47218_, new_n47215_ );
nor  ( new_n47220_, new_n47219_, new_n47214_ );
nor  ( new_n47221_, new_n47220_, new_n47206_ );
nor  ( new_n47222_, new_n47221_, new_n47205_ );
and  ( new_n47223_, new_n47111_, new_n47106_ );
and  ( new_n47224_, new_n47112_, new_n47099_ );
or   ( new_n47225_, new_n47224_, new_n47223_ );
and  ( new_n47226_, new_n46935_, new_n456_ );
and  ( new_n47227_, new_n46738_, new_n454_ );
nor  ( new_n47228_, new_n47227_, new_n47226_ );
nand ( new_n47229_, new_n46942_, new_n1741_ );
or   ( new_n47230_, new_n46743_, new_n1846_ );
and  ( new_n47231_, new_n47230_, new_n47229_ );
nand ( new_n47232_, new_n46759_, new_n660_ );
nand ( new_n47233_, new_n46891_, new_n662_ );
and  ( new_n47234_, new_n47233_, new_n47232_ );
xnor ( new_n47235_, new_n47234_, new_n47231_ );
xor  ( new_n47236_, new_n47235_, new_n47228_ );
xnor ( new_n47237_, new_n47236_, new_n47225_ );
xnor ( new_n47238_, new_n47237_, new_n47222_ );
and  ( new_n47239_, new_n47107_, new_n336_ );
nor  ( new_n47240_, new_n46772_, new_n340_ );
nor  ( new_n47241_, new_n47240_, new_n47239_ );
nand ( new_n47242_, new_n46928_, new_n373_ );
or   ( new_n47243_, new_n46734_, new_n411_ );
and  ( new_n47244_, new_n47243_, new_n47242_ );
xnor ( new_n47245_, new_n47244_, new_n47106_ );
xor  ( new_n47246_, new_n47245_, new_n47241_ );
and  ( new_n47247_, new_n46878_, new_n2930_ );
nor  ( new_n47248_, new_n46834_, new_n3119_ );
nor  ( new_n47249_, new_n47248_, new_n47247_ );
or   ( new_n47250_, new_n46885_, new_n2122_ );
nand ( new_n47251_, new_n46816_, new_n2000_ );
and  ( new_n47252_, new_n47251_, new_n47250_ );
or   ( new_n47253_, new_n47014_, new_n897_ );
or   ( new_n47254_, new_n46751_, new_n899_ );
and  ( new_n47255_, new_n47254_, new_n47253_ );
xnor ( new_n47256_, new_n47255_, new_n47252_ );
xor  ( new_n47257_, new_n47256_, new_n47249_ );
xor  ( new_n47258_, new_n47257_, new_n47246_ );
or   ( new_n47259_, new_n46996_, new_n1593_ );
nand ( new_n47260_, new_n46776_, new_n1474_ );
and  ( new_n47261_, new_n47260_, new_n47259_ );
nand ( new_n47262_, new_n46962_, new_n43880_ );
or   ( new_n47263_, new_n46767_, new_n320_ );
nand ( new_n47264_, new_n47002_, new_n316_ );
and  ( new_n47265_, new_n47264_, new_n47263_ );
xor  ( new_n47266_, new_n47265_, new_n47262_ );
xor  ( new_n47267_, new_n47266_, new_n47261_ );
xor  ( new_n47268_, new_n47267_, new_n47258_ );
xor  ( new_n47269_, new_n47268_, new_n47238_ );
xor  ( new_n47270_, new_n47269_, new_n47178_ );
or   ( new_n47271_, new_n47270_, new_n47044_ );
xor  ( new_n47272_, new_n47176_, new_n47175_ );
or   ( new_n47273_, new_n46933_, new_n526_ );
xor  ( new_n47274_, new_n45204_, RIbb2f070_13 );
nand ( new_n47275_, new_n47274_, new_n456_ );
and  ( new_n47276_, new_n47275_, new_n47273_ );
or   ( new_n47277_, new_n46930_, new_n411_ );
xor  ( new_n47278_, new_n45584_, new_n325_ );
or   ( new_n47279_, new_n47278_, new_n409_ );
and  ( new_n47280_, new_n47279_, new_n47277_ );
nor  ( new_n47281_, new_n47280_, new_n47276_ );
nor  ( new_n47282_, new_n46883_, new_n2124_ );
and  ( new_n47283_, new_n47139_, new_n2002_ );
nor  ( new_n47284_, new_n47283_, new_n47282_ );
and  ( new_n47285_, new_n47280_, new_n47276_ );
nor  ( new_n47286_, new_n47285_, new_n47284_ );
or   ( new_n47287_, new_n47286_, new_n47281_ );
xnor ( new_n47288_, new_n47016_, new_n47011_ );
xor  ( new_n47289_, new_n47288_, new_n47021_ );
xor  ( new_n47290_, new_n47289_, new_n47287_ );
xnor ( new_n47291_, new_n47033_, new_n47029_ );
xor  ( new_n47292_, new_n47291_, new_n47038_ );
xor  ( new_n47293_, new_n47292_, new_n47290_ );
and  ( new_n47294_, new_n47293_, new_n47272_ );
xor  ( new_n47295_, RIbb32838_168, RIbb2c5c8_104 );
xor  ( new_n47296_, new_n47295_, new_n46415_ );
and  ( new_n47297_, new_n47296_, new_n43880_ );
not  ( new_n47298_, new_n47297_ );
xor  ( new_n47299_, new_n47046_, new_n43945_ );
not  ( new_n47300_, new_n47299_ );
or   ( new_n47301_, new_n47300_, new_n43983_ );
xor  ( new_n47302_, RIbb32748_166, RIbb2c6b8_102 );
xor  ( new_n47303_, new_n47302_, new_n46955_ );
or   ( new_n47304_, new_n47303_, new_n43880_ );
and  ( new_n47305_, new_n47303_, new_n43880_ );
not  ( new_n47306_, new_n47305_ );
and  ( new_n47307_, new_n47306_, new_n43978_ );
nand ( new_n47308_, new_n47307_, new_n47304_ );
and  ( new_n47309_, new_n47308_, new_n47301_ );
nor  ( new_n47310_, new_n47309_, new_n47298_ );
nor  ( new_n47311_, new_n47049_, new_n302_ );
xor  ( new_n47312_, new_n46958_, new_n43945_ );
not  ( new_n47313_, new_n47312_ );
and  ( new_n47314_, new_n47313_, new_n43949_ );
nor  ( new_n47315_, new_n47314_, new_n47311_ );
xor  ( new_n47316_, new_n47309_, new_n47297_ );
nor  ( new_n47317_, new_n47316_, new_n47315_ );
nor  ( new_n47318_, new_n47317_, new_n47310_ );
nor  ( new_n47319_, new_n47055_, new_n286_ );
xor  ( new_n47320_, new_n46789_, new_n275_ );
nor  ( new_n47321_, new_n47320_, new_n283_ );
nor  ( new_n47322_, new_n47321_, new_n47319_ );
or   ( new_n47323_, new_n47162_, new_n320_ );
xor  ( new_n47324_, new_n46427_, new_n309_ );
or   ( new_n47325_, new_n47324_, new_n317_ );
and  ( new_n47326_, new_n47325_, new_n47323_ );
and  ( new_n47327_, new_n47326_, new_n4294_ );
or   ( new_n47328_, new_n47327_, new_n47322_ );
or   ( new_n47329_, new_n47326_, new_n4294_ );
and  ( new_n47330_, new_n47329_, new_n47328_ );
nor  ( new_n47331_, new_n47330_, new_n47318_ );
xor  ( new_n47332_, new_n47330_, new_n47318_ );
xor  ( new_n47333_, new_n47058_, new_n47057_ );
and  ( new_n47334_, new_n47333_, new_n47332_ );
or   ( new_n47335_, new_n47334_, new_n47331_ );
xor  ( new_n47336_, new_n47087_, new_n47086_ );
and  ( new_n47337_, new_n47336_, new_n47335_ );
and  ( new_n47338_, new_n47122_, new_n2928_ );
xor  ( new_n47339_, new_n43888_, RIbb2e710_33 );
and  ( new_n47340_, new_n47339_, new_n2930_ );
nor  ( new_n47341_, new_n47340_, new_n47338_ );
nand ( new_n47342_, new_n47126_, new_n1251_ );
xor  ( new_n47343_, new_n44600_, new_n1126_ );
or   ( new_n47344_, new_n47343_, new_n1364_ );
and  ( new_n47345_, new_n47344_, new_n47342_ );
nor  ( new_n47346_, new_n47345_, new_n47341_ );
and  ( new_n47347_, new_n47167_, new_n1474_ );
xor  ( new_n47348_, new_n44407_, RIbb2ebc0_23 );
and  ( new_n47349_, new_n47348_, new_n1476_ );
nor  ( new_n47350_, new_n47349_, new_n47347_ );
and  ( new_n47351_, new_n47345_, new_n47341_ );
nor  ( new_n47352_, new_n47351_, new_n47350_ );
nor  ( new_n47353_, new_n47352_, new_n47346_ );
xor  ( new_n47354_, new_n43787_, new_n3892_ );
or   ( new_n47355_, new_n47354_, new_n4302_ );
nand ( new_n47356_, new_n47064_, new_n4032_ );
and  ( new_n47357_, new_n47356_, new_n47355_ );
or   ( new_n47358_, new_n47081_, new_n3463_ );
xor  ( new_n47359_, new_n43803_, new_n3113_ );
or   ( new_n47360_, new_n47359_, new_n3461_ );
and  ( new_n47361_, new_n47360_, new_n47358_ );
or   ( new_n47362_, new_n47361_, new_n47357_ );
xor  ( new_n47363_, new_n44183_, RIbb2ead0_25 );
and  ( new_n47364_, new_n47363_, new_n1739_ );
xor  ( new_n47365_, new_n44218_, RIbb2ead0_25 );
and  ( new_n47366_, new_n47365_, new_n1741_ );
or   ( new_n47367_, new_n47366_, new_n47364_ );
xor  ( new_n47368_, new_n47361_, new_n47357_ );
nand ( new_n47369_, new_n47368_, new_n47367_ );
and  ( new_n47370_, new_n47369_, new_n47362_ );
nor  ( new_n47371_, new_n47370_, new_n47353_ );
xor  ( new_n47372_, new_n45597_, RIbb2f160_11 );
nand ( new_n47373_, new_n47372_, new_n373_ );
xor  ( new_n47374_, new_n45738_, new_n325_ );
or   ( new_n47375_, new_n47374_, new_n411_ );
and  ( new_n47376_, new_n47375_, new_n47373_ );
xor  ( new_n47377_, new_n43914_, RIbb2e9e0_27 );
nand ( new_n47378_, new_n47377_, new_n2002_ );
or   ( new_n47379_, new_n47141_, new_n2124_ );
and  ( new_n47380_, new_n47379_, new_n47378_ );
nor  ( new_n47381_, new_n47380_, new_n47376_ );
xor  ( new_n47382_, new_n46037_, new_n329_ );
nor  ( new_n47383_, new_n47382_, new_n337_ );
xor  ( new_n47384_, new_n45928_, new_n329_ );
nor  ( new_n47385_, new_n47384_, new_n340_ );
nor  ( new_n47386_, new_n47385_, new_n47383_ );
xnor ( new_n47387_, new_n47380_, new_n47376_ );
nor  ( new_n47388_, new_n47387_, new_n47386_ );
or   ( new_n47389_, new_n47388_, new_n47381_ );
xor  ( new_n47390_, new_n47370_, new_n47353_ );
and  ( new_n47391_, new_n47390_, new_n47389_ );
or   ( new_n47392_, new_n47391_, new_n47371_ );
xor  ( new_n47393_, new_n47336_, new_n47335_ );
and  ( new_n47394_, new_n47393_, new_n47392_ );
or   ( new_n47395_, new_n47394_, new_n47337_ );
xor  ( new_n47396_, new_n47293_, new_n47272_ );
and  ( new_n47397_, new_n47396_, new_n47395_ );
or   ( new_n47398_, new_n47397_, new_n47294_ );
xor  ( new_n47399_, new_n47270_, new_n47044_ );
nand ( new_n47400_, new_n47399_, new_n47398_ );
and  ( new_n47401_, new_n47400_, new_n47271_ );
or   ( new_n47402_, new_n46963_, new_n43977_ );
or   ( new_n47403_, new_n47313_, new_n43983_ );
and  ( new_n47404_, new_n47403_, new_n47402_ );
nor  ( new_n47405_, new_n47404_, new_n47306_ );
and  ( new_n47406_, new_n46940_, new_n1739_ );
xor  ( new_n47407_, new_n43914_, RIbb2ead0_25 );
and  ( new_n47408_, new_n47407_, new_n1741_ );
or   ( new_n47409_, new_n47408_, new_n47406_ );
xor  ( new_n47410_, new_n47404_, new_n47306_ );
and  ( new_n47411_, new_n47410_, new_n47409_ );
or   ( new_n47412_, new_n47411_, new_n47405_ );
xor  ( new_n47413_, new_n46974_, new_n46973_ );
and  ( new_n47414_, new_n47413_, new_n47412_ );
or   ( new_n47415_, new_n47068_, new_n2425_ );
or   ( new_n47416_, new_n47008_, new_n2427_ );
and  ( new_n47417_, new_n47416_, new_n47415_ );
nand ( new_n47418_, new_n46889_, new_n660_ );
nand ( new_n47419_, new_n47145_, new_n662_ );
and  ( new_n47420_, new_n47419_, new_n47418_ );
nor  ( new_n47421_, new_n47420_, new_n47417_ );
and  ( new_n47422_, new_n47012_, new_n820_ );
and  ( new_n47423_, new_n47134_, new_n822_ );
or   ( new_n47424_, new_n47423_, new_n47422_ );
xor  ( new_n47425_, new_n47420_, new_n47417_ );
and  ( new_n47426_, new_n47425_, new_n47424_ );
nor  ( new_n47427_, new_n47426_, new_n47421_ );
not  ( new_n47428_, new_n47427_ );
xor  ( new_n47429_, new_n47413_, new_n47412_ );
and  ( new_n47430_, new_n47429_, new_n47428_ );
nor  ( new_n47431_, new_n47430_, new_n47414_ );
nand ( new_n47432_, new_n47289_, new_n47287_ );
nand ( new_n47433_, new_n47292_, new_n47290_ );
and  ( new_n47434_, new_n47433_, new_n47432_ );
xor  ( new_n47435_, new_n47434_, new_n47431_ );
xnor ( new_n47436_, new_n46998_, new_n46993_ );
xor  ( new_n47437_, new_n47436_, new_n47004_ );
xor  ( new_n47438_, new_n46894_, new_n46893_ );
or   ( new_n47439_, new_n47438_, new_n47437_ );
xor  ( new_n47440_, new_n46937_, new_n46932_ );
not  ( new_n47441_, new_n47440_ );
and  ( new_n47442_, new_n47441_, new_n46944_ );
and  ( new_n47443_, new_n46946_, new_n46939_ );
nor  ( new_n47444_, new_n47443_, new_n47442_ );
and  ( new_n47445_, new_n47438_, new_n47437_ );
or   ( new_n47446_, new_n47445_, new_n47444_ );
and  ( new_n47447_, new_n47446_, new_n47439_ );
xnor ( new_n47448_, new_n47447_, new_n47435_ );
or   ( new_n47449_, new_n47374_, new_n409_ );
or   ( new_n47450_, new_n47278_, new_n411_ );
nand ( new_n47451_, new_n47450_, new_n47449_ );
and  ( new_n47452_, new_n47451_, new_n47066_ );
and  ( new_n47453_, new_n47274_, new_n454_ );
xor  ( new_n47454_, new_n45403_, new_n400_ );
nor  ( new_n47455_, new_n47454_, new_n524_ );
or   ( new_n47456_, new_n47455_, new_n47453_ );
xor  ( new_n47457_, new_n47451_, new_n47066_ );
and  ( new_n47458_, new_n47457_, new_n47456_ );
or   ( new_n47459_, new_n47458_, new_n47452_ );
xor  ( new_n47460_, new_n47425_, new_n47424_ );
nand ( new_n47461_, new_n47460_, new_n47459_ );
xor  ( new_n47462_, new_n47460_, new_n47459_ );
xnor ( new_n47463_, new_n47213_, new_n47209_ );
nand ( new_n47464_, new_n47463_, new_n47218_ );
not  ( new_n47465_, new_n47219_ );
or   ( new_n47466_, new_n47465_, new_n47214_ );
and  ( new_n47467_, new_n47466_, new_n47464_ );
nand ( new_n47468_, new_n47467_, new_n47462_ );
and  ( new_n47469_, new_n47468_, new_n47461_ );
xnor ( new_n47470_, new_n47184_, new_n47181_ );
nand ( new_n47471_, new_n47470_, new_n47188_ );
not  ( new_n47472_, new_n47190_ );
or   ( new_n47473_, new_n47472_, new_n47185_ );
and  ( new_n47474_, new_n47473_, new_n47471_ );
xnor ( new_n47475_, new_n47197_, new_n47194_ );
xor  ( new_n47476_, new_n47475_, new_n47201_ );
nand ( new_n47477_, new_n47476_, new_n47474_ );
xor  ( new_n47478_, new_n47476_, new_n47474_ );
xnor ( new_n47479_, new_n47280_, new_n47276_ );
nand ( new_n47480_, new_n47479_, new_n47284_ );
not  ( new_n47481_, new_n47281_ );
nand ( new_n47482_, new_n47286_, new_n47481_ );
and  ( new_n47483_, new_n47482_, new_n47480_ );
nand ( new_n47484_, new_n47483_, new_n47478_ );
and  ( new_n47485_, new_n47484_, new_n47477_ );
or   ( new_n47486_, new_n47485_, new_n47469_ );
or   ( new_n47487_, new_n47210_, new_n340_ );
or   ( new_n47488_, new_n47384_, new_n337_ );
and  ( new_n47489_, new_n47488_, new_n47487_ );
xor  ( new_n47490_, new_n47303_, new_n43945_ );
not  ( new_n47491_, new_n47490_ );
or   ( new_n47492_, new_n47491_, new_n43983_ );
nor  ( new_n47493_, new_n46958_, new_n43880_ );
or   ( new_n47494_, new_n46959_, new_n43977_ );
or   ( new_n47495_, new_n47494_, new_n47493_ );
and  ( new_n47496_, new_n47495_, new_n47492_ );
nor  ( new_n47497_, new_n47496_, new_n47489_ );
and  ( new_n47498_, new_n47407_, new_n1739_ );
and  ( new_n47499_, new_n47363_, new_n1741_ );
nor  ( new_n47500_, new_n47499_, new_n47498_ );
xnor ( new_n47501_, new_n47496_, new_n47489_ );
nor  ( new_n47502_, new_n47501_, new_n47500_ );
or   ( new_n47503_, new_n47502_, new_n47497_ );
xor  ( new_n47504_, new_n47097_, new_n47096_ );
and  ( new_n47505_, new_n47504_, new_n47503_ );
xor  ( new_n47506_, new_n47504_, new_n47503_ );
xor  ( new_n47507_, new_n47410_, new_n47409_ );
and  ( new_n47508_, new_n47507_, new_n47506_ );
nor  ( new_n47509_, new_n47508_, new_n47505_ );
and  ( new_n47510_, new_n47485_, new_n47469_ );
or   ( new_n47511_, new_n47510_, new_n47509_ );
and  ( new_n47512_, new_n47511_, new_n47486_ );
nor  ( new_n47513_, new_n47512_, new_n47448_ );
xor  ( new_n47514_, new_n47429_, new_n47428_ );
xnor ( new_n47515_, new_n47204_, new_n47191_ );
xor  ( new_n47516_, new_n47515_, new_n47220_ );
and  ( new_n47517_, new_n47516_, new_n47514_ );
xnor ( new_n47518_, new_n47516_, new_n47514_ );
xnor ( new_n47519_, new_n47438_, new_n47437_ );
xor  ( new_n47520_, new_n47519_, new_n47444_ );
nor  ( new_n47521_, new_n47520_, new_n47518_ );
nor  ( new_n47522_, new_n47521_, new_n47517_ );
xnor ( new_n47523_, new_n47512_, new_n47448_ );
nor  ( new_n47524_, new_n47523_, new_n47522_ );
nor  ( new_n47525_, new_n47524_, new_n47513_ );
nor  ( new_n47526_, new_n47434_, new_n47431_ );
and  ( new_n47527_, new_n47447_, new_n47435_ );
nor  ( new_n47528_, new_n47527_, new_n47526_ );
and  ( new_n47529_, new_n46987_, new_n46976_ );
nor  ( new_n47530_, new_n46987_, new_n46976_ );
nor  ( new_n47531_, new_n47530_, new_n46948_ );
nor  ( new_n47532_, new_n47531_, new_n47529_ );
or   ( new_n47533_, new_n47024_, new_n47007_ );
and  ( new_n47534_, new_n47024_, new_n47007_ );
or   ( new_n47535_, new_n47041_, new_n47534_ );
and  ( new_n47536_, new_n47535_, new_n47533_ );
xor  ( new_n47537_, new_n47536_, new_n47532_ );
xor  ( new_n47538_, new_n46774_, new_n46770_ );
xor  ( new_n47539_, new_n47538_, new_n46780_ );
or   ( new_n47540_, new_n47255_, new_n47252_ );
and  ( new_n47541_, new_n47255_, new_n47252_ );
or   ( new_n47542_, new_n47541_, new_n47249_ );
and  ( new_n47543_, new_n47542_, new_n47540_ );
or   ( new_n47544_, new_n47234_, new_n47231_ );
and  ( new_n47545_, new_n47234_, new_n47231_ );
or   ( new_n47546_, new_n47545_, new_n47228_ );
and  ( new_n47547_, new_n47546_, new_n47544_ );
xor  ( new_n47548_, new_n47547_, new_n47543_ );
xor  ( new_n47549_, new_n47548_, new_n47539_ );
xnor ( new_n47550_, new_n47549_, new_n47537_ );
nand ( new_n47551_, new_n47042_, new_n46989_ );
nor  ( new_n47552_, new_n47042_, new_n46989_ );
or   ( new_n47553_, new_n47552_, new_n46927_ );
and  ( new_n47554_, new_n47553_, new_n47551_ );
xnor ( new_n47555_, new_n47554_, new_n47550_ );
xnor ( new_n47556_, new_n47555_, new_n47528_ );
and  ( new_n47557_, new_n47236_, new_n47225_ );
nor  ( new_n47558_, new_n47237_, new_n47222_ );
nor  ( new_n47559_, new_n47558_, new_n47557_ );
not  ( new_n47560_, new_n47559_ );
not  ( new_n47561_, new_n46723_ );
or   ( new_n47562_, new_n46985_, new_n3459_ );
and  ( new_n47563_, new_n46985_, new_n3459_ );
or   ( new_n47564_, new_n47563_, new_n46979_ );
and  ( new_n47565_, new_n47564_, new_n47562_ );
xor  ( new_n47566_, new_n47565_, new_n47561_ );
xor  ( new_n47567_, new_n46804_, new_n46803_ );
xor  ( new_n47568_, new_n47567_, new_n47566_ );
xor  ( new_n47569_, new_n46741_, new_n46737_ );
xor  ( new_n47570_, new_n47569_, new_n46746_ );
or   ( new_n47571_, new_n47244_, new_n47106_ );
and  ( new_n47572_, new_n47244_, new_n47106_ );
or   ( new_n47573_, new_n47572_, new_n47241_ );
and  ( new_n47574_, new_n47573_, new_n47571_ );
xor  ( new_n47575_, new_n47574_, new_n47570_ );
xor  ( new_n47576_, new_n47575_, new_n47568_ );
xnor ( new_n47577_, new_n46757_, new_n46753_ );
nand ( new_n47578_, new_n47577_, new_n46762_ );
not  ( new_n47579_, new_n46764_ );
or   ( new_n47580_, new_n47579_, new_n46758_ );
and  ( new_n47581_, new_n47580_, new_n47578_ );
xnor ( new_n47582_, new_n46814_, new_n46810_ );
xor  ( new_n47583_, new_n47582_, new_n46819_ );
xnor ( new_n47584_, new_n46832_, new_n46828_ );
xor  ( new_n47585_, new_n47584_, new_n46837_ );
xor  ( new_n47586_, new_n47585_, new_n47583_ );
xor  ( new_n47587_, new_n47586_, new_n47581_ );
xor  ( new_n47588_, new_n47587_, new_n47576_ );
xor  ( new_n47589_, new_n47588_, new_n47560_ );
not  ( new_n47590_, new_n47589_ );
or   ( new_n47591_, new_n47268_, new_n47238_ );
and  ( new_n47592_, new_n47268_, new_n47238_ );
or   ( new_n47593_, new_n47592_, new_n47178_ );
and  ( new_n47594_, new_n47593_, new_n47591_ );
and  ( new_n47595_, new_n46911_, new_n46897_ );
and  ( new_n47596_, new_n46926_, new_n46912_ );
nor  ( new_n47597_, new_n47596_, new_n47595_ );
or   ( new_n47598_, new_n46909_, new_n46905_ );
and  ( new_n47599_, new_n46909_, new_n46905_ );
or   ( new_n47600_, new_n47599_, new_n46901_ );
and  ( new_n47601_, new_n47600_, new_n47598_ );
or   ( new_n47602_, new_n46924_, new_n46920_ );
and  ( new_n47603_, new_n46924_, new_n46920_ );
or   ( new_n47604_, new_n47603_, new_n46916_ );
and  ( new_n47605_, new_n47604_, new_n47602_ );
xor  ( new_n47606_, new_n47605_, new_n47601_ );
or   ( new_n47607_, new_n47265_, new_n47262_ );
and  ( new_n47608_, new_n47265_, new_n47262_ );
or   ( new_n47609_, new_n47608_, new_n47261_ );
and  ( new_n47610_, new_n47609_, new_n47607_ );
xor  ( new_n47611_, new_n47610_, new_n47606_ );
nand ( new_n47612_, new_n47257_, new_n47246_ );
nor  ( new_n47613_, new_n47257_, new_n47246_ );
or   ( new_n47614_, new_n47267_, new_n47613_ );
and  ( new_n47615_, new_n47614_, new_n47612_ );
xor  ( new_n47616_, new_n47615_, new_n47611_ );
xor  ( new_n47617_, new_n47616_, new_n47597_ );
xor  ( new_n47618_, new_n47617_, new_n47594_ );
xor  ( new_n47619_, new_n47618_, new_n47590_ );
xor  ( new_n47620_, new_n47619_, new_n47556_ );
xor  ( new_n47621_, new_n47620_, new_n47525_ );
nor  ( new_n47622_, new_n47621_, new_n47401_ );
nand ( new_n47623_, new_n47621_, new_n47401_ );
xnor ( new_n47624_, new_n47523_, new_n47522_ );
xor  ( new_n47625_, new_n47396_, new_n47395_ );
xnor ( new_n47626_, new_n47485_, new_n47469_ );
xor  ( new_n47627_, new_n47626_, new_n47509_ );
nand ( new_n47628_, new_n47627_, new_n47625_ );
nor  ( new_n47629_, new_n47627_, new_n47625_ );
xnor ( new_n47630_, new_n47333_, new_n47332_ );
xor  ( new_n47631_, RIbb328b0_169, RIbb2c550_105 );
and  ( new_n47632_, new_n46412_, new_n43561_ );
nor  ( new_n47633_, new_n47632_, new_n43643_ );
not  ( new_n47634_, new_n47633_ );
and  ( new_n47635_, new_n47634_, new_n43564_ );
nor  ( new_n47636_, new_n47635_, new_n43642_ );
not  ( new_n47637_, new_n47636_ );
and  ( new_n47638_, new_n47637_, new_n43566_ );
nor  ( new_n47639_, new_n47638_, new_n43641_ );
xnor ( new_n47640_, new_n47639_, new_n47631_ );
and  ( new_n47641_, new_n47640_, new_n43880_ );
not  ( new_n47642_, new_n47641_ );
or   ( new_n47643_, new_n47490_, new_n44007_ );
or   ( new_n47644_, new_n47312_, new_n302_ );
and  ( new_n47645_, new_n47644_, new_n47643_ );
nor  ( new_n47646_, new_n47645_, new_n47642_ );
xor  ( new_n47647_, new_n44183_, RIbb2e9e0_27 );
and  ( new_n47648_, new_n47647_, new_n2002_ );
and  ( new_n47649_, new_n47377_, new_n2000_ );
or   ( new_n47650_, new_n47649_, new_n47648_ );
xor  ( new_n47651_, new_n47645_, new_n47642_ );
and  ( new_n47652_, new_n47651_, new_n47650_ );
or   ( new_n47653_, new_n47652_, new_n47646_ );
xor  ( new_n47654_, new_n47326_, new_n4295_ );
xor  ( new_n47655_, new_n47654_, new_n47322_ );
nand ( new_n47656_, new_n47655_, new_n47653_ );
nor  ( new_n47657_, new_n47655_, new_n47653_ );
xnor ( new_n47658_, new_n47316_, new_n47315_ );
or   ( new_n47659_, new_n47658_, new_n47657_ );
and  ( new_n47660_, new_n47659_, new_n47656_ );
nor  ( new_n47661_, new_n47660_, new_n47630_ );
or   ( new_n47662_, new_n47359_, new_n3463_ );
xor  ( new_n47663_, new_n43884_, new_n3113_ );
or   ( new_n47664_, new_n47663_, new_n3461_ );
and  ( new_n47665_, new_n47664_, new_n47662_ );
nand ( new_n47666_, new_n47348_, new_n1474_ );
xor  ( new_n47667_, new_n44506_, new_n1355_ );
or   ( new_n47668_, new_n47667_, new_n1593_ );
and  ( new_n47669_, new_n47668_, new_n47666_ );
or   ( new_n47670_, new_n47669_, new_n47665_ );
and  ( new_n47671_, new_n47365_, new_n1739_ );
xor  ( new_n47672_, new_n44319_, RIbb2ead0_25 );
and  ( new_n47673_, new_n47672_, new_n1741_ );
or   ( new_n47674_, new_n47673_, new_n47671_ );
xor  ( new_n47675_, new_n47669_, new_n47665_ );
nand ( new_n47676_, new_n47675_, new_n47674_ );
and  ( new_n47677_, new_n47676_, new_n47670_ );
nand ( new_n47678_, new_n47339_, new_n2928_ );
xor  ( new_n47679_, new_n43937_, RIbb2e710_33 );
nand ( new_n47680_, new_n47679_, new_n2930_ );
and  ( new_n47681_, new_n47680_, new_n47678_ );
xor  ( new_n47682_, new_n44681_, RIbb2ecb0_21 );
nand ( new_n47683_, new_n47682_, new_n1253_ );
or   ( new_n47684_, new_n47343_, new_n1366_ );
and  ( new_n47685_, new_n47684_, new_n47683_ );
or   ( new_n47686_, new_n47685_, new_n47681_ );
xor  ( new_n47687_, new_n43894_, RIbb2e530_37 );
and  ( new_n47688_, new_n47687_, new_n3731_ );
xor  ( new_n47689_, new_n43799_, new_n3457_ );
nor  ( new_n47690_, new_n47689_, new_n3896_ );
nor  ( new_n47691_, new_n47690_, new_n47688_ );
and  ( new_n47692_, new_n47685_, new_n47681_ );
or   ( new_n47693_, new_n47692_, new_n47691_ );
and  ( new_n47694_, new_n47693_, new_n47686_ );
nor  ( new_n47695_, new_n47694_, new_n47677_ );
or   ( new_n47696_, new_n47354_, new_n4304_ );
xor  ( new_n47697_, new_n43898_, new_n3892_ );
or   ( new_n47698_, new_n47697_, new_n4302_ );
and  ( new_n47699_, new_n47698_, new_n47696_ );
or   ( new_n47700_, new_n47382_, new_n340_ );
xor  ( new_n47701_, new_n46137_, RIbb2f250_9 );
nand ( new_n47702_, new_n47701_, new_n336_ );
and  ( new_n47703_, new_n47702_, new_n47700_ );
nor  ( new_n47704_, new_n47703_, new_n47699_ );
and  ( new_n47705_, new_n47372_, new_n371_ );
xor  ( new_n47706_, new_n45928_, new_n325_ );
nor  ( new_n47707_, new_n47706_, new_n409_ );
nor  ( new_n47708_, new_n47707_, new_n47705_ );
xnor ( new_n47709_, new_n47703_, new_n47699_ );
nor  ( new_n47710_, new_n47709_, new_n47708_ );
or   ( new_n47711_, new_n47710_, new_n47704_ );
xor  ( new_n47712_, new_n47694_, new_n47677_ );
and  ( new_n47713_, new_n47712_, new_n47711_ );
or   ( new_n47714_, new_n47713_, new_n47695_ );
xor  ( new_n47715_, new_n47660_, new_n47630_ );
and  ( new_n47716_, new_n47715_, new_n47714_ );
or   ( new_n47717_, new_n47716_, new_n47661_ );
xor  ( new_n47718_, new_n47483_, new_n47478_ );
nand ( new_n47719_, new_n47718_, new_n47717_ );
xor  ( new_n47720_, new_n47718_, new_n47717_ );
xor  ( new_n47721_, new_n47393_, new_n47392_ );
nand ( new_n47722_, new_n47721_, new_n47720_ );
and  ( new_n47723_, new_n47722_, new_n47719_ );
or   ( new_n47724_, new_n47723_, new_n47629_ );
and  ( new_n47725_, new_n47724_, new_n47628_ );
nor  ( new_n47726_, new_n47725_, new_n47624_ );
or   ( new_n47727_, new_n47070_, new_n2427_ );
xor  ( new_n47728_, new_n43985_, new_n2118_ );
or   ( new_n47729_, new_n47728_, new_n2425_ );
and  ( new_n47730_, new_n47729_, new_n47727_ );
or   ( new_n47731_, new_n47147_, new_n757_ );
xor  ( new_n47732_, new_n45204_, RIbb2ef80_15 );
nand ( new_n47733_, new_n47732_, new_n662_ );
and  ( new_n47734_, new_n47733_, new_n47731_ );
or   ( new_n47735_, new_n47734_, new_n47730_ );
and  ( new_n47736_, new_n47136_, new_n820_ );
xor  ( new_n47737_, new_n44974_, RIbb2ee90_17 );
and  ( new_n47738_, new_n47737_, new_n822_ );
or   ( new_n47739_, new_n47738_, new_n47736_ );
xor  ( new_n47740_, new_n47734_, new_n47730_ );
nand ( new_n47741_, new_n47740_, new_n47739_ );
and  ( new_n47742_, new_n47741_, new_n47735_ );
or   ( new_n47743_, new_n47117_, new_n2809_ );
xor  ( new_n47744_, new_n43956_, new_n2421_ );
or   ( new_n47745_, new_n47744_, new_n2807_ );
and  ( new_n47746_, new_n47745_, new_n47743_ );
or   ( new_n47747_, new_n47075_, new_n1137_ );
xor  ( new_n47748_, new_n44785_, new_n893_ );
or   ( new_n47749_, new_n47748_, new_n1135_ );
and  ( new_n47750_, new_n47749_, new_n47747_ );
or   ( new_n47751_, new_n47750_, new_n47746_ );
and  ( new_n47752_, new_n47687_, new_n3733_ );
nor  ( new_n47753_, new_n47157_, new_n3898_ );
or   ( new_n47754_, new_n47753_, new_n47752_ );
xor  ( new_n47755_, new_n47750_, new_n47746_ );
nand ( new_n47756_, new_n47755_, new_n47754_ );
and  ( new_n47757_, new_n47756_, new_n47751_ );
nor  ( new_n47758_, new_n47757_, new_n47742_ );
xor  ( new_n47759_, new_n47757_, new_n47742_ );
xor  ( new_n47760_, new_n47457_, new_n47456_ );
and  ( new_n47761_, new_n47760_, new_n47759_ );
or   ( new_n47762_, new_n47761_, new_n47758_ );
xor  ( new_n47763_, new_n47507_, new_n47506_ );
nand ( new_n47764_, new_n47763_, new_n47762_ );
xor  ( new_n47765_, new_n47763_, new_n47762_ );
xor  ( new_n47766_, new_n47173_, new_n47154_ );
nand ( new_n47767_, new_n47766_, new_n47765_ );
and  ( new_n47768_, new_n47767_, new_n47764_ );
xor  ( new_n47769_, new_n47131_, new_n47130_ );
xnor ( new_n47770_, new_n47077_, new_n47072_ );
nand ( new_n47771_, new_n47770_, new_n47083_ );
not  ( new_n47772_, new_n47078_ );
nand ( new_n47773_, new_n47085_, new_n47772_ );
and  ( new_n47774_, new_n47773_, new_n47771_ );
nor  ( new_n47775_, new_n47774_, new_n47769_ );
nand ( new_n47776_, new_n47774_, new_n47769_ );
xnor ( new_n47777_, new_n47501_, new_n47500_ );
and  ( new_n47778_, new_n47777_, new_n47776_ );
or   ( new_n47779_, new_n47778_, new_n47775_ );
xor  ( new_n47780_, new_n47150_, new_n47149_ );
xnor ( new_n47781_, new_n47164_, new_n47159_ );
nand ( new_n47782_, new_n47781_, new_n47171_ );
not  ( new_n47783_, new_n47172_ );
or   ( new_n47784_, new_n47783_, new_n47165_ );
and  ( new_n47785_, new_n47784_, new_n47782_ );
nand ( new_n47786_, new_n47785_, new_n47780_ );
nor  ( new_n47787_, new_n47785_, new_n47780_ );
or   ( new_n47788_, new_n47454_, new_n526_ );
xor  ( new_n47789_, new_n45584_, new_n400_ );
or   ( new_n47790_, new_n47789_, new_n524_ );
and  ( new_n47791_, new_n47790_, new_n47788_ );
nor  ( new_n47792_, RIbb2e260_43, RIbb2e2d8_42 );
not  ( new_n47793_, new_n47792_ );
and  ( new_n47794_, new_n47793_, new_n4294_ );
xor  ( new_n47795_, new_n43793_, new_n4292_ );
and  ( new_n47796_, new_n47795_, new_n4543_ );
nor  ( new_n47797_, new_n47796_, new_n47794_ );
or   ( new_n47798_, new_n47797_, new_n47791_ );
or   ( new_n47799_, new_n47320_, new_n286_ );
xor  ( new_n47800_, new_n46962_, new_n275_ );
or   ( new_n47801_, new_n47800_, new_n283_ );
and  ( new_n47802_, new_n47801_, new_n47799_ );
or   ( new_n47803_, new_n47324_, new_n320_ );
xor  ( new_n47804_, new_n46619_, new_n309_ );
or   ( new_n47805_, new_n47804_, new_n317_ );
and  ( new_n47806_, new_n47805_, new_n47803_ );
nor  ( new_n47807_, new_n47806_, new_n47802_ );
nand ( new_n47808_, new_n47806_, new_n47802_ );
xor  ( new_n47809_, new_n47296_, new_n43945_ );
and  ( new_n47810_, new_n47809_, new_n43982_ );
or   ( new_n47811_, new_n47046_, new_n43880_ );
and  ( new_n47812_, new_n47047_, new_n43978_ );
and  ( new_n47813_, new_n47812_, new_n47811_ );
or   ( new_n47814_, new_n47813_, new_n47810_ );
and  ( new_n47815_, new_n47814_, new_n47808_ );
or   ( new_n47816_, new_n47815_, new_n47807_ );
xor  ( new_n47817_, new_n47797_, new_n47791_ );
nand ( new_n47818_, new_n47817_, new_n47816_ );
and  ( new_n47819_, new_n47818_, new_n47798_ );
or   ( new_n47820_, new_n47819_, new_n47787_ );
and  ( new_n47821_, new_n47820_, new_n47786_ );
or   ( new_n47822_, new_n47821_, new_n47779_ );
xor  ( new_n47823_, new_n47467_, new_n47462_ );
xor  ( new_n47824_, new_n47821_, new_n47779_ );
nand ( new_n47825_, new_n47824_, new_n47823_ );
and  ( new_n47826_, new_n47825_, new_n47822_ );
nand ( new_n47827_, new_n47826_, new_n47768_ );
nor  ( new_n47828_, new_n47826_, new_n47768_ );
xor  ( new_n47829_, new_n47520_, new_n47518_ );
or   ( new_n47830_, new_n47829_, new_n47828_ );
and  ( new_n47831_, new_n47830_, new_n47827_ );
nand ( new_n47832_, new_n47725_, new_n47624_ );
and  ( new_n47833_, new_n47832_, new_n47831_ );
or   ( new_n47834_, new_n47833_, new_n47726_ );
and  ( new_n47835_, new_n47834_, new_n47623_ );
or   ( new_n47836_, new_n47835_, new_n47622_ );
nor  ( new_n47837_, new_n47619_, new_n47556_ );
and  ( new_n47838_, new_n47619_, new_n47556_ );
nor  ( new_n47839_, new_n47838_, new_n47525_ );
nor  ( new_n47840_, new_n47839_, new_n47837_ );
and  ( new_n47841_, new_n47587_, new_n47576_ );
and  ( new_n47842_, new_n47588_, new_n47560_ );
or   ( new_n47843_, new_n47842_, new_n47841_ );
xor  ( new_n47844_, new_n46731_, new_n46729_ );
not  ( new_n47845_, new_n47844_ );
xnor ( new_n47846_, new_n46572_, new_n46568_ );
nand ( new_n47847_, new_n47846_, new_n46577_ );
not  ( new_n47848_, new_n46579_ );
or   ( new_n47849_, new_n47848_, new_n46573_ );
and  ( new_n47850_, new_n47849_, new_n47847_ );
xnor ( new_n47851_, new_n46588_, new_n46584_ );
nand ( new_n47852_, new_n47851_, new_n46593_ );
not  ( new_n47853_, new_n46595_ );
or   ( new_n47854_, new_n47853_, new_n46589_ );
and  ( new_n47855_, new_n47854_, new_n47852_ );
xor  ( new_n47856_, new_n47855_, new_n47850_ );
xor  ( new_n47857_, new_n47856_, new_n47845_ );
xnor ( new_n47858_, new_n46858_, new_n46856_ );
or   ( new_n47859_, new_n47574_, new_n47570_ );
nand ( new_n47860_, new_n47574_, new_n47570_ );
nand ( new_n47861_, new_n47860_, new_n47568_ );
and  ( new_n47862_, new_n47861_, new_n47859_ );
xnor ( new_n47863_, new_n47862_, new_n47858_ );
xor  ( new_n47864_, new_n47863_, new_n47857_ );
xor  ( new_n47865_, new_n46840_, new_n46825_ );
xor  ( new_n47866_, new_n46784_, new_n46783_ );
or   ( new_n47867_, new_n47585_, new_n47583_ );
and  ( new_n47868_, new_n47585_, new_n47583_ );
or   ( new_n47869_, new_n47868_, new_n47581_ );
and  ( new_n47870_, new_n47869_, new_n47867_ );
xor  ( new_n47871_, new_n47870_, new_n47866_ );
xor  ( new_n47872_, new_n47871_, new_n47865_ );
xor  ( new_n47873_, new_n47872_, new_n47864_ );
xor  ( new_n47874_, new_n47873_, new_n47843_ );
nor  ( new_n47875_, new_n47617_, new_n47594_ );
and  ( new_n47876_, new_n47617_, new_n47594_ );
nor  ( new_n47877_, new_n47876_, new_n47590_ );
nor  ( new_n47878_, new_n47877_, new_n47875_ );
nor  ( new_n47879_, new_n47554_, new_n47550_ );
nor  ( new_n47880_, new_n47555_, new_n47528_ );
or   ( new_n47881_, new_n47880_, new_n47879_ );
nor  ( new_n47882_, new_n47615_, new_n47611_ );
and  ( new_n47883_, new_n47615_, new_n47611_ );
nor  ( new_n47884_, new_n47883_, new_n47597_ );
nor  ( new_n47885_, new_n47884_, new_n47882_ );
nor  ( new_n47886_, new_n47536_, new_n47532_ );
and  ( new_n47887_, new_n47549_, new_n47537_ );
or   ( new_n47888_, new_n47887_, new_n47886_ );
nor  ( new_n47889_, new_n47605_, new_n47601_ );
and  ( new_n47890_, new_n47605_, new_n47601_ );
nor  ( new_n47891_, new_n47610_, new_n47890_ );
nor  ( new_n47892_, new_n47891_, new_n47889_ );
nor  ( new_n47893_, new_n47565_, new_n47561_ );
and  ( new_n47894_, new_n47567_, new_n47566_ );
nor  ( new_n47895_, new_n47894_, new_n47893_ );
nor  ( new_n47896_, new_n47547_, new_n47543_ );
and  ( new_n47897_, new_n47547_, new_n47543_ );
not  ( new_n47898_, new_n47897_ );
and  ( new_n47899_, new_n47898_, new_n47539_ );
nor  ( new_n47900_, new_n47899_, new_n47896_ );
xnor ( new_n47901_, new_n47900_, new_n47895_ );
nand ( new_n47902_, new_n47901_, new_n47892_ );
nor  ( new_n47903_, new_n47900_, new_n47895_ );
and  ( new_n47904_, new_n47900_, new_n47895_ );
nor  ( new_n47905_, new_n47904_, new_n47892_ );
not  ( new_n47906_, new_n47905_ );
or   ( new_n47907_, new_n47906_, new_n47903_ );
and  ( new_n47908_, new_n47907_, new_n47902_ );
xnor ( new_n47909_, new_n47908_, new_n47888_ );
xor  ( new_n47910_, new_n47909_, new_n47885_ );
xnor ( new_n47911_, new_n47910_, new_n47881_ );
xor  ( new_n47912_, new_n47911_, new_n47878_ );
xnor ( new_n47913_, new_n47912_, new_n47874_ );
xor  ( new_n47914_, new_n47913_, new_n47840_ );
nor  ( new_n47915_, new_n47914_, new_n47836_ );
xor  ( new_n47916_, new_n47399_, new_n47398_ );
xor  ( new_n47917_, new_n47725_, new_n47624_ );
xor  ( new_n47918_, new_n47917_, new_n47831_ );
or   ( new_n47919_, new_n47918_, new_n47916_ );
nand ( new_n47920_, new_n47918_, new_n47916_ );
xnor ( new_n47921_, new_n47387_, new_n47386_ );
xor  ( new_n47922_, new_n43952_, new_n2421_ );
or   ( new_n47923_, new_n47922_, new_n2807_ );
or   ( new_n47924_, new_n47744_, new_n2809_ );
and  ( new_n47925_, new_n47924_, new_n47923_ );
xor  ( new_n47926_, new_n44877_, new_n893_ );
or   ( new_n47927_, new_n47926_, new_n1135_ );
or   ( new_n47928_, new_n47748_, new_n1137_ );
and  ( new_n47929_, new_n47928_, new_n47927_ );
or   ( new_n47930_, new_n47929_, new_n47925_ );
xor  ( new_n47931_, new_n45119_, new_n745_ );
nor  ( new_n47932_, new_n47931_, new_n897_ );
and  ( new_n47933_, new_n47737_, new_n820_ );
nor  ( new_n47934_, new_n47933_, new_n47932_ );
and  ( new_n47935_, new_n47929_, new_n47925_ );
or   ( new_n47936_, new_n47935_, new_n47934_ );
and  ( new_n47937_, new_n47936_, new_n47930_ );
nor  ( new_n47938_, new_n47937_, new_n47921_ );
nand ( new_n47939_, new_n47937_, new_n47921_ );
xor  ( new_n47940_, new_n45738_, RIbb2f070_13 );
nand ( new_n47941_, new_n47940_, new_n456_ );
or   ( new_n47942_, new_n47789_, new_n526_ );
and  ( new_n47943_, new_n47942_, new_n47941_ );
or   ( new_n47944_, new_n47728_, new_n2427_ );
xor  ( new_n47945_, new_n43812_, new_n2118_ );
or   ( new_n47946_, new_n47945_, new_n2425_ );
and  ( new_n47947_, new_n47946_, new_n47944_ );
nor  ( new_n47948_, new_n47947_, new_n47943_ );
xor  ( new_n47949_, new_n45403_, new_n520_ );
nor  ( new_n47950_, new_n47949_, new_n755_ );
and  ( new_n47951_, new_n47732_, new_n660_ );
or   ( new_n47952_, new_n47951_, new_n47950_ );
nand ( new_n47953_, new_n47947_, new_n47943_ );
and  ( new_n47954_, new_n47953_, new_n47952_ );
or   ( new_n47955_, new_n47954_, new_n47948_ );
and  ( new_n47956_, new_n47955_, new_n47939_ );
or   ( new_n47957_, new_n47956_, new_n47938_ );
xor  ( new_n47958_, new_n47755_, new_n47754_ );
xor  ( new_n47959_, new_n47368_, new_n47367_ );
or   ( new_n47960_, new_n47959_, new_n47958_ );
and  ( new_n47961_, new_n47959_, new_n47958_ );
xor  ( new_n47962_, new_n47345_, new_n47341_ );
not  ( new_n47963_, new_n47962_ );
and  ( new_n47964_, new_n47963_, new_n47350_ );
not  ( new_n47965_, new_n47346_ );
and  ( new_n47966_, new_n47352_, new_n47965_ );
nor  ( new_n47967_, new_n47966_, new_n47964_ );
or   ( new_n47968_, new_n47967_, new_n47961_ );
and  ( new_n47969_, new_n47968_, new_n47960_ );
and  ( new_n47970_, new_n47969_, new_n47957_ );
xor  ( new_n47971_, new_n47760_, new_n47759_ );
xor  ( new_n47972_, new_n47969_, new_n47957_ );
and  ( new_n47973_, new_n47972_, new_n47971_ );
or   ( new_n47974_, new_n47973_, new_n47970_ );
xor  ( new_n47975_, new_n47766_, new_n47765_ );
and  ( new_n47976_, new_n47975_, new_n47974_ );
xor  ( new_n47977_, new_n47740_, new_n47739_ );
xor  ( new_n47978_, new_n47817_, new_n47816_ );
and  ( new_n47979_, new_n47978_, new_n47977_ );
and  ( new_n47980_, new_n47300_, new_n43949_ );
and  ( new_n47981_, new_n47491_, new_n295_ );
nor  ( new_n47982_, new_n47981_, new_n47980_ );
xor  ( new_n47983_, new_n47640_, new_n43945_ );
not  ( new_n47984_, new_n47983_ );
or   ( new_n47985_, new_n47984_, new_n43983_ );
not  ( new_n47986_, new_n47296_ );
and  ( new_n47987_, new_n47986_, new_n43879_ );
or   ( new_n47988_, new_n47297_, new_n43977_ );
or   ( new_n47989_, new_n47988_, new_n47987_ );
and  ( new_n47990_, new_n47989_, new_n47985_ );
nor  ( new_n47991_, new_n47990_, new_n47982_ );
and  ( new_n47992_, new_n47990_, new_n47982_ );
nor  ( new_n47993_, new_n47800_, new_n286_ );
xor  ( new_n47994_, new_n46958_, RIbb2f430_5 );
and  ( new_n47995_, new_n47994_, new_n282_ );
nor  ( new_n47996_, new_n47995_, new_n47993_ );
nor  ( new_n47997_, new_n47996_, new_n47992_ );
or   ( new_n47998_, new_n47997_, new_n47991_ );
and  ( new_n47999_, new_n47998_, new_n47797_ );
or   ( new_n48000_, new_n47804_, new_n320_ );
xor  ( new_n48001_, new_n46789_, new_n309_ );
or   ( new_n48002_, new_n48001_, new_n317_ );
and  ( new_n48003_, new_n48002_, new_n48000_ );
nor  ( new_n48004_, new_n48003_, new_n4707_ );
and  ( new_n48005_, new_n47701_, new_n334_ );
xor  ( new_n48006_, new_n46427_, RIbb2f250_9 );
and  ( new_n48007_, new_n48006_, new_n336_ );
nor  ( new_n48008_, new_n48007_, new_n48005_ );
xor  ( new_n48009_, new_n48003_, new_n4708_ );
nor  ( new_n48010_, new_n48009_, new_n48008_ );
or   ( new_n48011_, new_n48010_, new_n48004_ );
xor  ( new_n48012_, new_n47998_, new_n47797_ );
and  ( new_n48013_, new_n48012_, new_n48011_ );
or   ( new_n48014_, new_n48013_, new_n47999_ );
xor  ( new_n48015_, new_n47978_, new_n47977_ );
and  ( new_n48016_, new_n48015_, new_n48014_ );
nor  ( new_n48017_, new_n48016_, new_n47979_ );
xnor ( new_n48018_, new_n47390_, new_n47389_ );
nor  ( new_n48019_, new_n48018_, new_n48017_ );
xnor ( new_n48020_, new_n48018_, new_n48017_ );
xor  ( new_n48021_, new_n47785_, new_n47780_ );
xor  ( new_n48022_, new_n48021_, new_n47819_ );
nor  ( new_n48023_, new_n48022_, new_n48020_ );
or   ( new_n48024_, new_n48023_, new_n48019_ );
xor  ( new_n48025_, new_n47975_, new_n47974_ );
and  ( new_n48026_, new_n48025_, new_n48024_ );
or   ( new_n48027_, new_n48026_, new_n47976_ );
xor  ( new_n48028_, new_n47826_, new_n47768_ );
xor  ( new_n48029_, new_n48028_, new_n47829_ );
and  ( new_n48030_, new_n48029_, new_n48027_ );
xor  ( new_n48031_, new_n47774_, new_n47769_ );
xor  ( new_n48032_, new_n48031_, new_n47777_ );
xor  ( new_n48033_, new_n47651_, new_n47650_ );
xor  ( new_n48034_, new_n47806_, new_n47802_ );
xor  ( new_n48035_, new_n48034_, new_n47814_ );
nand ( new_n48036_, new_n48035_, new_n48033_ );
nor  ( new_n48037_, new_n48035_, new_n48033_ );
xor  ( new_n48038_, RIbb32928_170, RIbb2c4d8_106 );
xor  ( new_n48039_, new_n48038_, new_n47637_ );
not  ( new_n48040_, new_n48039_ );
or   ( new_n48041_, new_n48040_, new_n43879_ );
xor  ( new_n48042_, new_n43914_, new_n2118_ );
or   ( new_n48043_, new_n48042_, new_n2425_ );
or   ( new_n48044_, new_n47945_, new_n2427_ );
and  ( new_n48045_, new_n48044_, new_n48043_ );
nor  ( new_n48046_, new_n48045_, new_n48041_ );
and  ( new_n48047_, new_n48045_, new_n48041_ );
xor  ( new_n48048_, new_n45597_, RIbb2f070_13 );
and  ( new_n48049_, new_n48048_, new_n456_ );
and  ( new_n48050_, new_n47940_, new_n454_ );
nor  ( new_n48051_, new_n48050_, new_n48049_ );
nor  ( new_n48052_, new_n48051_, new_n48047_ );
nor  ( new_n48053_, new_n48052_, new_n48046_ );
or   ( new_n48054_, new_n48053_, new_n48037_ );
and  ( new_n48055_, new_n48054_, new_n48036_ );
xor  ( new_n48056_, new_n43956_, new_n2797_ );
nor  ( new_n48057_, new_n48056_, new_n3117_ );
and  ( new_n48058_, new_n47679_, new_n2928_ );
nor  ( new_n48059_, new_n48058_, new_n48057_ );
xor  ( new_n48060_, new_n44600_, RIbb2ebc0_23 );
nand ( new_n48061_, new_n48060_, new_n1476_ );
or   ( new_n48062_, new_n47667_, new_n1595_ );
and  ( new_n48063_, new_n48062_, new_n48061_ );
nor  ( new_n48064_, new_n48063_, new_n48059_ );
xor  ( new_n48065_, new_n43894_, RIbb2e440_39 );
and  ( new_n48066_, new_n48065_, new_n4034_ );
nor  ( new_n48067_, new_n47697_, new_n4304_ );
nor  ( new_n48068_, new_n48067_, new_n48066_ );
and  ( new_n48069_, new_n48063_, new_n48059_ );
nor  ( new_n48070_, new_n48069_, new_n48068_ );
nor  ( new_n48071_, new_n48070_, new_n48064_ );
or   ( new_n48072_, new_n47663_, new_n3463_ );
xor  ( new_n48073_, new_n43888_, new_n3113_ );
or   ( new_n48074_, new_n48073_, new_n3461_ );
and  ( new_n48075_, new_n48074_, new_n48072_ );
or   ( new_n48076_, new_n47689_, new_n3898_ );
xor  ( new_n48077_, new_n43803_, new_n3457_ );
or   ( new_n48078_, new_n48077_, new_n3896_ );
and  ( new_n48079_, new_n48078_, new_n48076_ );
nor  ( new_n48080_, new_n48079_, new_n48075_ );
xor  ( new_n48081_, new_n44407_, RIbb2ead0_25 );
and  ( new_n48082_, new_n48081_, new_n1741_ );
and  ( new_n48083_, new_n47672_, new_n1739_ );
nor  ( new_n48084_, new_n48083_, new_n48082_ );
and  ( new_n48085_, new_n48079_, new_n48075_ );
nor  ( new_n48086_, new_n48085_, new_n48084_ );
nor  ( new_n48087_, new_n48086_, new_n48080_ );
or   ( new_n48088_, new_n48087_, new_n48071_ );
and  ( new_n48089_, new_n48087_, new_n48071_ );
xor  ( new_n48090_, new_n46037_, new_n325_ );
or   ( new_n48091_, new_n48090_, new_n409_ );
or   ( new_n48092_, new_n47706_, new_n411_ );
and  ( new_n48093_, new_n48092_, new_n48091_ );
xor  ( new_n48094_, new_n43787_, new_n4292_ );
or   ( new_n48095_, new_n48094_, new_n4709_ );
nand ( new_n48096_, new_n47795_, new_n4541_ );
and  ( new_n48097_, new_n48096_, new_n48095_ );
nor  ( new_n48098_, new_n48097_, new_n48093_ );
and  ( new_n48099_, new_n47647_, new_n2000_ );
xor  ( new_n48100_, new_n44218_, RIbb2e9e0_27 );
and  ( new_n48101_, new_n48100_, new_n2002_ );
nor  ( new_n48102_, new_n48101_, new_n48099_ );
and  ( new_n48103_, new_n48097_, new_n48093_ );
nor  ( new_n48104_, new_n48103_, new_n48102_ );
nor  ( new_n48105_, new_n48104_, new_n48098_ );
or   ( new_n48106_, new_n48105_, new_n48089_ );
and  ( new_n48107_, new_n48106_, new_n48088_ );
or   ( new_n48108_, new_n48107_, new_n48055_ );
and  ( new_n48109_, new_n48107_, new_n48055_ );
xor  ( new_n48110_, new_n46619_, new_n329_ );
nor  ( new_n48111_, new_n48110_, new_n337_ );
and  ( new_n48112_, new_n48006_, new_n334_ );
nor  ( new_n48113_, new_n48112_, new_n48111_ );
or   ( new_n48114_, new_n47931_, new_n899_ );
xor  ( new_n48115_, new_n45204_, RIbb2ee90_17 );
nand ( new_n48116_, new_n48115_, new_n822_ );
and  ( new_n48117_, new_n48116_, new_n48114_ );
nor  ( new_n48118_, new_n48117_, new_n48113_ );
xor  ( new_n48119_, new_n45584_, RIbb2ef80_15 );
and  ( new_n48120_, new_n48119_, new_n662_ );
nor  ( new_n48121_, new_n47949_, new_n757_ );
or   ( new_n48122_, new_n48121_, new_n48120_ );
xor  ( new_n48123_, new_n48117_, new_n48113_ );
and  ( new_n48124_, new_n48123_, new_n48122_ );
or   ( new_n48125_, new_n48124_, new_n48118_ );
xor  ( new_n48126_, new_n47675_, new_n47674_ );
and  ( new_n48127_, new_n48126_, new_n48125_ );
nor  ( new_n48128_, new_n48126_, new_n48125_ );
not  ( new_n48129_, new_n48128_ );
xor  ( new_n48130_, new_n47929_, new_n47925_ );
xnor ( new_n48131_, new_n48130_, new_n47934_ );
and  ( new_n48132_, new_n48131_, new_n48129_ );
nor  ( new_n48133_, new_n48132_, new_n48127_ );
or   ( new_n48134_, new_n48133_, new_n48109_ );
and  ( new_n48135_, new_n48134_, new_n48108_ );
nor  ( new_n48136_, new_n48135_, new_n48032_ );
xor  ( new_n48137_, new_n47715_, new_n47714_ );
xor  ( new_n48138_, new_n48135_, new_n48032_ );
and  ( new_n48139_, new_n48138_, new_n48137_ );
or   ( new_n48140_, new_n48139_, new_n48136_ );
xor  ( new_n48141_, new_n47824_, new_n47823_ );
and  ( new_n48142_, new_n48141_, new_n48140_ );
xor  ( new_n48143_, new_n48141_, new_n48140_ );
xor  ( new_n48144_, new_n47721_, new_n47720_ );
and  ( new_n48145_, new_n48144_, new_n48143_ );
nor  ( new_n48146_, new_n48145_, new_n48142_ );
not  ( new_n48147_, new_n48146_ );
xor  ( new_n48148_, new_n48029_, new_n48027_ );
and  ( new_n48149_, new_n48148_, new_n48147_ );
nor  ( new_n48150_, new_n48149_, new_n48030_ );
nand ( new_n48151_, new_n48150_, new_n47920_ );
and  ( new_n48152_, new_n48151_, new_n47919_ );
xor  ( new_n48153_, new_n47621_, new_n47401_ );
xor  ( new_n48154_, new_n48153_, new_n47834_ );
and  ( new_n48155_, new_n48154_, new_n48152_ );
nor  ( new_n48156_, new_n48154_, new_n48152_ );
xor  ( new_n48157_, new_n48025_, new_n48024_ );
xor  ( new_n48158_, new_n47972_, new_n47971_ );
xor  ( new_n48159_, new_n48022_, new_n48020_ );
or   ( new_n48160_, new_n48159_, new_n48158_ );
and  ( new_n48161_, new_n48159_, new_n48158_ );
xnor ( new_n48162_, new_n47709_, new_n47708_ );
or   ( new_n48163_, new_n47926_, new_n1137_ );
xor  ( new_n48164_, new_n44974_, new_n893_ );
or   ( new_n48165_, new_n48164_, new_n1135_ );
and  ( new_n48166_, new_n48165_, new_n48163_ );
xor  ( new_n48167_, new_n43985_, new_n2421_ );
or   ( new_n48168_, new_n48167_, new_n2807_ );
or   ( new_n48169_, new_n47922_, new_n2809_ );
and  ( new_n48170_, new_n48169_, new_n48168_ );
nor  ( new_n48171_, new_n48170_, new_n48166_ );
and  ( new_n48172_, new_n48170_, new_n48166_ );
xor  ( new_n48173_, new_n44785_, RIbb2ecb0_21 );
and  ( new_n48174_, new_n48173_, new_n1253_ );
and  ( new_n48175_, new_n47682_, new_n1251_ );
nor  ( new_n48176_, new_n48175_, new_n48174_ );
nor  ( new_n48177_, new_n48176_, new_n48172_ );
nor  ( new_n48178_, new_n48177_, new_n48171_ );
nor  ( new_n48179_, new_n48178_, new_n48162_ );
nand ( new_n48180_, new_n48178_, new_n48162_ );
xnor ( new_n48181_, new_n47685_, new_n47681_ );
xor  ( new_n48182_, new_n48181_, new_n47691_ );
and  ( new_n48183_, new_n48182_, new_n48180_ );
or   ( new_n48184_, new_n48183_, new_n48179_ );
xor  ( new_n48185_, new_n47937_, new_n47921_ );
xor  ( new_n48186_, new_n48185_, new_n47955_ );
and  ( new_n48187_, new_n48186_, new_n48184_ );
or   ( new_n48188_, new_n48186_, new_n48184_ );
xor  ( new_n48189_, new_n47712_, new_n47711_ );
and  ( new_n48190_, new_n48189_, new_n48188_ );
or   ( new_n48191_, new_n48190_, new_n48187_ );
or   ( new_n48192_, new_n48191_, new_n48161_ );
and  ( new_n48193_, new_n48192_, new_n48160_ );
nand ( new_n48194_, new_n48193_, new_n48157_ );
xor  ( new_n48195_, new_n48193_, new_n48157_ );
xor  ( new_n48196_, new_n48144_, new_n48143_ );
nand ( new_n48197_, new_n48196_, new_n48195_ );
and  ( new_n48198_, new_n48197_, new_n48194_ );
xor  ( new_n48199_, new_n47627_, new_n47625_ );
xor  ( new_n48200_, new_n48199_, new_n47723_ );
or   ( new_n48201_, new_n48200_, new_n48198_ );
xor  ( new_n48202_, new_n48148_, new_n48147_ );
xor  ( new_n48203_, new_n48200_, new_n48198_ );
nand ( new_n48204_, new_n48203_, new_n48202_ );
and  ( new_n48205_, new_n48204_, new_n48201_ );
xor  ( new_n48206_, new_n47918_, new_n47916_ );
xor  ( new_n48207_, new_n48206_, new_n48150_ );
nor  ( new_n48208_, new_n48207_, new_n48205_ );
and  ( new_n48209_, new_n48207_, new_n48205_ );
xnor ( new_n48210_, new_n48203_, new_n48202_ );
xor  ( new_n48211_, new_n48196_, new_n48195_ );
xor  ( new_n48212_, new_n47655_, new_n47653_ );
xor  ( new_n48213_, new_n48212_, new_n47658_ );
xnor ( new_n48214_, new_n47959_, new_n47958_ );
xor  ( new_n48215_, new_n48214_, new_n47967_ );
nor  ( new_n48216_, new_n48215_, new_n48213_ );
xor  ( new_n48217_, new_n48012_, new_n48011_ );
xor  ( new_n48218_, new_n47947_, new_n47943_ );
xor  ( new_n48219_, new_n48218_, new_n47952_ );
and  ( new_n48220_, new_n48219_, new_n48217_ );
xnor ( new_n48221_, new_n48009_, new_n48008_ );
xor  ( new_n48222_, new_n43812_, new_n2421_ );
or   ( new_n48223_, new_n48222_, new_n2807_ );
or   ( new_n48224_, new_n48167_, new_n2809_ );
and  ( new_n48225_, new_n48224_, new_n48223_ );
xor  ( new_n48226_, new_n45119_, new_n893_ );
or   ( new_n48227_, new_n48226_, new_n1135_ );
or   ( new_n48228_, new_n48164_, new_n1137_ );
and  ( new_n48229_, new_n48228_, new_n48227_ );
or   ( new_n48230_, new_n48229_, new_n48225_ );
xor  ( new_n48231_, new_n45403_, new_n745_ );
nor  ( new_n48232_, new_n48231_, new_n897_ );
and  ( new_n48233_, new_n48115_, new_n820_ );
nor  ( new_n48234_, new_n48233_, new_n48232_ );
and  ( new_n48235_, new_n48229_, new_n48225_ );
or   ( new_n48236_, new_n48235_, new_n48234_ );
and  ( new_n48237_, new_n48236_, new_n48230_ );
nor  ( new_n48238_, new_n48237_, new_n48221_ );
or   ( new_n48239_, new_n48090_, new_n411_ );
xor  ( new_n48240_, new_n46137_, RIbb2f160_11 );
nand ( new_n48241_, new_n48240_, new_n373_ );
and  ( new_n48242_, new_n48241_, new_n48239_ );
xor  ( new_n48243_, new_n44183_, new_n2118_ );
or   ( new_n48244_, new_n48243_, new_n2425_ );
or   ( new_n48245_, new_n48042_, new_n2427_ );
and  ( new_n48246_, new_n48245_, new_n48244_ );
nor  ( new_n48247_, new_n48246_, new_n48242_ );
xor  ( new_n48248_, new_n45928_, new_n400_ );
nor  ( new_n48249_, new_n48248_, new_n524_ );
and  ( new_n48250_, new_n48048_, new_n454_ );
or   ( new_n48251_, new_n48250_, new_n48249_ );
xor  ( new_n48252_, new_n48246_, new_n48242_ );
and  ( new_n48253_, new_n48252_, new_n48251_ );
nor  ( new_n48254_, new_n48253_, new_n48247_ );
and  ( new_n48255_, new_n48237_, new_n48221_ );
nor  ( new_n48256_, new_n48255_, new_n48254_ );
nor  ( new_n48257_, new_n48256_, new_n48238_ );
not  ( new_n48258_, new_n48257_ );
xor  ( new_n48259_, new_n48219_, new_n48217_ );
and  ( new_n48260_, new_n48259_, new_n48258_ );
or   ( new_n48261_, new_n48260_, new_n48220_ );
xor  ( new_n48262_, new_n48215_, new_n48213_ );
and  ( new_n48263_, new_n48262_, new_n48261_ );
or   ( new_n48264_, new_n48263_, new_n48216_ );
xor  ( new_n48265_, new_n48138_, new_n48137_ );
or   ( new_n48266_, new_n48265_, new_n48264_ );
and  ( new_n48267_, new_n48265_, new_n48264_ );
xor  ( new_n48268_, new_n48015_, new_n48014_ );
xnor ( new_n48269_, new_n48107_, new_n48055_ );
xor  ( new_n48270_, new_n48269_, new_n48133_ );
nor  ( new_n48271_, new_n48270_, new_n48268_ );
and  ( new_n48272_, new_n48270_, new_n48268_ );
not  ( new_n48273_, new_n48272_ );
xor  ( new_n48274_, new_n47303_, new_n275_ );
or   ( new_n48275_, new_n48274_, new_n283_ );
nand ( new_n48276_, new_n47994_, new_n280_ );
and  ( new_n48277_, new_n48276_, new_n48275_ );
xor  ( new_n48278_, new_n46962_, new_n309_ );
or   ( new_n48279_, new_n48278_, new_n317_ );
or   ( new_n48280_, new_n48001_, new_n320_ );
and  ( new_n48281_, new_n48280_, new_n48279_ );
nor  ( new_n48282_, new_n48281_, new_n48277_ );
not  ( new_n48283_, new_n47809_ );
and  ( new_n48284_, new_n48283_, new_n43949_ );
and  ( new_n48285_, new_n47300_, new_n295_ );
nor  ( new_n48286_, new_n48285_, new_n48284_ );
and  ( new_n48287_, new_n48281_, new_n48277_ );
nor  ( new_n48288_, new_n48287_, new_n48286_ );
or   ( new_n48289_, new_n48288_, new_n48282_ );
xor  ( new_n48290_, RIbb329a0_171, RIbb2c460_107 );
xor  ( new_n48291_, new_n48290_, new_n47634_ );
and  ( new_n48292_, new_n48291_, new_n43880_ );
not  ( new_n48293_, new_n48292_ );
nor  ( new_n48294_, RIbb2e170_45, RIbb2e1e8_44 );
or   ( new_n48295_, new_n48294_, new_n4708_ );
xor  ( new_n48296_, new_n43793_, RIbb2e260_43 );
or   ( new_n48297_, new_n48296_, new_n5207_ );
and  ( new_n48298_, new_n48297_, new_n48295_ );
nand ( new_n48299_, new_n48298_, new_n48293_ );
xor  ( new_n48300_, new_n48298_, new_n48293_ );
xor  ( new_n48301_, new_n48039_, new_n43945_ );
not  ( new_n48302_, new_n48301_ );
or   ( new_n48303_, new_n48302_, new_n43983_ );
nor  ( new_n48304_, new_n47640_, new_n43880_ );
or   ( new_n48305_, new_n47641_, new_n43977_ );
or   ( new_n48306_, new_n48305_, new_n48304_ );
and  ( new_n48307_, new_n48306_, new_n48303_ );
nand ( new_n48308_, new_n48307_, new_n48300_ );
and  ( new_n48309_, new_n48308_, new_n48299_ );
nor  ( new_n48310_, new_n48309_, new_n48289_ );
and  ( new_n48311_, new_n48309_, new_n48289_ );
xor  ( new_n48312_, new_n47990_, new_n47982_ );
not  ( new_n48313_, new_n48312_ );
and  ( new_n48314_, new_n48313_, new_n47996_ );
not  ( new_n48315_, new_n47991_ );
and  ( new_n48316_, new_n47997_, new_n48315_ );
nor  ( new_n48317_, new_n48316_, new_n48314_ );
nor  ( new_n48318_, new_n48317_, new_n48311_ );
nor  ( new_n48319_, new_n48318_, new_n48310_ );
not  ( new_n48320_, new_n48319_ );
or   ( new_n48321_, new_n48077_, new_n3898_ );
xor  ( new_n48322_, new_n43884_, RIbb2e530_37 );
nand ( new_n48323_, new_n48322_, new_n3733_ );
and  ( new_n48324_, new_n48323_, new_n48321_ );
or   ( new_n48325_, new_n48094_, new_n4711_ );
xor  ( new_n48326_, new_n43898_, new_n4292_ );
or   ( new_n48327_, new_n48326_, new_n4709_ );
and  ( new_n48328_, new_n48327_, new_n48325_ );
nor  ( new_n48329_, new_n48328_, new_n48324_ );
and  ( new_n48330_, new_n48100_, new_n2000_ );
xor  ( new_n48331_, new_n44319_, RIbb2e9e0_27 );
and  ( new_n48332_, new_n48331_, new_n2002_ );
nor  ( new_n48333_, new_n48332_, new_n48330_ );
and  ( new_n48334_, new_n48328_, new_n48324_ );
nor  ( new_n48335_, new_n48334_, new_n48333_ );
nor  ( new_n48336_, new_n48335_, new_n48329_ );
xor  ( new_n48337_, new_n43799_, new_n3892_ );
or   ( new_n48338_, new_n48337_, new_n4302_ );
nand ( new_n48339_, new_n48065_, new_n4032_ );
and  ( new_n48340_, new_n48339_, new_n48338_ );
xor  ( new_n48341_, new_n43952_, new_n2797_ );
or   ( new_n48342_, new_n48341_, new_n3117_ );
or   ( new_n48343_, new_n48056_, new_n3119_ );
and  ( new_n48344_, new_n48343_, new_n48342_ );
or   ( new_n48345_, new_n48344_, new_n48340_ );
and  ( new_n48346_, new_n48173_, new_n1251_ );
xor  ( new_n48347_, new_n44877_, RIbb2ecb0_21 );
and  ( new_n48348_, new_n48347_, new_n1253_ );
nor  ( new_n48349_, new_n48348_, new_n48346_ );
and  ( new_n48350_, new_n48344_, new_n48340_ );
or   ( new_n48351_, new_n48350_, new_n48349_ );
and  ( new_n48352_, new_n48351_, new_n48345_ );
or   ( new_n48353_, new_n48352_, new_n48336_ );
and  ( new_n48354_, new_n48352_, new_n48336_ );
or   ( new_n48355_, new_n48073_, new_n3463_ );
xor  ( new_n48356_, new_n43937_, RIbb2e620_35 );
nand ( new_n48357_, new_n48356_, new_n3293_ );
and  ( new_n48358_, new_n48357_, new_n48355_ );
xor  ( new_n48359_, new_n44506_, new_n1583_ );
or   ( new_n48360_, new_n48359_, new_n1844_ );
nand ( new_n48361_, new_n48081_, new_n1739_ );
and  ( new_n48362_, new_n48361_, new_n48360_ );
or   ( new_n48363_, new_n48362_, new_n48358_ );
xor  ( new_n48364_, new_n44681_, RIbb2ebc0_23 );
and  ( new_n48365_, new_n48364_, new_n1476_ );
and  ( new_n48366_, new_n48060_, new_n1474_ );
nor  ( new_n48367_, new_n48366_, new_n48365_ );
and  ( new_n48368_, new_n48362_, new_n48358_ );
or   ( new_n48369_, new_n48368_, new_n48367_ );
and  ( new_n48370_, new_n48369_, new_n48363_ );
or   ( new_n48371_, new_n48370_, new_n48354_ );
and  ( new_n48372_, new_n48371_, new_n48353_ );
nor  ( new_n48373_, new_n48372_, new_n48320_ );
xor  ( new_n48374_, new_n48372_, new_n48320_ );
xnor ( new_n48375_, new_n48087_, new_n48071_ );
xor  ( new_n48376_, new_n48375_, new_n48105_ );
and  ( new_n48377_, new_n48376_, new_n48374_ );
nor  ( new_n48378_, new_n48377_, new_n48373_ );
and  ( new_n48379_, new_n48378_, new_n48273_ );
nor  ( new_n48380_, new_n48379_, new_n48271_ );
or   ( new_n48381_, new_n48380_, new_n48267_ );
and  ( new_n48382_, new_n48381_, new_n48266_ );
nand ( new_n48383_, new_n48382_, new_n48211_ );
nor  ( new_n48384_, new_n48382_, new_n48211_ );
xor  ( new_n48385_, new_n48123_, new_n48122_ );
xnor ( new_n48386_, new_n48079_, new_n48075_ );
nand ( new_n48387_, new_n48386_, new_n48084_ );
not  ( new_n48388_, new_n48086_ );
or   ( new_n48389_, new_n48388_, new_n48080_ );
and  ( new_n48390_, new_n48389_, new_n48387_ );
and  ( new_n48391_, new_n48390_, new_n48385_ );
or   ( new_n48392_, new_n48390_, new_n48385_ );
xnor ( new_n48393_, new_n48045_, new_n48041_ );
xor  ( new_n48394_, new_n48393_, new_n48051_ );
and  ( new_n48395_, new_n48394_, new_n48392_ );
or   ( new_n48396_, new_n48395_, new_n48391_ );
xnor ( new_n48397_, new_n48035_, new_n48033_ );
xor  ( new_n48398_, new_n48397_, new_n48053_ );
and  ( new_n48399_, new_n48398_, new_n48396_ );
xor  ( new_n48400_, new_n48063_, new_n48059_ );
not  ( new_n48401_, new_n48400_ );
and  ( new_n48402_, new_n48401_, new_n48068_ );
not  ( new_n48403_, new_n48064_ );
and  ( new_n48404_, new_n48070_, new_n48403_ );
nor  ( new_n48405_, new_n48404_, new_n48402_ );
xnor ( new_n48406_, new_n48097_, new_n48093_ );
xor  ( new_n48407_, new_n48406_, new_n48102_ );
and  ( new_n48408_, new_n48407_, new_n48405_ );
xor  ( new_n48409_, new_n48407_, new_n48405_ );
xnor ( new_n48410_, new_n48170_, new_n48166_ );
nand ( new_n48411_, new_n48410_, new_n48176_ );
not  ( new_n48412_, new_n48177_ );
or   ( new_n48413_, new_n48412_, new_n48171_ );
and  ( new_n48414_, new_n48413_, new_n48411_ );
and  ( new_n48415_, new_n48414_, new_n48409_ );
nor  ( new_n48416_, new_n48415_, new_n48408_ );
xnor ( new_n48417_, new_n48398_, new_n48396_ );
nor  ( new_n48418_, new_n48417_, new_n48416_ );
or   ( new_n48419_, new_n48418_, new_n48399_ );
xor  ( new_n48420_, new_n48186_, new_n48184_ );
xor  ( new_n48421_, new_n48420_, new_n48189_ );
and  ( new_n48422_, new_n48421_, new_n48419_ );
or   ( new_n48423_, new_n48421_, new_n48419_ );
xor  ( new_n48424_, new_n48262_, new_n48261_ );
and  ( new_n48425_, new_n48424_, new_n48423_ );
or   ( new_n48426_, new_n48425_, new_n48422_ );
xor  ( new_n48427_, new_n48159_, new_n48158_ );
xor  ( new_n48428_, new_n48427_, new_n48191_ );
and  ( new_n48429_, new_n48428_, new_n48426_ );
nor  ( new_n48430_, new_n48428_, new_n48426_ );
xor  ( new_n48431_, new_n48178_, new_n48162_ );
xor  ( new_n48432_, new_n48431_, new_n48182_ );
xor  ( new_n48433_, new_n48126_, new_n48125_ );
xor  ( new_n48434_, new_n48433_, new_n48131_ );
nor  ( new_n48435_, new_n48434_, new_n48432_ );
nand ( new_n48436_, new_n48434_, new_n48432_ );
not  ( new_n48437_, new_n48113_ );
xor  ( new_n48438_, new_n45738_, RIbb2ef80_15 );
nand ( new_n48439_, new_n48438_, new_n662_ );
nand ( new_n48440_, new_n48119_, new_n660_ );
and  ( new_n48441_, new_n48440_, new_n48439_ );
nor  ( new_n48442_, new_n48441_, new_n48437_ );
or   ( new_n48443_, new_n48110_, new_n340_ );
xor  ( new_n48444_, new_n46789_, new_n329_ );
or   ( new_n48445_, new_n48444_, new_n337_ );
and  ( new_n48446_, new_n48445_, new_n48443_ );
nor  ( new_n48447_, new_n48446_, new_n5205_ );
and  ( new_n48448_, new_n48240_, new_n371_ );
xor  ( new_n48449_, new_n46427_, RIbb2f160_11 );
and  ( new_n48450_, new_n48449_, new_n373_ );
nor  ( new_n48451_, new_n48450_, new_n48448_ );
xor  ( new_n48452_, new_n48446_, new_n5206_ );
nor  ( new_n48453_, new_n48452_, new_n48451_ );
or   ( new_n48454_, new_n48453_, new_n48447_ );
xor  ( new_n48455_, new_n48441_, new_n48437_ );
and  ( new_n48456_, new_n48455_, new_n48454_ );
nor  ( new_n48457_, new_n48456_, new_n48442_ );
or   ( new_n48458_, new_n48278_, new_n320_ );
xor  ( new_n48459_, new_n46958_, new_n309_ );
or   ( new_n48460_, new_n48459_, new_n317_ );
and  ( new_n48461_, new_n48460_, new_n48458_ );
or   ( new_n48462_, new_n48274_, new_n286_ );
xor  ( new_n48463_, new_n47046_, new_n275_ );
or   ( new_n48464_, new_n48463_, new_n283_ );
and  ( new_n48465_, new_n48464_, new_n48462_ );
or   ( new_n48466_, new_n48465_, new_n48461_ );
and  ( new_n48467_, new_n47984_, new_n43949_ );
and  ( new_n48468_, new_n48283_, new_n295_ );
nor  ( new_n48469_, new_n48468_, new_n48467_ );
xnor ( new_n48470_, new_n48465_, new_n48461_ );
or   ( new_n48471_, new_n48470_, new_n48469_ );
and  ( new_n48472_, new_n48471_, new_n48466_ );
xor  ( new_n48473_, new_n48307_, new_n48300_ );
or   ( new_n48474_, new_n48473_, new_n48472_ );
xor  ( new_n48475_, new_n43985_, RIbb2e710_33 );
nand ( new_n48476_, new_n48475_, new_n2930_ );
or   ( new_n48477_, new_n48341_, new_n3119_ );
and  ( new_n48478_, new_n48477_, new_n48476_ );
or   ( new_n48479_, new_n48231_, new_n899_ );
xor  ( new_n48480_, new_n45584_, new_n745_ );
or   ( new_n48481_, new_n48480_, new_n897_ );
and  ( new_n48482_, new_n48481_, new_n48479_ );
or   ( new_n48483_, new_n48482_, new_n48478_ );
nor  ( new_n48484_, new_n48226_, new_n1137_ );
xor  ( new_n48485_, new_n45204_, RIbb2eda0_19 );
and  ( new_n48486_, new_n48485_, new_n1042_ );
or   ( new_n48487_, new_n48486_, new_n48484_ );
xor  ( new_n48488_, new_n48482_, new_n48478_ );
nand ( new_n48489_, new_n48488_, new_n48487_ );
and  ( new_n48490_, new_n48489_, new_n48483_ );
and  ( new_n48491_, new_n48473_, new_n48472_ );
or   ( new_n48492_, new_n48491_, new_n48490_ );
and  ( new_n48493_, new_n48492_, new_n48474_ );
nor  ( new_n48494_, new_n48493_, new_n48457_ );
xor  ( new_n48495_, new_n48493_, new_n48457_ );
not  ( new_n48496_, new_n48495_ );
xor  ( new_n48497_, new_n48281_, new_n48277_ );
xor  ( new_n48498_, new_n48497_, new_n48286_ );
xor  ( new_n48499_, new_n44785_, RIbb2ebc0_23 );
nand ( new_n48500_, new_n48499_, new_n1476_ );
nand ( new_n48501_, new_n48364_, new_n1474_ );
and  ( new_n48502_, new_n48501_, new_n48500_ );
nand ( new_n48503_, new_n48347_, new_n1251_ );
xor  ( new_n48504_, new_n44974_, new_n1126_ );
or   ( new_n48505_, new_n48504_, new_n1364_ );
and  ( new_n48506_, new_n48505_, new_n48503_ );
or   ( new_n48507_, new_n48506_, new_n48502_ );
and  ( new_n48508_, new_n48356_, new_n3291_ );
xor  ( new_n48509_, new_n43956_, new_n3113_ );
nor  ( new_n48510_, new_n48509_, new_n3461_ );
nor  ( new_n48511_, new_n48510_, new_n48508_ );
and  ( new_n48512_, new_n48506_, new_n48502_ );
or   ( new_n48513_, new_n48512_, new_n48511_ );
and  ( new_n48514_, new_n48513_, new_n48507_ );
or   ( new_n48515_, new_n48514_, new_n48498_ );
and  ( new_n48516_, new_n48514_, new_n48498_ );
xor  ( new_n48517_, RIbb32a18_172, RIbb2c3e8_108 );
xor  ( new_n48518_, new_n48517_, new_n46412_ );
not  ( new_n48519_, new_n48518_ );
or   ( new_n48520_, new_n48519_, new_n43879_ );
or   ( new_n48521_, new_n48222_, new_n2809_ );
xor  ( new_n48522_, new_n43914_, new_n2421_ );
or   ( new_n48523_, new_n48522_, new_n2807_ );
and  ( new_n48524_, new_n48523_, new_n48521_ );
nor  ( new_n48525_, new_n48524_, new_n48520_ );
and  ( new_n48526_, new_n48524_, new_n48520_ );
xor  ( new_n48527_, new_n48291_, new_n43945_ );
and  ( new_n48528_, new_n48527_, new_n43982_ );
and  ( new_n48529_, new_n48040_, new_n43879_ );
not  ( new_n48530_, new_n48529_ );
and  ( new_n48531_, new_n48041_, new_n43978_ );
and  ( new_n48532_, new_n48531_, new_n48530_ );
nor  ( new_n48533_, new_n48532_, new_n48528_ );
nor  ( new_n48534_, new_n48533_, new_n48526_ );
nor  ( new_n48535_, new_n48534_, new_n48525_ );
or   ( new_n48536_, new_n48535_, new_n48516_ );
and  ( new_n48537_, new_n48536_, new_n48515_ );
nor  ( new_n48538_, new_n48537_, new_n48496_ );
nor  ( new_n48539_, new_n48538_, new_n48494_ );
and  ( new_n48540_, new_n48539_, new_n48436_ );
or   ( new_n48541_, new_n48540_, new_n48435_ );
xor  ( new_n48542_, new_n48270_, new_n48268_ );
xor  ( new_n48543_, new_n48542_, new_n48378_ );
nor  ( new_n48544_, new_n48543_, new_n48541_ );
and  ( new_n48545_, new_n48543_, new_n48541_ );
xnor ( new_n48546_, new_n48376_, new_n48374_ );
xor  ( new_n48547_, new_n43894_, new_n4292_ );
or   ( new_n48548_, new_n48547_, new_n4709_ );
or   ( new_n48549_, new_n48326_, new_n4711_ );
and  ( new_n48550_, new_n48549_, new_n48548_ );
or   ( new_n48551_, new_n48359_, new_n1846_ );
xor  ( new_n48552_, new_n44600_, new_n1583_ );
or   ( new_n48553_, new_n48552_, new_n1844_ );
and  ( new_n48554_, new_n48553_, new_n48551_ );
nor  ( new_n48555_, new_n48554_, new_n48550_ );
xor  ( new_n48556_, new_n43888_, RIbb2e530_37 );
and  ( new_n48557_, new_n48556_, new_n3733_ );
and  ( new_n48558_, new_n48322_, new_n3731_ );
nor  ( new_n48559_, new_n48558_, new_n48557_ );
and  ( new_n48560_, new_n48554_, new_n48550_ );
nor  ( new_n48561_, new_n48560_, new_n48559_ );
nor  ( new_n48562_, new_n48561_, new_n48555_ );
or   ( new_n48563_, new_n48243_, new_n2427_ );
xor  ( new_n48564_, new_n44218_, new_n2118_ );
or   ( new_n48565_, new_n48564_, new_n2425_ );
and  ( new_n48566_, new_n48565_, new_n48563_ );
xor  ( new_n48567_, new_n43803_, new_n3892_ );
or   ( new_n48568_, new_n48567_, new_n4302_ );
or   ( new_n48569_, new_n48337_, new_n4304_ );
and  ( new_n48570_, new_n48569_, new_n48568_ );
or   ( new_n48571_, new_n48570_, new_n48566_ );
xor  ( new_n48572_, new_n44407_, RIbb2e9e0_27 );
and  ( new_n48573_, new_n48572_, new_n2002_ );
and  ( new_n48574_, new_n48331_, new_n2000_ );
nor  ( new_n48575_, new_n48574_, new_n48573_ );
and  ( new_n48576_, new_n48570_, new_n48566_ );
or   ( new_n48577_, new_n48576_, new_n48575_ );
and  ( new_n48578_, new_n48577_, new_n48571_ );
nor  ( new_n48579_, new_n48578_, new_n48562_ );
xor  ( new_n48580_, new_n43787_, RIbb2e260_43 );
nand ( new_n48581_, new_n48580_, new_n4960_ );
or   ( new_n48582_, new_n48296_, new_n5209_ );
and  ( new_n48583_, new_n48582_, new_n48581_ );
xor  ( new_n48584_, new_n46037_, new_n400_ );
or   ( new_n48585_, new_n48584_, new_n524_ );
or   ( new_n48586_, new_n48248_, new_n526_ );
and  ( new_n48587_, new_n48586_, new_n48585_ );
nor  ( new_n48588_, new_n48587_, new_n48583_ );
xor  ( new_n48589_, new_n45597_, RIbb2ef80_15 );
and  ( new_n48590_, new_n48589_, new_n662_ );
and  ( new_n48591_, new_n48438_, new_n660_ );
nor  ( new_n48592_, new_n48591_, new_n48590_ );
and  ( new_n48593_, new_n48587_, new_n48583_ );
nor  ( new_n48594_, new_n48593_, new_n48592_ );
or   ( new_n48595_, new_n48594_, new_n48588_ );
xor  ( new_n48596_, new_n48578_, new_n48562_ );
and  ( new_n48597_, new_n48596_, new_n48595_ );
or   ( new_n48598_, new_n48597_, new_n48579_ );
xor  ( new_n48599_, new_n48309_, new_n48289_ );
xor  ( new_n48600_, new_n48599_, new_n48317_ );
nand ( new_n48601_, new_n48600_, new_n48598_ );
nor  ( new_n48602_, new_n48600_, new_n48598_ );
xnor ( new_n48603_, new_n48328_, new_n48324_ );
nand ( new_n48604_, new_n48603_, new_n48333_ );
not  ( new_n48605_, new_n48335_ );
or   ( new_n48606_, new_n48605_, new_n48329_ );
and  ( new_n48607_, new_n48606_, new_n48604_ );
xnor ( new_n48608_, new_n48344_, new_n48340_ );
xor  ( new_n48609_, new_n48608_, new_n48349_ );
and  ( new_n48610_, new_n48609_, new_n48607_ );
nor  ( new_n48611_, new_n48609_, new_n48607_ );
not  ( new_n48612_, new_n48611_ );
xor  ( new_n48613_, new_n48229_, new_n48225_ );
xnor ( new_n48614_, new_n48613_, new_n48234_ );
and  ( new_n48615_, new_n48614_, new_n48612_ );
nor  ( new_n48616_, new_n48615_, new_n48610_ );
or   ( new_n48617_, new_n48616_, new_n48602_ );
and  ( new_n48618_, new_n48617_, new_n48601_ );
nor  ( new_n48619_, new_n48618_, new_n48546_ );
and  ( new_n48620_, new_n48618_, new_n48546_ );
not  ( new_n48621_, new_n48620_ );
xor  ( new_n48622_, new_n48259_, new_n48258_ );
and  ( new_n48623_, new_n48622_, new_n48621_ );
nor  ( new_n48624_, new_n48623_, new_n48619_ );
nor  ( new_n48625_, new_n48624_, new_n48545_ );
nor  ( new_n48626_, new_n48625_, new_n48544_ );
nor  ( new_n48627_, new_n48626_, new_n48430_ );
nor  ( new_n48628_, new_n48627_, new_n48429_ );
or   ( new_n48629_, new_n48628_, new_n48384_ );
and  ( new_n48630_, new_n48629_, new_n48383_ );
nor  ( new_n48631_, new_n48630_, new_n48210_ );
and  ( new_n48632_, new_n48630_, new_n48210_ );
xor  ( new_n48633_, new_n48428_, new_n48426_ );
xor  ( new_n48634_, new_n48633_, new_n48626_ );
xnor ( new_n48635_, new_n48265_, new_n48264_ );
xor  ( new_n48636_, new_n48635_, new_n48380_ );
and  ( new_n48637_, new_n48636_, new_n48634_ );
xnor ( new_n48638_, new_n48417_, new_n48416_ );
xor  ( new_n48639_, new_n48352_, new_n48336_ );
xor  ( new_n48640_, new_n48639_, new_n48370_ );
xor  ( new_n48641_, new_n48237_, new_n48221_ );
xor  ( new_n48642_, new_n48641_, new_n48254_ );
or   ( new_n48643_, new_n48642_, new_n48640_ );
and  ( new_n48644_, new_n48642_, new_n48640_ );
xor  ( new_n48645_, new_n48252_, new_n48251_ );
xnor ( new_n48646_, new_n48362_, new_n48358_ );
xor  ( new_n48647_, new_n48646_, new_n48367_ );
nand ( new_n48648_, new_n48647_, new_n48645_ );
nor  ( new_n48649_, new_n48647_, new_n48645_ );
and  ( new_n48650_, new_n48449_, new_n371_ );
xor  ( new_n48651_, new_n46619_, new_n325_ );
nor  ( new_n48652_, new_n48651_, new_n409_ );
nor  ( new_n48653_, new_n48652_, new_n48650_ );
xor  ( new_n48654_, new_n47303_, new_n309_ );
or   ( new_n48655_, new_n48654_, new_n317_ );
or   ( new_n48656_, new_n48459_, new_n320_ );
and  ( new_n48657_, new_n48656_, new_n48655_ );
or   ( new_n48658_, new_n48444_, new_n340_ );
xor  ( new_n48659_, new_n46962_, new_n329_ );
or   ( new_n48660_, new_n48659_, new_n337_ );
and  ( new_n48661_, new_n48660_, new_n48658_ );
or   ( new_n48662_, new_n48661_, new_n48657_ );
xor  ( new_n48663_, new_n47296_, RIbb2f430_5 );
and  ( new_n48664_, new_n48663_, new_n282_ );
nor  ( new_n48665_, new_n48463_, new_n286_ );
nor  ( new_n48666_, new_n48665_, new_n48664_ );
xnor ( new_n48667_, new_n48661_, new_n48657_ );
or   ( new_n48668_, new_n48667_, new_n48666_ );
and  ( new_n48669_, new_n48668_, new_n48662_ );
or   ( new_n48670_, new_n48669_, new_n48653_ );
nor  ( new_n48671_, RIbb2e080_47, RIbb2e0f8_46 );
or   ( new_n48672_, new_n48671_, new_n5206_ );
xor  ( new_n48673_, new_n43793_, RIbb2e170_45 );
or   ( new_n48674_, new_n48673_, new_n5604_ );
and  ( new_n48675_, new_n48674_, new_n48672_ );
xor  ( new_n48676_, new_n48518_, new_n43945_ );
not  ( new_n48677_, new_n48676_ );
or   ( new_n48678_, new_n48677_, new_n43983_ );
nor  ( new_n48679_, new_n48291_, new_n43880_ );
or   ( new_n48680_, new_n48292_, new_n43977_ );
or   ( new_n48681_, new_n48680_, new_n48679_ );
and  ( new_n48682_, new_n48681_, new_n48678_ );
nor  ( new_n48683_, new_n48682_, new_n48675_ );
and  ( new_n48684_, new_n47984_, new_n295_ );
and  ( new_n48685_, new_n48302_, new_n43949_ );
nor  ( new_n48686_, new_n48685_, new_n48684_ );
xnor ( new_n48687_, new_n48682_, new_n48675_ );
nor  ( new_n48688_, new_n48687_, new_n48686_ );
or   ( new_n48689_, new_n48688_, new_n48683_ );
xor  ( new_n48690_, new_n48669_, new_n48653_ );
nand ( new_n48691_, new_n48690_, new_n48689_ );
and  ( new_n48692_, new_n48691_, new_n48670_ );
or   ( new_n48693_, new_n48692_, new_n48649_ );
and  ( new_n48694_, new_n48693_, new_n48648_ );
or   ( new_n48695_, new_n48694_, new_n48644_ );
and  ( new_n48696_, new_n48695_, new_n48643_ );
nor  ( new_n48697_, new_n48696_, new_n48638_ );
and  ( new_n48698_, new_n48696_, new_n48638_ );
xor  ( new_n48699_, new_n48414_, new_n48409_ );
xor  ( new_n48700_, new_n48390_, new_n48385_ );
xor  ( new_n48701_, new_n48700_, new_n48394_ );
and  ( new_n48702_, new_n48701_, new_n48699_ );
xor  ( new_n48703_, new_n48701_, new_n48699_ );
xor  ( new_n48704_, new_n48455_, new_n48454_ );
xnor ( new_n48705_, new_n48470_, new_n48469_ );
xor  ( new_n48706_, new_n45119_, new_n1126_ );
or   ( new_n48707_, new_n48706_, new_n1364_ );
or   ( new_n48708_, new_n48504_, new_n1366_ );
and  ( new_n48709_, new_n48708_, new_n48707_ );
xor  ( new_n48710_, new_n43952_, new_n3113_ );
or   ( new_n48711_, new_n48710_, new_n3461_ );
or   ( new_n48712_, new_n48509_, new_n3463_ );
and  ( new_n48713_, new_n48712_, new_n48711_ );
nor  ( new_n48714_, new_n48713_, new_n48709_ );
and  ( new_n48715_, new_n48713_, new_n48709_ );
and  ( new_n48716_, new_n48475_, new_n2928_ );
xor  ( new_n48717_, new_n43812_, RIbb2e710_33 );
and  ( new_n48718_, new_n48717_, new_n2930_ );
nor  ( new_n48719_, new_n48718_, new_n48716_ );
nor  ( new_n48720_, new_n48719_, new_n48715_ );
nor  ( new_n48721_, new_n48720_, new_n48714_ );
nand ( new_n48722_, new_n48721_, new_n48705_ );
nor  ( new_n48723_, new_n48721_, new_n48705_ );
xor  ( new_n48724_, new_n48524_, new_n48520_ );
xnor ( new_n48725_, new_n48724_, new_n48533_ );
or   ( new_n48726_, new_n48725_, new_n48723_ );
and  ( new_n48727_, new_n48726_, new_n48722_ );
or   ( new_n48728_, new_n48727_, new_n48704_ );
nand ( new_n48729_, new_n48727_, new_n48704_ );
xnor ( new_n48730_, new_n48452_, new_n48451_ );
or   ( new_n48731_, new_n48547_, new_n4711_ );
xor  ( new_n48732_, new_n43799_, new_n4292_ );
or   ( new_n48733_, new_n48732_, new_n4709_ );
and  ( new_n48734_, new_n48733_, new_n48731_ );
xor  ( new_n48735_, new_n44681_, RIbb2ead0_25 );
nand ( new_n48736_, new_n48735_, new_n1741_ );
or   ( new_n48737_, new_n48552_, new_n1846_ );
and  ( new_n48738_, new_n48737_, new_n48736_ );
or   ( new_n48739_, new_n48738_, new_n48734_ );
xor  ( new_n48740_, new_n44877_, RIbb2ebc0_23 );
and  ( new_n48741_, new_n48740_, new_n1476_ );
and  ( new_n48742_, new_n48499_, new_n1474_ );
nor  ( new_n48743_, new_n48742_, new_n48741_ );
and  ( new_n48744_, new_n48738_, new_n48734_ );
or   ( new_n48745_, new_n48744_, new_n48743_ );
and  ( new_n48746_, new_n48745_, new_n48739_ );
nor  ( new_n48747_, new_n48746_, new_n48730_ );
xor  ( new_n48748_, RIbb32a90_173, RIbb2c370_109 );
and  ( new_n48749_, new_n46409_, new_n43555_ );
nor  ( new_n48750_, new_n48749_, new_n43597_ );
not  ( new_n48751_, new_n48750_ );
and  ( new_n48752_, new_n48751_, new_n43553_ );
nor  ( new_n48753_, new_n48752_, new_n43600_ );
nor  ( new_n48754_, new_n48753_, new_n43549_ );
nor  ( new_n48755_, new_n48754_, new_n43601_ );
xnor ( new_n48756_, new_n48755_, new_n48748_ );
and  ( new_n48757_, new_n48756_, new_n43880_ );
not  ( new_n48758_, new_n48757_ );
xor  ( new_n48759_, new_n44183_, new_n2421_ );
or   ( new_n48760_, new_n48759_, new_n2807_ );
or   ( new_n48761_, new_n48522_, new_n2809_ );
and  ( new_n48762_, new_n48761_, new_n48760_ );
nor  ( new_n48763_, new_n48762_, new_n48758_ );
and  ( new_n48764_, new_n48589_, new_n660_ );
xor  ( new_n48765_, new_n45928_, new_n520_ );
nor  ( new_n48766_, new_n48765_, new_n755_ );
or   ( new_n48767_, new_n48766_, new_n48764_ );
xor  ( new_n48768_, new_n48762_, new_n48758_ );
and  ( new_n48769_, new_n48768_, new_n48767_ );
nor  ( new_n48770_, new_n48769_, new_n48763_ );
and  ( new_n48771_, new_n48746_, new_n48730_ );
nor  ( new_n48772_, new_n48771_, new_n48770_ );
nor  ( new_n48773_, new_n48772_, new_n48747_ );
nand ( new_n48774_, new_n48773_, new_n48729_ );
and  ( new_n48775_, new_n48774_, new_n48728_ );
and  ( new_n48776_, new_n48775_, new_n48703_ );
nor  ( new_n48777_, new_n48776_, new_n48702_ );
nor  ( new_n48778_, new_n48777_, new_n48698_ );
nor  ( new_n48779_, new_n48778_, new_n48697_ );
xor  ( new_n48780_, new_n48421_, new_n48419_ );
xnor ( new_n48781_, new_n48780_, new_n48424_ );
and  ( new_n48782_, new_n48781_, new_n48779_ );
xnor ( new_n48783_, new_n48781_, new_n48779_ );
xnor ( new_n48784_, new_n48543_, new_n48541_ );
xor  ( new_n48785_, new_n48784_, new_n48624_ );
nor  ( new_n48786_, new_n48785_, new_n48783_ );
or   ( new_n48787_, new_n48786_, new_n48782_ );
xor  ( new_n48788_, new_n48636_, new_n48634_ );
and  ( new_n48789_, new_n48788_, new_n48787_ );
nor  ( new_n48790_, new_n48789_, new_n48637_ );
xor  ( new_n48791_, new_n48382_, new_n48211_ );
xnor ( new_n48792_, new_n48791_, new_n48628_ );
and  ( new_n48793_, new_n48792_, new_n48790_ );
nor  ( new_n48794_, new_n48792_, new_n48790_ );
xor  ( new_n48795_, new_n48537_, new_n48496_ );
xnor ( new_n48796_, new_n48600_, new_n48598_ );
xor  ( new_n48797_, new_n48796_, new_n48616_ );
and  ( new_n48798_, new_n48797_, new_n48795_ );
xor  ( new_n48799_, new_n48797_, new_n48795_ );
xor  ( new_n48800_, new_n48473_, new_n48472_ );
xor  ( new_n48801_, new_n48800_, new_n48490_ );
or   ( new_n48802_, new_n48567_, new_n4304_ );
xor  ( new_n48803_, new_n43884_, new_n3892_ );
or   ( new_n48804_, new_n48803_, new_n4302_ );
and  ( new_n48805_, new_n48804_, new_n48802_ );
nand ( new_n48806_, new_n48556_, new_n3731_ );
xor  ( new_n48807_, new_n43937_, new_n3457_ );
or   ( new_n48808_, new_n48807_, new_n3896_ );
and  ( new_n48809_, new_n48808_, new_n48806_ );
or   ( new_n48810_, new_n48809_, new_n48805_ );
and  ( new_n48811_, new_n48572_, new_n2000_ );
xor  ( new_n48812_, new_n44506_, RIbb2e9e0_27 );
and  ( new_n48813_, new_n48812_, new_n2002_ );
or   ( new_n48814_, new_n48813_, new_n48811_ );
xor  ( new_n48815_, new_n48809_, new_n48805_ );
nand ( new_n48816_, new_n48815_, new_n48814_ );
and  ( new_n48817_, new_n48816_, new_n48810_ );
not  ( new_n48818_, new_n48653_ );
xor  ( new_n48819_, new_n45738_, new_n745_ );
or   ( new_n48820_, new_n48819_, new_n897_ );
or   ( new_n48821_, new_n48480_, new_n899_ );
and  ( new_n48822_, new_n48821_, new_n48820_ );
or   ( new_n48823_, new_n48822_, new_n48818_ );
and  ( new_n48824_, new_n48485_, new_n1040_ );
xor  ( new_n48825_, new_n45403_, new_n893_ );
nor  ( new_n48826_, new_n48825_, new_n1135_ );
or   ( new_n48827_, new_n48826_, new_n48824_ );
xor  ( new_n48828_, new_n48822_, new_n48818_ );
nand ( new_n48829_, new_n48828_, new_n48827_ );
and  ( new_n48830_, new_n48829_, new_n48823_ );
or   ( new_n48831_, new_n48830_, new_n48817_ );
and  ( new_n48832_, new_n48830_, new_n48817_ );
or   ( new_n48833_, new_n48584_, new_n526_ );
xor  ( new_n48834_, new_n46137_, RIbb2f070_13 );
nand ( new_n48835_, new_n48834_, new_n456_ );
and  ( new_n48836_, new_n48835_, new_n48833_ );
xor  ( new_n48837_, new_n44319_, RIbb2e8f0_29 );
nand ( new_n48838_, new_n48837_, new_n2244_ );
or   ( new_n48839_, new_n48564_, new_n2427_ );
and  ( new_n48840_, new_n48839_, new_n48838_ );
or   ( new_n48841_, new_n48840_, new_n48836_ );
and  ( new_n48842_, new_n48580_, new_n4958_ );
xor  ( new_n48843_, new_n43898_, new_n4705_ );
nor  ( new_n48844_, new_n48843_, new_n5207_ );
nor  ( new_n48845_, new_n48844_, new_n48842_ );
and  ( new_n48846_, new_n48840_, new_n48836_ );
or   ( new_n48847_, new_n48846_, new_n48845_ );
and  ( new_n48848_, new_n48847_, new_n48841_ );
or   ( new_n48849_, new_n48848_, new_n48832_ );
and  ( new_n48850_, new_n48849_, new_n48831_ );
nand ( new_n48851_, new_n48850_, new_n48801_ );
xor  ( new_n48852_, new_n48596_, new_n48595_ );
nor  ( new_n48853_, new_n48850_, new_n48801_ );
or   ( new_n48854_, new_n48853_, new_n48852_ );
and  ( new_n48855_, new_n48854_, new_n48851_ );
and  ( new_n48856_, new_n48855_, new_n48799_ );
or   ( new_n48857_, new_n48856_, new_n48798_ );
xor  ( new_n48858_, new_n48618_, new_n48546_ );
xor  ( new_n48859_, new_n48858_, new_n48622_ );
nor  ( new_n48860_, new_n48859_, new_n48857_ );
xor  ( new_n48861_, new_n48434_, new_n48432_ );
xnor ( new_n48862_, new_n48861_, new_n48539_ );
and  ( new_n48863_, new_n48859_, new_n48857_ );
nor  ( new_n48864_, new_n48863_, new_n48862_ );
nor  ( new_n48865_, new_n48864_, new_n48860_ );
not  ( new_n48866_, new_n48865_ );
xor  ( new_n48867_, new_n48696_, new_n48638_ );
xor  ( new_n48868_, new_n48867_, new_n48777_ );
xnor ( new_n48869_, new_n48775_, new_n48703_ );
xor  ( new_n48870_, new_n48609_, new_n48607_ );
xor  ( new_n48871_, new_n48870_, new_n48614_ );
xnor ( new_n48872_, new_n48514_, new_n48498_ );
xor  ( new_n48873_, new_n48872_, new_n48535_ );
nand ( new_n48874_, new_n48873_, new_n48871_ );
nor  ( new_n48875_, new_n48873_, new_n48871_ );
xor  ( new_n48876_, new_n48488_, new_n48487_ );
xnor ( new_n48877_, new_n48570_, new_n48566_ );
xor  ( new_n48878_, new_n48877_, new_n48575_ );
and  ( new_n48879_, new_n48878_, new_n48876_ );
nor  ( new_n48880_, new_n48878_, new_n48876_ );
xor  ( new_n48881_, new_n48506_, new_n48502_ );
xnor ( new_n48882_, new_n48881_, new_n48511_ );
not  ( new_n48883_, new_n48882_ );
nor  ( new_n48884_, new_n48883_, new_n48880_ );
nor  ( new_n48885_, new_n48884_, new_n48879_ );
or   ( new_n48886_, new_n48885_, new_n48875_ );
and  ( new_n48887_, new_n48886_, new_n48874_ );
or   ( new_n48888_, new_n48887_, new_n48869_ );
and  ( new_n48889_, new_n48887_, new_n48869_ );
xor  ( new_n48890_, new_n48642_, new_n48640_ );
xor  ( new_n48891_, new_n48890_, new_n48694_ );
or   ( new_n48892_, new_n48891_, new_n48889_ );
and  ( new_n48893_, new_n48892_, new_n48888_ );
or   ( new_n48894_, new_n48893_, new_n48868_ );
and  ( new_n48895_, new_n48893_, new_n48868_ );
xnor ( new_n48896_, new_n48554_, new_n48550_ );
nand ( new_n48897_, new_n48896_, new_n48559_ );
not  ( new_n48898_, new_n48561_ );
or   ( new_n48899_, new_n48898_, new_n48555_ );
and  ( new_n48900_, new_n48899_, new_n48897_ );
xnor ( new_n48901_, new_n48587_, new_n48583_ );
nand ( new_n48902_, new_n48901_, new_n48592_ );
not  ( new_n48903_, new_n48588_ );
nand ( new_n48904_, new_n48594_, new_n48903_ );
and  ( new_n48905_, new_n48904_, new_n48902_ );
nand ( new_n48906_, new_n48905_, new_n48900_ );
xor  ( new_n48907_, RIbb32b08_174, RIbb2c2f8_110 );
xnor ( new_n48908_, new_n48907_, new_n48753_ );
and  ( new_n48909_, new_n48908_, new_n43880_ );
not  ( new_n48910_, new_n48909_ );
xor  ( new_n48911_, new_n48756_, new_n43945_ );
not  ( new_n48912_, new_n48911_ );
or   ( new_n48913_, new_n48912_, new_n43983_ );
and  ( new_n48914_, new_n48519_, new_n43879_ );
nand ( new_n48915_, new_n48520_, new_n43978_ );
or   ( new_n48916_, new_n48915_, new_n48914_ );
and  ( new_n48917_, new_n48916_, new_n48913_ );
or   ( new_n48918_, new_n48917_, new_n48910_ );
not  ( new_n48919_, new_n48527_ );
and  ( new_n48920_, new_n48919_, new_n43949_ );
and  ( new_n48921_, new_n48302_, new_n295_ );
or   ( new_n48922_, new_n48921_, new_n48920_ );
xor  ( new_n48923_, new_n48917_, new_n48910_ );
nand ( new_n48924_, new_n48923_, new_n48922_ );
and  ( new_n48925_, new_n48924_, new_n48918_ );
xor  ( new_n48926_, new_n46789_, new_n325_ );
or   ( new_n48927_, new_n48926_, new_n409_ );
or   ( new_n48928_, new_n48651_, new_n411_ );
and  ( new_n48929_, new_n48928_, new_n48927_ );
or   ( new_n48930_, new_n48929_, new_n5596_ );
and  ( new_n48931_, new_n48834_, new_n454_ );
xor  ( new_n48932_, new_n46427_, RIbb2f070_13 );
and  ( new_n48933_, new_n48932_, new_n456_ );
or   ( new_n48934_, new_n48933_, new_n48931_ );
xor  ( new_n48935_, new_n48929_, new_n5596_ );
nand ( new_n48936_, new_n48935_, new_n48934_ );
and  ( new_n48937_, new_n48936_, new_n48930_ );
nor  ( new_n48938_, new_n48937_, new_n48925_ );
nand ( new_n48939_, new_n48663_, new_n280_ );
xor  ( new_n48940_, new_n47640_, new_n275_ );
or   ( new_n48941_, new_n48940_, new_n283_ );
and  ( new_n48942_, new_n48941_, new_n48939_ );
or   ( new_n48943_, new_n48659_, new_n340_ );
xor  ( new_n48944_, new_n46958_, new_n329_ );
or   ( new_n48945_, new_n48944_, new_n337_ );
and  ( new_n48946_, new_n48945_, new_n48943_ );
nor  ( new_n48947_, new_n48946_, new_n48942_ );
nor  ( new_n48948_, new_n48654_, new_n320_ );
xor  ( new_n48949_, new_n47046_, new_n309_ );
nor  ( new_n48950_, new_n48949_, new_n317_ );
nor  ( new_n48951_, new_n48950_, new_n48948_ );
xnor ( new_n48952_, new_n48946_, new_n48942_ );
nor  ( new_n48953_, new_n48952_, new_n48951_ );
or   ( new_n48954_, new_n48953_, new_n48947_ );
xor  ( new_n48955_, new_n48937_, new_n48925_ );
and  ( new_n48956_, new_n48955_, new_n48954_ );
nor  ( new_n48957_, new_n48956_, new_n48938_ );
xnor ( new_n48958_, new_n48905_, new_n48900_ );
or   ( new_n48959_, new_n48958_, new_n48957_ );
and  ( new_n48960_, new_n48959_, new_n48906_ );
xor  ( new_n48961_, new_n48647_, new_n48645_ );
xor  ( new_n48962_, new_n48961_, new_n48692_ );
or   ( new_n48963_, new_n48962_, new_n48960_ );
xnor ( new_n48964_, new_n48687_, new_n48686_ );
xor  ( new_n48965_, new_n43888_, new_n3892_ );
or   ( new_n48966_, new_n48965_, new_n4302_ );
or   ( new_n48967_, new_n48803_, new_n4304_ );
and  ( new_n48968_, new_n48967_, new_n48966_ );
nand ( new_n48969_, new_n48812_, new_n2000_ );
xor  ( new_n48970_, new_n44600_, RIbb2e9e0_27 );
nand ( new_n48971_, new_n48970_, new_n2002_ );
and  ( new_n48972_, new_n48971_, new_n48969_ );
nor  ( new_n48973_, new_n48972_, new_n48968_ );
and  ( new_n48974_, new_n48837_, new_n2242_ );
xor  ( new_n48975_, new_n44407_, RIbb2e8f0_29 );
and  ( new_n48976_, new_n48975_, new_n2244_ );
nor  ( new_n48977_, new_n48976_, new_n48974_ );
and  ( new_n48978_, new_n48972_, new_n48968_ );
nor  ( new_n48979_, new_n48978_, new_n48977_ );
nor  ( new_n48980_, new_n48979_, new_n48973_ );
nor  ( new_n48981_, new_n48980_, new_n48964_ );
xor  ( new_n48982_, new_n43914_, RIbb2e710_33 );
nand ( new_n48983_, new_n48982_, new_n2930_ );
nand ( new_n48984_, new_n48717_, new_n2928_ );
and  ( new_n48985_, new_n48984_, new_n48983_ );
or   ( new_n48986_, new_n48819_, new_n899_ );
xor  ( new_n48987_, new_n45597_, RIbb2ee90_17 );
nand ( new_n48988_, new_n48987_, new_n822_ );
and  ( new_n48989_, new_n48988_, new_n48986_ );
nor  ( new_n48990_, new_n48989_, new_n48985_ );
nor  ( new_n48991_, new_n48765_, new_n757_ );
xor  ( new_n48992_, new_n46037_, new_n520_ );
nor  ( new_n48993_, new_n48992_, new_n755_ );
or   ( new_n48994_, new_n48993_, new_n48991_ );
xor  ( new_n48995_, new_n48989_, new_n48985_ );
and  ( new_n48996_, new_n48995_, new_n48994_ );
or   ( new_n48997_, new_n48996_, new_n48990_ );
xor  ( new_n48998_, new_n48980_, new_n48964_ );
and  ( new_n48999_, new_n48998_, new_n48997_ );
or   ( new_n49000_, new_n48999_, new_n48981_ );
xor  ( new_n49001_, new_n48690_, new_n48689_ );
and  ( new_n49002_, new_n49001_, new_n49000_ );
xnor ( new_n49003_, new_n48667_, new_n48666_ );
or   ( new_n49004_, new_n48710_, new_n3463_ );
xor  ( new_n49005_, new_n43985_, new_n3113_ );
or   ( new_n49006_, new_n49005_, new_n3461_ );
and  ( new_n49007_, new_n49006_, new_n49004_ );
nand ( new_n49008_, new_n48740_, new_n1474_ );
xor  ( new_n49009_, new_n44974_, RIbb2ebc0_23 );
nand ( new_n49010_, new_n49009_, new_n1476_ );
and  ( new_n49011_, new_n49010_, new_n49008_ );
or   ( new_n49012_, new_n49011_, new_n49007_ );
nor  ( new_n49013_, new_n48706_, new_n1366_ );
xor  ( new_n49014_, new_n45204_, RIbb2ecb0_21 );
and  ( new_n49015_, new_n49014_, new_n1253_ );
nor  ( new_n49016_, new_n49015_, new_n49013_ );
and  ( new_n49017_, new_n49011_, new_n49007_ );
or   ( new_n49018_, new_n49017_, new_n49016_ );
and  ( new_n49019_, new_n49018_, new_n49012_ );
nor  ( new_n49020_, new_n49019_, new_n49003_ );
xor  ( new_n49021_, new_n43956_, new_n3457_ );
or   ( new_n49022_, new_n49021_, new_n3896_ );
or   ( new_n49023_, new_n48807_, new_n3898_ );
and  ( new_n49024_, new_n49023_, new_n49022_ );
or   ( new_n49025_, new_n48843_, new_n5209_ );
xor  ( new_n49026_, new_n43894_, new_n4705_ );
or   ( new_n49027_, new_n49026_, new_n5207_ );
and  ( new_n49028_, new_n49027_, new_n49025_ );
nor  ( new_n49029_, new_n49028_, new_n49024_ );
and  ( new_n49030_, new_n48735_, new_n1739_ );
xor  ( new_n49031_, new_n44785_, RIbb2ead0_25 );
and  ( new_n49032_, new_n49031_, new_n1741_ );
or   ( new_n49033_, new_n49032_, new_n49030_ );
xor  ( new_n49034_, new_n49028_, new_n49024_ );
and  ( new_n49035_, new_n49034_, new_n49033_ );
nor  ( new_n49036_, new_n49035_, new_n49029_ );
not  ( new_n49037_, new_n49036_ );
xor  ( new_n49038_, new_n49019_, new_n49003_ );
and  ( new_n49039_, new_n49038_, new_n49037_ );
or   ( new_n49040_, new_n49039_, new_n49020_ );
xor  ( new_n49041_, new_n49001_, new_n49000_ );
and  ( new_n49042_, new_n49041_, new_n49040_ );
nor  ( new_n49043_, new_n49042_, new_n49002_ );
not  ( new_n49044_, new_n49043_ );
xor  ( new_n49045_, new_n48962_, new_n48960_ );
nand ( new_n49046_, new_n49045_, new_n49044_ );
and  ( new_n49047_, new_n49046_, new_n48963_ );
xor  ( new_n49048_, new_n48830_, new_n48817_ );
xor  ( new_n49049_, new_n49048_, new_n48848_ );
xnor ( new_n49050_, new_n48721_, new_n48705_ );
xor  ( new_n49051_, new_n49050_, new_n48725_ );
or   ( new_n49052_, new_n49051_, new_n49049_ );
nand ( new_n49053_, new_n49051_, new_n49049_ );
xor  ( new_n49054_, new_n48878_, new_n48876_ );
xor  ( new_n49055_, new_n49054_, new_n48882_ );
nand ( new_n49056_, new_n49055_, new_n49053_ );
and  ( new_n49057_, new_n49056_, new_n49052_ );
xor  ( new_n49058_, new_n48727_, new_n48704_ );
xor  ( new_n49059_, new_n49058_, new_n48773_ );
or   ( new_n49060_, new_n49059_, new_n49057_ );
and  ( new_n49061_, new_n49059_, new_n49057_ );
or   ( new_n49062_, new_n48759_, new_n2809_ );
xor  ( new_n49063_, new_n44218_, RIbb2e800_31 );
nand ( new_n49064_, new_n49063_, new_n2615_ );
and  ( new_n49065_, new_n49064_, new_n49062_ );
xor  ( new_n49066_, new_n43787_, new_n5203_ );
or   ( new_n49067_, new_n49066_, new_n5604_ );
or   ( new_n49068_, new_n48673_, new_n5606_ );
and  ( new_n49069_, new_n49068_, new_n49067_ );
nor  ( new_n49070_, new_n49069_, new_n49065_ );
nor  ( new_n49071_, new_n48732_, new_n4711_ );
xor  ( new_n49072_, new_n43803_, RIbb2e350_41 );
and  ( new_n49073_, new_n49072_, new_n4543_ );
or   ( new_n49074_, new_n49073_, new_n49071_ );
xor  ( new_n49075_, new_n49069_, new_n49065_ );
and  ( new_n49076_, new_n49075_, new_n49074_ );
or   ( new_n49077_, new_n49076_, new_n49070_ );
xor  ( new_n49078_, new_n48815_, new_n48814_ );
nand ( new_n49079_, new_n49078_, new_n49077_ );
xor  ( new_n49080_, new_n49078_, new_n49077_ );
xor  ( new_n49081_, new_n48828_, new_n48827_ );
nand ( new_n49082_, new_n49081_, new_n49080_ );
and  ( new_n49083_, new_n49082_, new_n49079_ );
xor  ( new_n49084_, new_n48746_, new_n48730_ );
xor  ( new_n49085_, new_n49084_, new_n48770_ );
nor  ( new_n49086_, new_n49085_, new_n49083_ );
and  ( new_n49087_, new_n49085_, new_n49083_ );
xor  ( new_n49088_, new_n48768_, new_n48767_ );
xnor ( new_n49089_, new_n48738_, new_n48734_ );
xor  ( new_n49090_, new_n49089_, new_n48743_ );
and  ( new_n49091_, new_n49090_, new_n49088_ );
xor  ( new_n49092_, new_n49090_, new_n49088_ );
xnor ( new_n49093_, new_n48840_, new_n48836_ );
xor  ( new_n49094_, new_n49093_, new_n48845_ );
and  ( new_n49095_, new_n49094_, new_n49092_ );
nor  ( new_n49096_, new_n49095_, new_n49091_ );
nor  ( new_n49097_, new_n49096_, new_n49087_ );
nor  ( new_n49098_, new_n49097_, new_n49086_ );
or   ( new_n49099_, new_n49098_, new_n49061_ );
and  ( new_n49100_, new_n49099_, new_n49060_ );
or   ( new_n49101_, new_n49100_, new_n49047_ );
nand ( new_n49102_, new_n49100_, new_n49047_ );
xor  ( new_n49103_, new_n48855_, new_n48799_ );
nand ( new_n49104_, new_n49103_, new_n49102_ );
and  ( new_n49105_, new_n49104_, new_n49101_ );
or   ( new_n49106_, new_n49105_, new_n48895_ );
and  ( new_n49107_, new_n49106_, new_n48894_ );
and  ( new_n49108_, new_n49107_, new_n48866_ );
xor  ( new_n49109_, new_n49107_, new_n48866_ );
xor  ( new_n49110_, new_n48785_, new_n48783_ );
and  ( new_n49111_, new_n49110_, new_n49109_ );
or   ( new_n49112_, new_n49111_, new_n49108_ );
xor  ( new_n49113_, new_n48788_, new_n48787_ );
nor  ( new_n49114_, new_n49113_, new_n49112_ );
and  ( new_n49115_, new_n49113_, new_n49112_ );
xor  ( new_n49116_, new_n49110_, new_n49109_ );
xor  ( new_n49117_, new_n48893_, new_n48868_ );
xor  ( new_n49118_, new_n49117_, new_n49105_ );
xnor ( new_n49119_, new_n48859_, new_n48857_ );
xor  ( new_n49120_, new_n49119_, new_n48862_ );
or   ( new_n49121_, new_n49120_, new_n49118_ );
and  ( new_n49122_, new_n49120_, new_n49118_ );
xor  ( new_n49123_, new_n48850_, new_n48801_ );
xor  ( new_n49124_, new_n49123_, new_n48852_ );
xnor ( new_n49125_, new_n48873_, new_n48871_ );
xor  ( new_n49126_, new_n49125_, new_n48885_ );
nand ( new_n49127_, new_n49126_, new_n49124_ );
or   ( new_n49128_, new_n49126_, new_n49124_ );
xor  ( new_n49129_, new_n49045_, new_n49044_ );
nand ( new_n49130_, new_n49129_, new_n49128_ );
and  ( new_n49131_, new_n49130_, new_n49127_ );
xor  ( new_n49132_, new_n48887_, new_n48869_ );
xor  ( new_n49133_, new_n49132_, new_n48891_ );
nor  ( new_n49134_, new_n49133_, new_n49131_ );
and  ( new_n49135_, new_n49133_, new_n49131_ );
not  ( new_n49136_, new_n49135_ );
nand ( new_n49137_, new_n49072_, new_n4541_ );
xor  ( new_n49138_, new_n43884_, new_n4292_ );
or   ( new_n49139_, new_n49138_, new_n4709_ );
and  ( new_n49140_, new_n49139_, new_n49137_ );
xor  ( new_n49141_, new_n44506_, new_n2118_ );
or   ( new_n49142_, new_n49141_, new_n2425_ );
nand ( new_n49143_, new_n48975_, new_n2242_ );
and  ( new_n49144_, new_n49143_, new_n49142_ );
nor  ( new_n49145_, new_n49144_, new_n49140_ );
and  ( new_n49146_, new_n49063_, new_n2613_ );
xor  ( new_n49147_, new_n44319_, RIbb2e800_31 );
and  ( new_n49148_, new_n49147_, new_n2615_ );
nor  ( new_n49149_, new_n49148_, new_n49146_ );
not  ( new_n49150_, new_n49149_ );
xor  ( new_n49151_, new_n49144_, new_n49140_ );
and  ( new_n49152_, new_n49151_, new_n49150_ );
nor  ( new_n49153_, new_n49152_, new_n49145_ );
not  ( new_n49154_, new_n49153_ );
xor  ( new_n49155_, new_n49034_, new_n49033_ );
and  ( new_n49156_, new_n49155_, new_n49154_ );
xor  ( new_n49157_, new_n49155_, new_n49154_ );
xnor ( new_n49158_, new_n49011_, new_n49007_ );
xor  ( new_n49159_, new_n49158_, new_n49016_ );
and  ( new_n49160_, new_n49159_, new_n49157_ );
nor  ( new_n49161_, new_n49160_, new_n49156_ );
not  ( new_n49162_, new_n49161_ );
xor  ( new_n49163_, new_n48998_, new_n48997_ );
and  ( new_n49164_, new_n49163_, new_n49162_ );
xor  ( new_n49165_, new_n49163_, new_n49162_ );
xor  ( new_n49166_, new_n49075_, new_n49074_ );
xnor ( new_n49167_, new_n48972_, new_n48968_ );
nand ( new_n49168_, new_n49167_, new_n48977_ );
not  ( new_n49169_, new_n48979_ );
or   ( new_n49170_, new_n49169_, new_n48973_ );
and  ( new_n49171_, new_n49170_, new_n49168_ );
or   ( new_n49172_, new_n49171_, new_n49166_ );
and  ( new_n49173_, new_n49171_, new_n49166_ );
xor  ( new_n49174_, new_n48995_, new_n48994_ );
or   ( new_n49175_, new_n49174_, new_n49173_ );
and  ( new_n49176_, new_n49175_, new_n49172_ );
and  ( new_n49177_, new_n49176_, new_n49165_ );
or   ( new_n49178_, new_n49177_, new_n49164_ );
xor  ( new_n49179_, new_n49041_, new_n49040_ );
and  ( new_n49180_, new_n49179_, new_n49178_ );
xor  ( new_n49181_, new_n49179_, new_n49178_ );
xnor ( new_n49182_, new_n49085_, new_n49083_ );
xor  ( new_n49183_, new_n49182_, new_n49096_ );
and  ( new_n49184_, new_n49183_, new_n49181_ );
nor  ( new_n49185_, new_n49184_, new_n49180_ );
xnor ( new_n49186_, new_n48958_, new_n48957_ );
xor  ( new_n49187_, new_n48955_, new_n48954_ );
xnor ( new_n49188_, new_n48713_, new_n48709_ );
nand ( new_n49189_, new_n49188_, new_n48719_ );
not  ( new_n49190_, new_n48720_ );
or   ( new_n49191_, new_n49190_, new_n48714_ );
and  ( new_n49192_, new_n49191_, new_n49189_ );
nand ( new_n49193_, new_n49192_, new_n49187_ );
nor  ( new_n49194_, new_n49192_, new_n49187_ );
and  ( new_n49195_, new_n48932_, new_n454_ );
xor  ( new_n49196_, new_n46619_, new_n400_ );
nor  ( new_n49197_, new_n49196_, new_n524_ );
nor  ( new_n49198_, new_n49197_, new_n49195_ );
or   ( new_n49199_, new_n48825_, new_n1137_ );
xor  ( new_n49200_, new_n45584_, RIbb2eda0_19 );
nand ( new_n49201_, new_n49200_, new_n1042_ );
and  ( new_n49202_, new_n49201_, new_n49199_ );
or   ( new_n49203_, new_n49202_, new_n49198_ );
or   ( new_n49204_, new_n48949_, new_n320_ );
xor  ( new_n49205_, new_n47296_, new_n309_ );
or   ( new_n49206_, new_n49205_, new_n317_ );
and  ( new_n49207_, new_n49206_, new_n49204_ );
or   ( new_n49208_, new_n48944_, new_n340_ );
xor  ( new_n49209_, new_n47303_, new_n329_ );
or   ( new_n49210_, new_n49209_, new_n337_ );
and  ( new_n49211_, new_n49210_, new_n49208_ );
nor  ( new_n49212_, new_n49211_, new_n49207_ );
nor  ( new_n49213_, new_n48926_, new_n411_ );
xor  ( new_n49214_, new_n46962_, new_n325_ );
nor  ( new_n49215_, new_n49214_, new_n409_ );
nor  ( new_n49216_, new_n49215_, new_n49213_ );
and  ( new_n49217_, new_n49211_, new_n49207_ );
nor  ( new_n49218_, new_n49217_, new_n49216_ );
or   ( new_n49219_, new_n49218_, new_n49212_ );
xor  ( new_n49220_, new_n49202_, new_n49198_ );
nand ( new_n49221_, new_n49220_, new_n49219_ );
and  ( new_n49222_, new_n49221_, new_n49203_ );
or   ( new_n49223_, new_n49222_, new_n49194_ );
and  ( new_n49224_, new_n49223_, new_n49193_ );
nor  ( new_n49225_, new_n49224_, new_n49186_ );
xor  ( new_n49226_, new_n48935_, new_n48934_ );
xor  ( new_n49227_, new_n48923_, new_n48922_ );
nand ( new_n49228_, new_n49227_, new_n49226_ );
or   ( new_n49229_, new_n49005_, new_n3463_ );
xor  ( new_n49230_, new_n43812_, new_n3113_ );
or   ( new_n49231_, new_n49230_, new_n3461_ );
and  ( new_n49232_, new_n49231_, new_n49229_ );
nand ( new_n49233_, new_n49014_, new_n1251_ );
xor  ( new_n49234_, new_n45403_, new_n1126_ );
or   ( new_n49235_, new_n49234_, new_n1364_ );
and  ( new_n49236_, new_n49235_, new_n49233_ );
nor  ( new_n49237_, new_n49236_, new_n49232_ );
xor  ( new_n49238_, new_n45738_, RIbb2eda0_19 );
and  ( new_n49239_, new_n49238_, new_n1042_ );
and  ( new_n49240_, new_n49200_, new_n1040_ );
or   ( new_n49241_, new_n49240_, new_n49239_ );
xor  ( new_n49242_, new_n49236_, new_n49232_ );
and  ( new_n49243_, new_n49242_, new_n49241_ );
or   ( new_n49244_, new_n49243_, new_n49237_ );
xor  ( new_n49245_, new_n49227_, new_n49226_ );
nand ( new_n49246_, new_n49245_, new_n49244_ );
and  ( new_n49247_, new_n49246_, new_n49228_ );
or   ( new_n49248_, new_n49066_, new_n5606_ );
xor  ( new_n49249_, new_n43898_, new_n5203_ );
or   ( new_n49250_, new_n49249_, new_n5604_ );
and  ( new_n49251_, new_n49250_, new_n49248_ );
or   ( new_n49252_, new_n48992_, new_n757_ );
xor  ( new_n49253_, new_n46137_, RIbb2ef80_15 );
nand ( new_n49254_, new_n49253_, new_n662_ );
and  ( new_n49255_, new_n49254_, new_n49252_ );
or   ( new_n49256_, new_n49255_, new_n49251_ );
and  ( new_n49257_, new_n48987_, new_n820_ );
xor  ( new_n49258_, new_n45928_, new_n745_ );
nor  ( new_n49259_, new_n49258_, new_n897_ );
or   ( new_n49260_, new_n49259_, new_n49257_ );
xor  ( new_n49261_, new_n49255_, new_n49251_ );
nand ( new_n49262_, new_n49261_, new_n49260_ );
and  ( new_n49263_, new_n49262_, new_n49256_ );
xor  ( new_n49264_, RIbb32b80_175, RIbb2c280_111 );
xor  ( new_n49265_, new_n49264_, new_n48751_ );
not  ( new_n49266_, new_n49265_ );
or   ( new_n49267_, new_n49266_, new_n43879_ );
xor  ( new_n49268_, new_n48908_, new_n43945_ );
not  ( new_n49269_, new_n49268_ );
or   ( new_n49270_, new_n49269_, new_n43983_ );
not  ( new_n49271_, new_n48756_ );
and  ( new_n49272_, new_n49271_, new_n43879_ );
or   ( new_n49273_, new_n48757_, new_n43977_ );
or   ( new_n49274_, new_n49273_, new_n49272_ );
and  ( new_n49275_, new_n49274_, new_n49270_ );
or   ( new_n49276_, new_n49275_, new_n49267_ );
and  ( new_n49277_, new_n49275_, new_n49267_ );
and  ( new_n49278_, new_n48982_, new_n2928_ );
xor  ( new_n49279_, new_n44183_, RIbb2e710_33 );
and  ( new_n49280_, new_n49279_, new_n2930_ );
nor  ( new_n49281_, new_n49280_, new_n49278_ );
or   ( new_n49282_, new_n49281_, new_n49277_ );
and  ( new_n49283_, new_n49282_, new_n49276_ );
or   ( new_n49284_, new_n49283_, new_n49263_ );
and  ( new_n49285_, new_n49283_, new_n49263_ );
xnor ( new_n49286_, new_n48952_, new_n48951_ );
or   ( new_n49287_, new_n49286_, new_n49285_ );
and  ( new_n49288_, new_n49287_, new_n49284_ );
nor  ( new_n49289_, new_n49288_, new_n49247_ );
or   ( new_n49290_, new_n48940_, new_n286_ );
xor  ( new_n49291_, new_n48039_, new_n275_ );
or   ( new_n49292_, new_n49291_, new_n283_ );
and  ( new_n49293_, new_n49292_, new_n49290_ );
nor  ( new_n49294_, RIbb2df90_49, RIbb2e008_48 );
or   ( new_n49295_, new_n49294_, new_n5597_ );
xor  ( new_n49296_, new_n43793_, RIbb2e080_47 );
or   ( new_n49297_, new_n49296_, new_n6173_ );
and  ( new_n49298_, new_n49297_, new_n49295_ );
or   ( new_n49299_, new_n49298_, new_n49293_ );
and  ( new_n49300_, new_n48919_, new_n295_ );
and  ( new_n49301_, new_n48677_, new_n43949_ );
or   ( new_n49302_, new_n49301_, new_n49300_ );
xor  ( new_n49303_, new_n49298_, new_n49293_ );
nand ( new_n49304_, new_n49303_, new_n49302_ );
and  ( new_n49305_, new_n49304_, new_n49299_ );
or   ( new_n49306_, new_n48965_, new_n4304_ );
xor  ( new_n49307_, new_n43937_, new_n3892_ );
or   ( new_n49308_, new_n49307_, new_n4302_ );
and  ( new_n49309_, new_n49308_, new_n49306_ );
or   ( new_n49310_, new_n49026_, new_n5209_ );
xor  ( new_n49311_, new_n43799_, new_n4705_ );
or   ( new_n49312_, new_n49311_, new_n5207_ );
and  ( new_n49313_, new_n49312_, new_n49310_ );
or   ( new_n49314_, new_n49313_, new_n49309_ );
xor  ( new_n49315_, new_n44681_, RIbb2e9e0_27 );
and  ( new_n49316_, new_n49315_, new_n2002_ );
and  ( new_n49317_, new_n48970_, new_n2000_ );
nor  ( new_n49318_, new_n49317_, new_n49316_ );
xnor ( new_n49319_, new_n49313_, new_n49309_ );
or   ( new_n49320_, new_n49319_, new_n49318_ );
and  ( new_n49321_, new_n49320_, new_n49314_ );
nor  ( new_n49322_, new_n49321_, new_n49305_ );
nand ( new_n49323_, new_n49031_, new_n1739_ );
xor  ( new_n49324_, new_n44877_, RIbb2ead0_25 );
nand ( new_n49325_, new_n49324_, new_n1741_ );
and  ( new_n49326_, new_n49325_, new_n49323_ );
or   ( new_n49327_, new_n49021_, new_n3898_ );
xor  ( new_n49328_, new_n43952_, new_n3457_ );
or   ( new_n49329_, new_n49328_, new_n3896_ );
and  ( new_n49330_, new_n49329_, new_n49327_ );
nor  ( new_n49331_, new_n49330_, new_n49326_ );
and  ( new_n49332_, new_n49009_, new_n1474_ );
xor  ( new_n49333_, new_n45119_, new_n1355_ );
nor  ( new_n49334_, new_n49333_, new_n1593_ );
nor  ( new_n49335_, new_n49334_, new_n49332_ );
not  ( new_n49336_, new_n49335_ );
xor  ( new_n49337_, new_n49330_, new_n49326_ );
and  ( new_n49338_, new_n49337_, new_n49336_ );
or   ( new_n49339_, new_n49338_, new_n49331_ );
xor  ( new_n49340_, new_n49321_, new_n49305_ );
and  ( new_n49341_, new_n49340_, new_n49339_ );
nor  ( new_n49342_, new_n49341_, new_n49322_ );
xnor ( new_n49343_, new_n49288_, new_n49247_ );
nor  ( new_n49344_, new_n49343_, new_n49342_ );
or   ( new_n49345_, new_n49344_, new_n49289_ );
xor  ( new_n49346_, new_n49224_, new_n49186_ );
and  ( new_n49347_, new_n49346_, new_n49345_ );
or   ( new_n49348_, new_n49347_, new_n49225_ );
xnor ( new_n49349_, new_n49059_, new_n49057_ );
xor  ( new_n49350_, new_n49349_, new_n49098_ );
and  ( new_n49351_, new_n49350_, new_n49348_ );
not  ( new_n49352_, new_n49351_ );
and  ( new_n49353_, new_n49352_, new_n49185_ );
nor  ( new_n49354_, new_n49350_, new_n49348_ );
nor  ( new_n49355_, new_n49354_, new_n49353_ );
and  ( new_n49356_, new_n49355_, new_n49136_ );
nor  ( new_n49357_, new_n49356_, new_n49134_ );
or   ( new_n49358_, new_n49357_, new_n49122_ );
and  ( new_n49359_, new_n49358_, new_n49121_ );
nor  ( new_n49360_, new_n49359_, new_n49116_ );
and  ( new_n49361_, new_n49359_, new_n49116_ );
xor  ( new_n49362_, new_n49100_, new_n49047_ );
xor  ( new_n49363_, new_n49362_, new_n49103_ );
xor  ( new_n49364_, new_n49133_, new_n49131_ );
xor  ( new_n49365_, new_n49364_, new_n49355_ );
and  ( new_n49366_, new_n49365_, new_n49363_ );
nor  ( new_n49367_, new_n49365_, new_n49363_ );
xnor ( new_n49368_, new_n49343_, new_n49342_ );
xnor ( new_n49369_, new_n49319_, new_n49318_ );
xor  ( new_n49370_, new_n43787_, new_n5594_ );
or   ( new_n49371_, new_n49370_, new_n6173_ );
or   ( new_n49372_, new_n49296_, new_n6175_ );
and  ( new_n49373_, new_n49372_, new_n49371_ );
nand ( new_n49374_, new_n49279_, new_n2928_ );
xor  ( new_n49375_, new_n44218_, new_n2797_ );
or   ( new_n49376_, new_n49375_, new_n3117_ );
and  ( new_n49377_, new_n49376_, new_n49374_ );
or   ( new_n49378_, new_n49377_, new_n49373_ );
nor  ( new_n49379_, new_n49258_, new_n899_ );
xor  ( new_n49380_, new_n46037_, new_n745_ );
nor  ( new_n49381_, new_n49380_, new_n897_ );
or   ( new_n49382_, new_n49381_, new_n49379_ );
xor  ( new_n49383_, new_n49377_, new_n49373_ );
nand ( new_n49384_, new_n49383_, new_n49382_ );
and  ( new_n49385_, new_n49384_, new_n49378_ );
and  ( new_n49386_, new_n49385_, new_n49369_ );
xor  ( new_n49387_, new_n49337_, new_n49336_ );
nor  ( new_n49388_, new_n49385_, new_n49369_ );
nor  ( new_n49389_, new_n49388_, new_n49387_ );
or   ( new_n49390_, new_n49389_, new_n49386_ );
xor  ( new_n49391_, new_n49283_, new_n49263_ );
xor  ( new_n49392_, new_n49391_, new_n49286_ );
or   ( new_n49393_, new_n49392_, new_n49390_ );
and  ( new_n49394_, new_n49392_, new_n49390_ );
xor  ( new_n49395_, new_n49261_, new_n49260_ );
xor  ( new_n49396_, new_n49242_, new_n49241_ );
nor  ( new_n49397_, new_n49396_, new_n49395_ );
xor  ( new_n49398_, new_n49151_, new_n49150_ );
and  ( new_n49399_, new_n49396_, new_n49395_ );
nor  ( new_n49400_, new_n49399_, new_n49398_ );
or   ( new_n49401_, new_n49400_, new_n49397_ );
or   ( new_n49402_, new_n49401_, new_n49394_ );
and  ( new_n49403_, new_n49402_, new_n49393_ );
nor  ( new_n49404_, new_n49403_, new_n49368_ );
xor  ( new_n49405_, new_n49176_, new_n49165_ );
xor  ( new_n49406_, new_n49403_, new_n49368_ );
and  ( new_n49407_, new_n49406_, new_n49405_ );
or   ( new_n49408_, new_n49407_, new_n49404_ );
xor  ( new_n49409_, new_n49346_, new_n49345_ );
and  ( new_n49410_, new_n49409_, new_n49408_ );
xor  ( new_n49411_, new_n49183_, new_n49181_ );
xor  ( new_n49412_, new_n49409_, new_n49408_ );
and  ( new_n49413_, new_n49412_, new_n49411_ );
or   ( new_n49414_, new_n49413_, new_n49410_ );
xor  ( new_n49415_, new_n49126_, new_n49124_ );
xor  ( new_n49416_, new_n49415_, new_n49129_ );
and  ( new_n49417_, new_n49416_, new_n49414_ );
nor  ( new_n49418_, new_n49416_, new_n49414_ );
xor  ( new_n49419_, new_n49038_, new_n49037_ );
xor  ( new_n49420_, new_n49081_, new_n49080_ );
and  ( new_n49421_, new_n49420_, new_n49419_ );
xor  ( new_n49422_, new_n49420_, new_n49419_ );
xor  ( new_n49423_, new_n49094_, new_n49092_ );
and  ( new_n49424_, new_n49423_, new_n49422_ );
nor  ( new_n49425_, new_n49424_, new_n49421_ );
xor  ( new_n49426_, RIbb32bf8_176, RIbb2c208_112 );
xor  ( new_n49427_, new_n49426_, new_n46409_ );
and  ( new_n49428_, new_n49427_, new_n43880_ );
nand ( new_n49429_, new_n49428_, new_n6166_ );
and  ( new_n49430_, new_n49253_, new_n660_ );
xor  ( new_n49431_, new_n46427_, RIbb2ef80_15 );
and  ( new_n49432_, new_n49431_, new_n662_ );
nor  ( new_n49433_, new_n49432_, new_n49430_ );
xor  ( new_n49434_, new_n49428_, new_n6165_ );
or   ( new_n49435_, new_n49434_, new_n49433_ );
nand ( new_n49436_, new_n49435_, new_n49429_ );
and  ( new_n49437_, new_n49436_, new_n49198_ );
xnor ( new_n49438_, new_n49436_, new_n49198_ );
or   ( new_n49439_, new_n49214_, new_n411_ );
xor  ( new_n49440_, new_n46958_, new_n325_ );
or   ( new_n49441_, new_n49440_, new_n409_ );
and  ( new_n49442_, new_n49441_, new_n49439_ );
or   ( new_n49443_, new_n49196_, new_n526_ );
xor  ( new_n49444_, new_n46789_, new_n400_ );
or   ( new_n49445_, new_n49444_, new_n524_ );
and  ( new_n49446_, new_n49445_, new_n49443_ );
nor  ( new_n49447_, new_n49446_, new_n49442_ );
and  ( new_n49448_, new_n49446_, new_n49442_ );
nor  ( new_n49449_, new_n49209_, new_n340_ );
xor  ( new_n49450_, new_n47046_, new_n329_ );
nor  ( new_n49451_, new_n49450_, new_n337_ );
nor  ( new_n49452_, new_n49451_, new_n49449_ );
nor  ( new_n49453_, new_n49452_, new_n49448_ );
nor  ( new_n49454_, new_n49453_, new_n49447_ );
nor  ( new_n49455_, new_n49454_, new_n49438_ );
or   ( new_n49456_, new_n49455_, new_n49437_ );
xor  ( new_n49457_, new_n49220_, new_n49219_ );
nand ( new_n49458_, new_n49457_, new_n49456_ );
xor  ( new_n49459_, new_n48291_, RIbb2f430_5 );
nand ( new_n49460_, new_n49459_, new_n282_ );
or   ( new_n49461_, new_n49291_, new_n286_ );
and  ( new_n49462_, new_n49461_, new_n49460_ );
or   ( new_n49463_, new_n49205_, new_n320_ );
xor  ( new_n49464_, new_n47640_, new_n309_ );
or   ( new_n49465_, new_n49464_, new_n317_ );
and  ( new_n49466_, new_n49465_, new_n49463_ );
nor  ( new_n49467_, new_n49466_, new_n49462_ );
and  ( new_n49468_, new_n48912_, new_n43949_ );
and  ( new_n49469_, new_n48677_, new_n295_ );
nor  ( new_n49470_, new_n49469_, new_n49468_ );
and  ( new_n49471_, new_n49466_, new_n49462_ );
nor  ( new_n49472_, new_n49471_, new_n49470_ );
nor  ( new_n49473_, new_n49472_, new_n49467_ );
xor  ( new_n49474_, RIbb32c70_177, RIbb2c190_113 );
nor  ( new_n49475_, new_n43618_, new_n43534_ );
not  ( new_n49476_, new_n49475_ );
and  ( new_n49477_, new_n49476_, new_n43512_ );
nor  ( new_n49478_, new_n49477_, new_n43546_ );
not  ( new_n49479_, new_n49478_ );
and  ( new_n49480_, new_n49479_, new_n43497_ );
nor  ( new_n49481_, new_n49480_, new_n43625_ );
not  ( new_n49482_, new_n49481_ );
and  ( new_n49483_, new_n49482_, new_n43500_ );
nor  ( new_n49484_, new_n49483_, new_n43624_ );
not  ( new_n49485_, new_n49484_ );
and  ( new_n49486_, new_n49485_, new_n43502_ );
nor  ( new_n49487_, new_n49486_, new_n43623_ );
xnor ( new_n49488_, new_n49487_, new_n49474_ );
and  ( new_n49489_, new_n49488_, new_n43880_ );
not  ( new_n49490_, new_n49489_ );
xor  ( new_n49491_, new_n43956_, new_n3892_ );
or   ( new_n49492_, new_n49491_, new_n4302_ );
or   ( new_n49493_, new_n49307_, new_n4304_ );
and  ( new_n49494_, new_n49493_, new_n49492_ );
or   ( new_n49495_, new_n49494_, new_n49490_ );
and  ( new_n49496_, new_n49324_, new_n1739_ );
xor  ( new_n49497_, new_n44974_, RIbb2ead0_25 );
and  ( new_n49498_, new_n49497_, new_n1741_ );
nor  ( new_n49499_, new_n49498_, new_n49496_ );
xor  ( new_n49500_, new_n49494_, new_n49489_ );
or   ( new_n49501_, new_n49500_, new_n49499_ );
and  ( new_n49502_, new_n49501_, new_n49495_ );
nor  ( new_n49503_, new_n49502_, new_n49473_ );
or   ( new_n49504_, new_n49138_, new_n4711_ );
xor  ( new_n49505_, new_n43888_, new_n4292_ );
or   ( new_n49506_, new_n49505_, new_n4709_ );
and  ( new_n49507_, new_n49506_, new_n49504_ );
or   ( new_n49508_, new_n49311_, new_n5209_ );
xor  ( new_n49509_, new_n43803_, RIbb2e260_43 );
nand ( new_n49510_, new_n49509_, new_n4960_ );
and  ( new_n49511_, new_n49510_, new_n49508_ );
nor  ( new_n49512_, new_n49511_, new_n49507_ );
and  ( new_n49513_, new_n49147_, new_n2613_ );
xor  ( new_n49514_, new_n44407_, RIbb2e800_31 );
and  ( new_n49515_, new_n49514_, new_n2615_ );
or   ( new_n49516_, new_n49515_, new_n49513_ );
xor  ( new_n49517_, new_n49511_, new_n49507_ );
and  ( new_n49518_, new_n49517_, new_n49516_ );
nor  ( new_n49519_, new_n49518_, new_n49512_ );
and  ( new_n49520_, new_n49502_, new_n49473_ );
nor  ( new_n49521_, new_n49520_, new_n49519_ );
or   ( new_n49522_, new_n49521_, new_n49503_ );
xor  ( new_n49523_, new_n49457_, new_n49456_ );
nand ( new_n49524_, new_n49523_, new_n49522_ );
and  ( new_n49525_, new_n49524_, new_n49458_ );
xor  ( new_n49526_, new_n49192_, new_n49187_ );
xor  ( new_n49527_, new_n49526_, new_n49222_ );
or   ( new_n49528_, new_n49527_, new_n49525_ );
and  ( new_n49529_, new_n49527_, new_n49525_ );
or   ( new_n49530_, new_n49230_, new_n3463_ );
xor  ( new_n49531_, new_n43914_, new_n3113_ );
or   ( new_n49532_, new_n49531_, new_n3461_ );
and  ( new_n49533_, new_n49532_, new_n49530_ );
xor  ( new_n49534_, new_n49265_, new_n43945_ );
nand ( new_n49535_, new_n49534_, new_n43982_ );
nor  ( new_n49536_, new_n48908_, new_n43880_ );
or   ( new_n49537_, new_n48909_, new_n43977_ );
or   ( new_n49538_, new_n49537_, new_n49536_ );
and  ( new_n49539_, new_n49538_, new_n49535_ );
nor  ( new_n49540_, new_n49539_, new_n49533_ );
xor  ( new_n49541_, new_n45597_, RIbb2eda0_19 );
and  ( new_n49542_, new_n49541_, new_n1042_ );
and  ( new_n49543_, new_n49238_, new_n1040_ );
nor  ( new_n49544_, new_n49543_, new_n49542_ );
not  ( new_n49545_, new_n49544_ );
xor  ( new_n49546_, new_n49539_, new_n49533_ );
and  ( new_n49547_, new_n49546_, new_n49545_ );
or   ( new_n49548_, new_n49547_, new_n49540_ );
xor  ( new_n49549_, new_n49303_, new_n49302_ );
and  ( new_n49550_, new_n49549_, new_n49548_ );
or   ( new_n49551_, new_n49549_, new_n49548_ );
or   ( new_n49552_, new_n49328_, new_n3898_ );
xor  ( new_n49553_, new_n43985_, new_n3457_ );
or   ( new_n49554_, new_n49553_, new_n3896_ );
and  ( new_n49555_, new_n49554_, new_n49552_ );
or   ( new_n49556_, new_n49333_, new_n1595_ );
xor  ( new_n49557_, new_n45204_, RIbb2ebc0_23 );
nand ( new_n49558_, new_n49557_, new_n1476_ );
and  ( new_n49559_, new_n49558_, new_n49556_ );
nor  ( new_n49560_, new_n49559_, new_n49555_ );
xor  ( new_n49561_, new_n45584_, RIbb2ecb0_21 );
and  ( new_n49562_, new_n49561_, new_n1253_ );
nor  ( new_n49563_, new_n49234_, new_n1366_ );
or   ( new_n49564_, new_n49563_, new_n49562_ );
xor  ( new_n49565_, new_n49559_, new_n49555_ );
and  ( new_n49566_, new_n49565_, new_n49564_ );
or   ( new_n49567_, new_n49566_, new_n49560_ );
and  ( new_n49568_, new_n49567_, new_n49551_ );
or   ( new_n49569_, new_n49568_, new_n49550_ );
or   ( new_n49570_, new_n49249_, new_n5606_ );
xor  ( new_n49571_, new_n43894_, new_n5203_ );
or   ( new_n49572_, new_n49571_, new_n5604_ );
and  ( new_n49573_, new_n49572_, new_n49570_ );
or   ( new_n49574_, new_n49141_, new_n2427_ );
xor  ( new_n49575_, new_n44600_, RIbb2e8f0_29 );
nand ( new_n49576_, new_n49575_, new_n2244_ );
and  ( new_n49577_, new_n49576_, new_n49574_ );
nor  ( new_n49578_, new_n49577_, new_n49573_ );
and  ( new_n49579_, new_n49315_, new_n2000_ );
xor  ( new_n49580_, new_n44785_, RIbb2e9e0_27 );
and  ( new_n49581_, new_n49580_, new_n2002_ );
nor  ( new_n49582_, new_n49581_, new_n49579_ );
and  ( new_n49583_, new_n49577_, new_n49573_ );
nor  ( new_n49584_, new_n49583_, new_n49582_ );
nor  ( new_n49585_, new_n49584_, new_n49578_ );
not  ( new_n49586_, new_n49585_ );
xnor ( new_n49587_, new_n49211_, new_n49207_ );
nand ( new_n49588_, new_n49587_, new_n49216_ );
not  ( new_n49589_, new_n49212_ );
nand ( new_n49590_, new_n49218_, new_n49589_ );
and  ( new_n49591_, new_n49590_, new_n49588_ );
xnor ( new_n49592_, new_n49275_, new_n49267_ );
xor  ( new_n49593_, new_n49592_, new_n49281_ );
and  ( new_n49594_, new_n49593_, new_n49591_ );
or   ( new_n49595_, new_n49594_, new_n49586_ );
or   ( new_n49596_, new_n49593_, new_n49591_ );
and  ( new_n49597_, new_n49596_, new_n49595_ );
and  ( new_n49598_, new_n49597_, new_n49569_ );
xor  ( new_n49599_, new_n49340_, new_n49339_ );
xor  ( new_n49600_, new_n49597_, new_n49569_ );
and  ( new_n49601_, new_n49600_, new_n49599_ );
nor  ( new_n49602_, new_n49601_, new_n49598_ );
or   ( new_n49603_, new_n49602_, new_n49529_ );
and  ( new_n49604_, new_n49603_, new_n49528_ );
nor  ( new_n49605_, new_n49604_, new_n49425_ );
xor  ( new_n49606_, new_n49604_, new_n49425_ );
xor  ( new_n49607_, new_n49051_, new_n49049_ );
xor  ( new_n49608_, new_n49607_, new_n49055_ );
and  ( new_n49609_, new_n49608_, new_n49606_ );
nor  ( new_n49610_, new_n49609_, new_n49605_ );
nor  ( new_n49611_, new_n49610_, new_n49418_ );
nor  ( new_n49612_, new_n49611_, new_n49417_ );
nor  ( new_n49613_, new_n49612_, new_n49367_ );
nor  ( new_n49614_, new_n49613_, new_n49366_ );
not  ( new_n49615_, new_n49614_ );
xnor ( new_n49616_, new_n49120_, new_n49118_ );
xor  ( new_n49617_, new_n49616_, new_n49357_ );
nor  ( new_n49618_, new_n49617_, new_n49615_ );
and  ( new_n49619_, new_n49617_, new_n49615_ );
xor  ( new_n49620_, new_n49608_, new_n49606_ );
not  ( new_n49621_, new_n49620_ );
xnor ( new_n49622_, new_n49423_, new_n49422_ );
xor  ( new_n49623_, new_n49245_, new_n49244_ );
xor  ( new_n49624_, new_n49171_, new_n49166_ );
xor  ( new_n49625_, new_n49624_, new_n49174_ );
nand ( new_n49626_, new_n49625_, new_n49623_ );
or   ( new_n49627_, new_n49625_, new_n49623_ );
xor  ( new_n49628_, new_n49159_, new_n49157_ );
nand ( new_n49629_, new_n49628_, new_n49627_ );
and  ( new_n49630_, new_n49629_, new_n49626_ );
or   ( new_n49631_, new_n49630_, new_n49622_ );
and  ( new_n49632_, new_n49630_, new_n49622_ );
xnor ( new_n49633_, new_n49434_, new_n49433_ );
or   ( new_n49634_, new_n49444_, new_n526_ );
xor  ( new_n49635_, new_n46962_, new_n400_ );
or   ( new_n49636_, new_n49635_, new_n524_ );
and  ( new_n49637_, new_n49636_, new_n49634_ );
xor  ( new_n49638_, new_n47303_, new_n325_ );
or   ( new_n49639_, new_n49638_, new_n409_ );
or   ( new_n49640_, new_n49440_, new_n411_ );
and  ( new_n49641_, new_n49640_, new_n49639_ );
or   ( new_n49642_, new_n49641_, new_n49637_ );
xor  ( new_n49643_, new_n46619_, new_n520_ );
nor  ( new_n49644_, new_n49643_, new_n755_ );
and  ( new_n49645_, new_n49431_, new_n660_ );
nor  ( new_n49646_, new_n49645_, new_n49644_ );
and  ( new_n49647_, new_n49641_, new_n49637_ );
or   ( new_n49648_, new_n49647_, new_n49646_ );
and  ( new_n49649_, new_n49648_, new_n49642_ );
nor  ( new_n49650_, new_n49649_, new_n49633_ );
xor  ( new_n49651_, new_n48039_, new_n309_ );
or   ( new_n49652_, new_n49651_, new_n317_ );
or   ( new_n49653_, new_n49464_, new_n320_ );
and  ( new_n49654_, new_n49653_, new_n49652_ );
or   ( new_n49655_, new_n49450_, new_n340_ );
xor  ( new_n49656_, new_n47296_, new_n329_ );
or   ( new_n49657_, new_n49656_, new_n337_ );
and  ( new_n49658_, new_n49657_, new_n49655_ );
nor  ( new_n49659_, new_n49658_, new_n49654_ );
and  ( new_n49660_, new_n49459_, new_n280_ );
xor  ( new_n49661_, new_n48518_, RIbb2f430_5 );
and  ( new_n49662_, new_n49661_, new_n282_ );
or   ( new_n49663_, new_n49662_, new_n49660_ );
xor  ( new_n49664_, new_n49658_, new_n49654_ );
and  ( new_n49665_, new_n49664_, new_n49663_ );
or   ( new_n49666_, new_n49665_, new_n49659_ );
xor  ( new_n49667_, new_n49649_, new_n49633_ );
and  ( new_n49668_, new_n49667_, new_n49666_ );
or   ( new_n49669_, new_n49668_, new_n49650_ );
xor  ( new_n49670_, new_n49454_, new_n49438_ );
and  ( new_n49671_, new_n49670_, new_n49669_ );
and  ( new_n49672_, new_n48912_, new_n295_ );
and  ( new_n49673_, new_n49269_, new_n43949_ );
nor  ( new_n49674_, new_n49673_, new_n49672_ );
xor  ( new_n49675_, new_n49427_, new_n43945_ );
not  ( new_n49676_, new_n49675_ );
or   ( new_n49677_, new_n49676_, new_n43983_ );
and  ( new_n49678_, new_n49266_, new_n43879_ );
nand ( new_n49679_, new_n49267_, new_n43978_ );
or   ( new_n49680_, new_n49679_, new_n49678_ );
and  ( new_n49681_, new_n49680_, new_n49677_ );
nor  ( new_n49682_, new_n49681_, new_n49674_ );
xnor ( new_n49683_, new_n49681_, new_n49674_ );
not  ( new_n49684_, RIbb2df18_50 );
and  ( new_n49685_, new_n6635_, new_n49684_ );
or   ( new_n49686_, new_n49685_, new_n6166_ );
xor  ( new_n49687_, new_n43793_, RIbb2df90_49 );
or   ( new_n49688_, new_n49687_, new_n6645_ );
and  ( new_n49689_, new_n49688_, new_n49686_ );
nor  ( new_n49690_, new_n49689_, new_n49683_ );
or   ( new_n49691_, new_n49690_, new_n49682_ );
xnor ( new_n49692_, new_n49466_, new_n49462_ );
nand ( new_n49693_, new_n49692_, new_n49470_ );
not  ( new_n49694_, new_n49472_ );
or   ( new_n49695_, new_n49694_, new_n49467_ );
and  ( new_n49696_, new_n49695_, new_n49693_ );
and  ( new_n49697_, new_n49696_, new_n49691_ );
xor  ( new_n49698_, new_n43799_, new_n5203_ );
or   ( new_n49699_, new_n49698_, new_n5604_ );
or   ( new_n49700_, new_n49571_, new_n5606_ );
and  ( new_n49701_, new_n49700_, new_n49699_ );
nand ( new_n49702_, new_n49580_, new_n2000_ );
xor  ( new_n49703_, new_n44877_, new_n1840_ );
or   ( new_n49704_, new_n49703_, new_n2122_ );
and  ( new_n49705_, new_n49704_, new_n49702_ );
nor  ( new_n49706_, new_n49705_, new_n49701_ );
xor  ( new_n49707_, new_n44681_, RIbb2e8f0_29 );
and  ( new_n49708_, new_n49707_, new_n2244_ );
and  ( new_n49709_, new_n49575_, new_n2242_ );
or   ( new_n49710_, new_n49709_, new_n49708_ );
xor  ( new_n49711_, new_n49705_, new_n49701_ );
and  ( new_n49712_, new_n49711_, new_n49710_ );
or   ( new_n49713_, new_n49712_, new_n49706_ );
xor  ( new_n49714_, new_n49696_, new_n49691_ );
and  ( new_n49715_, new_n49714_, new_n49713_ );
or   ( new_n49716_, new_n49715_, new_n49697_ );
xor  ( new_n49717_, new_n49670_, new_n49669_ );
and  ( new_n49718_, new_n49717_, new_n49716_ );
or   ( new_n49719_, new_n49718_, new_n49671_ );
xor  ( new_n49720_, new_n49523_, new_n49522_ );
nand ( new_n49721_, new_n49720_, new_n49719_ );
or   ( new_n49722_, new_n49531_, new_n3463_ );
xor  ( new_n49723_, new_n44183_, RIbb2e620_35 );
nand ( new_n49724_, new_n49723_, new_n3293_ );
and  ( new_n49725_, new_n49724_, new_n49722_ );
or   ( new_n49726_, new_n49380_, new_n899_ );
xor  ( new_n49727_, new_n46137_, RIbb2ee90_17 );
nand ( new_n49728_, new_n49727_, new_n822_ );
and  ( new_n49729_, new_n49728_, new_n49726_ );
nor  ( new_n49730_, new_n49729_, new_n49725_ );
and  ( new_n49731_, new_n49541_, new_n1040_ );
xor  ( new_n49732_, new_n45928_, new_n893_ );
nor  ( new_n49733_, new_n49732_, new_n1135_ );
or   ( new_n49734_, new_n49733_, new_n49731_ );
xor  ( new_n49735_, new_n49729_, new_n49725_ );
and  ( new_n49736_, new_n49735_, new_n49734_ );
nor  ( new_n49737_, new_n49736_, new_n49730_ );
not  ( new_n49738_, new_n49737_ );
xor  ( new_n49739_, new_n43952_, new_n3892_ );
or   ( new_n49740_, new_n49739_, new_n4302_ );
or   ( new_n49741_, new_n49491_, new_n4304_ );
and  ( new_n49742_, new_n49741_, new_n49740_ );
xor  ( new_n49743_, new_n43812_, RIbb2e530_37 );
nand ( new_n49744_, new_n49743_, new_n3733_ );
or   ( new_n49745_, new_n49553_, new_n3898_ );
and  ( new_n49746_, new_n49745_, new_n49744_ );
nor  ( new_n49747_, new_n49746_, new_n49742_ );
and  ( new_n49748_, new_n49497_, new_n1739_ );
xor  ( new_n49749_, new_n45119_, new_n1583_ );
nor  ( new_n49750_, new_n49749_, new_n1844_ );
or   ( new_n49751_, new_n49750_, new_n49748_ );
xor  ( new_n49752_, new_n49746_, new_n49742_ );
and  ( new_n49753_, new_n49752_, new_n49751_ );
nor  ( new_n49754_, new_n49753_, new_n49747_ );
not  ( new_n49755_, new_n49754_ );
and  ( new_n49756_, new_n49755_, new_n49738_ );
xor  ( new_n49757_, RIbb32ce8_178, RIbb2c118_114 );
xor  ( new_n49758_, new_n49757_, new_n49485_ );
and  ( new_n49759_, new_n49758_, new_n43880_ );
nand ( new_n49760_, new_n49759_, new_n6638_ );
xor  ( new_n49761_, new_n49759_, new_n6637_ );
xor  ( new_n49762_, new_n49488_, new_n43945_ );
not  ( new_n49763_, new_n49762_ );
or   ( new_n49764_, new_n49763_, new_n43983_ );
nor  ( new_n49765_, new_n49427_, new_n43880_ );
or   ( new_n49766_, new_n49428_, new_n43977_ );
or   ( new_n49767_, new_n49766_, new_n49765_ );
and  ( new_n49768_, new_n49767_, new_n49764_ );
or   ( new_n49769_, new_n49768_, new_n49761_ );
and  ( new_n49770_, new_n49769_, new_n49760_ );
nand ( new_n49771_, new_n49561_, new_n1251_ );
xor  ( new_n49772_, new_n45738_, RIbb2ecb0_21 );
nand ( new_n49773_, new_n49772_, new_n1253_ );
and  ( new_n49774_, new_n49773_, new_n49771_ );
nor  ( new_n49775_, new_n49774_, new_n49770_ );
and  ( new_n49776_, new_n49557_, new_n1474_ );
xor  ( new_n49777_, new_n45403_, new_n1355_ );
nor  ( new_n49778_, new_n49777_, new_n1593_ );
or   ( new_n49779_, new_n49778_, new_n49776_ );
xor  ( new_n49780_, new_n49774_, new_n49770_ );
and  ( new_n49781_, new_n49780_, new_n49779_ );
nor  ( new_n49782_, new_n49781_, new_n49775_ );
and  ( new_n49783_, new_n49754_, new_n49737_ );
nor  ( new_n49784_, new_n49783_, new_n49782_ );
nor  ( new_n49785_, new_n49784_, new_n49756_ );
xor  ( new_n49786_, new_n49546_, new_n49545_ );
xor  ( new_n49787_, new_n49517_, new_n49516_ );
nand ( new_n49788_, new_n49787_, new_n49786_ );
xor  ( new_n49789_, new_n49787_, new_n49786_ );
xor  ( new_n49790_, new_n49565_, new_n49564_ );
nand ( new_n49791_, new_n49790_, new_n49789_ );
and  ( new_n49792_, new_n49791_, new_n49788_ );
nor  ( new_n49793_, new_n49792_, new_n49785_ );
xor  ( new_n49794_, new_n49792_, new_n49785_ );
xor  ( new_n49795_, new_n49549_, new_n49548_ );
xor  ( new_n49796_, new_n49795_, new_n49567_ );
and  ( new_n49797_, new_n49796_, new_n49794_ );
or   ( new_n49798_, new_n49797_, new_n49793_ );
xor  ( new_n49799_, new_n49720_, new_n49719_ );
nand ( new_n49800_, new_n49799_, new_n49798_ );
and  ( new_n49801_, new_n49800_, new_n49721_ );
or   ( new_n49802_, new_n49801_, new_n49632_ );
and  ( new_n49803_, new_n49802_, new_n49631_ );
nor  ( new_n49804_, new_n49803_, new_n49621_ );
xor  ( new_n49805_, new_n49803_, new_n49621_ );
not  ( new_n49806_, new_n49805_ );
xor  ( new_n49807_, new_n43937_, RIbb2e350_41 );
nand ( new_n49808_, new_n49807_, new_n4543_ );
or   ( new_n49809_, new_n49505_, new_n4711_ );
and  ( new_n49810_, new_n49809_, new_n49808_ );
nor  ( new_n49811_, new_n49810_, new_n49489_ );
xor  ( new_n49812_, new_n44506_, RIbb2e800_31 );
and  ( new_n49813_, new_n49812_, new_n2615_ );
and  ( new_n49814_, new_n49514_, new_n2613_ );
or   ( new_n49815_, new_n49814_, new_n49813_ );
xor  ( new_n49816_, new_n49810_, new_n49489_ );
and  ( new_n49817_, new_n49816_, new_n49815_ );
or   ( new_n49818_, new_n49817_, new_n49811_ );
xnor ( new_n49819_, new_n49446_, new_n49442_ );
nand ( new_n49820_, new_n49819_, new_n49452_ );
not  ( new_n49821_, new_n49453_ );
or   ( new_n49822_, new_n49821_, new_n49447_ );
and  ( new_n49823_, new_n49822_, new_n49820_ );
and  ( new_n49824_, new_n49823_, new_n49818_ );
xor  ( new_n49825_, new_n43898_, new_n5594_ );
or   ( new_n49826_, new_n49825_, new_n6173_ );
or   ( new_n49827_, new_n49370_, new_n6175_ );
and  ( new_n49828_, new_n49827_, new_n49826_ );
or   ( new_n49829_, new_n49375_, new_n3119_ );
xor  ( new_n49830_, new_n44319_, new_n2797_ );
or   ( new_n49831_, new_n49830_, new_n3117_ );
and  ( new_n49832_, new_n49831_, new_n49829_ );
nor  ( new_n49833_, new_n49832_, new_n49828_ );
xor  ( new_n49834_, new_n43884_, RIbb2e260_43 );
and  ( new_n49835_, new_n49834_, new_n4960_ );
and  ( new_n49836_, new_n49509_, new_n4958_ );
or   ( new_n49837_, new_n49836_, new_n49835_ );
xor  ( new_n49838_, new_n49832_, new_n49828_ );
and  ( new_n49839_, new_n49838_, new_n49837_ );
or   ( new_n49840_, new_n49839_, new_n49833_ );
xor  ( new_n49841_, new_n49823_, new_n49818_ );
and  ( new_n49842_, new_n49841_, new_n49840_ );
or   ( new_n49843_, new_n49842_, new_n49824_ );
xnor ( new_n49844_, new_n49502_, new_n49473_ );
nand ( new_n49845_, new_n49844_, new_n49519_ );
not  ( new_n49846_, new_n49503_ );
nand ( new_n49847_, new_n49521_, new_n49846_ );
and  ( new_n49848_, new_n49847_, new_n49845_ );
nor  ( new_n49849_, new_n49848_, new_n49843_ );
nand ( new_n49850_, new_n49848_, new_n49843_ );
xor  ( new_n49851_, new_n49383_, new_n49382_ );
xnor ( new_n49852_, new_n49577_, new_n49573_ );
xor  ( new_n49853_, new_n49852_, new_n49582_ );
nor  ( new_n49854_, new_n49853_, new_n49851_ );
nand ( new_n49855_, new_n49853_, new_n49851_ );
xnor ( new_n49856_, new_n49500_, new_n49499_ );
and  ( new_n49857_, new_n49856_, new_n49855_ );
or   ( new_n49858_, new_n49857_, new_n49854_ );
and  ( new_n49859_, new_n49858_, new_n49850_ );
or   ( new_n49860_, new_n49859_, new_n49849_ );
xor  ( new_n49861_, new_n49392_, new_n49390_ );
xor  ( new_n49862_, new_n49861_, new_n49401_ );
nand ( new_n49863_, new_n49862_, new_n49860_ );
nor  ( new_n49864_, new_n49862_, new_n49860_ );
xor  ( new_n49865_, new_n49600_, new_n49599_ );
or   ( new_n49866_, new_n49865_, new_n49864_ );
and  ( new_n49867_, new_n49866_, new_n49863_ );
xnor ( new_n49868_, new_n49527_, new_n49525_ );
xor  ( new_n49869_, new_n49868_, new_n49602_ );
nand ( new_n49870_, new_n49869_, new_n49867_ );
nor  ( new_n49871_, new_n49869_, new_n49867_ );
xnor ( new_n49872_, new_n49406_, new_n49405_ );
or   ( new_n49873_, new_n49872_, new_n49871_ );
and  ( new_n49874_, new_n49873_, new_n49870_ );
nor  ( new_n49875_, new_n49874_, new_n49806_ );
nor  ( new_n49876_, new_n49875_, new_n49804_ );
xor  ( new_n49877_, new_n49350_, new_n49348_ );
xor  ( new_n49878_, new_n49877_, new_n49185_ );
and  ( new_n49879_, new_n49878_, new_n49876_ );
xnor ( new_n49880_, new_n49878_, new_n49876_ );
xnor ( new_n49881_, new_n49416_, new_n49414_ );
xor  ( new_n49882_, new_n49881_, new_n49610_ );
nor  ( new_n49883_, new_n49882_, new_n49880_ );
nor  ( new_n49884_, new_n49883_, new_n49879_ );
xor  ( new_n49885_, new_n49365_, new_n49363_ );
xnor ( new_n49886_, new_n49885_, new_n49612_ );
nor  ( new_n49887_, new_n49886_, new_n49884_ );
and  ( new_n49888_, new_n49886_, new_n49884_ );
xor  ( new_n49889_, new_n49874_, new_n49806_ );
xor  ( new_n49890_, new_n49412_, new_n49411_ );
and  ( new_n49891_, new_n49890_, new_n49889_ );
xor  ( new_n49892_, new_n49890_, new_n49889_ );
not  ( new_n49893_, new_n49892_ );
xor  ( new_n49894_, new_n49385_, new_n49369_ );
xor  ( new_n49895_, new_n49894_, new_n49387_ );
xor  ( new_n49896_, new_n49396_, new_n49395_ );
xor  ( new_n49897_, new_n49896_, new_n49398_ );
or   ( new_n49898_, new_n49897_, new_n49895_ );
and  ( new_n49899_, new_n49897_, new_n49895_ );
xor  ( new_n49900_, new_n49593_, new_n49591_ );
xor  ( new_n49901_, new_n49900_, new_n49586_ );
or   ( new_n49902_, new_n49901_, new_n49899_ );
and  ( new_n49903_, new_n49902_, new_n49898_ );
xor  ( new_n49904_, new_n49625_, new_n49623_ );
xor  ( new_n49905_, new_n49904_, new_n49628_ );
nand ( new_n49906_, new_n49905_, new_n49903_ );
xor  ( new_n49907_, new_n49905_, new_n49903_ );
xor  ( new_n49908_, new_n49799_, new_n49798_ );
nand ( new_n49909_, new_n49908_, new_n49907_ );
and  ( new_n49910_, new_n49909_, new_n49906_ );
xor  ( new_n49911_, new_n49630_, new_n49622_ );
xor  ( new_n49912_, new_n49911_, new_n49801_ );
or   ( new_n49913_, new_n49912_, new_n49910_ );
and  ( new_n49914_, new_n49912_, new_n49910_ );
xor  ( new_n49915_, new_n43888_, new_n4705_ );
or   ( new_n49916_, new_n49915_, new_n5207_ );
nand ( new_n49917_, new_n49834_, new_n4958_ );
and  ( new_n49918_, new_n49917_, new_n49916_ );
xor  ( new_n49919_, new_n44600_, new_n2421_ );
or   ( new_n49920_, new_n49919_, new_n2807_ );
nand ( new_n49921_, new_n49812_, new_n2613_ );
and  ( new_n49922_, new_n49921_, new_n49920_ );
nor  ( new_n49923_, new_n49922_, new_n49918_ );
and  ( new_n49924_, new_n49922_, new_n49918_ );
xor  ( new_n49925_, new_n43894_, RIbb2e080_47 );
and  ( new_n49926_, new_n49925_, new_n5917_ );
nor  ( new_n49927_, new_n49825_, new_n6175_ );
nor  ( new_n49928_, new_n49927_, new_n49926_ );
nor  ( new_n49929_, new_n49928_, new_n49924_ );
nor  ( new_n49930_, new_n49929_, new_n49923_ );
xor  ( new_n49931_, new_n44974_, RIbb2e9e0_27 );
nand ( new_n49932_, new_n49931_, new_n2002_ );
or   ( new_n49933_, new_n49703_, new_n2124_ );
and  ( new_n49934_, new_n49933_, new_n49932_ );
xor  ( new_n49935_, new_n44785_, RIbb2e8f0_29 );
nand ( new_n49936_, new_n49935_, new_n2244_ );
nand ( new_n49937_, new_n49707_, new_n2242_ );
and  ( new_n49938_, new_n49937_, new_n49936_ );
nor  ( new_n49939_, new_n49938_, new_n49934_ );
and  ( new_n49940_, new_n49938_, new_n49934_ );
xor  ( new_n49941_, new_n43956_, new_n4292_ );
nor  ( new_n49942_, new_n49941_, new_n4709_ );
and  ( new_n49943_, new_n49807_, new_n4541_ );
nor  ( new_n49944_, new_n49943_, new_n49942_ );
nor  ( new_n49945_, new_n49944_, new_n49940_ );
nor  ( new_n49946_, new_n49945_, new_n49939_ );
nor  ( new_n49947_, new_n49946_, new_n49930_ );
xor  ( new_n49948_, new_n43803_, new_n5203_ );
or   ( new_n49949_, new_n49948_, new_n5604_ );
or   ( new_n49950_, new_n49698_, new_n5606_ );
and  ( new_n49951_, new_n49950_, new_n49949_ );
xor  ( new_n49952_, new_n44407_, RIbb2e710_33 );
nand ( new_n49953_, new_n49952_, new_n2930_ );
or   ( new_n49954_, new_n49830_, new_n3119_ );
and  ( new_n49955_, new_n49954_, new_n49953_ );
nor  ( new_n49956_, new_n49955_, new_n49951_ );
and  ( new_n49957_, new_n49723_, new_n3291_ );
xor  ( new_n49958_, new_n44218_, RIbb2e620_35 );
and  ( new_n49959_, new_n49958_, new_n3293_ );
or   ( new_n49960_, new_n49959_, new_n49957_ );
xor  ( new_n49961_, new_n49955_, new_n49951_ );
and  ( new_n49962_, new_n49961_, new_n49960_ );
nor  ( new_n49963_, new_n49962_, new_n49956_ );
and  ( new_n49964_, new_n49946_, new_n49930_ );
nor  ( new_n49965_, new_n49964_, new_n49963_ );
or   ( new_n49966_, new_n49965_, new_n49947_ );
xor  ( new_n49967_, new_n49667_, new_n49666_ );
and  ( new_n49968_, new_n49967_, new_n49966_ );
xor  ( new_n49969_, new_n49689_, new_n49683_ );
xnor ( new_n49970_, new_n49641_, new_n49637_ );
xor  ( new_n49971_, new_n49970_, new_n49646_ );
and  ( new_n49972_, new_n49971_, new_n49969_ );
or   ( new_n49973_, new_n49739_, new_n4304_ );
xor  ( new_n49974_, new_n43985_, new_n3892_ );
or   ( new_n49975_, new_n49974_, new_n4302_ );
and  ( new_n49976_, new_n49975_, new_n49973_ );
xor  ( new_n49977_, new_n49758_, new_n43945_ );
and  ( new_n49978_, new_n49977_, new_n43982_ );
not  ( new_n49979_, new_n49488_ );
and  ( new_n49980_, new_n49979_, new_n43879_ );
not  ( new_n49981_, new_n49980_ );
and  ( new_n49982_, new_n49490_, new_n43978_ );
and  ( new_n49983_, new_n49982_, new_n49981_ );
nor  ( new_n49984_, new_n49983_, new_n49978_ );
nor  ( new_n49985_, new_n49984_, new_n49976_ );
nor  ( new_n49986_, new_n49749_, new_n1846_ );
xor  ( new_n49987_, new_n45204_, RIbb2ead0_25 );
and  ( new_n49988_, new_n49987_, new_n1741_ );
or   ( new_n49989_, new_n49988_, new_n49986_ );
xor  ( new_n49990_, new_n49984_, new_n49976_ );
and  ( new_n49991_, new_n49990_, new_n49989_ );
nor  ( new_n49992_, new_n49991_, new_n49985_ );
not  ( new_n49993_, new_n49992_ );
xor  ( new_n49994_, new_n49971_, new_n49969_ );
and  ( new_n49995_, new_n49994_, new_n49993_ );
or   ( new_n49996_, new_n49995_, new_n49972_ );
xor  ( new_n49997_, new_n49967_, new_n49966_ );
and  ( new_n49998_, new_n49997_, new_n49996_ );
or   ( new_n49999_, new_n49998_, new_n49968_ );
xor  ( new_n50000_, new_n49717_, new_n49716_ );
nand ( new_n50001_, new_n50000_, new_n49999_ );
xor  ( new_n50002_, new_n48291_, new_n309_ );
or   ( new_n50003_, new_n50002_, new_n317_ );
or   ( new_n50004_, new_n49651_, new_n320_ );
and  ( new_n50005_, new_n50004_, new_n50003_ );
xor  ( new_n50006_, new_n47640_, new_n329_ );
or   ( new_n50007_, new_n50006_, new_n337_ );
or   ( new_n50008_, new_n49656_, new_n340_ );
and  ( new_n50009_, new_n50008_, new_n50007_ );
or   ( new_n50010_, new_n50009_, new_n50005_ );
nor  ( new_n50011_, new_n49638_, new_n411_ );
xor  ( new_n50012_, new_n47046_, new_n325_ );
nor  ( new_n50013_, new_n50012_, new_n409_ );
or   ( new_n50014_, new_n50013_, new_n50011_ );
xor  ( new_n50015_, new_n50009_, new_n50005_ );
nand ( new_n50016_, new_n50015_, new_n50014_ );
and  ( new_n50017_, new_n50016_, new_n50010_ );
xor  ( new_n50018_, new_n46958_, new_n400_ );
or   ( new_n50019_, new_n50018_, new_n524_ );
or   ( new_n50020_, new_n49635_, new_n526_ );
and  ( new_n50021_, new_n50020_, new_n50019_ );
xor  ( new_n50022_, new_n46789_, new_n520_ );
or   ( new_n50023_, new_n50022_, new_n755_ );
or   ( new_n50024_, new_n49643_, new_n757_ );
and  ( new_n50025_, new_n50024_, new_n50023_ );
or   ( new_n50026_, new_n50025_, new_n50021_ );
and  ( new_n50027_, new_n49727_, new_n820_ );
xor  ( new_n50028_, new_n46427_, RIbb2ee90_17 );
and  ( new_n50029_, new_n50028_, new_n822_ );
or   ( new_n50030_, new_n50029_, new_n50027_ );
xor  ( new_n50031_, new_n50025_, new_n50021_ );
nand ( new_n50032_, new_n50031_, new_n50030_ );
and  ( new_n50033_, new_n50032_, new_n50026_ );
nor  ( new_n50034_, new_n50033_, new_n50017_ );
xor  ( new_n50035_, new_n43787_, new_n6163_ );
or   ( new_n50036_, new_n50035_, new_n6645_ );
or   ( new_n50037_, new_n49687_, new_n6647_ );
and  ( new_n50038_, new_n50037_, new_n50036_ );
or   ( new_n50039_, new_n49732_, new_n1137_ );
xor  ( new_n50040_, new_n46037_, new_n893_ );
or   ( new_n50041_, new_n50040_, new_n1135_ );
and  ( new_n50042_, new_n50041_, new_n50039_ );
nor  ( new_n50043_, new_n50042_, new_n50038_ );
and  ( new_n50044_, new_n49772_, new_n1251_ );
xor  ( new_n50045_, new_n45597_, RIbb2ecb0_21 );
and  ( new_n50046_, new_n50045_, new_n1253_ );
or   ( new_n50047_, new_n50046_, new_n50044_ );
xor  ( new_n50048_, new_n50042_, new_n50038_ );
and  ( new_n50049_, new_n50048_, new_n50047_ );
nor  ( new_n50050_, new_n50049_, new_n50043_ );
xnor ( new_n50051_, new_n50033_, new_n50017_ );
nor  ( new_n50052_, new_n50051_, new_n50050_ );
or   ( new_n50053_, new_n50052_, new_n50034_ );
xor  ( new_n50054_, new_n49714_, new_n49713_ );
and  ( new_n50055_, new_n50054_, new_n50053_ );
xor  ( new_n50056_, new_n50054_, new_n50053_ );
xor  ( new_n50057_, new_n49754_, new_n49738_ );
nand ( new_n50058_, new_n50057_, new_n49782_ );
or   ( new_n50059_, new_n49783_, new_n49782_ );
or   ( new_n50060_, new_n50059_, new_n49756_ );
and  ( new_n50061_, new_n50060_, new_n50058_ );
and  ( new_n50062_, new_n50061_, new_n50056_ );
or   ( new_n50063_, new_n50062_, new_n50055_ );
xor  ( new_n50064_, new_n50000_, new_n49999_ );
nand ( new_n50065_, new_n50064_, new_n50063_ );
and  ( new_n50066_, new_n50065_, new_n50001_ );
xor  ( new_n50067_, new_n48756_, new_n275_ );
or   ( new_n50068_, new_n50067_, new_n283_ );
nand ( new_n50069_, new_n49661_, new_n280_ );
and  ( new_n50070_, new_n50069_, new_n50068_ );
or   ( new_n50071_, new_n49534_, new_n44007_ );
or   ( new_n50072_, new_n49268_, new_n302_ );
and  ( new_n50073_, new_n50072_, new_n50071_ );
nor  ( new_n50074_, new_n50073_, new_n50070_ );
nand ( new_n50075_, new_n50073_, new_n50070_ );
xor  ( new_n50076_, new_n43914_, RIbb2e530_37 );
and  ( new_n50077_, new_n50076_, new_n3733_ );
and  ( new_n50078_, new_n49743_, new_n3731_ );
or   ( new_n50079_, new_n50078_, new_n50077_ );
and  ( new_n50080_, new_n50079_, new_n50075_ );
or   ( new_n50081_, new_n50080_, new_n50074_ );
xor  ( new_n50082_, new_n49664_, new_n49663_ );
nand ( new_n50083_, new_n50082_, new_n50081_ );
xor  ( new_n50084_, new_n50082_, new_n50081_ );
xor  ( new_n50085_, new_n49752_, new_n49751_ );
nand ( new_n50086_, new_n50085_, new_n50084_ );
and  ( new_n50087_, new_n50086_, new_n50083_ );
xor  ( new_n50088_, new_n49816_, new_n49815_ );
xor  ( new_n50089_, new_n49711_, new_n49710_ );
nand ( new_n50090_, new_n50089_, new_n50088_ );
xor  ( new_n50091_, new_n50089_, new_n50088_ );
xor  ( new_n50092_, new_n49838_, new_n49837_ );
nand ( new_n50093_, new_n50092_, new_n50091_ );
and  ( new_n50094_, new_n50093_, new_n50090_ );
nor  ( new_n50095_, new_n50094_, new_n50087_ );
xor  ( new_n50096_, new_n49841_, new_n49840_ );
xor  ( new_n50097_, new_n50094_, new_n50087_ );
and  ( new_n50098_, new_n50097_, new_n50096_ );
or   ( new_n50099_, new_n50098_, new_n50095_ );
xor  ( new_n50100_, new_n49796_, new_n49794_ );
nand ( new_n50101_, new_n50100_, new_n50099_ );
nor  ( new_n50102_, new_n50100_, new_n50099_ );
xnor ( new_n50103_, new_n49790_, new_n49789_ );
xor  ( new_n50104_, new_n49853_, new_n49851_ );
xor  ( new_n50105_, new_n50104_, new_n49856_ );
nor  ( new_n50106_, new_n50105_, new_n50103_ );
and  ( new_n50107_, new_n50105_, new_n50103_ );
nor  ( new_n50108_, new_n49777_, new_n1595_ );
xor  ( new_n50109_, new_n45584_, RIbb2ebc0_23 );
and  ( new_n50110_, new_n50109_, new_n1476_ );
or   ( new_n50111_, new_n50110_, new_n50108_ );
xor  ( new_n50112_, new_n49768_, new_n49761_ );
and  ( new_n50113_, new_n50112_, new_n50111_ );
xor  ( new_n50114_, RIbb32d60_179, RIbb2c0a0_115 );
xor  ( new_n50115_, new_n50114_, new_n49482_ );
and  ( new_n50116_, new_n50115_, new_n43880_ );
not  ( new_n50117_, new_n50116_ );
nand ( new_n50118_, new_n50028_, new_n820_ );
xor  ( new_n50119_, new_n46619_, new_n745_ );
or   ( new_n50120_, new_n50119_, new_n897_ );
and  ( new_n50121_, new_n50120_, new_n50118_ );
nor  ( new_n50122_, new_n50121_, new_n50117_ );
nor  ( new_n50123_, new_n50022_, new_n757_ );
xor  ( new_n50124_, new_n46962_, new_n520_ );
nor  ( new_n50125_, new_n50124_, new_n755_ );
or   ( new_n50126_, new_n50125_, new_n50123_ );
xor  ( new_n50127_, new_n50121_, new_n50117_ );
and  ( new_n50128_, new_n50127_, new_n50126_ );
or   ( new_n50129_, new_n50128_, new_n50122_ );
xor  ( new_n50130_, new_n50112_, new_n50111_ );
and  ( new_n50131_, new_n50130_, new_n50129_ );
or   ( new_n50132_, new_n50131_, new_n50113_ );
xor  ( new_n50133_, new_n49780_, new_n49779_ );
and  ( new_n50134_, new_n50133_, new_n50132_ );
xor  ( new_n50135_, new_n50133_, new_n50132_ );
xor  ( new_n50136_, new_n49735_, new_n49734_ );
and  ( new_n50137_, new_n50136_, new_n50135_ );
nor  ( new_n50138_, new_n50137_, new_n50134_ );
nor  ( new_n50139_, new_n50138_, new_n50107_ );
nor  ( new_n50140_, new_n50139_, new_n50106_ );
or   ( new_n50141_, new_n50140_, new_n50102_ );
and  ( new_n50142_, new_n50141_, new_n50101_ );
or   ( new_n50143_, new_n50142_, new_n50066_ );
xor  ( new_n50144_, new_n50142_, new_n50066_ );
xor  ( new_n50145_, new_n49862_, new_n49860_ );
xor  ( new_n50146_, new_n50145_, new_n49865_ );
nand ( new_n50147_, new_n50146_, new_n50144_ );
and  ( new_n50148_, new_n50147_, new_n50143_ );
or   ( new_n50149_, new_n50148_, new_n49914_ );
and  ( new_n50150_, new_n50149_, new_n49913_ );
nor  ( new_n50151_, new_n50150_, new_n49893_ );
nor  ( new_n50152_, new_n50151_, new_n49891_ );
xor  ( new_n50153_, new_n49882_, new_n49880_ );
and  ( new_n50154_, new_n50153_, new_n50152_ );
nor  ( new_n50155_, new_n50153_, new_n50152_ );
xor  ( new_n50156_, new_n50150_, new_n49893_ );
not  ( new_n50157_, new_n50156_ );
xor  ( new_n50158_, new_n49912_, new_n49910_ );
xor  ( new_n50159_, new_n50158_, new_n50148_ );
xor  ( new_n50160_, new_n49869_, new_n49867_ );
xor  ( new_n50161_, new_n50160_, new_n49872_ );
or   ( new_n50162_, new_n50161_, new_n50159_ );
and  ( new_n50163_, new_n50161_, new_n50159_ );
xor  ( new_n50164_, new_n49848_, new_n49843_ );
xor  ( new_n50165_, new_n50164_, new_n49858_ );
xnor ( new_n50166_, new_n49897_, new_n49895_ );
xor  ( new_n50167_, new_n50166_, new_n49901_ );
nor  ( new_n50168_, new_n50167_, new_n50165_ );
xnor ( new_n50169_, new_n50051_, new_n50050_ );
nand ( new_n50170_, new_n49987_, new_n1739_ );
xor  ( new_n50171_, new_n45403_, new_n1583_ );
or   ( new_n50172_, new_n50171_, new_n1844_ );
and  ( new_n50173_, new_n50172_, new_n50170_ );
xor  ( new_n50174_, new_n43812_, new_n3892_ );
or   ( new_n50175_, new_n50174_, new_n4302_ );
or   ( new_n50176_, new_n49974_, new_n4304_ );
and  ( new_n50177_, new_n50176_, new_n50175_ );
nor  ( new_n50178_, new_n50177_, new_n50173_ );
xor  ( new_n50179_, new_n45738_, RIbb2ebc0_23 );
and  ( new_n50180_, new_n50179_, new_n1476_ );
and  ( new_n50181_, new_n50109_, new_n1474_ );
or   ( new_n50182_, new_n50181_, new_n50180_ );
xor  ( new_n50183_, new_n50177_, new_n50173_ );
and  ( new_n50184_, new_n50183_, new_n50182_ );
or   ( new_n50185_, new_n50184_, new_n50178_ );
xor  ( new_n50186_, new_n50031_, new_n50030_ );
nand ( new_n50187_, new_n50186_, new_n50185_ );
nor  ( new_n50188_, new_n50186_, new_n50185_ );
xor  ( new_n50189_, new_n43952_, new_n4292_ );
or   ( new_n50190_, new_n50189_, new_n4709_ );
or   ( new_n50191_, new_n49941_, new_n4711_ );
nand ( new_n50192_, new_n50191_, new_n50190_ );
and  ( new_n50193_, new_n50192_, new_n49984_ );
xor  ( new_n50194_, new_n45119_, new_n1840_ );
nor  ( new_n50195_, new_n50194_, new_n2122_ );
and  ( new_n50196_, new_n49931_, new_n2000_ );
or   ( new_n50197_, new_n50196_, new_n50195_ );
xor  ( new_n50198_, new_n50192_, new_n49984_ );
and  ( new_n50199_, new_n50198_, new_n50197_ );
nor  ( new_n50200_, new_n50199_, new_n50193_ );
or   ( new_n50201_, new_n50200_, new_n50188_ );
and  ( new_n50202_, new_n50201_, new_n50187_ );
nor  ( new_n50203_, new_n50202_, new_n50169_ );
xor  ( new_n50204_, new_n43898_, new_n6163_ );
or   ( new_n50205_, new_n50204_, new_n6645_ );
or   ( new_n50206_, new_n50035_, new_n6647_ );
and  ( new_n50207_, new_n50206_, new_n50205_ );
or   ( new_n50208_, new_n50040_, new_n1137_ );
xor  ( new_n50209_, new_n46137_, new_n893_ );
or   ( new_n50210_, new_n50209_, new_n1135_ );
and  ( new_n50211_, new_n50210_, new_n50208_ );
or   ( new_n50212_, new_n50211_, new_n50207_ );
xor  ( new_n50213_, new_n44319_, RIbb2e620_35 );
and  ( new_n50214_, new_n50213_, new_n3293_ );
and  ( new_n50215_, new_n49958_, new_n3291_ );
or   ( new_n50216_, new_n50215_, new_n50214_ );
xor  ( new_n50217_, new_n50211_, new_n50207_ );
nand ( new_n50218_, new_n50217_, new_n50216_ );
and  ( new_n50219_, new_n50218_, new_n50212_ );
xor  ( new_n50220_, new_n44681_, new_n2421_ );
or   ( new_n50221_, new_n50220_, new_n2807_ );
or   ( new_n50222_, new_n49919_, new_n2809_ );
and  ( new_n50223_, new_n50222_, new_n50221_ );
xor  ( new_n50224_, new_n43799_, new_n5594_ );
or   ( new_n50225_, new_n50224_, new_n6173_ );
nand ( new_n50226_, new_n49925_, new_n5915_ );
and  ( new_n50227_, new_n50226_, new_n50225_ );
or   ( new_n50228_, new_n50227_, new_n50223_ );
xor  ( new_n50229_, new_n44877_, RIbb2e8f0_29 );
and  ( new_n50230_, new_n50229_, new_n2244_ );
and  ( new_n50231_, new_n49935_, new_n2242_ );
or   ( new_n50232_, new_n50231_, new_n50230_ );
xor  ( new_n50233_, new_n50227_, new_n50223_ );
nand ( new_n50234_, new_n50233_, new_n50232_ );
and  ( new_n50235_, new_n50234_, new_n50228_ );
nor  ( new_n50236_, new_n50235_, new_n50219_ );
xor  ( new_n50237_, new_n43937_, RIbb2e260_43 );
nand ( new_n50238_, new_n50237_, new_n4960_ );
or   ( new_n50239_, new_n49915_, new_n5209_ );
and  ( new_n50240_, new_n50239_, new_n50238_ );
or   ( new_n50241_, new_n49948_, new_n5606_ );
xor  ( new_n50242_, new_n43884_, RIbb2e170_45 );
nand ( new_n50243_, new_n50242_, new_n5373_ );
and  ( new_n50244_, new_n50243_, new_n50241_ );
nor  ( new_n50245_, new_n50244_, new_n50240_ );
and  ( new_n50246_, new_n49952_, new_n2928_ );
xor  ( new_n50247_, new_n44506_, RIbb2e710_33 );
and  ( new_n50248_, new_n50247_, new_n2930_ );
or   ( new_n50249_, new_n50248_, new_n50246_ );
xor  ( new_n50250_, new_n50244_, new_n50240_ );
and  ( new_n50251_, new_n50250_, new_n50249_ );
or   ( new_n50252_, new_n50251_, new_n50245_ );
xor  ( new_n50253_, new_n50235_, new_n50219_ );
and  ( new_n50254_, new_n50253_, new_n50252_ );
or   ( new_n50255_, new_n50254_, new_n50236_ );
xor  ( new_n50256_, new_n50202_, new_n50169_ );
and  ( new_n50257_, new_n50256_, new_n50255_ );
or   ( new_n50258_, new_n50257_, new_n50203_ );
xor  ( new_n50259_, new_n49997_, new_n49996_ );
and  ( new_n50260_, new_n50259_, new_n50258_ );
xor  ( new_n50261_, new_n49946_, new_n49930_ );
xor  ( new_n50262_, new_n50261_, new_n49963_ );
xor  ( new_n50263_, new_n49961_, new_n49960_ );
xor  ( new_n50264_, new_n50048_, new_n50047_ );
nand ( new_n50265_, new_n50264_, new_n50263_ );
xor  ( new_n50266_, new_n50264_, new_n50263_ );
xnor ( new_n50267_, new_n49922_, new_n49918_ );
nand ( new_n50268_, new_n50267_, new_n49928_ );
not  ( new_n50269_, new_n49929_ );
or   ( new_n50270_, new_n50269_, new_n49923_ );
and  ( new_n50271_, new_n50270_, new_n50268_ );
nand ( new_n50272_, new_n50271_, new_n50266_ );
and  ( new_n50273_, new_n50272_, new_n50265_ );
nor  ( new_n50274_, new_n50273_, new_n50262_ );
xor  ( new_n50275_, new_n49994_, new_n49993_ );
xor  ( new_n50276_, new_n50273_, new_n50262_ );
and  ( new_n50277_, new_n50276_, new_n50275_ );
nor  ( new_n50278_, new_n50277_, new_n50274_ );
xnor ( new_n50279_, new_n50259_, new_n50258_ );
nor  ( new_n50280_, new_n50279_, new_n50278_ );
or   ( new_n50281_, new_n50280_, new_n50260_ );
xor  ( new_n50282_, new_n50167_, new_n50165_ );
and  ( new_n50283_, new_n50282_, new_n50281_ );
or   ( new_n50284_, new_n50283_, new_n50168_ );
xor  ( new_n50285_, new_n49908_, new_n49907_ );
and  ( new_n50286_, new_n50285_, new_n50284_ );
xor  ( new_n50287_, new_n50285_, new_n50284_ );
xor  ( new_n50288_, new_n50146_, new_n50144_ );
and  ( new_n50289_, new_n50288_, new_n50287_ );
nor  ( new_n50290_, new_n50289_, new_n50286_ );
or   ( new_n50291_, new_n50290_, new_n50163_ );
and  ( new_n50292_, new_n50291_, new_n50162_ );
and  ( new_n50293_, new_n50292_, new_n50157_ );
nor  ( new_n50294_, new_n50292_, new_n50157_ );
or   ( new_n50295_, new_n50002_, new_n320_ );
xor  ( new_n50296_, new_n48518_, new_n309_ );
or   ( new_n50297_, new_n50296_, new_n317_ );
and  ( new_n50298_, new_n50297_, new_n50295_ );
xor  ( new_n50299_, new_n48908_, new_n275_ );
or   ( new_n50300_, new_n50299_, new_n283_ );
or   ( new_n50301_, new_n50067_, new_n286_ );
and  ( new_n50302_, new_n50301_, new_n50300_ );
or   ( new_n50303_, new_n50302_, new_n50298_ );
and  ( new_n50304_, new_n50302_, new_n50298_ );
nor  ( new_n50305_, RIbb2ddb0_53, RIbb2de28_52 );
not  ( new_n50306_, new_n50305_ );
and  ( new_n50307_, new_n50306_, new_n6637_ );
xor  ( new_n50308_, new_n43793_, new_n6635_ );
and  ( new_n50309_, new_n50308_, new_n6910_ );
nor  ( new_n50310_, new_n50309_, new_n50307_ );
or   ( new_n50311_, new_n50310_, new_n50304_ );
and  ( new_n50312_, new_n50311_, new_n50303_ );
xor  ( new_n50313_, new_n47296_, new_n325_ );
or   ( new_n50314_, new_n50313_, new_n409_ );
or   ( new_n50315_, new_n50012_, new_n411_ );
and  ( new_n50316_, new_n50315_, new_n50314_ );
xor  ( new_n50317_, new_n47303_, new_n400_ );
or   ( new_n50318_, new_n50317_, new_n524_ );
or   ( new_n50319_, new_n50018_, new_n526_ );
and  ( new_n50320_, new_n50319_, new_n50318_ );
or   ( new_n50321_, new_n50320_, new_n50316_ );
nor  ( new_n50322_, new_n50006_, new_n340_ );
xor  ( new_n50323_, new_n48039_, RIbb2f250_9 );
and  ( new_n50324_, new_n50323_, new_n336_ );
nor  ( new_n50325_, new_n50324_, new_n50322_ );
and  ( new_n50326_, new_n50320_, new_n50316_ );
or   ( new_n50327_, new_n50326_, new_n50325_ );
and  ( new_n50328_, new_n50327_, new_n50321_ );
nor  ( new_n50329_, new_n50328_, new_n50312_ );
or   ( new_n50330_, new_n49534_, new_n302_ );
or   ( new_n50331_, new_n49675_, new_n44007_ );
and  ( new_n50332_, new_n50331_, new_n50330_ );
xor  ( new_n50333_, new_n44183_, RIbb2e530_37 );
nand ( new_n50334_, new_n50333_, new_n3733_ );
nand ( new_n50335_, new_n50076_, new_n3731_ );
and  ( new_n50336_, new_n50335_, new_n50334_ );
nor  ( new_n50337_, new_n50336_, new_n50332_ );
xor  ( new_n50338_, new_n45928_, new_n1126_ );
nor  ( new_n50339_, new_n50338_, new_n1364_ );
and  ( new_n50340_, new_n50045_, new_n1251_ );
or   ( new_n50341_, new_n50340_, new_n50339_ );
xor  ( new_n50342_, new_n50336_, new_n50332_ );
and  ( new_n50343_, new_n50342_, new_n50341_ );
or   ( new_n50344_, new_n50343_, new_n50337_ );
xor  ( new_n50345_, new_n50328_, new_n50312_ );
and  ( new_n50346_, new_n50345_, new_n50344_ );
or   ( new_n50347_, new_n50346_, new_n50329_ );
xor  ( new_n50348_, new_n50015_, new_n50014_ );
xor  ( new_n50349_, new_n50073_, new_n50070_ );
xor  ( new_n50350_, new_n50349_, new_n50079_ );
or   ( new_n50351_, new_n50350_, new_n50348_ );
and  ( new_n50352_, new_n50350_, new_n50348_ );
xnor ( new_n50353_, new_n49938_, new_n49934_ );
nand ( new_n50354_, new_n50353_, new_n49944_ );
not  ( new_n50355_, new_n49945_ );
or   ( new_n50356_, new_n50355_, new_n49939_ );
and  ( new_n50357_, new_n50356_, new_n50354_ );
or   ( new_n50358_, new_n50357_, new_n50352_ );
and  ( new_n50359_, new_n50358_, new_n50351_ );
and  ( new_n50360_, new_n50359_, new_n50347_ );
xor  ( new_n50361_, new_n50085_, new_n50084_ );
xor  ( new_n50362_, new_n50359_, new_n50347_ );
and  ( new_n50363_, new_n50362_, new_n50361_ );
or   ( new_n50364_, new_n50363_, new_n50360_ );
xor  ( new_n50365_, new_n50097_, new_n50096_ );
and  ( new_n50366_, new_n50365_, new_n50364_ );
xor  ( new_n50367_, new_n50061_, new_n50056_ );
xor  ( new_n50368_, new_n50365_, new_n50364_ );
and  ( new_n50369_, new_n50368_, new_n50367_ );
or   ( new_n50370_, new_n50369_, new_n50366_ );
xor  ( new_n50371_, new_n50064_, new_n50063_ );
and  ( new_n50372_, new_n50371_, new_n50370_ );
xor  ( new_n50373_, new_n50371_, new_n50370_ );
xnor ( new_n50374_, new_n50100_, new_n50099_ );
xor  ( new_n50375_, new_n50374_, new_n50140_ );
and  ( new_n50376_, new_n50375_, new_n50373_ );
or   ( new_n50377_, new_n50376_, new_n50372_ );
xor  ( new_n50378_, new_n50288_, new_n50287_ );
and  ( new_n50379_, new_n50378_, new_n50377_ );
xor  ( new_n50380_, new_n50105_, new_n50103_ );
xor  ( new_n50381_, new_n50380_, new_n50138_ );
xor  ( new_n50382_, new_n50092_, new_n50091_ );
xor  ( new_n50383_, new_n50136_, new_n50135_ );
nand ( new_n50384_, new_n50383_, new_n50382_ );
nor  ( new_n50385_, new_n50383_, new_n50382_ );
xor  ( new_n50386_, new_n50127_, new_n50126_ );
xnor ( new_n50387_, new_n50302_, new_n50298_ );
xor  ( new_n50388_, new_n50387_, new_n50310_ );
and  ( new_n50389_, new_n50388_, new_n50386_ );
xor  ( new_n50390_, new_n50388_, new_n50386_ );
xnor ( new_n50391_, new_n50320_, new_n50316_ );
xor  ( new_n50392_, new_n50391_, new_n50325_ );
and  ( new_n50393_, new_n50392_, new_n50390_ );
or   ( new_n50394_, new_n50393_, new_n50389_ );
xor  ( new_n50395_, new_n50130_, new_n50129_ );
and  ( new_n50396_, new_n50395_, new_n50394_ );
or   ( new_n50397_, new_n50220_, new_n2809_ );
xor  ( new_n50398_, new_n44785_, new_n2421_ );
or   ( new_n50399_, new_n50398_, new_n2807_ );
and  ( new_n50400_, new_n50399_, new_n50397_ );
xor  ( new_n50401_, new_n43894_, RIbb2df90_49 );
nand ( new_n50402_, new_n50401_, new_n6510_ );
or   ( new_n50403_, new_n50204_, new_n6647_ );
and  ( new_n50404_, new_n50403_, new_n50402_ );
or   ( new_n50405_, new_n50404_, new_n50400_ );
and  ( new_n50406_, new_n50237_, new_n4958_ );
xor  ( new_n50407_, new_n43956_, new_n4705_ );
nor  ( new_n50408_, new_n50407_, new_n5207_ );
or   ( new_n50409_, new_n50408_, new_n50406_ );
xor  ( new_n50410_, new_n50404_, new_n50400_ );
nand ( new_n50411_, new_n50410_, new_n50409_ );
and  ( new_n50412_, new_n50411_, new_n50405_ );
xor  ( new_n50413_, new_n44407_, new_n3113_ );
or   ( new_n50414_, new_n50413_, new_n3461_ );
nand ( new_n50415_, new_n50213_, new_n3291_ );
and  ( new_n50416_, new_n50415_, new_n50414_ );
xor  ( new_n50417_, new_n44600_, new_n2797_ );
or   ( new_n50418_, new_n50417_, new_n3117_ );
nand ( new_n50419_, new_n50247_, new_n2928_ );
and  ( new_n50420_, new_n50419_, new_n50418_ );
or   ( new_n50421_, new_n50420_, new_n50416_ );
xor  ( new_n50422_, new_n43888_, RIbb2e170_45 );
and  ( new_n50423_, new_n50422_, new_n5373_ );
and  ( new_n50424_, new_n50242_, new_n5371_ );
nor  ( new_n50425_, new_n50424_, new_n50423_ );
and  ( new_n50426_, new_n50420_, new_n50416_ );
or   ( new_n50427_, new_n50426_, new_n50425_ );
and  ( new_n50428_, new_n50427_, new_n50421_ );
nor  ( new_n50429_, new_n50428_, new_n50412_ );
or   ( new_n50430_, new_n50189_, new_n4711_ );
xor  ( new_n50431_, new_n43985_, new_n4292_ );
or   ( new_n50432_, new_n50431_, new_n4709_ );
and  ( new_n50433_, new_n50432_, new_n50430_ );
nand ( new_n50434_, new_n50229_, new_n2242_ );
xor  ( new_n50435_, new_n44974_, RIbb2e8f0_29 );
nand ( new_n50436_, new_n50435_, new_n2244_ );
and  ( new_n50437_, new_n50436_, new_n50434_ );
nor  ( new_n50438_, new_n50437_, new_n50433_ );
nor  ( new_n50439_, new_n50194_, new_n2124_ );
xor  ( new_n50440_, new_n45204_, RIbb2e9e0_27 );
and  ( new_n50441_, new_n50440_, new_n2002_ );
or   ( new_n50442_, new_n50441_, new_n50439_ );
xor  ( new_n50443_, new_n50437_, new_n50433_ );
and  ( new_n50444_, new_n50443_, new_n50442_ );
or   ( new_n50445_, new_n50444_, new_n50438_ );
xor  ( new_n50446_, new_n50428_, new_n50412_ );
and  ( new_n50447_, new_n50446_, new_n50445_ );
or   ( new_n50448_, new_n50447_, new_n50429_ );
xor  ( new_n50449_, new_n50395_, new_n50394_ );
and  ( new_n50450_, new_n50449_, new_n50448_ );
nor  ( new_n50451_, new_n50450_, new_n50396_ );
or   ( new_n50452_, new_n50451_, new_n50385_ );
and  ( new_n50453_, new_n50452_, new_n50384_ );
nor  ( new_n50454_, new_n50453_, new_n50381_ );
xor  ( new_n50455_, new_n50115_, new_n43945_ );
not  ( new_n50456_, new_n50455_ );
or   ( new_n50457_, new_n50456_, new_n43983_ );
nor  ( new_n50458_, new_n49758_, new_n43880_ );
or   ( new_n50459_, new_n49759_, new_n43977_ );
or   ( new_n50460_, new_n50459_, new_n50458_ );
and  ( new_n50461_, new_n50460_, new_n50457_ );
or   ( new_n50462_, new_n50461_, new_n7176_ );
and  ( new_n50463_, new_n49676_, new_n295_ );
and  ( new_n50464_, new_n49763_, new_n43949_ );
or   ( new_n50465_, new_n50464_, new_n50463_ );
xor  ( new_n50466_, new_n50461_, new_n7176_ );
nand ( new_n50467_, new_n50466_, new_n50465_ );
and  ( new_n50468_, new_n50467_, new_n50462_ );
or   ( new_n50469_, new_n50299_, new_n286_ );
xor  ( new_n50470_, new_n49265_, new_n275_ );
or   ( new_n50471_, new_n50470_, new_n283_ );
and  ( new_n50472_, new_n50471_, new_n50469_ );
nand ( new_n50473_, new_n50323_, new_n334_ );
xor  ( new_n50474_, new_n48291_, new_n329_ );
or   ( new_n50475_, new_n50474_, new_n337_ );
and  ( new_n50476_, new_n50475_, new_n50473_ );
or   ( new_n50477_, new_n50476_, new_n50472_ );
or   ( new_n50478_, new_n50296_, new_n320_ );
xor  ( new_n50479_, new_n48756_, new_n309_ );
or   ( new_n50480_, new_n50479_, new_n317_ );
and  ( new_n50481_, new_n50480_, new_n50478_ );
and  ( new_n50482_, new_n50476_, new_n50472_ );
or   ( new_n50483_, new_n50482_, new_n50481_ );
and  ( new_n50484_, new_n50483_, new_n50477_ );
nor  ( new_n50485_, new_n50484_, new_n50468_ );
xor  ( new_n50486_, RIbb32dd8_180, RIbb2c028_116 );
xor  ( new_n50487_, new_n50486_, new_n49479_ );
and  ( new_n50488_, new_n50487_, new_n43880_ );
not  ( new_n50489_, new_n50488_ );
or   ( new_n50490_, new_n50209_, new_n1137_ );
xor  ( new_n50491_, new_n46427_, RIbb2eda0_19 );
nand ( new_n50492_, new_n50491_, new_n1042_ );
and  ( new_n50493_, new_n50492_, new_n50490_ );
nor  ( new_n50494_, new_n50493_, new_n50489_ );
xor  ( new_n50495_, new_n46789_, new_n745_ );
nor  ( new_n50496_, new_n50495_, new_n897_ );
nor  ( new_n50497_, new_n50119_, new_n899_ );
or   ( new_n50498_, new_n50497_, new_n50496_ );
xor  ( new_n50499_, new_n50493_, new_n50489_ );
and  ( new_n50500_, new_n50499_, new_n50498_ );
or   ( new_n50501_, new_n50500_, new_n50494_ );
xor  ( new_n50502_, new_n50484_, new_n50468_ );
and  ( new_n50503_, new_n50502_, new_n50501_ );
nor  ( new_n50504_, new_n50503_, new_n50485_ );
not  ( new_n50505_, new_n50504_ );
xor  ( new_n50506_, new_n49990_, new_n49989_ );
and  ( new_n50507_, new_n50506_, new_n50505_ );
xor  ( new_n50508_, new_n50506_, new_n50505_ );
xor  ( new_n50509_, new_n50345_, new_n50344_ );
and  ( new_n50510_, new_n50509_, new_n50508_ );
or   ( new_n50511_, new_n50510_, new_n50507_ );
xor  ( new_n50512_, new_n50253_, new_n50252_ );
xor  ( new_n50513_, new_n50350_, new_n50348_ );
xor  ( new_n50514_, new_n50513_, new_n50357_ );
or   ( new_n50515_, new_n50514_, new_n50512_ );
and  ( new_n50516_, new_n50514_, new_n50512_ );
xor  ( new_n50517_, new_n50186_, new_n50185_ );
xnor ( new_n50518_, new_n50517_, new_n50200_ );
or   ( new_n50519_, new_n50518_, new_n50516_ );
and  ( new_n50520_, new_n50519_, new_n50515_ );
and  ( new_n50521_, new_n50520_, new_n50511_ );
or   ( new_n50522_, new_n50317_, new_n526_ );
xor  ( new_n50523_, new_n47046_, new_n400_ );
or   ( new_n50524_, new_n50523_, new_n524_ );
and  ( new_n50525_, new_n50524_, new_n50522_ );
or   ( new_n50526_, new_n50313_, new_n411_ );
xor  ( new_n50527_, new_n47640_, new_n325_ );
or   ( new_n50528_, new_n50527_, new_n409_ );
and  ( new_n50529_, new_n50528_, new_n50526_ );
or   ( new_n50530_, new_n50529_, new_n50525_ );
nor  ( new_n50531_, new_n50124_, new_n757_ );
xor  ( new_n50532_, new_n46958_, RIbb2ef80_15 );
and  ( new_n50533_, new_n50532_, new_n662_ );
or   ( new_n50534_, new_n50533_, new_n50531_ );
xor  ( new_n50535_, new_n50529_, new_n50525_ );
nand ( new_n50536_, new_n50535_, new_n50534_ );
and  ( new_n50537_, new_n50536_, new_n50530_ );
xor  ( new_n50538_, new_n43787_, new_n6635_ );
or   ( new_n50539_, new_n50538_, new_n7184_ );
nand ( new_n50540_, new_n50308_, new_n6908_ );
and  ( new_n50541_, new_n50540_, new_n50539_ );
or   ( new_n50542_, new_n50224_, new_n6175_ );
xor  ( new_n50543_, new_n43803_, RIbb2e080_47 );
nand ( new_n50544_, new_n50543_, new_n5917_ );
and  ( new_n50545_, new_n50544_, new_n50542_ );
or   ( new_n50546_, new_n50545_, new_n50541_ );
and  ( new_n50547_, new_n50333_, new_n3731_ );
xor  ( new_n50548_, new_n44218_, RIbb2e530_37 );
and  ( new_n50549_, new_n50548_, new_n3733_ );
or   ( new_n50550_, new_n50549_, new_n50547_ );
xor  ( new_n50551_, new_n50545_, new_n50541_ );
nand ( new_n50552_, new_n50551_, new_n50550_ );
and  ( new_n50553_, new_n50552_, new_n50546_ );
or   ( new_n50554_, new_n50553_, new_n50537_ );
or   ( new_n50555_, new_n50174_, new_n4304_ );
xor  ( new_n50556_, new_n43914_, RIbb2e440_39 );
nand ( new_n50557_, new_n50556_, new_n4034_ );
and  ( new_n50558_, new_n50557_, new_n50555_ );
nand ( new_n50559_, new_n50179_, new_n1474_ );
xor  ( new_n50560_, new_n45597_, new_n1355_ );
or   ( new_n50561_, new_n50560_, new_n1593_ );
and  ( new_n50562_, new_n50561_, new_n50559_ );
nor  ( new_n50563_, new_n50562_, new_n50558_ );
nor  ( new_n50564_, new_n50338_, new_n1366_ );
xor  ( new_n50565_, new_n46037_, new_n1126_ );
nor  ( new_n50566_, new_n50565_, new_n1364_ );
or   ( new_n50567_, new_n50566_, new_n50564_ );
xor  ( new_n50568_, new_n50562_, new_n50558_ );
and  ( new_n50569_, new_n50568_, new_n50567_ );
or   ( new_n50570_, new_n50569_, new_n50563_ );
xor  ( new_n50571_, new_n50553_, new_n50537_ );
nand ( new_n50572_, new_n50571_, new_n50570_ );
and  ( new_n50573_, new_n50572_, new_n50554_ );
xor  ( new_n50574_, new_n50250_, new_n50249_ );
xor  ( new_n50575_, new_n50198_, new_n50197_ );
nand ( new_n50576_, new_n50575_, new_n50574_ );
xor  ( new_n50577_, new_n50183_, new_n50182_ );
xor  ( new_n50578_, new_n50575_, new_n50574_ );
nand ( new_n50579_, new_n50578_, new_n50577_ );
and  ( new_n50580_, new_n50579_, new_n50576_ );
nor  ( new_n50581_, new_n50580_, new_n50573_ );
xor  ( new_n50582_, new_n50217_, new_n50216_ );
xor  ( new_n50583_, new_n50233_, new_n50232_ );
and  ( new_n50584_, new_n50583_, new_n50582_ );
xor  ( new_n50585_, new_n50583_, new_n50582_ );
xor  ( new_n50586_, new_n50342_, new_n50341_ );
and  ( new_n50587_, new_n50586_, new_n50585_ );
or   ( new_n50588_, new_n50587_, new_n50584_ );
xor  ( new_n50589_, new_n50580_, new_n50573_ );
and  ( new_n50590_, new_n50589_, new_n50588_ );
or   ( new_n50591_, new_n50590_, new_n50581_ );
xor  ( new_n50592_, new_n50520_, new_n50511_ );
and  ( new_n50593_, new_n50592_, new_n50591_ );
nor  ( new_n50594_, new_n50593_, new_n50521_ );
xnor ( new_n50595_, new_n50453_, new_n50381_ );
nor  ( new_n50596_, new_n50595_, new_n50594_ );
or   ( new_n50597_, new_n50596_, new_n50454_ );
xor  ( new_n50598_, new_n50282_, new_n50281_ );
and  ( new_n50599_, new_n50598_, new_n50597_ );
xnor ( new_n50600_, new_n50279_, new_n50278_ );
xor  ( new_n50601_, new_n50256_, new_n50255_ );
xor  ( new_n50602_, new_n50362_, new_n50361_ );
nand ( new_n50603_, new_n50602_, new_n50601_ );
or   ( new_n50604_, new_n50602_, new_n50601_ );
xor  ( new_n50605_, new_n50276_, new_n50275_ );
nand ( new_n50606_, new_n50605_, new_n50604_ );
and  ( new_n50607_, new_n50606_, new_n50603_ );
nor  ( new_n50608_, new_n50607_, new_n50600_ );
xor  ( new_n50609_, new_n50607_, new_n50600_ );
xor  ( new_n50610_, new_n50368_, new_n50367_ );
and  ( new_n50611_, new_n50610_, new_n50609_ );
or   ( new_n50612_, new_n50611_, new_n50608_ );
xor  ( new_n50613_, new_n50598_, new_n50597_ );
and  ( new_n50614_, new_n50613_, new_n50612_ );
or   ( new_n50615_, new_n50614_, new_n50599_ );
xor  ( new_n50616_, new_n50378_, new_n50377_ );
and  ( new_n50617_, new_n50616_, new_n50615_ );
nor  ( new_n50618_, new_n50617_, new_n50379_ );
xor  ( new_n50619_, new_n50161_, new_n50159_ );
xnor ( new_n50620_, new_n50619_, new_n50290_ );
not  ( new_n50621_, new_n50620_ );
and  ( new_n50622_, new_n50621_, new_n50618_ );
nor  ( new_n50623_, new_n50621_, new_n50618_ );
xnor ( new_n50624_, new_n50595_, new_n50594_ );
xor  ( new_n50625_, new_n50509_, new_n50508_ );
xor  ( new_n50626_, new_n50271_, new_n50266_ );
and  ( new_n50627_, new_n50626_, new_n50625_ );
xnor ( new_n50628_, new_n50626_, new_n50625_ );
nor  ( new_n50629_, new_n49977_, new_n44007_ );
and  ( new_n50630_, new_n49763_, new_n295_ );
nor  ( new_n50631_, new_n50630_, new_n50629_ );
not  ( new_n50632_, new_n50631_ );
or   ( new_n50633_, new_n50431_, new_n4711_ );
xor  ( new_n50634_, new_n43812_, new_n4292_ );
or   ( new_n50635_, new_n50634_, new_n4709_ );
and  ( new_n50636_, new_n50635_, new_n50633_ );
nor  ( new_n50637_, new_n50636_, new_n50632_ );
and  ( new_n50638_, new_n50440_, new_n2000_ );
xor  ( new_n50639_, new_n45403_, new_n1840_ );
nor  ( new_n50640_, new_n50639_, new_n2122_ );
or   ( new_n50641_, new_n50640_, new_n50638_ );
xor  ( new_n50642_, new_n50636_, new_n50632_ );
and  ( new_n50643_, new_n50642_, new_n50641_ );
or   ( new_n50644_, new_n50643_, new_n50637_ );
xor  ( new_n50645_, new_n50499_, new_n50498_ );
and  ( new_n50646_, new_n50645_, new_n50644_ );
xor  ( new_n50647_, new_n50645_, new_n50644_ );
xor  ( new_n50648_, new_n50535_, new_n50534_ );
and  ( new_n50649_, new_n50648_, new_n50647_ );
nor  ( new_n50650_, new_n50649_, new_n50646_ );
not  ( new_n50651_, new_n50650_ );
xor  ( new_n50652_, new_n50476_, new_n50472_ );
xor  ( new_n50653_, new_n50652_, new_n50481_ );
xor  ( new_n50654_, new_n44319_, RIbb2e530_37 );
nand ( new_n50655_, new_n50654_, new_n3733_ );
nand ( new_n50656_, new_n50548_, new_n3731_ );
and  ( new_n50657_, new_n50656_, new_n50655_ );
or   ( new_n50658_, new_n50413_, new_n3463_ );
xor  ( new_n50659_, new_n44506_, new_n3113_ );
or   ( new_n50660_, new_n50659_, new_n3461_ );
and  ( new_n50661_, new_n50660_, new_n50658_ );
nor  ( new_n50662_, new_n50661_, new_n50657_ );
and  ( new_n50663_, new_n50661_, new_n50657_ );
and  ( new_n50664_, new_n50543_, new_n5915_ );
xor  ( new_n50665_, new_n43884_, RIbb2e080_47 );
and  ( new_n50666_, new_n50665_, new_n5917_ );
nor  ( new_n50667_, new_n50666_, new_n50664_ );
nor  ( new_n50668_, new_n50667_, new_n50663_ );
nor  ( new_n50669_, new_n50668_, new_n50662_ );
nor  ( new_n50670_, new_n50669_, new_n50653_ );
or   ( new_n50671_, new_n50417_, new_n3119_ );
xor  ( new_n50672_, new_n44681_, new_n2797_ );
or   ( new_n50673_, new_n50672_, new_n3117_ );
and  ( new_n50674_, new_n50673_, new_n50671_ );
nand ( new_n50675_, new_n50422_, new_n5371_ );
xor  ( new_n50676_, new_n43937_, RIbb2e170_45 );
nand ( new_n50677_, new_n50676_, new_n5373_ );
and  ( new_n50678_, new_n50677_, new_n50675_ );
nor  ( new_n50679_, new_n50678_, new_n50674_ );
and  ( new_n50680_, new_n50401_, new_n6508_ );
xor  ( new_n50681_, new_n43799_, new_n6163_ );
nor  ( new_n50682_, new_n50681_, new_n6645_ );
or   ( new_n50683_, new_n50682_, new_n50680_ );
xor  ( new_n50684_, new_n50678_, new_n50674_ );
and  ( new_n50685_, new_n50684_, new_n50683_ );
or   ( new_n50686_, new_n50685_, new_n50679_ );
xor  ( new_n50687_, new_n50669_, new_n50653_ );
and  ( new_n50688_, new_n50687_, new_n50686_ );
nor  ( new_n50689_, new_n50688_, new_n50670_ );
not  ( new_n50690_, new_n50689_ );
and  ( new_n50691_, new_n50690_, new_n50651_ );
and  ( new_n50692_, new_n50689_, new_n50650_ );
or   ( new_n50693_, new_n50470_, new_n286_ );
xor  ( new_n50694_, new_n49427_, RIbb2f430_5 );
nand ( new_n50695_, new_n50694_, new_n282_ );
and  ( new_n50696_, new_n50695_, new_n50693_ );
or   ( new_n50697_, new_n50479_, new_n320_ );
xor  ( new_n50698_, new_n48908_, new_n309_ );
or   ( new_n50699_, new_n50698_, new_n317_ );
and  ( new_n50700_, new_n50699_, new_n50697_ );
or   ( new_n50701_, new_n50700_, new_n50696_ );
xor  ( new_n50702_, new_n44183_, RIbb2e440_39 );
and  ( new_n50703_, new_n50702_, new_n4034_ );
and  ( new_n50704_, new_n50556_, new_n4032_ );
nor  ( new_n50705_, new_n50704_, new_n50703_ );
not  ( new_n50706_, new_n50705_ );
xor  ( new_n50707_, new_n50700_, new_n50696_ );
nand ( new_n50708_, new_n50707_, new_n50706_ );
and  ( new_n50709_, new_n50708_, new_n50701_ );
or   ( new_n50710_, new_n50538_, new_n7186_ );
xor  ( new_n50711_, new_n43898_, new_n6635_ );
or   ( new_n50712_, new_n50711_, new_n7184_ );
and  ( new_n50713_, new_n50712_, new_n50710_ );
xor  ( new_n50714_, new_n45928_, new_n1355_ );
or   ( new_n50715_, new_n50714_, new_n1593_ );
or   ( new_n50716_, new_n50560_, new_n1595_ );
and  ( new_n50717_, new_n50716_, new_n50715_ );
or   ( new_n50718_, new_n50717_, new_n50713_ );
nor  ( new_n50719_, new_n50565_, new_n1366_ );
xor  ( new_n50720_, new_n46137_, RIbb2ecb0_21 );
and  ( new_n50721_, new_n50720_, new_n1253_ );
or   ( new_n50722_, new_n50721_, new_n50719_ );
xor  ( new_n50723_, new_n50717_, new_n50713_ );
nand ( new_n50724_, new_n50723_, new_n50722_ );
and  ( new_n50725_, new_n50724_, new_n50718_ );
nor  ( new_n50726_, new_n50725_, new_n50709_ );
or   ( new_n50727_, new_n50407_, new_n5209_ );
xor  ( new_n50728_, new_n43952_, new_n4705_ );
or   ( new_n50729_, new_n50728_, new_n5207_ );
and  ( new_n50730_, new_n50729_, new_n50727_ );
or   ( new_n50731_, new_n50398_, new_n2809_ );
xor  ( new_n50732_, new_n44877_, new_n2421_ );
or   ( new_n50733_, new_n50732_, new_n2807_ );
and  ( new_n50734_, new_n50733_, new_n50731_ );
nor  ( new_n50735_, new_n50734_, new_n50730_ );
and  ( new_n50736_, new_n50435_, new_n2242_ );
xor  ( new_n50737_, new_n45119_, new_n2118_ );
nor  ( new_n50738_, new_n50737_, new_n2425_ );
nor  ( new_n50739_, new_n50738_, new_n50736_ );
not  ( new_n50740_, new_n50739_ );
xor  ( new_n50741_, new_n50734_, new_n50730_ );
and  ( new_n50742_, new_n50741_, new_n50740_ );
nor  ( new_n50743_, new_n50742_, new_n50735_ );
not  ( new_n50744_, new_n50743_ );
xor  ( new_n50745_, new_n50725_, new_n50709_ );
and  ( new_n50746_, new_n50745_, new_n50744_ );
nor  ( new_n50747_, new_n50746_, new_n50726_ );
nor  ( new_n50748_, new_n50747_, new_n50692_ );
nor  ( new_n50749_, new_n50748_, new_n50691_ );
nor  ( new_n50750_, new_n50749_, new_n50628_ );
or   ( new_n50751_, new_n50750_, new_n50627_ );
xnor ( new_n50752_, new_n50383_, new_n50382_ );
xor  ( new_n50753_, new_n50752_, new_n50451_ );
nand ( new_n50754_, new_n50753_, new_n50751_ );
xor  ( new_n50755_, new_n45584_, new_n1583_ );
or   ( new_n50756_, new_n50755_, new_n1844_ );
or   ( new_n50757_, new_n50171_, new_n1846_ );
and  ( new_n50758_, new_n50757_, new_n50756_ );
or   ( new_n50759_, new_n50758_, new_n50631_ );
or   ( new_n50760_, new_n50474_, new_n340_ );
xor  ( new_n50761_, new_n48518_, new_n329_ );
or   ( new_n50762_, new_n50761_, new_n337_ );
and  ( new_n50763_, new_n50762_, new_n50760_ );
not  ( new_n50764_, RIbb2dd38_54 );
and  ( new_n50765_, new_n7722_, new_n50764_ );
or   ( new_n50766_, new_n50765_, new_n7177_ );
xor  ( new_n50767_, new_n43793_, RIbb2ddb0_53 );
or   ( new_n50768_, new_n50767_, new_n7732_ );
and  ( new_n50769_, new_n50768_, new_n50766_ );
nor  ( new_n50770_, new_n50769_, new_n50763_ );
nor  ( new_n50771_, new_n50527_, new_n411_ );
xor  ( new_n50772_, new_n48039_, RIbb2f160_11 );
and  ( new_n50773_, new_n50772_, new_n373_ );
or   ( new_n50774_, new_n50773_, new_n50771_ );
nand ( new_n50775_, new_n50769_, new_n50763_ );
and  ( new_n50776_, new_n50775_, new_n50774_ );
or   ( new_n50777_, new_n50776_, new_n50770_ );
xor  ( new_n50778_, new_n50758_, new_n50631_ );
nand ( new_n50779_, new_n50778_, new_n50777_ );
and  ( new_n50780_, new_n50779_, new_n50759_ );
xor  ( new_n50781_, RIbb32e50_181, RIbb2bfb0_117 );
nor  ( new_n50782_, new_n49475_, new_n43510_ );
nor  ( new_n50783_, new_n50782_, new_n43537_ );
nor  ( new_n50784_, new_n50783_, new_n43507_ );
nor  ( new_n50785_, new_n50784_, new_n43536_ );
nor  ( new_n50786_, new_n50785_, new_n43506_ );
nor  ( new_n50787_, new_n50786_, new_n43542_ );
xnor ( new_n50788_, new_n50787_, new_n50781_ );
and  ( new_n50789_, new_n50788_, new_n43880_ );
not  ( new_n50790_, new_n50789_ );
xor  ( new_n50791_, new_n50487_, new_n43945_ );
not  ( new_n50792_, new_n50791_ );
or   ( new_n50793_, new_n50792_, new_n43983_ );
nor  ( new_n50794_, new_n50115_, new_n43880_ );
or   ( new_n50795_, new_n50116_, new_n43977_ );
or   ( new_n50796_, new_n50795_, new_n50794_ );
and  ( new_n50797_, new_n50796_, new_n50793_ );
nor  ( new_n50798_, new_n50797_, new_n50790_ );
and  ( new_n50799_, new_n50491_, new_n1040_ );
xor  ( new_n50800_, new_n46619_, new_n893_ );
nor  ( new_n50801_, new_n50800_, new_n1135_ );
or   ( new_n50802_, new_n50801_, new_n50799_ );
xor  ( new_n50803_, new_n50797_, new_n50790_ );
and  ( new_n50804_, new_n50803_, new_n50802_ );
or   ( new_n50805_, new_n50804_, new_n50798_ );
xor  ( new_n50806_, new_n50466_, new_n50465_ );
nand ( new_n50807_, new_n50806_, new_n50805_ );
xor  ( new_n50808_, new_n47303_, new_n520_ );
or   ( new_n50809_, new_n50808_, new_n755_ );
nand ( new_n50810_, new_n50532_, new_n660_ );
and  ( new_n50811_, new_n50810_, new_n50809_ );
xor  ( new_n50812_, new_n47296_, RIbb2f070_13 );
nand ( new_n50813_, new_n50812_, new_n456_ );
or   ( new_n50814_, new_n50523_, new_n526_ );
and  ( new_n50815_, new_n50814_, new_n50813_ );
nor  ( new_n50816_, new_n50815_, new_n50811_ );
nor  ( new_n50817_, new_n50495_, new_n899_ );
xor  ( new_n50818_, new_n46962_, new_n745_ );
nor  ( new_n50819_, new_n50818_, new_n897_ );
nor  ( new_n50820_, new_n50819_, new_n50817_ );
and  ( new_n50821_, new_n50815_, new_n50811_ );
nor  ( new_n50822_, new_n50821_, new_n50820_ );
or   ( new_n50823_, new_n50822_, new_n50816_ );
xor  ( new_n50824_, new_n50806_, new_n50805_ );
nand ( new_n50825_, new_n50824_, new_n50823_ );
and  ( new_n50826_, new_n50825_, new_n50807_ );
nor  ( new_n50827_, new_n50826_, new_n50780_ );
xor  ( new_n50828_, new_n50502_, new_n50501_ );
xor  ( new_n50829_, new_n50826_, new_n50780_ );
and  ( new_n50830_, new_n50829_, new_n50828_ );
or   ( new_n50831_, new_n50830_, new_n50827_ );
xor  ( new_n50832_, new_n50449_, new_n50448_ );
nand ( new_n50833_, new_n50832_, new_n50831_ );
xor  ( new_n50834_, new_n50571_, new_n50570_ );
xor  ( new_n50835_, new_n50392_, new_n50390_ );
and  ( new_n50836_, new_n50835_, new_n50834_ );
xor  ( new_n50837_, new_n50410_, new_n50409_ );
xor  ( new_n50838_, new_n50568_, new_n50567_ );
and  ( new_n50839_, new_n50838_, new_n50837_ );
xor  ( new_n50840_, new_n50838_, new_n50837_ );
xnor ( new_n50841_, new_n50420_, new_n50416_ );
xor  ( new_n50842_, new_n50841_, new_n50425_ );
and  ( new_n50843_, new_n50842_, new_n50840_ );
or   ( new_n50844_, new_n50843_, new_n50839_ );
xor  ( new_n50845_, new_n50835_, new_n50834_ );
and  ( new_n50846_, new_n50845_, new_n50844_ );
nor  ( new_n50847_, new_n50846_, new_n50836_ );
not  ( new_n50848_, new_n50847_ );
xor  ( new_n50849_, new_n50832_, new_n50831_ );
nand ( new_n50850_, new_n50849_, new_n50848_ );
and  ( new_n50851_, new_n50850_, new_n50833_ );
nor  ( new_n50852_, new_n50753_, new_n50751_ );
or   ( new_n50853_, new_n50852_, new_n50851_ );
and  ( new_n50854_, new_n50853_, new_n50754_ );
nor  ( new_n50855_, new_n50854_, new_n50624_ );
xor  ( new_n50856_, new_n50854_, new_n50624_ );
xor  ( new_n50857_, new_n50610_, new_n50609_ );
and  ( new_n50858_, new_n50857_, new_n50856_ );
or   ( new_n50859_, new_n50858_, new_n50855_ );
xor  ( new_n50860_, new_n50375_, new_n50373_ );
and  ( new_n50861_, new_n50860_, new_n50859_ );
xor  ( new_n50862_, new_n50613_, new_n50612_ );
xor  ( new_n50863_, new_n50860_, new_n50859_ );
and  ( new_n50864_, new_n50863_, new_n50862_ );
or   ( new_n50865_, new_n50864_, new_n50861_ );
xor  ( new_n50866_, new_n50616_, new_n50615_ );
nor  ( new_n50867_, new_n50866_, new_n50865_ );
and  ( new_n50868_, new_n50866_, new_n50865_ );
xor  ( new_n50869_, new_n50592_, new_n50591_ );
xor  ( new_n50870_, new_n50602_, new_n50601_ );
xor  ( new_n50871_, new_n50870_, new_n50605_ );
and  ( new_n50872_, new_n50871_, new_n50869_ );
xor  ( new_n50873_, new_n50446_, new_n50445_ );
xor  ( new_n50874_, new_n50586_, new_n50585_ );
and  ( new_n50875_, new_n50874_, new_n50873_ );
xor  ( new_n50876_, new_n50874_, new_n50873_ );
xor  ( new_n50877_, new_n50578_, new_n50577_ );
and  ( new_n50878_, new_n50877_, new_n50876_ );
nor  ( new_n50879_, new_n50878_, new_n50875_ );
xnor ( new_n50880_, new_n50589_, new_n50588_ );
nor  ( new_n50881_, new_n50880_, new_n50879_ );
xnor ( new_n50882_, new_n50880_, new_n50879_ );
xnor ( new_n50883_, new_n50514_, new_n50512_ );
xor  ( new_n50884_, new_n50883_, new_n50518_ );
nor  ( new_n50885_, new_n50884_, new_n50882_ );
nor  ( new_n50886_, new_n50885_, new_n50881_ );
xnor ( new_n50887_, new_n50871_, new_n50869_ );
nor  ( new_n50888_, new_n50887_, new_n50886_ );
nor  ( new_n50889_, new_n50888_, new_n50872_ );
xor  ( new_n50890_, new_n50551_, new_n50550_ );
xor  ( new_n50891_, new_n50443_, new_n50442_ );
and  ( new_n50892_, new_n50891_, new_n50890_ );
xor  ( new_n50893_, RIbb32ec8_182, RIbb2bf38_118 );
xnor ( new_n50894_, new_n50893_, new_n50785_ );
not  ( new_n50895_, new_n50894_ );
or   ( new_n50896_, new_n50895_, new_n43879_ );
nor  ( new_n50897_, new_n50487_, new_n43880_ );
or   ( new_n50898_, new_n50488_, new_n43977_ );
or   ( new_n50899_, new_n50898_, new_n50897_ );
xor  ( new_n50900_, new_n50788_, new_n43945_ );
nand ( new_n50901_, new_n50900_, new_n43982_ );
and  ( new_n50902_, new_n50901_, new_n50899_ );
or   ( new_n50903_, new_n50902_, new_n50896_ );
and  ( new_n50904_, new_n50902_, new_n50896_ );
and  ( new_n50905_, new_n50720_, new_n1251_ );
xor  ( new_n50906_, new_n46427_, RIbb2ecb0_21 );
and  ( new_n50907_, new_n50906_, new_n1253_ );
nor  ( new_n50908_, new_n50907_, new_n50905_ );
or   ( new_n50909_, new_n50908_, new_n50904_ );
and  ( new_n50910_, new_n50909_, new_n50903_ );
xor  ( new_n50911_, new_n48756_, RIbb2f250_9 );
nand ( new_n50912_, new_n50911_, new_n336_ );
or   ( new_n50913_, new_n50761_, new_n340_ );
and  ( new_n50914_, new_n50913_, new_n50912_ );
xor  ( new_n50915_, new_n48291_, new_n325_ );
or   ( new_n50916_, new_n50915_, new_n409_ );
nand ( new_n50917_, new_n50772_, new_n371_ );
and  ( new_n50918_, new_n50917_, new_n50916_ );
or   ( new_n50919_, new_n50918_, new_n50914_ );
and  ( new_n50920_, new_n50812_, new_n454_ );
xor  ( new_n50921_, new_n47640_, new_n400_ );
nor  ( new_n50922_, new_n50921_, new_n524_ );
nor  ( new_n50923_, new_n50922_, new_n50920_ );
and  ( new_n50924_, new_n50918_, new_n50914_ );
or   ( new_n50925_, new_n50924_, new_n50923_ );
and  ( new_n50926_, new_n50925_, new_n50919_ );
nor  ( new_n50927_, new_n50926_, new_n50910_ );
xor  ( new_n50928_, new_n50926_, new_n50910_ );
xor  ( new_n50929_, new_n50803_, new_n50802_ );
and  ( new_n50930_, new_n50929_, new_n50928_ );
or   ( new_n50931_, new_n50930_, new_n50927_ );
xor  ( new_n50932_, new_n50891_, new_n50890_ );
and  ( new_n50933_, new_n50932_, new_n50931_ );
nor  ( new_n50934_, new_n50933_, new_n50892_ );
or   ( new_n50935_, new_n49977_, new_n302_ );
or   ( new_n50936_, new_n50455_, new_n44007_ );
and  ( new_n50937_, new_n50936_, new_n50935_ );
nor  ( new_n50938_, new_n50937_, new_n7724_ );
and  ( new_n50939_, new_n50694_, new_n280_ );
xor  ( new_n50940_, new_n49488_, RIbb2f430_5 );
and  ( new_n50941_, new_n50940_, new_n282_ );
or   ( new_n50942_, new_n50941_, new_n50939_ );
xor  ( new_n50943_, new_n50937_, new_n7724_ );
and  ( new_n50944_, new_n50943_, new_n50942_ );
nor  ( new_n50945_, new_n50944_, new_n50938_ );
or   ( new_n50946_, new_n50755_, new_n1846_ );
xor  ( new_n50947_, new_n45738_, RIbb2ead0_25 );
nand ( new_n50948_, new_n50947_, new_n1741_ );
and  ( new_n50949_, new_n50948_, new_n50946_ );
nor  ( new_n50950_, new_n50949_, new_n50945_ );
xnor ( new_n50951_, new_n50949_, new_n50945_ );
xor  ( new_n50952_, new_n46958_, new_n745_ );
or   ( new_n50953_, new_n50952_, new_n897_ );
or   ( new_n50954_, new_n50818_, new_n899_ );
and  ( new_n50955_, new_n50954_, new_n50953_ );
or   ( new_n50956_, new_n50800_, new_n1137_ );
xor  ( new_n50957_, new_n46789_, new_n893_ );
or   ( new_n50958_, new_n50957_, new_n1135_ );
and  ( new_n50959_, new_n50958_, new_n50956_ );
nor  ( new_n50960_, new_n50959_, new_n50955_ );
and  ( new_n50961_, new_n50959_, new_n50955_ );
nor  ( new_n50962_, new_n50808_, new_n757_ );
xor  ( new_n50963_, new_n47046_, new_n520_ );
nor  ( new_n50964_, new_n50963_, new_n755_ );
nor  ( new_n50965_, new_n50964_, new_n50962_ );
nor  ( new_n50966_, new_n50965_, new_n50961_ );
nor  ( new_n50967_, new_n50966_, new_n50960_ );
nor  ( new_n50968_, new_n50967_, new_n50951_ );
or   ( new_n50969_, new_n50968_, new_n50950_ );
xor  ( new_n50970_, new_n50778_, new_n50777_ );
nand ( new_n50971_, new_n50970_, new_n50969_ );
xor  ( new_n50972_, new_n50970_, new_n50969_ );
xor  ( new_n50973_, new_n50824_, new_n50823_ );
nand ( new_n50974_, new_n50973_, new_n50972_ );
and  ( new_n50975_, new_n50974_, new_n50971_ );
nor  ( new_n50976_, new_n50975_, new_n50934_ );
xor  ( new_n50977_, new_n50975_, new_n50934_ );
xor  ( new_n50978_, new_n50829_, new_n50828_ );
and  ( new_n50979_, new_n50978_, new_n50977_ );
or   ( new_n50980_, new_n50979_, new_n50976_ );
xor  ( new_n50981_, new_n50749_, new_n50628_ );
and  ( new_n50982_, new_n50981_, new_n50980_ );
and  ( new_n50983_, new_n50940_, new_n280_ );
xor  ( new_n50984_, new_n49758_, new_n275_ );
nor  ( new_n50985_, new_n50984_, new_n283_ );
nor  ( new_n50986_, new_n50985_, new_n50983_ );
xor  ( new_n50987_, new_n43985_, new_n4705_ );
or   ( new_n50988_, new_n50987_, new_n5207_ );
or   ( new_n50989_, new_n50728_, new_n5209_ );
and  ( new_n50990_, new_n50989_, new_n50988_ );
nor  ( new_n50991_, new_n50990_, new_n50986_ );
nor  ( new_n50992_, new_n50639_, new_n2124_ );
xor  ( new_n50993_, new_n45584_, RIbb2e9e0_27 );
and  ( new_n50994_, new_n50993_, new_n2002_ );
nor  ( new_n50995_, new_n50994_, new_n50992_ );
and  ( new_n50996_, new_n50990_, new_n50986_ );
nor  ( new_n50997_, new_n50996_, new_n50995_ );
or   ( new_n50998_, new_n50997_, new_n50991_ );
xor  ( new_n50999_, new_n50769_, new_n50763_ );
xor  ( new_n51000_, new_n50999_, new_n50774_ );
nand ( new_n51001_, new_n51000_, new_n50998_ );
or   ( new_n51002_, new_n51000_, new_n50998_ );
xor  ( new_n51003_, new_n50707_, new_n50706_ );
nand ( new_n51004_, new_n51003_, new_n51002_ );
and  ( new_n51005_, new_n51004_, new_n51001_ );
xor  ( new_n51006_, new_n43803_, new_n6163_ );
or   ( new_n51007_, new_n51006_, new_n6645_ );
or   ( new_n51008_, new_n50681_, new_n6647_ );
and  ( new_n51009_, new_n51008_, new_n51007_ );
xor  ( new_n51010_, new_n43888_, RIbb2e080_47 );
nand ( new_n51011_, new_n51010_, new_n5917_ );
nand ( new_n51012_, new_n50665_, new_n5915_ );
and  ( new_n51013_, new_n51012_, new_n51011_ );
nor  ( new_n51014_, new_n51013_, new_n51009_ );
and  ( new_n51015_, new_n50654_, new_n3731_ );
xor  ( new_n51016_, new_n44407_, RIbb2e530_37 );
and  ( new_n51017_, new_n51016_, new_n3733_ );
nor  ( new_n51018_, new_n51017_, new_n51015_ );
and  ( new_n51019_, new_n51013_, new_n51009_ );
nor  ( new_n51020_, new_n51019_, new_n51018_ );
nor  ( new_n51021_, new_n51020_, new_n51014_ );
xor  ( new_n51022_, new_n44785_, new_n2797_ );
or   ( new_n51023_, new_n51022_, new_n3117_ );
or   ( new_n51024_, new_n50672_, new_n3119_ );
and  ( new_n51025_, new_n51024_, new_n51023_ );
or   ( new_n51026_, new_n50659_, new_n3463_ );
xor  ( new_n51027_, new_n44600_, new_n3113_ );
or   ( new_n51028_, new_n51027_, new_n3461_ );
and  ( new_n51029_, new_n51028_, new_n51026_ );
or   ( new_n51030_, new_n51029_, new_n51025_ );
xor  ( new_n51031_, new_n43894_, RIbb2dea0_51 );
and  ( new_n51032_, new_n51031_, new_n6910_ );
nor  ( new_n51033_, new_n50711_, new_n7186_ );
or   ( new_n51034_, new_n51033_, new_n51032_ );
xor  ( new_n51035_, new_n51029_, new_n51025_ );
nand ( new_n51036_, new_n51035_, new_n51034_ );
and  ( new_n51037_, new_n51036_, new_n51030_ );
nor  ( new_n51038_, new_n51037_, new_n51021_ );
and  ( new_n51039_, new_n51037_, new_n51021_ );
xor  ( new_n51040_, new_n45204_, RIbb2e8f0_29 );
nand ( new_n51041_, new_n51040_, new_n2244_ );
or   ( new_n51042_, new_n50737_, new_n2427_ );
and  ( new_n51043_, new_n51042_, new_n51041_ );
xor  ( new_n51044_, new_n44974_, new_n2421_ );
or   ( new_n51045_, new_n51044_, new_n2807_ );
or   ( new_n51046_, new_n50732_, new_n2809_ );
and  ( new_n51047_, new_n51046_, new_n51045_ );
nor  ( new_n51048_, new_n51047_, new_n51043_ );
and  ( new_n51049_, new_n50676_, new_n5371_ );
xor  ( new_n51050_, new_n43956_, new_n5203_ );
nor  ( new_n51051_, new_n51050_, new_n5604_ );
nor  ( new_n51052_, new_n51051_, new_n51049_ );
and  ( new_n51053_, new_n51047_, new_n51043_ );
nor  ( new_n51054_, new_n51053_, new_n51052_ );
nor  ( new_n51055_, new_n51054_, new_n51048_ );
nor  ( new_n51056_, new_n51055_, new_n51039_ );
nor  ( new_n51057_, new_n51056_, new_n51038_ );
or   ( new_n51058_, new_n51057_, new_n51005_ );
xor  ( new_n51059_, new_n49265_, new_n309_ );
or   ( new_n51060_, new_n51059_, new_n317_ );
or   ( new_n51061_, new_n50698_, new_n320_ );
and  ( new_n51062_, new_n51061_, new_n51060_ );
xor  ( new_n51063_, new_n43914_, new_n4292_ );
or   ( new_n51064_, new_n51063_, new_n4709_ );
or   ( new_n51065_, new_n50634_, new_n4711_ );
and  ( new_n51066_, new_n51065_, new_n51064_ );
nor  ( new_n51067_, new_n51066_, new_n51062_ );
and  ( new_n51068_, new_n50947_, new_n1739_ );
xor  ( new_n51069_, new_n45597_, RIbb2ead0_25 );
and  ( new_n51070_, new_n51069_, new_n1741_ );
or   ( new_n51071_, new_n51070_, new_n51068_ );
xor  ( new_n51072_, new_n51066_, new_n51062_ );
and  ( new_n51073_, new_n51072_, new_n51071_ );
nor  ( new_n51074_, new_n51073_, new_n51067_ );
xor  ( new_n51075_, new_n43787_, RIbb2ddb0_53 );
nand ( new_n51076_, new_n51075_, new_n7489_ );
or   ( new_n51077_, new_n50767_, new_n7734_ );
and  ( new_n51078_, new_n51077_, new_n51076_ );
nand ( new_n51079_, new_n50702_, new_n4032_ );
xor  ( new_n51080_, new_n44218_, new_n3892_ );
or   ( new_n51081_, new_n51080_, new_n4302_ );
and  ( new_n51082_, new_n51081_, new_n51079_ );
or   ( new_n51083_, new_n51082_, new_n51078_ );
xor  ( new_n51084_, new_n46037_, new_n1355_ );
nor  ( new_n51085_, new_n51084_, new_n1593_ );
nor  ( new_n51086_, new_n50714_, new_n1595_ );
nor  ( new_n51087_, new_n51086_, new_n51085_ );
not  ( new_n51088_, new_n51087_ );
xor  ( new_n51089_, new_n51082_, new_n51078_ );
nand ( new_n51090_, new_n51089_, new_n51088_ );
and  ( new_n51091_, new_n51090_, new_n51083_ );
nor  ( new_n51092_, new_n51091_, new_n51074_ );
xor  ( new_n51093_, new_n51091_, new_n51074_ );
xnor ( new_n51094_, new_n50815_, new_n50811_ );
nand ( new_n51095_, new_n51094_, new_n50820_ );
not  ( new_n51096_, new_n50816_ );
nand ( new_n51097_, new_n50822_, new_n51096_ );
and  ( new_n51098_, new_n51097_, new_n51095_ );
and  ( new_n51099_, new_n51098_, new_n51093_ );
nor  ( new_n51100_, new_n51099_, new_n51092_ );
xnor ( new_n51101_, new_n51057_, new_n51005_ );
or   ( new_n51102_, new_n51101_, new_n51100_ );
and  ( new_n51103_, new_n51102_, new_n51058_ );
xor  ( new_n51104_, new_n50745_, new_n50744_ );
xor  ( new_n51105_, new_n50648_, new_n50647_ );
nand ( new_n51106_, new_n51105_, new_n51104_ );
xor  ( new_n51107_, new_n51105_, new_n51104_ );
xor  ( new_n51108_, new_n50723_, new_n50722_ );
xor  ( new_n51109_, new_n50684_, new_n50683_ );
or   ( new_n51110_, new_n51109_, new_n51108_ );
xor  ( new_n51111_, new_n50741_, new_n50740_ );
and  ( new_n51112_, new_n51109_, new_n51108_ );
or   ( new_n51113_, new_n51112_, new_n51111_ );
and  ( new_n51114_, new_n51113_, new_n51110_ );
nand ( new_n51115_, new_n51114_, new_n51107_ );
and  ( new_n51116_, new_n51115_, new_n51106_ );
nor  ( new_n51117_, new_n51116_, new_n51103_ );
xor  ( new_n51118_, new_n51116_, new_n51103_ );
xor  ( new_n51119_, new_n50689_, new_n50651_ );
nand ( new_n51120_, new_n51119_, new_n50747_ );
or   ( new_n51121_, new_n50747_, new_n50692_ );
or   ( new_n51122_, new_n51121_, new_n50691_ );
and  ( new_n51123_, new_n51122_, new_n51120_ );
and  ( new_n51124_, new_n51123_, new_n51118_ );
or   ( new_n51125_, new_n51124_, new_n51117_ );
xor  ( new_n51126_, new_n50981_, new_n50980_ );
and  ( new_n51127_, new_n51126_, new_n51125_ );
nor  ( new_n51128_, new_n51127_, new_n50982_ );
xor  ( new_n51129_, new_n50753_, new_n50751_ );
xor  ( new_n51130_, new_n51129_, new_n50851_ );
or   ( new_n51131_, new_n51130_, new_n51128_ );
xor  ( new_n51132_, new_n51130_, new_n51128_ );
not  ( new_n51133_, new_n51132_ );
xor  ( new_n51134_, new_n50642_, new_n50641_ );
xnor ( new_n51135_, new_n50661_, new_n50657_ );
nand ( new_n51136_, new_n51135_, new_n50667_ );
not  ( new_n51137_, new_n50668_ );
or   ( new_n51138_, new_n51137_, new_n50662_ );
and  ( new_n51139_, new_n51138_, new_n51136_ );
and  ( new_n51140_, new_n51139_, new_n51134_ );
xor  ( new_n51141_, RIbb32f40_183, RIbb2bec0_119 );
xnor ( new_n51142_, new_n51141_, new_n50783_ );
and  ( new_n51143_, new_n51142_, new_n43880_ );
xor  ( new_n51144_, new_n50894_, new_n43945_ );
not  ( new_n51145_, new_n51144_ );
or   ( new_n51146_, new_n51145_, new_n43983_ );
nor  ( new_n51147_, new_n50788_, new_n43880_ );
or   ( new_n51148_, new_n50789_, new_n43977_ );
or   ( new_n51149_, new_n51148_, new_n51147_ );
nand ( new_n51150_, new_n51149_, new_n51146_ );
nand ( new_n51151_, new_n51150_, new_n51143_ );
and  ( new_n51152_, new_n50456_, new_n295_ );
and  ( new_n51153_, new_n50792_, new_n43949_ );
nor  ( new_n51154_, new_n51153_, new_n51152_ );
xnor ( new_n51155_, new_n51150_, new_n51143_ );
or   ( new_n51156_, new_n51155_, new_n51154_ );
and  ( new_n51157_, new_n51156_, new_n51151_ );
or   ( new_n51158_, new_n50952_, new_n899_ );
xor  ( new_n51159_, new_n47303_, new_n745_ );
or   ( new_n51160_, new_n51159_, new_n897_ );
and  ( new_n51161_, new_n51160_, new_n51158_ );
xor  ( new_n51162_, new_n46619_, new_n1126_ );
or   ( new_n51163_, new_n51162_, new_n1364_ );
nand ( new_n51164_, new_n50906_, new_n1251_ );
and  ( new_n51165_, new_n51164_, new_n51163_ );
nor  ( new_n51166_, new_n51165_, new_n51161_ );
nor  ( new_n51167_, new_n50957_, new_n1137_ );
xor  ( new_n51168_, new_n46962_, new_n893_ );
nor  ( new_n51169_, new_n51168_, new_n1135_ );
nor  ( new_n51170_, new_n51169_, new_n51167_ );
and  ( new_n51171_, new_n51165_, new_n51161_ );
nor  ( new_n51172_, new_n51171_, new_n51170_ );
nor  ( new_n51173_, new_n51172_, new_n51166_ );
nor  ( new_n51174_, new_n51173_, new_n51157_ );
xor  ( new_n51175_, new_n48518_, RIbb2f160_11 );
nand ( new_n51176_, new_n51175_, new_n373_ );
or   ( new_n51177_, new_n50915_, new_n411_ );
and  ( new_n51178_, new_n51177_, new_n51176_ );
or   ( new_n51179_, new_n50963_, new_n757_ );
xor  ( new_n51180_, new_n47296_, new_n520_ );
or   ( new_n51181_, new_n51180_, new_n755_ );
and  ( new_n51182_, new_n51181_, new_n51179_ );
nor  ( new_n51183_, new_n51182_, new_n51178_ );
xor  ( new_n51184_, new_n48039_, RIbb2f070_13 );
and  ( new_n51185_, new_n51184_, new_n456_ );
nor  ( new_n51186_, new_n50921_, new_n526_ );
or   ( new_n51187_, new_n51186_, new_n51185_ );
xor  ( new_n51188_, new_n51182_, new_n51178_ );
and  ( new_n51189_, new_n51188_, new_n51187_ );
or   ( new_n51190_, new_n51189_, new_n51183_ );
xor  ( new_n51191_, new_n51173_, new_n51157_ );
and  ( new_n51192_, new_n51191_, new_n51190_ );
or   ( new_n51193_, new_n51192_, new_n51174_ );
xor  ( new_n51194_, new_n51139_, new_n51134_ );
and  ( new_n51195_, new_n51194_, new_n51193_ );
nor  ( new_n51196_, new_n51195_, new_n51140_ );
not  ( new_n51197_, new_n51196_ );
xor  ( new_n51198_, new_n50687_, new_n50686_ );
and  ( new_n51199_, new_n51198_, new_n51197_ );
xor  ( new_n51200_, new_n51198_, new_n51197_ );
xor  ( new_n51201_, new_n50932_, new_n50931_ );
and  ( new_n51202_, new_n51201_, new_n51200_ );
or   ( new_n51203_, new_n51202_, new_n51199_ );
xor  ( new_n51204_, new_n50845_, new_n50844_ );
and  ( new_n51205_, new_n51204_, new_n51203_ );
xor  ( new_n51206_, new_n50973_, new_n50972_ );
xor  ( new_n51207_, new_n50842_, new_n50840_ );
and  ( new_n51208_, new_n51207_, new_n51206_ );
xor  ( new_n51209_, new_n50943_, new_n50942_ );
xnor ( new_n51210_, new_n50902_, new_n50896_ );
xor  ( new_n51211_, new_n51210_, new_n50908_ );
and  ( new_n51212_, new_n51211_, new_n51209_ );
or   ( new_n51213_, new_n51059_, new_n320_ );
xor  ( new_n51214_, new_n49427_, RIbb2f340_7 );
nand ( new_n51215_, new_n51214_, new_n316_ );
and  ( new_n51216_, new_n51215_, new_n51213_ );
nor  ( new_n51217_, RIbb2dbd0_57, RIbb2dc48_56 );
or   ( new_n51218_, new_n51217_, new_n7725_ );
xor  ( new_n51219_, new_n43793_, new_n7722_ );
nand ( new_n51220_, new_n51219_, new_n8042_ );
and  ( new_n51221_, new_n51220_, new_n51218_ );
nor  ( new_n51222_, new_n51221_, new_n51216_ );
xor  ( new_n51223_, new_n48908_, new_n329_ );
nor  ( new_n51224_, new_n51223_, new_n337_ );
and  ( new_n51225_, new_n50911_, new_n334_ );
or   ( new_n51226_, new_n51225_, new_n51224_ );
xor  ( new_n51227_, new_n51221_, new_n51216_ );
and  ( new_n51228_, new_n51227_, new_n51226_ );
or   ( new_n51229_, new_n51228_, new_n51222_ );
xor  ( new_n51230_, new_n51211_, new_n51209_ );
and  ( new_n51231_, new_n51230_, new_n51229_ );
or   ( new_n51232_, new_n51231_, new_n51212_ );
xor  ( new_n51233_, new_n50967_, new_n50951_ );
and  ( new_n51234_, new_n51233_, new_n51232_ );
xor  ( new_n51235_, new_n50929_, new_n50928_ );
xor  ( new_n51236_, new_n51233_, new_n51232_ );
and  ( new_n51237_, new_n51236_, new_n51235_ );
nor  ( new_n51238_, new_n51237_, new_n51234_ );
xnor ( new_n51239_, new_n51207_, new_n51206_ );
nor  ( new_n51240_, new_n51239_, new_n51238_ );
or   ( new_n51241_, new_n51240_, new_n51208_ );
xor  ( new_n51242_, new_n51204_, new_n51203_ );
and  ( new_n51243_, new_n51242_, new_n51241_ );
or   ( new_n51244_, new_n51243_, new_n51205_ );
xor  ( new_n51245_, new_n50884_, new_n50882_ );
nand ( new_n51246_, new_n51245_, new_n51244_ );
or   ( new_n51247_, new_n51245_, new_n51244_ );
xor  ( new_n51248_, new_n50849_, new_n50848_ );
nand ( new_n51249_, new_n51248_, new_n51247_ );
and  ( new_n51250_, new_n51249_, new_n51246_ );
or   ( new_n51251_, new_n51250_, new_n51133_ );
and  ( new_n51252_, new_n51251_, new_n51131_ );
nor  ( new_n51253_, new_n51252_, new_n50889_ );
xor  ( new_n51254_, new_n51252_, new_n50889_ );
xor  ( new_n51255_, new_n50857_, new_n50856_ );
and  ( new_n51256_, new_n51255_, new_n51254_ );
nor  ( new_n51257_, new_n51256_, new_n51253_ );
not  ( new_n51258_, new_n51257_ );
xor  ( new_n51259_, new_n50863_, new_n50862_ );
nor  ( new_n51260_, new_n51259_, new_n51258_ );
and  ( new_n51261_, new_n51259_, new_n51258_ );
xor  ( new_n51262_, new_n51255_, new_n51254_ );
not  ( new_n51263_, new_n51262_ );
xnor ( new_n51264_, new_n50887_, new_n50886_ );
xor  ( new_n51265_, new_n50978_, new_n50977_ );
xor  ( new_n51266_, new_n50877_, new_n50876_ );
and  ( new_n51267_, new_n51266_, new_n51265_ );
xor  ( new_n51268_, new_n51266_, new_n51265_ );
not  ( new_n51269_, new_n51268_ );
xnor ( new_n51270_, new_n51101_, new_n51100_ );
xor  ( new_n51271_, new_n51035_, new_n51034_ );
xnor ( new_n51272_, new_n51047_, new_n51043_ );
xor  ( new_n51273_, new_n51272_, new_n51052_ );
or   ( new_n51274_, new_n51273_, new_n51271_ );
and  ( new_n51275_, new_n51273_, new_n51271_ );
xor  ( new_n51276_, new_n51089_, new_n51088_ );
or   ( new_n51277_, new_n51276_, new_n51275_ );
and  ( new_n51278_, new_n51277_, new_n51274_ );
xor  ( new_n51279_, new_n51000_, new_n50998_ );
xor  ( new_n51280_, new_n51279_, new_n51003_ );
nand ( new_n51281_, new_n51280_, new_n51278_ );
nor  ( new_n51282_, new_n51280_, new_n51278_ );
not  ( new_n51283_, new_n50986_ );
xor  ( new_n51284_, new_n45119_, new_n2421_ );
or   ( new_n51285_, new_n51284_, new_n2807_ );
or   ( new_n51286_, new_n51044_, new_n2809_ );
and  ( new_n51287_, new_n51286_, new_n51285_ );
nor  ( new_n51288_, new_n51287_, new_n51283_ );
xor  ( new_n51289_, new_n45403_, new_n2118_ );
nor  ( new_n51290_, new_n51289_, new_n2425_ );
and  ( new_n51291_, new_n51040_, new_n2242_ );
or   ( new_n51292_, new_n51291_, new_n51290_ );
nand ( new_n51293_, new_n51287_, new_n51283_ );
and  ( new_n51294_, new_n51293_, new_n51292_ );
or   ( new_n51295_, new_n51294_, new_n51288_ );
xor  ( new_n51296_, new_n50990_, new_n51283_ );
nand ( new_n51297_, new_n51296_, new_n50995_ );
not  ( new_n51298_, new_n50991_ );
nand ( new_n51299_, new_n50997_, new_n51298_ );
and  ( new_n51300_, new_n51299_, new_n51297_ );
and  ( new_n51301_, new_n51300_, new_n51295_ );
nor  ( new_n51302_, new_n51300_, new_n51295_ );
xor  ( new_n51303_, new_n43812_, RIbb2e260_43 );
nand ( new_n51304_, new_n51303_, new_n4960_ );
or   ( new_n51305_, new_n50987_, new_n5209_ );
and  ( new_n51306_, new_n51305_, new_n51304_ );
xor  ( new_n51307_, new_n45738_, new_n1840_ );
or   ( new_n51308_, new_n51307_, new_n2122_ );
nand ( new_n51309_, new_n50993_, new_n2000_ );
and  ( new_n51310_, new_n51309_, new_n51308_ );
nor  ( new_n51311_, new_n51310_, new_n51306_ );
or   ( new_n51312_, new_n50900_, new_n44007_ );
or   ( new_n51313_, new_n50791_, new_n302_ );
and  ( new_n51314_, new_n51313_, new_n51312_ );
xor  ( new_n51315_, new_n51142_, new_n43945_ );
not  ( new_n51316_, new_n51315_ );
or   ( new_n51317_, new_n51316_, new_n43983_ );
and  ( new_n51318_, new_n50895_, new_n43879_ );
nand ( new_n51319_, new_n50896_, new_n43978_ );
or   ( new_n51320_, new_n51319_, new_n51318_ );
and  ( new_n51321_, new_n51320_, new_n51317_ );
nor  ( new_n51322_, new_n51321_, new_n51314_ );
and  ( new_n51323_, new_n51214_, new_n314_ );
xor  ( new_n51324_, new_n49488_, RIbb2f340_7 );
and  ( new_n51325_, new_n51324_, new_n316_ );
or   ( new_n51326_, new_n51325_, new_n51323_ );
xor  ( new_n51327_, new_n51321_, new_n51314_ );
and  ( new_n51328_, new_n51327_, new_n51326_ );
nor  ( new_n51329_, new_n51328_, new_n51322_ );
and  ( new_n51330_, new_n51310_, new_n51306_ );
nor  ( new_n51331_, new_n51330_, new_n51329_ );
nor  ( new_n51332_, new_n51331_, new_n51311_ );
nor  ( new_n51333_, new_n51332_, new_n51302_ );
nor  ( new_n51334_, new_n51333_, new_n51301_ );
or   ( new_n51335_, new_n51334_, new_n51282_ );
and  ( new_n51336_, new_n51335_, new_n51281_ );
or   ( new_n51337_, new_n51336_, new_n51270_ );
and  ( new_n51338_, new_n51336_, new_n51270_ );
xnor ( new_n51339_, new_n51098_, new_n51093_ );
xnor ( new_n51340_, new_n50959_, new_n50955_ );
nand ( new_n51341_, new_n51340_, new_n50965_ );
not  ( new_n51342_, new_n50966_ );
or   ( new_n51343_, new_n51342_, new_n50960_ );
and  ( new_n51344_, new_n51343_, new_n51341_ );
xnor ( new_n51345_, new_n50918_, new_n50914_ );
xor  ( new_n51346_, new_n51345_, new_n50923_ );
nand ( new_n51347_, new_n51346_, new_n51344_ );
nor  ( new_n51348_, new_n51346_, new_n51344_ );
xor  ( new_n51349_, new_n43952_, new_n5203_ );
or   ( new_n51350_, new_n51349_, new_n5604_ );
or   ( new_n51351_, new_n51050_, new_n5606_ );
and  ( new_n51352_, new_n51351_, new_n51350_ );
xor  ( new_n51353_, new_n44877_, RIbb2e710_33 );
nand ( new_n51354_, new_n51353_, new_n2930_ );
or   ( new_n51355_, new_n51022_, new_n3119_ );
and  ( new_n51356_, new_n51355_, new_n51354_ );
nor  ( new_n51357_, new_n51356_, new_n51352_ );
xor  ( new_n51358_, new_n43799_, new_n6635_ );
nor  ( new_n51359_, new_n51358_, new_n7184_ );
and  ( new_n51360_, new_n51031_, new_n6908_ );
nor  ( new_n51361_, new_n51360_, new_n51359_ );
not  ( new_n51362_, new_n51361_ );
xor  ( new_n51363_, new_n51356_, new_n51352_ );
and  ( new_n51364_, new_n51363_, new_n51362_ );
nor  ( new_n51365_, new_n51364_, new_n51357_ );
or   ( new_n51366_, new_n51365_, new_n51348_ );
and  ( new_n51367_, new_n51366_, new_n51347_ );
nor  ( new_n51368_, new_n51367_, new_n51339_ );
and  ( new_n51369_, new_n51367_, new_n51339_ );
xor  ( new_n51370_, new_n43884_, RIbb2df90_49 );
nand ( new_n51371_, new_n51370_, new_n6510_ );
or   ( new_n51372_, new_n51006_, new_n6647_ );
and  ( new_n51373_, new_n51372_, new_n51371_ );
xor  ( new_n51374_, new_n44319_, new_n3892_ );
or   ( new_n51375_, new_n51374_, new_n4302_ );
or   ( new_n51376_, new_n51080_, new_n4304_ );
and  ( new_n51377_, new_n51376_, new_n51375_ );
or   ( new_n51378_, new_n51377_, new_n51373_ );
xor  ( new_n51379_, new_n43898_, new_n7174_ );
nor  ( new_n51380_, new_n51379_, new_n7732_ );
and  ( new_n51381_, new_n51075_, new_n7487_ );
nor  ( new_n51382_, new_n51381_, new_n51380_ );
and  ( new_n51383_, new_n51377_, new_n51373_ );
or   ( new_n51384_, new_n51383_, new_n51382_ );
and  ( new_n51385_, new_n51384_, new_n51378_ );
or   ( new_n51386_, new_n51084_, new_n1595_ );
xor  ( new_n51387_, new_n46137_, new_n1355_ );
or   ( new_n51388_, new_n51387_, new_n1593_ );
and  ( new_n51389_, new_n51388_, new_n51386_ );
xor  ( new_n51390_, new_n44183_, new_n4292_ );
or   ( new_n51391_, new_n51390_, new_n4709_ );
or   ( new_n51392_, new_n51063_, new_n4711_ );
and  ( new_n51393_, new_n51392_, new_n51391_ );
or   ( new_n51394_, new_n51393_, new_n51389_ );
xor  ( new_n51395_, new_n45928_, new_n1583_ );
nor  ( new_n51396_, new_n51395_, new_n1844_ );
and  ( new_n51397_, new_n51069_, new_n1739_ );
nor  ( new_n51398_, new_n51397_, new_n51396_ );
and  ( new_n51399_, new_n51393_, new_n51389_ );
or   ( new_n51400_, new_n51399_, new_n51398_ );
and  ( new_n51401_, new_n51400_, new_n51394_ );
nor  ( new_n51402_, new_n51401_, new_n51385_ );
and  ( new_n51403_, new_n51401_, new_n51385_ );
nand ( new_n51404_, new_n51016_, new_n3731_ );
xor  ( new_n51405_, new_n44506_, new_n3457_ );
or   ( new_n51406_, new_n51405_, new_n3896_ );
and  ( new_n51407_, new_n51406_, new_n51404_ );
xor  ( new_n51408_, new_n44681_, new_n3113_ );
or   ( new_n51409_, new_n51408_, new_n3461_ );
or   ( new_n51410_, new_n51027_, new_n3463_ );
and  ( new_n51411_, new_n51410_, new_n51409_ );
nor  ( new_n51412_, new_n51411_, new_n51407_ );
and  ( new_n51413_, new_n51411_, new_n51407_ );
xor  ( new_n51414_, new_n43937_, RIbb2e080_47 );
and  ( new_n51415_, new_n51414_, new_n5917_ );
and  ( new_n51416_, new_n51010_, new_n5915_ );
nor  ( new_n51417_, new_n51416_, new_n51415_ );
nor  ( new_n51418_, new_n51417_, new_n51413_ );
nor  ( new_n51419_, new_n51418_, new_n51412_ );
nor  ( new_n51420_, new_n51419_, new_n51403_ );
nor  ( new_n51421_, new_n51420_, new_n51402_ );
nor  ( new_n51422_, new_n51421_, new_n51369_ );
nor  ( new_n51423_, new_n51422_, new_n51368_ );
or   ( new_n51424_, new_n51423_, new_n51338_ );
and  ( new_n51425_, new_n51424_, new_n51337_ );
nor  ( new_n51426_, new_n51425_, new_n51269_ );
or   ( new_n51427_, new_n51426_, new_n51267_ );
xor  ( new_n51428_, new_n51126_, new_n51125_ );
nand ( new_n51429_, new_n51428_, new_n51427_ );
nor  ( new_n51430_, new_n51428_, new_n51427_ );
xnor ( new_n51431_, new_n51114_, new_n51107_ );
xnor ( new_n51432_, new_n51037_, new_n51021_ );
and  ( new_n51433_, new_n51432_, new_n51055_ );
not  ( new_n51434_, new_n51038_ );
and  ( new_n51435_, new_n51056_, new_n51434_ );
or   ( new_n51436_, new_n51435_, new_n51433_ );
xor  ( new_n51437_, new_n51072_, new_n51071_ );
xnor ( new_n51438_, new_n51013_, new_n51009_ );
nand ( new_n51439_, new_n51438_, new_n51018_ );
not  ( new_n51440_, new_n51020_ );
or   ( new_n51441_, new_n51440_, new_n51014_ );
and  ( new_n51442_, new_n51441_, new_n51439_ );
nand ( new_n51443_, new_n51442_, new_n51437_ );
nor  ( new_n51444_, new_n51442_, new_n51437_ );
xor  ( new_n51445_, RIbb32fb8_184, RIbb2be48_120 );
xor  ( new_n51446_, new_n51445_, new_n49476_ );
and  ( new_n51447_, new_n51446_, new_n43880_ );
nand ( new_n51448_, new_n51447_, new_n8257_ );
xor  ( new_n51449_, new_n50115_, new_n275_ );
nor  ( new_n51450_, new_n51449_, new_n283_ );
nor  ( new_n51451_, new_n50984_, new_n286_ );
or   ( new_n51452_, new_n51451_, new_n51450_ );
xor  ( new_n51453_, new_n51447_, new_n8257_ );
nand ( new_n51454_, new_n51453_, new_n51452_ );
and  ( new_n51455_, new_n51454_, new_n51448_ );
xor  ( new_n51456_, new_n46958_, new_n893_ );
or   ( new_n51457_, new_n51456_, new_n1135_ );
or   ( new_n51458_, new_n51168_, new_n1137_ );
and  ( new_n51459_, new_n51458_, new_n51457_ );
or   ( new_n51460_, new_n51180_, new_n757_ );
xor  ( new_n51461_, new_n47640_, new_n520_ );
or   ( new_n51462_, new_n51461_, new_n755_ );
and  ( new_n51463_, new_n51462_, new_n51460_ );
nor  ( new_n51464_, new_n51463_, new_n51459_ );
and  ( new_n51465_, new_n51463_, new_n51459_ );
xor  ( new_n51466_, new_n47046_, new_n745_ );
nor  ( new_n51467_, new_n51466_, new_n897_ );
nor  ( new_n51468_, new_n51159_, new_n899_ );
nor  ( new_n51469_, new_n51468_, new_n51467_ );
nor  ( new_n51470_, new_n51469_, new_n51465_ );
nor  ( new_n51471_, new_n51470_, new_n51464_ );
or   ( new_n51472_, new_n51471_, new_n51455_ );
xor  ( new_n51473_, RIbb33030_185, RIbb2bdd0_121 );
nor  ( new_n51474_, new_n43613_, new_n43533_ );
nor  ( new_n51475_, new_n51474_, new_n43513_ );
nor  ( new_n51476_, new_n51475_, new_n43609_ );
xnor ( new_n51477_, new_n51476_, new_n51473_ );
and  ( new_n51478_, new_n51477_, new_n43880_ );
not  ( new_n51479_, new_n51478_ );
or   ( new_n51480_, new_n51387_, new_n1595_ );
xor  ( new_n51481_, new_n46427_, RIbb2ebc0_23 );
nand ( new_n51482_, new_n51481_, new_n1476_ );
and  ( new_n51483_, new_n51482_, new_n51480_ );
nor  ( new_n51484_, new_n51483_, new_n51479_ );
xor  ( new_n51485_, new_n46789_, new_n1126_ );
nor  ( new_n51486_, new_n51485_, new_n1364_ );
nor  ( new_n51487_, new_n51162_, new_n1366_ );
or   ( new_n51488_, new_n51487_, new_n51486_ );
xor  ( new_n51489_, new_n51483_, new_n51479_ );
and  ( new_n51490_, new_n51489_, new_n51488_ );
or   ( new_n51491_, new_n51490_, new_n51484_ );
xor  ( new_n51492_, new_n51471_, new_n51455_ );
nand ( new_n51493_, new_n51492_, new_n51491_ );
and  ( new_n51494_, new_n51493_, new_n51472_ );
or   ( new_n51495_, new_n51494_, new_n51444_ );
and  ( new_n51496_, new_n51495_, new_n51443_ );
or   ( new_n51497_, new_n51496_, new_n51436_ );
nand ( new_n51498_, new_n51496_, new_n51436_ );
xor  ( new_n51499_, new_n51109_, new_n51108_ );
xor  ( new_n51500_, new_n51499_, new_n51111_ );
nand ( new_n51501_, new_n51500_, new_n51498_ );
and  ( new_n51502_, new_n51501_, new_n51497_ );
nor  ( new_n51503_, new_n51502_, new_n51431_ );
xor  ( new_n51504_, new_n51201_, new_n51200_ );
xor  ( new_n51505_, new_n51502_, new_n51431_ );
and  ( new_n51506_, new_n51505_, new_n51504_ );
or   ( new_n51507_, new_n51506_, new_n51503_ );
xor  ( new_n51508_, new_n51123_, new_n51118_ );
and  ( new_n51509_, new_n51508_, new_n51507_ );
xor  ( new_n51510_, new_n51508_, new_n51507_ );
xor  ( new_n51511_, new_n51242_, new_n51241_ );
and  ( new_n51512_, new_n51511_, new_n51510_ );
nor  ( new_n51513_, new_n51512_, new_n51509_ );
or   ( new_n51514_, new_n51513_, new_n51430_ );
and  ( new_n51515_, new_n51514_, new_n51429_ );
or   ( new_n51516_, new_n51515_, new_n51264_ );
nand ( new_n51517_, new_n51515_, new_n51264_ );
xor  ( new_n51518_, new_n51250_, new_n51133_ );
nand ( new_n51519_, new_n51518_, new_n51517_ );
and  ( new_n51520_, new_n51519_, new_n51516_ );
and  ( new_n51521_, new_n51520_, new_n51263_ );
nor  ( new_n51522_, new_n51520_, new_n51263_ );
xor  ( new_n51523_, new_n51425_, new_n51269_ );
xnor ( new_n51524_, new_n51239_, new_n51238_ );
xor  ( new_n51525_, new_n43803_, new_n6635_ );
or   ( new_n51526_, new_n51525_, new_n7184_ );
or   ( new_n51527_, new_n51358_, new_n7186_ );
and  ( new_n51528_, new_n51527_, new_n51526_ );
xor  ( new_n51529_, new_n44218_, RIbb2e350_41 );
nand ( new_n51530_, new_n51529_, new_n4543_ );
or   ( new_n51531_, new_n51390_, new_n4711_ );
and  ( new_n51532_, new_n51531_, new_n51530_ );
or   ( new_n51533_, new_n51532_, new_n51528_ );
xor  ( new_n51534_, new_n43787_, RIbb2dcc0_55 );
and  ( new_n51535_, new_n51534_, new_n8042_ );
and  ( new_n51536_, new_n51219_, new_n8040_ );
nor  ( new_n51537_, new_n51536_, new_n51535_ );
and  ( new_n51538_, new_n51532_, new_n51528_ );
or   ( new_n51539_, new_n51538_, new_n51537_ );
and  ( new_n51540_, new_n51539_, new_n51533_ );
or   ( new_n51541_, new_n51405_, new_n3898_ );
xor  ( new_n51542_, new_n44600_, RIbb2e530_37 );
nand ( new_n51543_, new_n51542_, new_n3733_ );
and  ( new_n51544_, new_n51543_, new_n51541_ );
xor  ( new_n51545_, new_n44407_, new_n3892_ );
or   ( new_n51546_, new_n51545_, new_n4302_ );
or   ( new_n51547_, new_n51374_, new_n4304_ );
and  ( new_n51548_, new_n51547_, new_n51546_ );
or   ( new_n51549_, new_n51548_, new_n51544_ );
xor  ( new_n51550_, new_n43888_, RIbb2df90_49 );
and  ( new_n51551_, new_n51550_, new_n6510_ );
and  ( new_n51552_, new_n51370_, new_n6508_ );
nor  ( new_n51553_, new_n51552_, new_n51551_ );
and  ( new_n51554_, new_n51548_, new_n51544_ );
or   ( new_n51555_, new_n51554_, new_n51553_ );
and  ( new_n51556_, new_n51555_, new_n51549_ );
nor  ( new_n51557_, new_n51556_, new_n51540_ );
nand ( new_n51558_, new_n51556_, new_n51540_ );
xor  ( new_n51559_, new_n45597_, RIbb2e9e0_27 );
nand ( new_n51560_, new_n51559_, new_n2002_ );
or   ( new_n51561_, new_n51307_, new_n2124_ );
and  ( new_n51562_, new_n51561_, new_n51560_ );
xor  ( new_n51563_, new_n46037_, new_n1583_ );
or   ( new_n51564_, new_n51563_, new_n1844_ );
or   ( new_n51565_, new_n51395_, new_n1846_ );
and  ( new_n51566_, new_n51565_, new_n51564_ );
nor  ( new_n51567_, new_n51566_, new_n51562_ );
xor  ( new_n51568_, new_n43914_, RIbb2e260_43 );
and  ( new_n51569_, new_n51568_, new_n4960_ );
and  ( new_n51570_, new_n51303_, new_n4958_ );
or   ( new_n51571_, new_n51570_, new_n51569_ );
nand ( new_n51572_, new_n51566_, new_n51562_ );
and  ( new_n51573_, new_n51572_, new_n51571_ );
or   ( new_n51574_, new_n51573_, new_n51567_ );
and  ( new_n51575_, new_n51574_, new_n51558_ );
or   ( new_n51576_, new_n51575_, new_n51557_ );
xnor ( new_n51577_, new_n51401_, new_n51385_ );
xor  ( new_n51578_, new_n51577_, new_n51419_ );
and  ( new_n51579_, new_n51578_, new_n51576_ );
or   ( new_n51580_, new_n51578_, new_n51576_ );
xnor ( new_n51581_, new_n51155_, new_n51154_ );
xor  ( new_n51582_, new_n48291_, new_n400_ );
or   ( new_n51583_, new_n51582_, new_n524_ );
nand ( new_n51584_, new_n51184_, new_n454_ );
and  ( new_n51585_, new_n51584_, new_n51583_ );
or   ( new_n51586_, new_n51223_, new_n340_ );
xor  ( new_n51587_, new_n49265_, new_n329_ );
or   ( new_n51588_, new_n51587_, new_n337_ );
and  ( new_n51589_, new_n51588_, new_n51586_ );
or   ( new_n51590_, new_n51589_, new_n51585_ );
xor  ( new_n51591_, new_n48756_, RIbb2f160_11 );
and  ( new_n51592_, new_n51591_, new_n373_ );
and  ( new_n51593_, new_n51175_, new_n371_ );
nor  ( new_n51594_, new_n51593_, new_n51592_ );
and  ( new_n51595_, new_n51589_, new_n51585_ );
or   ( new_n51596_, new_n51595_, new_n51594_ );
and  ( new_n51597_, new_n51596_, new_n51590_ );
nor  ( new_n51598_, new_n51597_, new_n51581_ );
xor  ( new_n51599_, new_n43956_, new_n5594_ );
or   ( new_n51600_, new_n51599_, new_n6173_ );
nand ( new_n51601_, new_n51414_, new_n5915_ );
and  ( new_n51602_, new_n51601_, new_n51600_ );
xor  ( new_n51603_, new_n44785_, RIbb2e620_35 );
nand ( new_n51604_, new_n51603_, new_n3293_ );
or   ( new_n51605_, new_n51408_, new_n3463_ );
and  ( new_n51606_, new_n51605_, new_n51604_ );
nor  ( new_n51607_, new_n51606_, new_n51602_ );
xor  ( new_n51608_, new_n43894_, RIbb2ddb0_53 );
and  ( new_n51609_, new_n51608_, new_n7489_ );
nor  ( new_n51610_, new_n51379_, new_n7734_ );
nor  ( new_n51611_, new_n51610_, new_n51609_ );
and  ( new_n51612_, new_n51606_, new_n51602_ );
nor  ( new_n51613_, new_n51612_, new_n51611_ );
or   ( new_n51614_, new_n51613_, new_n51607_ );
xor  ( new_n51615_, new_n51597_, new_n51581_ );
and  ( new_n51616_, new_n51615_, new_n51614_ );
or   ( new_n51617_, new_n51616_, new_n51598_ );
and  ( new_n51618_, new_n51617_, new_n51580_ );
or   ( new_n51619_, new_n51618_, new_n51579_ );
xnor ( new_n51620_, new_n51367_, new_n51339_ );
xor  ( new_n51621_, new_n51620_, new_n51421_ );
nand ( new_n51622_, new_n51621_, new_n51619_ );
nor  ( new_n51623_, new_n51621_, new_n51619_ );
xnor ( new_n51624_, new_n51346_, new_n51344_ );
xor  ( new_n51625_, new_n51624_, new_n51365_ );
xnor ( new_n51626_, new_n51377_, new_n51373_ );
xor  ( new_n51627_, new_n51626_, new_n51382_ );
xor  ( new_n51628_, new_n51287_, new_n51283_ );
xor  ( new_n51629_, new_n51628_, new_n51292_ );
or   ( new_n51630_, new_n51629_, new_n51627_ );
xor  ( new_n51631_, new_n51363_, new_n51362_ );
and  ( new_n51632_, new_n51629_, new_n51627_ );
or   ( new_n51633_, new_n51632_, new_n51631_ );
and  ( new_n51634_, new_n51633_, new_n51630_ );
and  ( new_n51635_, new_n51634_, new_n51625_ );
xor  ( new_n51636_, new_n50487_, new_n275_ );
or   ( new_n51637_, new_n51636_, new_n283_ );
or   ( new_n51638_, new_n51449_, new_n286_ );
and  ( new_n51639_, new_n51638_, new_n51637_ );
xor  ( new_n51640_, new_n51446_, new_n43950_ );
or   ( new_n51641_, new_n51640_, new_n43983_ );
nor  ( new_n51642_, new_n51142_, new_n43880_ );
or   ( new_n51643_, new_n51143_, new_n43977_ );
or   ( new_n51644_, new_n51643_, new_n51642_ );
and  ( new_n51645_, new_n51644_, new_n51641_ );
nor  ( new_n51646_, new_n51645_, new_n51639_ );
and  ( new_n51647_, new_n51324_, new_n314_ );
xor  ( new_n51648_, new_n49758_, new_n309_ );
nor  ( new_n51649_, new_n51648_, new_n317_ );
or   ( new_n51650_, new_n51649_, new_n51647_ );
xor  ( new_n51651_, new_n51645_, new_n51639_ );
and  ( new_n51652_, new_n51651_, new_n51650_ );
or   ( new_n51653_, new_n51652_, new_n51646_ );
xor  ( new_n51654_, new_n51453_, new_n51452_ );
and  ( new_n51655_, new_n51654_, new_n51653_ );
xor  ( new_n51656_, new_n45584_, RIbb2e8f0_29 );
and  ( new_n51657_, new_n51656_, new_n2244_ );
nor  ( new_n51658_, new_n51289_, new_n2427_ );
or   ( new_n51659_, new_n51658_, new_n51657_ );
xor  ( new_n51660_, new_n51654_, new_n51653_ );
and  ( new_n51661_, new_n51660_, new_n51659_ );
or   ( new_n51662_, new_n51661_, new_n51655_ );
xnor ( new_n51663_, new_n51165_, new_n51161_ );
nand ( new_n51664_, new_n51663_, new_n51170_ );
not  ( new_n51665_, new_n51172_ );
or   ( new_n51666_, new_n51665_, new_n51166_ );
and  ( new_n51667_, new_n51666_, new_n51664_ );
and  ( new_n51668_, new_n51667_, new_n51662_ );
xor  ( new_n51669_, new_n51667_, new_n51662_ );
xnor ( new_n51670_, new_n51310_, new_n51306_ );
nand ( new_n51671_, new_n51670_, new_n51329_ );
not  ( new_n51672_, new_n51331_ );
or   ( new_n51673_, new_n51672_, new_n51311_ );
and  ( new_n51674_, new_n51673_, new_n51671_ );
and  ( new_n51675_, new_n51674_, new_n51669_ );
or   ( new_n51676_, new_n51675_, new_n51668_ );
xor  ( new_n51677_, new_n51634_, new_n51625_ );
and  ( new_n51678_, new_n51677_, new_n51676_ );
nor  ( new_n51679_, new_n51678_, new_n51635_ );
or   ( new_n51680_, new_n51679_, new_n51623_ );
and  ( new_n51681_, new_n51680_, new_n51622_ );
or   ( new_n51682_, new_n51681_, new_n51524_ );
and  ( new_n51683_, new_n51681_, new_n51524_ );
xor  ( new_n51684_, new_n51194_, new_n51193_ );
xor  ( new_n51685_, new_n51236_, new_n51235_ );
nand ( new_n51686_, new_n51685_, new_n51684_ );
xor  ( new_n51687_, new_n51191_, new_n51190_ );
xor  ( new_n51688_, new_n51230_, new_n51229_ );
and  ( new_n51689_, new_n51688_, new_n51687_ );
xor  ( new_n51690_, new_n51227_, new_n51226_ );
xor  ( new_n51691_, new_n51188_, new_n51187_ );
and  ( new_n51692_, new_n51691_, new_n51690_ );
or   ( new_n51693_, new_n51284_, new_n2809_ );
xor  ( new_n51694_, new_n45204_, RIbb2e800_31 );
nand ( new_n51695_, new_n51694_, new_n2615_ );
and  ( new_n51696_, new_n51695_, new_n51693_ );
xor  ( new_n51697_, new_n43985_, new_n5203_ );
or   ( new_n51698_, new_n51697_, new_n5604_ );
or   ( new_n51699_, new_n51349_, new_n5606_ );
and  ( new_n51700_, new_n51699_, new_n51698_ );
nor  ( new_n51701_, new_n51700_, new_n51696_ );
and  ( new_n51702_, new_n51353_, new_n2928_ );
xor  ( new_n51703_, new_n44974_, RIbb2e710_33 );
and  ( new_n51704_, new_n51703_, new_n2930_ );
or   ( new_n51705_, new_n51704_, new_n51702_ );
xor  ( new_n51706_, new_n51700_, new_n51696_ );
and  ( new_n51707_, new_n51706_, new_n51705_ );
or   ( new_n51708_, new_n51707_, new_n51701_ );
xor  ( new_n51709_, new_n51691_, new_n51690_ );
and  ( new_n51710_, new_n51709_, new_n51708_ );
or   ( new_n51711_, new_n51710_, new_n51692_ );
xor  ( new_n51712_, new_n51688_, new_n51687_ );
and  ( new_n51713_, new_n51712_, new_n51711_ );
or   ( new_n51714_, new_n51713_, new_n51689_ );
xor  ( new_n51715_, new_n51685_, new_n51684_ );
nand ( new_n51716_, new_n51715_, new_n51714_ );
and  ( new_n51717_, new_n51716_, new_n51686_ );
or   ( new_n51718_, new_n51717_, new_n51683_ );
nand ( new_n51719_, new_n51718_, new_n51682_ );
and  ( new_n51720_, new_n51719_, new_n51523_ );
xnor ( new_n51721_, new_n51719_, new_n51523_ );
xor  ( new_n51722_, new_n51496_, new_n51436_ );
xor  ( new_n51723_, new_n51722_, new_n51500_ );
xnor ( new_n51724_, new_n51280_, new_n51278_ );
xor  ( new_n51725_, new_n51724_, new_n51334_ );
and  ( new_n51726_, new_n51725_, new_n51723_ );
or   ( new_n51727_, new_n51725_, new_n51723_ );
xnor ( new_n51728_, new_n51273_, new_n51271_ );
xor  ( new_n51729_, new_n51728_, new_n51276_ );
xor  ( new_n51730_, new_n51442_, new_n51437_ );
xor  ( new_n51731_, new_n51730_, new_n51494_ );
nor  ( new_n51732_, new_n51731_, new_n51729_ );
nand ( new_n51733_, new_n51731_, new_n51729_ );
xnor ( new_n51734_, new_n51411_, new_n51407_ );
nand ( new_n51735_, new_n51734_, new_n51417_ );
not  ( new_n51736_, new_n51418_ );
or   ( new_n51737_, new_n51736_, new_n51412_ );
and  ( new_n51738_, new_n51737_, new_n51735_ );
xnor ( new_n51739_, new_n51393_, new_n51389_ );
xor  ( new_n51740_, new_n51739_, new_n51398_ );
and  ( new_n51741_, new_n51740_, new_n51738_ );
or   ( new_n51742_, new_n51144_, new_n44007_ );
or   ( new_n51743_, new_n50900_, new_n302_ );
and  ( new_n51744_, new_n51743_, new_n51742_ );
nor  ( new_n51745_, new_n51744_, new_n51478_ );
xor  ( new_n51746_, new_n46619_, new_n1355_ );
nor  ( new_n51747_, new_n51746_, new_n1593_ );
and  ( new_n51748_, new_n51481_, new_n1474_ );
nor  ( new_n51749_, new_n51748_, new_n51747_ );
and  ( new_n51750_, new_n51744_, new_n51478_ );
nor  ( new_n51751_, new_n51750_, new_n51749_ );
nor  ( new_n51752_, new_n51751_, new_n51745_ );
xor  ( new_n51753_, RIbb330a8_186, RIbb2bd58_122 );
not  ( new_n51754_, new_n51753_ );
and  ( new_n51755_, new_n51754_, new_n51474_ );
not  ( new_n51756_, new_n43609_ );
and  ( new_n51757_, new_n51475_, new_n51756_ );
nor  ( new_n51758_, new_n51757_, new_n51755_ );
and  ( new_n51759_, new_n51758_, new_n43880_ );
nand ( new_n51760_, new_n51759_, new_n8873_ );
xor  ( new_n51761_, new_n51759_, new_n8872_ );
xor  ( new_n51762_, new_n51477_, new_n43945_ );
not  ( new_n51763_, new_n51762_ );
or   ( new_n51764_, new_n51763_, new_n43983_ );
nor  ( new_n51765_, new_n51446_, new_n43880_ );
or   ( new_n51766_, new_n51447_, new_n43977_ );
or   ( new_n51767_, new_n51766_, new_n51765_ );
and  ( new_n51768_, new_n51767_, new_n51764_ );
or   ( new_n51769_, new_n51768_, new_n51761_ );
and  ( new_n51770_, new_n51769_, new_n51760_ );
xor  ( new_n51771_, new_n47303_, new_n893_ );
or   ( new_n51772_, new_n51771_, new_n1135_ );
or   ( new_n51773_, new_n51456_, new_n1137_ );
and  ( new_n51774_, new_n51773_, new_n51772_ );
or   ( new_n51775_, new_n51774_, new_n51770_ );
xor  ( new_n51776_, new_n46962_, new_n1126_ );
nor  ( new_n51777_, new_n51776_, new_n1364_ );
nor  ( new_n51778_, new_n51485_, new_n1366_ );
or   ( new_n51779_, new_n51778_, new_n51777_ );
xor  ( new_n51780_, new_n51774_, new_n51770_ );
nand ( new_n51781_, new_n51780_, new_n51779_ );
and  ( new_n51782_, new_n51781_, new_n51775_ );
nor  ( new_n51783_, new_n51782_, new_n51752_ );
xnor ( new_n51784_, new_n51782_, new_n51752_ );
or   ( new_n51785_, new_n51582_, new_n526_ );
xor  ( new_n51786_, new_n48518_, RIbb2f070_13 );
nand ( new_n51787_, new_n51786_, new_n456_ );
and  ( new_n51788_, new_n51787_, new_n51785_ );
xor  ( new_n51789_, new_n47296_, new_n745_ );
or   ( new_n51790_, new_n51789_, new_n897_ );
or   ( new_n51791_, new_n51466_, new_n899_ );
and  ( new_n51792_, new_n51791_, new_n51790_ );
or   ( new_n51793_, new_n51792_, new_n51788_ );
xor  ( new_n51794_, new_n48039_, RIbb2ef80_15 );
and  ( new_n51795_, new_n51794_, new_n662_ );
nor  ( new_n51796_, new_n51461_, new_n757_ );
nor  ( new_n51797_, new_n51796_, new_n51795_ );
and  ( new_n51798_, new_n51792_, new_n51788_ );
or   ( new_n51799_, new_n51798_, new_n51797_ );
and  ( new_n51800_, new_n51799_, new_n51793_ );
nor  ( new_n51801_, new_n51800_, new_n51784_ );
or   ( new_n51802_, new_n51801_, new_n51783_ );
xor  ( new_n51803_, new_n51740_, new_n51738_ );
and  ( new_n51804_, new_n51803_, new_n51802_ );
or   ( new_n51805_, new_n51804_, new_n51741_ );
and  ( new_n51806_, new_n51805_, new_n51733_ );
or   ( new_n51807_, new_n51806_, new_n51732_ );
and  ( new_n51808_, new_n51807_, new_n51727_ );
or   ( new_n51809_, new_n51808_, new_n51726_ );
xnor ( new_n51810_, new_n51336_, new_n51270_ );
xor  ( new_n51811_, new_n51810_, new_n51423_ );
nand ( new_n51812_, new_n51811_, new_n51809_ );
or   ( new_n51813_, new_n51811_, new_n51809_ );
xor  ( new_n51814_, new_n51505_, new_n51504_ );
nand ( new_n51815_, new_n51814_, new_n51813_ );
and  ( new_n51816_, new_n51815_, new_n51812_ );
nor  ( new_n51817_, new_n51816_, new_n51721_ );
nor  ( new_n51818_, new_n51817_, new_n51720_ );
not  ( new_n51819_, new_n51818_ );
xor  ( new_n51820_, new_n51245_, new_n51244_ );
xor  ( new_n51821_, new_n51820_, new_n51248_ );
nor  ( new_n51822_, new_n51821_, new_n51819_ );
xor  ( new_n51823_, new_n51821_, new_n51819_ );
not  ( new_n51824_, new_n51823_ );
xnor ( new_n51825_, new_n51428_, new_n51427_ );
xor  ( new_n51826_, new_n51825_, new_n51513_ );
nor  ( new_n51827_, new_n51826_, new_n51824_ );
nor  ( new_n51828_, new_n51827_, new_n51822_ );
xor  ( new_n51829_, new_n51515_, new_n51264_ );
xor  ( new_n51830_, new_n51829_, new_n51518_ );
nor  ( new_n51831_, new_n51830_, new_n51828_ );
and  ( new_n51832_, new_n51830_, new_n51828_ );
xor  ( new_n51833_, new_n51826_, new_n51824_ );
xor  ( new_n51834_, new_n51511_, new_n51510_ );
xor  ( new_n51835_, new_n51816_, new_n51721_ );
nor  ( new_n51836_, new_n51835_, new_n51834_ );
xor  ( new_n51837_, new_n51492_, new_n51491_ );
xor  ( new_n51838_, new_n51615_, new_n51614_ );
and  ( new_n51839_, new_n51838_, new_n51837_ );
nand ( new_n51840_, new_n51534_, new_n8040_ );
xor  ( new_n51841_, new_n43898_, new_n7722_ );
or   ( new_n51842_, new_n51841_, new_n8264_ );
and  ( new_n51843_, new_n51842_, new_n51840_ );
or   ( new_n51844_, new_n51525_, new_n7186_ );
xor  ( new_n51845_, new_n43884_, RIbb2dea0_51 );
nand ( new_n51846_, new_n51845_, new_n6910_ );
and  ( new_n51847_, new_n51846_, new_n51844_ );
nor  ( new_n51848_, new_n51847_, new_n51843_ );
and  ( new_n51849_, new_n51847_, new_n51843_ );
xor  ( new_n51850_, new_n44319_, RIbb2e350_41 );
and  ( new_n51851_, new_n51850_, new_n4543_ );
and  ( new_n51852_, new_n51529_, new_n4541_ );
nor  ( new_n51853_, new_n51852_, new_n51851_ );
nor  ( new_n51854_, new_n51853_, new_n51849_ );
nor  ( new_n51855_, new_n51854_, new_n51848_ );
xor  ( new_n51856_, new_n43799_, new_n7174_ );
or   ( new_n51857_, new_n51856_, new_n7732_ );
nand ( new_n51858_, new_n51608_, new_n7487_ );
and  ( new_n51859_, new_n51858_, new_n51857_ );
xor  ( new_n51860_, new_n43952_, new_n5594_ );
or   ( new_n51861_, new_n51860_, new_n6173_ );
or   ( new_n51862_, new_n51599_, new_n6175_ );
and  ( new_n51863_, new_n51862_, new_n51861_ );
or   ( new_n51864_, new_n51863_, new_n51859_ );
xor  ( new_n51865_, new_n44877_, RIbb2e620_35 );
and  ( new_n51866_, new_n51865_, new_n3293_ );
and  ( new_n51867_, new_n51603_, new_n3291_ );
nor  ( new_n51868_, new_n51867_, new_n51866_ );
and  ( new_n51869_, new_n51863_, new_n51859_ );
or   ( new_n51870_, new_n51869_, new_n51868_ );
and  ( new_n51871_, new_n51870_, new_n51864_ );
nor  ( new_n51872_, new_n51871_, new_n51855_ );
nand ( new_n51873_, new_n51871_, new_n51855_ );
xor  ( new_n51874_, new_n43812_, RIbb2e170_45 );
nand ( new_n51875_, new_n51874_, new_n5373_ );
or   ( new_n51876_, new_n51697_, new_n5606_ );
and  ( new_n51877_, new_n51876_, new_n51875_ );
xor  ( new_n51878_, new_n45119_, new_n2797_ );
or   ( new_n51879_, new_n51878_, new_n3117_ );
nand ( new_n51880_, new_n51703_, new_n2928_ );
and  ( new_n51881_, new_n51880_, new_n51879_ );
nor  ( new_n51882_, new_n51881_, new_n51877_ );
and  ( new_n51883_, new_n51881_, new_n51877_ );
xor  ( new_n51884_, new_n45403_, new_n2421_ );
nor  ( new_n51885_, new_n51884_, new_n2807_ );
and  ( new_n51886_, new_n51694_, new_n2613_ );
nor  ( new_n51887_, new_n51886_, new_n51885_ );
nor  ( new_n51888_, new_n51887_, new_n51883_ );
or   ( new_n51889_, new_n51888_, new_n51882_ );
and  ( new_n51890_, new_n51889_, new_n51873_ );
or   ( new_n51891_, new_n51890_, new_n51872_ );
xor  ( new_n51892_, new_n51838_, new_n51837_ );
and  ( new_n51893_, new_n51892_, new_n51891_ );
or   ( new_n51894_, new_n51893_, new_n51839_ );
xnor ( new_n51895_, new_n51300_, new_n51295_ );
xor  ( new_n51896_, new_n51895_, new_n51332_ );
and  ( new_n51897_, new_n51896_, new_n51894_ );
xor  ( new_n51898_, new_n51896_, new_n51894_ );
xor  ( new_n51899_, new_n51709_, new_n51708_ );
xnor ( new_n51900_, new_n51548_, new_n51544_ );
xor  ( new_n51901_, new_n51900_, new_n51553_ );
xor  ( new_n51902_, new_n51566_, new_n51562_ );
xor  ( new_n51903_, new_n51902_, new_n51571_ );
or   ( new_n51904_, new_n51903_, new_n51901_ );
and  ( new_n51905_, new_n51903_, new_n51901_ );
xnor ( new_n51906_, new_n51532_, new_n51528_ );
xor  ( new_n51907_, new_n51906_, new_n51537_ );
or   ( new_n51908_, new_n51907_, new_n51905_ );
and  ( new_n51909_, new_n51908_, new_n51904_ );
or   ( new_n51910_, new_n51909_, new_n51899_ );
xor  ( new_n51911_, new_n43937_, new_n6163_ );
or   ( new_n51912_, new_n51911_, new_n6645_ );
nand ( new_n51913_, new_n51550_, new_n6508_ );
and  ( new_n51914_, new_n51913_, new_n51912_ );
or   ( new_n51915_, new_n51545_, new_n4304_ );
xor  ( new_n51916_, new_n44506_, new_n3892_ );
or   ( new_n51917_, new_n51916_, new_n4302_ );
and  ( new_n51918_, new_n51917_, new_n51915_ );
nor  ( new_n51919_, new_n51918_, new_n51914_ );
xor  ( new_n51920_, new_n44681_, RIbb2e530_37 );
and  ( new_n51921_, new_n51920_, new_n3733_ );
and  ( new_n51922_, new_n51542_, new_n3731_ );
nor  ( new_n51923_, new_n51922_, new_n51921_ );
not  ( new_n51924_, new_n51923_ );
nand ( new_n51925_, new_n51918_, new_n51914_ );
and  ( new_n51926_, new_n51925_, new_n51924_ );
or   ( new_n51927_, new_n51926_, new_n51919_ );
xor  ( new_n51928_, new_n51706_, new_n51705_ );
or   ( new_n51929_, new_n51928_, new_n51927_ );
and  ( new_n51930_, new_n51928_, new_n51927_ );
xnor ( new_n51931_, new_n51606_, new_n51602_ );
nand ( new_n51932_, new_n51931_, new_n51611_ );
not  ( new_n51933_, new_n51607_ );
nand ( new_n51934_, new_n51613_, new_n51933_ );
and  ( new_n51935_, new_n51934_, new_n51932_ );
or   ( new_n51936_, new_n51935_, new_n51930_ );
and  ( new_n51937_, new_n51936_, new_n51929_ );
and  ( new_n51938_, new_n51909_, new_n51899_ );
or   ( new_n51939_, new_n51938_, new_n51937_ );
and  ( new_n51940_, new_n51939_, new_n51910_ );
and  ( new_n51941_, new_n51940_, new_n51898_ );
or   ( new_n51942_, new_n51941_, new_n51897_ );
xor  ( new_n51943_, new_n51715_, new_n51714_ );
and  ( new_n51944_, new_n51943_, new_n51942_ );
xor  ( new_n51945_, new_n51489_, new_n51488_ );
xnor ( new_n51946_, new_n51463_, new_n51459_ );
nand ( new_n51947_, new_n51946_, new_n51469_ );
not  ( new_n51948_, new_n51470_ );
or   ( new_n51949_, new_n51948_, new_n51464_ );
and  ( new_n51950_, new_n51949_, new_n51947_ );
and  ( new_n51951_, new_n51950_, new_n51945_ );
xor  ( new_n51952_, new_n51950_, new_n51945_ );
xnor ( new_n51953_, new_n51589_, new_n51585_ );
xor  ( new_n51954_, new_n51953_, new_n51594_ );
and  ( new_n51955_, new_n51954_, new_n51952_ );
or   ( new_n51956_, new_n51955_, new_n51951_ );
or   ( new_n51957_, new_n51587_, new_n340_ );
xor  ( new_n51958_, new_n49427_, new_n329_ );
or   ( new_n51959_, new_n51958_, new_n337_ );
and  ( new_n51960_, new_n51959_, new_n51957_ );
not  ( new_n51961_, RIbb2db58_58 );
and  ( new_n51962_, new_n8870_, new_n51961_ );
or   ( new_n51963_, new_n51962_, new_n8257_ );
xor  ( new_n51964_, new_n43793_, RIbb2dbd0_57 );
or   ( new_n51965_, new_n51964_, new_n8874_ );
and  ( new_n51966_, new_n51965_, new_n51963_ );
or   ( new_n51967_, new_n51966_, new_n51960_ );
and  ( new_n51968_, new_n51591_, new_n371_ );
xor  ( new_n51969_, new_n48908_, new_n325_ );
nor  ( new_n51970_, new_n51969_, new_n409_ );
or   ( new_n51971_, new_n51970_, new_n51968_ );
xor  ( new_n51972_, new_n51966_, new_n51960_ );
nand ( new_n51973_, new_n51972_, new_n51971_ );
and  ( new_n51974_, new_n51973_, new_n51967_ );
or   ( new_n51975_, new_n51563_, new_n1846_ );
xor  ( new_n51976_, new_n46137_, RIbb2ead0_25 );
nand ( new_n51977_, new_n51976_, new_n1741_ );
and  ( new_n51978_, new_n51977_, new_n51975_ );
xor  ( new_n51979_, new_n44183_, new_n4705_ );
or   ( new_n51980_, new_n51979_, new_n5207_ );
nand ( new_n51981_, new_n51568_, new_n4958_ );
and  ( new_n51982_, new_n51981_, new_n51980_ );
or   ( new_n51983_, new_n51982_, new_n51978_ );
xor  ( new_n51984_, new_n45928_, new_n1840_ );
nor  ( new_n51985_, new_n51984_, new_n2122_ );
and  ( new_n51986_, new_n51559_, new_n2000_ );
nor  ( new_n51987_, new_n51986_, new_n51985_ );
and  ( new_n51988_, new_n51982_, new_n51978_ );
or   ( new_n51989_, new_n51988_, new_n51987_ );
and  ( new_n51990_, new_n51989_, new_n51983_ );
nand ( new_n51991_, new_n51990_, new_n51974_ );
nor  ( new_n51992_, new_n51990_, new_n51974_ );
xor  ( new_n51993_, new_n51327_, new_n51326_ );
or   ( new_n51994_, new_n51993_, new_n51992_ );
and  ( new_n51995_, new_n51994_, new_n51991_ );
and  ( new_n51996_, new_n51995_, new_n51956_ );
xor  ( new_n51997_, new_n51995_, new_n51956_ );
xor  ( new_n51998_, new_n51556_, new_n51540_ );
xor  ( new_n51999_, new_n51998_, new_n51574_ );
and  ( new_n52000_, new_n51999_, new_n51997_ );
nor  ( new_n52001_, new_n52000_, new_n51996_ );
not  ( new_n52002_, new_n52001_ );
xor  ( new_n52003_, new_n51712_, new_n51711_ );
and  ( new_n52004_, new_n52003_, new_n52002_ );
xor  ( new_n52005_, new_n52003_, new_n52002_ );
xor  ( new_n52006_, new_n51578_, new_n51576_ );
xor  ( new_n52007_, new_n52006_, new_n51617_ );
and  ( new_n52008_, new_n52007_, new_n52005_ );
nor  ( new_n52009_, new_n52008_, new_n52004_ );
not  ( new_n52010_, new_n52009_ );
xor  ( new_n52011_, new_n51943_, new_n51942_ );
and  ( new_n52012_, new_n52011_, new_n52010_ );
nor  ( new_n52013_, new_n52012_, new_n51944_ );
xor  ( new_n52014_, new_n51681_, new_n51524_ );
xor  ( new_n52015_, new_n52014_, new_n51717_ );
nor  ( new_n52016_, new_n52015_, new_n52013_ );
xnor ( new_n52017_, new_n52015_, new_n52013_ );
xnor ( new_n52018_, new_n51621_, new_n51619_ );
xor  ( new_n52019_, new_n52018_, new_n51679_ );
xor  ( new_n52020_, new_n51725_, new_n51723_ );
xor  ( new_n52021_, new_n52020_, new_n51807_ );
nand ( new_n52022_, new_n52021_, new_n52019_ );
xor  ( new_n52023_, new_n51677_, new_n51676_ );
xor  ( new_n52024_, new_n51731_, new_n51729_ );
xor  ( new_n52025_, new_n52024_, new_n51805_ );
nor  ( new_n52026_, new_n52025_, new_n52023_ );
xor  ( new_n52027_, new_n51803_, new_n51802_ );
xor  ( new_n52028_, new_n51674_, new_n51669_ );
nand ( new_n52029_, new_n52028_, new_n52027_ );
or   ( new_n52030_, new_n51648_, new_n320_ );
xor  ( new_n52031_, new_n50115_, new_n309_ );
or   ( new_n52032_, new_n52031_, new_n317_ );
and  ( new_n52033_, new_n52032_, new_n52030_ );
xor  ( new_n52034_, new_n51758_, new_n43950_ );
or   ( new_n52035_, new_n52034_, new_n43983_ );
nor  ( new_n52036_, new_n51477_, new_n43880_ );
or   ( new_n52037_, new_n51478_, new_n43977_ );
or   ( new_n52038_, new_n52037_, new_n52036_ );
and  ( new_n52039_, new_n52038_, new_n52035_ );
or   ( new_n52040_, new_n52039_, new_n52033_ );
and  ( new_n52041_, new_n51316_, new_n43949_ );
and  ( new_n52042_, new_n51145_, new_n295_ );
nor  ( new_n52043_, new_n52042_, new_n52041_ );
xnor ( new_n52044_, new_n52039_, new_n52033_ );
or   ( new_n52045_, new_n52044_, new_n52043_ );
and  ( new_n52046_, new_n52045_, new_n52040_ );
nand ( new_n52047_, new_n51656_, new_n2242_ );
xor  ( new_n52048_, new_n45738_, new_n2118_ );
or   ( new_n52049_, new_n52048_, new_n2425_ );
and  ( new_n52050_, new_n52049_, new_n52047_ );
nor  ( new_n52051_, new_n52050_, new_n52046_ );
or   ( new_n52052_, new_n51636_, new_n286_ );
xor  ( new_n52053_, new_n50788_, new_n275_ );
or   ( new_n52054_, new_n52053_, new_n283_ );
and  ( new_n52055_, new_n52054_, new_n52052_ );
or   ( new_n52056_, new_n51958_, new_n340_ );
xor  ( new_n52057_, new_n49488_, RIbb2f250_9 );
nand ( new_n52058_, new_n52057_, new_n336_ );
and  ( new_n52059_, new_n52058_, new_n52056_ );
nor  ( new_n52060_, new_n52059_, new_n52055_ );
and  ( new_n52061_, new_n51976_, new_n1739_ );
xor  ( new_n52062_, new_n46427_, RIbb2ead0_25 );
and  ( new_n52063_, new_n52062_, new_n1741_ );
or   ( new_n52064_, new_n52063_, new_n52061_ );
xor  ( new_n52065_, new_n52059_, new_n52055_ );
and  ( new_n52066_, new_n52065_, new_n52064_ );
nor  ( new_n52067_, new_n52066_, new_n52060_ );
xnor ( new_n52068_, new_n52050_, new_n52046_ );
nor  ( new_n52069_, new_n52068_, new_n52067_ );
or   ( new_n52070_, new_n52069_, new_n52051_ );
xor  ( new_n52071_, new_n51660_, new_n51659_ );
and  ( new_n52072_, new_n52071_, new_n52070_ );
or   ( new_n52073_, new_n51789_, new_n899_ );
xor  ( new_n52074_, new_n47640_, new_n745_ );
or   ( new_n52075_, new_n52074_, new_n897_ );
and  ( new_n52076_, new_n52075_, new_n52073_ );
nand ( new_n52077_, new_n51794_, new_n660_ );
xor  ( new_n52078_, new_n48291_, new_n520_ );
or   ( new_n52079_, new_n52078_, new_n755_ );
and  ( new_n52080_, new_n52079_, new_n52077_ );
nor  ( new_n52081_, new_n52080_, new_n52076_ );
and  ( new_n52082_, new_n52080_, new_n52076_ );
xor  ( new_n52083_, new_n48756_, RIbb2f070_13 );
and  ( new_n52084_, new_n52083_, new_n456_ );
and  ( new_n52085_, new_n51786_, new_n454_ );
nor  ( new_n52086_, new_n52085_, new_n52084_ );
nor  ( new_n52087_, new_n52086_, new_n52082_ );
nor  ( new_n52088_, new_n52087_, new_n52081_ );
xor  ( new_n52089_, new_n51744_, new_n51479_ );
nand ( new_n52090_, new_n52089_, new_n51749_ );
not  ( new_n52091_, new_n51751_ );
or   ( new_n52092_, new_n52091_, new_n51745_ );
nand ( new_n52093_, new_n52092_, new_n52090_ );
nor  ( new_n52094_, new_n52093_, new_n52088_ );
xnor ( new_n52095_, new_n52093_, new_n52088_ );
or   ( new_n52096_, new_n51776_, new_n1366_ );
xor  ( new_n52097_, new_n46958_, new_n1126_ );
or   ( new_n52098_, new_n52097_, new_n1364_ );
and  ( new_n52099_, new_n52098_, new_n52096_ );
or   ( new_n52100_, new_n51771_, new_n1137_ );
xor  ( new_n52101_, new_n47046_, new_n893_ );
or   ( new_n52102_, new_n52101_, new_n1135_ );
and  ( new_n52103_, new_n52102_, new_n52100_ );
or   ( new_n52104_, new_n52103_, new_n52099_ );
and  ( new_n52105_, new_n52103_, new_n52099_ );
xor  ( new_n52106_, new_n46789_, new_n1355_ );
nor  ( new_n52107_, new_n52106_, new_n1593_ );
nor  ( new_n52108_, new_n51746_, new_n1595_ );
nor  ( new_n52109_, new_n52108_, new_n52107_ );
or   ( new_n52110_, new_n52109_, new_n52105_ );
and  ( new_n52111_, new_n52110_, new_n52104_ );
nor  ( new_n52112_, new_n52111_, new_n52095_ );
or   ( new_n52113_, new_n52112_, new_n52094_ );
xor  ( new_n52114_, new_n52071_, new_n52070_ );
and  ( new_n52115_, new_n52114_, new_n52113_ );
or   ( new_n52116_, new_n52115_, new_n52072_ );
xor  ( new_n52117_, new_n52028_, new_n52027_ );
nand ( new_n52118_, new_n52117_, new_n52116_ );
and  ( new_n52119_, new_n52118_, new_n52029_ );
nand ( new_n52120_, new_n52025_, new_n52023_ );
and  ( new_n52121_, new_n52120_, new_n52119_ );
or   ( new_n52122_, new_n52121_, new_n52026_ );
nor  ( new_n52123_, new_n52021_, new_n52019_ );
or   ( new_n52124_, new_n52123_, new_n52122_ );
and  ( new_n52125_, new_n52124_, new_n52022_ );
nor  ( new_n52126_, new_n52125_, new_n52017_ );
nor  ( new_n52127_, new_n52126_, new_n52016_ );
not  ( new_n52128_, new_n52127_ );
and  ( new_n52129_, new_n51835_, new_n51834_ );
nor  ( new_n52130_, new_n52129_, new_n52128_ );
nor  ( new_n52131_, new_n52130_, new_n51836_ );
not  ( new_n52132_, new_n52131_ );
and  ( new_n52133_, new_n52132_, new_n51833_ );
xor  ( new_n52134_, new_n49265_, new_n325_ );
or   ( new_n52135_, new_n52134_, new_n409_ );
or   ( new_n52136_, new_n51969_, new_n411_ );
and  ( new_n52137_, new_n52136_, new_n52135_ );
or   ( new_n52138_, new_n52048_, new_n2427_ );
xor  ( new_n52139_, new_n45597_, new_n2118_ );
or   ( new_n52140_, new_n52139_, new_n2425_ );
and  ( new_n52141_, new_n52140_, new_n52138_ );
nor  ( new_n52142_, new_n52141_, new_n52137_ );
and  ( new_n52143_, new_n51874_, new_n5371_ );
xor  ( new_n52144_, new_n43914_, RIbb2e170_45 );
and  ( new_n52145_, new_n52144_, new_n5373_ );
or   ( new_n52146_, new_n52145_, new_n52143_ );
xor  ( new_n52147_, new_n52141_, new_n52137_ );
and  ( new_n52148_, new_n52147_, new_n52146_ );
nor  ( new_n52149_, new_n52148_, new_n52142_ );
not  ( new_n52150_, new_n52149_ );
xor  ( new_n52151_, new_n51651_, new_n51650_ );
nand ( new_n52152_, new_n52151_, new_n52150_ );
xor  ( new_n52153_, new_n52151_, new_n52150_ );
or   ( new_n52154_, new_n51856_, new_n7734_ );
xor  ( new_n52155_, new_n43803_, new_n7174_ );
or   ( new_n52156_, new_n52155_, new_n7732_ );
and  ( new_n52157_, new_n52156_, new_n52154_ );
xor  ( new_n52158_, new_n44407_, new_n4292_ );
or   ( new_n52159_, new_n52158_, new_n4709_ );
nand ( new_n52160_, new_n51850_, new_n4541_ );
and  ( new_n52161_, new_n52160_, new_n52159_ );
or   ( new_n52162_, new_n52161_, new_n52157_ );
and  ( new_n52163_, new_n51845_, new_n6908_ );
xor  ( new_n52164_, new_n43888_, RIbb2dea0_51 );
and  ( new_n52165_, new_n52164_, new_n6910_ );
nor  ( new_n52166_, new_n52165_, new_n52163_ );
and  ( new_n52167_, new_n52161_, new_n52157_ );
or   ( new_n52168_, new_n52167_, new_n52166_ );
nand ( new_n52169_, new_n52168_, new_n52162_ );
nand ( new_n52170_, new_n52169_, new_n52153_ );
and  ( new_n52171_, new_n52170_, new_n52152_ );
or   ( new_n52172_, new_n51911_, new_n6647_ );
xor  ( new_n52173_, new_n43956_, new_n6163_ );
or   ( new_n52174_, new_n52173_, new_n6645_ );
and  ( new_n52175_, new_n52174_, new_n52172_ );
xor  ( new_n52176_, new_n44974_, new_n3113_ );
or   ( new_n52177_, new_n52176_, new_n3461_ );
nand ( new_n52178_, new_n51865_, new_n3291_ );
and  ( new_n52179_, new_n52178_, new_n52177_ );
or   ( new_n52180_, new_n52179_, new_n52175_ );
and  ( new_n52181_, new_n52179_, new_n52175_ );
xor  ( new_n52182_, new_n45204_, RIbb2e710_33 );
and  ( new_n52183_, new_n52182_, new_n2930_ );
nor  ( new_n52184_, new_n51878_, new_n3119_ );
nor  ( new_n52185_, new_n52184_, new_n52183_ );
or   ( new_n52186_, new_n52185_, new_n52181_ );
and  ( new_n52187_, new_n52186_, new_n52180_ );
xor  ( new_n52188_, new_n44785_, new_n3457_ );
or   ( new_n52189_, new_n52188_, new_n3896_ );
nand ( new_n52190_, new_n51920_, new_n3731_ );
and  ( new_n52191_, new_n52190_, new_n52189_ );
or   ( new_n52192_, new_n51916_, new_n4304_ );
xor  ( new_n52193_, new_n44600_, RIbb2e440_39 );
nand ( new_n52194_, new_n52193_, new_n4034_ );
and  ( new_n52195_, new_n52194_, new_n52192_ );
or   ( new_n52196_, new_n52195_, new_n52191_ );
xor  ( new_n52197_, new_n43894_, RIbb2dcc0_55 );
and  ( new_n52198_, new_n52197_, new_n8042_ );
nor  ( new_n52199_, new_n51841_, new_n8266_ );
nor  ( new_n52200_, new_n52199_, new_n52198_ );
and  ( new_n52201_, new_n52195_, new_n52191_ );
or   ( new_n52202_, new_n52201_, new_n52200_ );
and  ( new_n52203_, new_n52202_, new_n52196_ );
or   ( new_n52204_, new_n52203_, new_n52187_ );
and  ( new_n52205_, new_n52203_, new_n52187_ );
xor  ( new_n52206_, new_n43787_, RIbb2dbd0_57 );
nand ( new_n52207_, new_n52206_, new_n8651_ );
or   ( new_n52208_, new_n51964_, new_n8876_ );
and  ( new_n52209_, new_n52208_, new_n52207_ );
or   ( new_n52210_, new_n51979_, new_n5209_ );
xor  ( new_n52211_, new_n44218_, new_n4705_ );
or   ( new_n52212_, new_n52211_, new_n5207_ );
and  ( new_n52213_, new_n52212_, new_n52210_ );
nor  ( new_n52214_, new_n52213_, new_n52209_ );
nor  ( new_n52215_, new_n51984_, new_n2124_ );
xor  ( new_n52216_, new_n46037_, new_n1840_ );
nor  ( new_n52217_, new_n52216_, new_n2122_ );
or   ( new_n52218_, new_n52217_, new_n52215_ );
xor  ( new_n52219_, new_n52213_, new_n52209_ );
and  ( new_n52220_, new_n52219_, new_n52218_ );
nor  ( new_n52221_, new_n52220_, new_n52214_ );
or   ( new_n52222_, new_n52221_, new_n52205_ );
and  ( new_n52223_, new_n52222_, new_n52204_ );
nor  ( new_n52224_, new_n52223_, new_n52171_ );
xor  ( new_n52225_, new_n51918_, new_n51914_ );
xor  ( new_n52226_, new_n52225_, new_n51924_ );
xnor ( new_n52227_, new_n51863_, new_n51859_ );
xor  ( new_n52228_, new_n52227_, new_n51868_ );
and  ( new_n52229_, new_n52228_, new_n52226_ );
xor  ( new_n52230_, new_n52228_, new_n52226_ );
xnor ( new_n52231_, new_n51982_, new_n51978_ );
xor  ( new_n52232_, new_n52231_, new_n51987_ );
and  ( new_n52233_, new_n52232_, new_n52230_ );
or   ( new_n52234_, new_n52233_, new_n52229_ );
xor  ( new_n52235_, new_n52223_, new_n52171_ );
and  ( new_n52236_, new_n52235_, new_n52234_ );
or   ( new_n52237_, new_n52236_, new_n52224_ );
xor  ( new_n52238_, new_n51892_, new_n51891_ );
xor  ( new_n52239_, new_n51999_, new_n51997_ );
xor  ( new_n52240_, new_n52239_, new_n52238_ );
xor  ( new_n52241_, new_n52240_, new_n52237_ );
xor  ( new_n52242_, new_n51954_, new_n51952_ );
xor  ( new_n52243_, new_n51780_, new_n51779_ );
xnor ( new_n52244_, new_n51847_, new_n51843_ );
nand ( new_n52245_, new_n52244_, new_n51853_ );
not  ( new_n52246_, new_n51854_ );
or   ( new_n52247_, new_n52246_, new_n51848_ );
and  ( new_n52248_, new_n52247_, new_n52245_ );
or   ( new_n52249_, new_n52248_, new_n52243_ );
and  ( new_n52250_, new_n52248_, new_n52243_ );
xnor ( new_n52251_, new_n51881_, new_n51877_ );
nand ( new_n52252_, new_n52251_, new_n51887_ );
not  ( new_n52253_, new_n51882_ );
nand ( new_n52254_, new_n51888_, new_n52253_ );
and  ( new_n52255_, new_n52254_, new_n52252_ );
or   ( new_n52256_, new_n52255_, new_n52250_ );
and  ( new_n52257_, new_n52256_, new_n52249_ );
xor  ( new_n52258_, new_n52257_, new_n52242_ );
xor  ( new_n52259_, new_n51871_, new_n51855_ );
xor  ( new_n52260_, new_n52259_, new_n51889_ );
xor  ( new_n52261_, new_n52260_, new_n52258_ );
xnor ( new_n52262_, new_n52068_, new_n52067_ );
or   ( new_n52263_, new_n52031_, new_n320_ );
xor  ( new_n52264_, new_n50487_, new_n309_ );
or   ( new_n52265_, new_n52264_, new_n317_ );
and  ( new_n52266_, new_n52265_, new_n52263_ );
or   ( new_n52267_, new_n52053_, new_n286_ );
xor  ( new_n52268_, new_n50894_, new_n275_ );
or   ( new_n52269_, new_n52268_, new_n283_ );
and  ( new_n52270_, new_n52269_, new_n52267_ );
nor  ( new_n52271_, new_n52270_, new_n52266_ );
and  ( new_n52272_, new_n51316_, new_n295_ );
and  ( new_n52273_, new_n51640_, new_n43949_ );
or   ( new_n52274_, new_n52273_, new_n52272_ );
xor  ( new_n52275_, new_n52270_, new_n52266_ );
and  ( new_n52276_, new_n52275_, new_n52274_ );
or   ( new_n52277_, new_n52276_, new_n52271_ );
nor  ( new_n52278_, new_n43611_, new_n43532_ );
xor  ( new_n52279_, RIbb33120_187, RIbb2bce0_123 );
xnor ( new_n52280_, new_n52279_, new_n52278_ );
and  ( new_n52281_, new_n52280_, new_n43880_ );
or   ( new_n52282_, new_n52281_, new_n52039_ );
and  ( new_n52283_, new_n52281_, new_n52039_ );
and  ( new_n52284_, new_n52057_, new_n334_ );
xor  ( new_n52285_, new_n49758_, new_n329_ );
nor  ( new_n52286_, new_n52285_, new_n337_ );
or   ( new_n52287_, new_n52286_, new_n52284_ );
or   ( new_n52288_, new_n52287_, new_n52283_ );
and  ( new_n52289_, new_n52288_, new_n52282_ );
nand ( new_n52290_, new_n52289_, new_n52277_ );
nor  ( new_n52291_, new_n52289_, new_n52277_ );
xor  ( new_n52292_, RIbb33198_188, RIbb2bc68_124 );
xor  ( new_n52293_, new_n52292_, new_n43531_ );
nor  ( new_n52294_, new_n52293_, new_n43879_ );
nand ( new_n52295_, new_n52294_, new_n9421_ );
and  ( new_n52296_, new_n51640_, new_n295_ );
and  ( new_n52297_, new_n51763_, new_n43949_ );
or   ( new_n52298_, new_n52297_, new_n52296_ );
xor  ( new_n52299_, new_n52294_, new_n9421_ );
nand ( new_n52300_, new_n52299_, new_n52298_ );
and  ( new_n52301_, new_n52300_, new_n52295_ );
or   ( new_n52302_, new_n52106_, new_n1595_ );
xor  ( new_n52303_, new_n46962_, new_n1355_ );
or   ( new_n52304_, new_n52303_, new_n1593_ );
and  ( new_n52305_, new_n52304_, new_n52302_ );
nor  ( new_n52306_, new_n52305_, new_n52301_ );
and  ( new_n52307_, new_n52062_, new_n1739_ );
xor  ( new_n52308_, new_n46619_, new_n1583_ );
nor  ( new_n52309_, new_n52308_, new_n1844_ );
nor  ( new_n52310_, new_n52309_, new_n52307_ );
xnor ( new_n52311_, new_n52305_, new_n52301_ );
nor  ( new_n52312_, new_n52311_, new_n52310_ );
nor  ( new_n52313_, new_n52312_, new_n52306_ );
or   ( new_n52314_, new_n52313_, new_n52291_ );
and  ( new_n52315_, new_n52314_, new_n52290_ );
nor  ( new_n52316_, new_n52315_, new_n52262_ );
xor  ( new_n52317_, new_n47303_, new_n1126_ );
or   ( new_n52318_, new_n52317_, new_n1364_ );
or   ( new_n52319_, new_n52097_, new_n1366_ );
and  ( new_n52320_, new_n52319_, new_n52318_ );
or   ( new_n52321_, new_n52101_, new_n1137_ );
xor  ( new_n52322_, new_n47296_, RIbb2eda0_19 );
nand ( new_n52323_, new_n52322_, new_n1042_ );
and  ( new_n52324_, new_n52323_, new_n52321_ );
nor  ( new_n52325_, new_n52324_, new_n52320_ );
nor  ( new_n52326_, new_n52074_, new_n899_ );
xor  ( new_n52327_, new_n48039_, RIbb2ee90_17 );
and  ( new_n52328_, new_n52327_, new_n822_ );
or   ( new_n52329_, new_n52328_, new_n52326_ );
xor  ( new_n52330_, new_n52324_, new_n52320_ );
and  ( new_n52331_, new_n52330_, new_n52329_ );
nor  ( new_n52332_, new_n52331_, new_n52325_ );
not  ( new_n52333_, new_n52332_ );
xor  ( new_n52334_, new_n52065_, new_n52064_ );
and  ( new_n52335_, new_n52334_, new_n52333_ );
xor  ( new_n52336_, new_n52334_, new_n52333_ );
not  ( new_n52337_, new_n52336_ );
or   ( new_n52338_, new_n52078_, new_n757_ );
xor  ( new_n52339_, new_n48518_, RIbb2ef80_15 );
nand ( new_n52340_, new_n52339_, new_n662_ );
and  ( new_n52341_, new_n52340_, new_n52338_ );
xor  ( new_n52342_, new_n48908_, new_n400_ );
or   ( new_n52343_, new_n52342_, new_n524_ );
nand ( new_n52344_, new_n52083_, new_n454_ );
and  ( new_n52345_, new_n52344_, new_n52343_ );
nor  ( new_n52346_, new_n52345_, new_n52341_ );
and  ( new_n52347_, new_n52345_, new_n52341_ );
nor  ( new_n52348_, RIbb2d9f0_61, RIbb2da68_60 );
not  ( new_n52349_, new_n52348_ );
and  ( new_n52350_, new_n52349_, new_n8872_ );
xor  ( new_n52351_, new_n43793_, new_n8870_ );
and  ( new_n52352_, new_n52351_, new_n9187_ );
nor  ( new_n52353_, new_n52352_, new_n52350_ );
nor  ( new_n52354_, new_n52353_, new_n52347_ );
nor  ( new_n52355_, new_n52354_, new_n52346_ );
nor  ( new_n52356_, new_n52355_, new_n52337_ );
or   ( new_n52357_, new_n52356_, new_n52335_ );
xor  ( new_n52358_, new_n52315_, new_n52262_ );
and  ( new_n52359_, new_n52358_, new_n52357_ );
or   ( new_n52360_, new_n52359_, new_n52316_ );
xor  ( new_n52361_, new_n51903_, new_n51901_ );
xor  ( new_n52362_, new_n52361_, new_n51907_ );
xor  ( new_n52363_, new_n51928_, new_n51927_ );
xor  ( new_n52364_, new_n52363_, new_n51935_ );
xor  ( new_n52365_, new_n52364_, new_n52362_ );
xor  ( new_n52366_, new_n52365_, new_n52360_ );
or   ( new_n52367_, new_n52366_, new_n52261_ );
nand ( new_n52368_, new_n52366_, new_n52261_ );
xor  ( new_n52369_, new_n52232_, new_n52230_ );
xor  ( new_n52370_, new_n52248_, new_n52243_ );
xor  ( new_n52371_, new_n52370_, new_n52255_ );
and  ( new_n52372_, new_n52371_, new_n52369_ );
xnor ( new_n52373_, new_n52371_, new_n52369_ );
xor  ( new_n52374_, new_n43803_, new_n7722_ );
or   ( new_n52375_, new_n52374_, new_n8264_ );
xor  ( new_n52376_, new_n43799_, new_n7722_ );
or   ( new_n52377_, new_n52376_, new_n8266_ );
and  ( new_n52378_, new_n52377_, new_n52375_ );
xor  ( new_n52379_, new_n43787_, new_n8870_ );
or   ( new_n52380_, new_n52379_, new_n9422_ );
nand ( new_n52381_, new_n52351_, new_n9185_ );
and  ( new_n52382_, new_n52381_, new_n52380_ );
nor  ( new_n52383_, new_n52382_, new_n52378_ );
xor  ( new_n52384_, new_n44183_, RIbb2e170_45 );
and  ( new_n52385_, new_n52384_, new_n5371_ );
xor  ( new_n52386_, new_n44218_, RIbb2e170_45 );
and  ( new_n52387_, new_n52386_, new_n5373_ );
nor  ( new_n52388_, new_n52387_, new_n52385_ );
and  ( new_n52389_, new_n52382_, new_n52378_ );
nor  ( new_n52390_, new_n52389_, new_n52388_ );
nor  ( new_n52391_, new_n52390_, new_n52383_ );
xor  ( new_n52392_, new_n45928_, new_n2118_ );
or   ( new_n52393_, new_n52392_, new_n2427_ );
xor  ( new_n52394_, new_n46037_, new_n2118_ );
or   ( new_n52395_, new_n52394_, new_n2425_ );
and  ( new_n52396_, new_n52395_, new_n52393_ );
xor  ( new_n52397_, new_n43914_, new_n5594_ );
or   ( new_n52398_, new_n52397_, new_n6173_ );
xor  ( new_n52399_, new_n43812_, new_n5594_ );
or   ( new_n52400_, new_n52399_, new_n6175_ );
and  ( new_n52401_, new_n52400_, new_n52398_ );
or   ( new_n52402_, new_n52401_, new_n52396_ );
xor  ( new_n52403_, new_n45597_, RIbb2e800_31 );
and  ( new_n52404_, new_n52403_, new_n2615_ );
xor  ( new_n52405_, new_n45738_, RIbb2e800_31 );
and  ( new_n52406_, new_n52405_, new_n2613_ );
nor  ( new_n52407_, new_n52406_, new_n52404_ );
and  ( new_n52408_, new_n52401_, new_n52396_ );
or   ( new_n52409_, new_n52408_, new_n52407_ );
and  ( new_n52410_, new_n52409_, new_n52402_ );
nor  ( new_n52411_, new_n52410_, new_n52391_ );
xor  ( new_n52412_, new_n44506_, new_n4292_ );
or   ( new_n52413_, new_n52412_, new_n4711_ );
xor  ( new_n52414_, new_n44600_, RIbb2e350_41 );
nand ( new_n52415_, new_n52414_, new_n4543_ );
and  ( new_n52416_, new_n52415_, new_n52413_ );
xor  ( new_n52417_, new_n43884_, new_n7174_ );
or   ( new_n52418_, new_n52417_, new_n7734_ );
xor  ( new_n52419_, new_n43888_, new_n7174_ );
or   ( new_n52420_, new_n52419_, new_n7732_ );
and  ( new_n52421_, new_n52420_, new_n52418_ );
nor  ( new_n52422_, new_n52421_, new_n52416_ );
xor  ( new_n52423_, new_n44319_, RIbb2e260_43 );
and  ( new_n52424_, new_n52423_, new_n4958_ );
xor  ( new_n52425_, new_n44407_, RIbb2e260_43 );
and  ( new_n52426_, new_n52425_, new_n4960_ );
nor  ( new_n52427_, new_n52426_, new_n52424_ );
and  ( new_n52428_, new_n52421_, new_n52416_ );
nor  ( new_n52429_, new_n52428_, new_n52427_ );
nor  ( new_n52430_, new_n52429_, new_n52422_ );
xnor ( new_n52431_, new_n52410_, new_n52391_ );
nor  ( new_n52432_, new_n52431_, new_n52430_ );
or   ( new_n52433_, new_n52432_, new_n52411_ );
xor  ( new_n52434_, new_n43894_, new_n8254_ );
or   ( new_n52435_, new_n52434_, new_n8874_ );
xor  ( new_n52436_, new_n43898_, new_n8254_ );
or   ( new_n52437_, new_n52436_, new_n8876_ );
and  ( new_n52438_, new_n52437_, new_n52435_ );
xor  ( new_n52439_, new_n43956_, new_n6635_ );
or   ( new_n52440_, new_n52439_, new_n7184_ );
xor  ( new_n52441_, new_n43937_, RIbb2dea0_51 );
nand ( new_n52442_, new_n52441_, new_n6908_ );
and  ( new_n52443_, new_n52442_, new_n52440_ );
nor  ( new_n52444_, new_n52443_, new_n52438_ );
xor  ( new_n52445_, new_n44681_, RIbb2e440_39 );
and  ( new_n52446_, new_n52445_, new_n4032_ );
xor  ( new_n52447_, new_n44785_, RIbb2e440_39 );
and  ( new_n52448_, new_n52447_, new_n4034_ );
or   ( new_n52449_, new_n52448_, new_n52446_ );
xor  ( new_n52450_, new_n52443_, new_n52438_ );
and  ( new_n52451_, new_n52450_, new_n52449_ );
or   ( new_n52452_, new_n52451_, new_n52444_ );
xor  ( new_n52453_, new_n52330_, new_n52329_ );
or   ( new_n52454_, new_n52453_, new_n52452_ );
and  ( new_n52455_, new_n52453_, new_n52452_ );
xnor ( new_n52456_, new_n52345_, new_n52341_ );
nand ( new_n52457_, new_n52456_, new_n52353_ );
not  ( new_n52458_, new_n52354_ );
or   ( new_n52459_, new_n52458_, new_n52346_ );
and  ( new_n52460_, new_n52459_, new_n52457_ );
or   ( new_n52461_, new_n52460_, new_n52455_ );
and  ( new_n52462_, new_n52461_, new_n52454_ );
nand ( new_n52463_, new_n52462_, new_n52433_ );
nor  ( new_n52464_, new_n52462_, new_n52433_ );
xor  ( new_n52465_, new_n52275_, new_n52274_ );
xor  ( new_n52466_, new_n52281_, new_n52039_ );
xor  ( new_n52467_, new_n52466_, new_n52287_ );
and  ( new_n52468_, new_n52467_, new_n52465_ );
nor  ( new_n52469_, new_n52467_, new_n52465_ );
and  ( new_n52470_, new_n52339_, new_n660_ );
xor  ( new_n52471_, new_n48756_, RIbb2ef80_15 );
and  ( new_n52472_, new_n52471_, new_n662_ );
or   ( new_n52473_, new_n52472_, new_n52470_ );
xor  ( new_n52474_, new_n52299_, new_n52298_ );
and  ( new_n52475_, new_n52474_, new_n52473_ );
nor  ( new_n52476_, new_n52342_, new_n526_ );
xor  ( new_n52477_, new_n49265_, new_n400_ );
nor  ( new_n52478_, new_n52477_, new_n524_ );
nor  ( new_n52479_, new_n52478_, new_n52476_ );
not  ( new_n52480_, new_n52479_ );
xor  ( new_n52481_, new_n52474_, new_n52473_ );
and  ( new_n52482_, new_n52481_, new_n52480_ );
nor  ( new_n52483_, new_n52482_, new_n52475_ );
nor  ( new_n52484_, new_n52483_, new_n52469_ );
nor  ( new_n52485_, new_n52484_, new_n52468_ );
or   ( new_n52486_, new_n52485_, new_n52464_ );
and  ( new_n52487_, new_n52486_, new_n52463_ );
nor  ( new_n52488_, new_n52487_, new_n52373_ );
nor  ( new_n52489_, new_n52488_, new_n52372_ );
nand ( new_n52490_, new_n52489_, new_n52368_ );
and  ( new_n52491_, new_n52490_, new_n52367_ );
nand ( new_n52492_, new_n52491_, new_n52241_ );
xor  ( new_n52493_, new_n52491_, new_n52241_ );
xor  ( new_n52494_, new_n52117_, new_n52116_ );
or   ( new_n52495_, new_n52364_, new_n52362_ );
and  ( new_n52496_, new_n52364_, new_n52362_ );
or   ( new_n52497_, new_n52496_, new_n52360_ );
and  ( new_n52498_, new_n52497_, new_n52495_ );
xor  ( new_n52499_, new_n51909_, new_n51899_ );
xor  ( new_n52500_, new_n52499_, new_n51937_ );
xor  ( new_n52501_, new_n52500_, new_n52498_ );
xor  ( new_n52502_, new_n52501_, new_n52494_ );
nand ( new_n52503_, new_n52502_, new_n52493_ );
and  ( new_n52504_, new_n52503_, new_n52492_ );
xnor ( new_n52505_, new_n52044_, new_n52043_ );
nand ( new_n52506_, new_n52423_, new_n4960_ );
or   ( new_n52507_, new_n52211_, new_n5209_ );
and  ( new_n52508_, new_n52507_, new_n52506_ );
or   ( new_n52509_, new_n52216_, new_n2124_ );
xor  ( new_n52510_, new_n46137_, new_n1840_ );
or   ( new_n52511_, new_n52510_, new_n2122_ );
and  ( new_n52512_, new_n52511_, new_n52509_ );
or   ( new_n52513_, new_n52512_, new_n52508_ );
and  ( new_n52514_, new_n52206_, new_n8649_ );
nor  ( new_n52515_, new_n52436_, new_n8874_ );
nor  ( new_n52516_, new_n52515_, new_n52514_ );
and  ( new_n52517_, new_n52512_, new_n52508_ );
or   ( new_n52518_, new_n52517_, new_n52516_ );
and  ( new_n52519_, new_n52518_, new_n52513_ );
nor  ( new_n52520_, new_n52519_, new_n52505_ );
or   ( new_n52521_, new_n52134_, new_n411_ );
xor  ( new_n52522_, new_n49427_, RIbb2f160_11 );
nand ( new_n52523_, new_n52522_, new_n373_ );
and  ( new_n52524_, new_n52523_, new_n52521_ );
or   ( new_n52525_, new_n52392_, new_n2425_ );
or   ( new_n52526_, new_n52139_, new_n2427_ );
and  ( new_n52527_, new_n52526_, new_n52525_ );
nor  ( new_n52528_, new_n52527_, new_n52524_ );
and  ( new_n52529_, new_n52384_, new_n5373_ );
and  ( new_n52530_, new_n52144_, new_n5371_ );
or   ( new_n52531_, new_n52530_, new_n52529_ );
xor  ( new_n52532_, new_n52527_, new_n52524_ );
and  ( new_n52533_, new_n52532_, new_n52531_ );
nor  ( new_n52534_, new_n52533_, new_n52528_ );
not  ( new_n52535_, new_n52534_ );
xor  ( new_n52536_, new_n52519_, new_n52505_ );
and  ( new_n52537_, new_n52536_, new_n52535_ );
nor  ( new_n52538_, new_n52537_, new_n52520_ );
xnor ( new_n52539_, new_n52111_, new_n52095_ );
nor  ( new_n52540_, new_n52539_, new_n52538_ );
xnor ( new_n52541_, new_n52539_, new_n52538_ );
nand ( new_n52542_, new_n52197_, new_n8040_ );
or   ( new_n52543_, new_n52376_, new_n8264_ );
and  ( new_n52544_, new_n52543_, new_n52542_ );
or   ( new_n52545_, new_n52188_, new_n3898_ );
xor  ( new_n52546_, new_n44877_, new_n3457_ );
or   ( new_n52547_, new_n52546_, new_n3896_ );
and  ( new_n52548_, new_n52547_, new_n52545_ );
nor  ( new_n52549_, new_n52548_, new_n52544_ );
and  ( new_n52550_, new_n52193_, new_n4032_ );
and  ( new_n52551_, new_n52445_, new_n4034_ );
nor  ( new_n52552_, new_n52551_, new_n52550_ );
and  ( new_n52553_, new_n52548_, new_n52544_ );
nor  ( new_n52554_, new_n52553_, new_n52552_ );
nor  ( new_n52555_, new_n52554_, new_n52549_ );
or   ( new_n52556_, new_n52176_, new_n3463_ );
xor  ( new_n52557_, new_n45119_, new_n3113_ );
or   ( new_n52558_, new_n52557_, new_n3461_ );
and  ( new_n52559_, new_n52558_, new_n52556_ );
xor  ( new_n52560_, new_n43952_, new_n6163_ );
or   ( new_n52561_, new_n52560_, new_n6645_ );
or   ( new_n52562_, new_n52173_, new_n6647_ );
and  ( new_n52563_, new_n52562_, new_n52561_ );
or   ( new_n52564_, new_n52563_, new_n52559_ );
and  ( new_n52565_, new_n52182_, new_n2928_ );
xor  ( new_n52566_, new_n45403_, new_n2797_ );
nor  ( new_n52567_, new_n52566_, new_n3117_ );
or   ( new_n52568_, new_n52567_, new_n52565_ );
xor  ( new_n52569_, new_n52563_, new_n52559_ );
nand ( new_n52570_, new_n52569_, new_n52568_ );
and  ( new_n52571_, new_n52570_, new_n52564_ );
nor  ( new_n52572_, new_n52571_, new_n52555_ );
and  ( new_n52573_, new_n52571_, new_n52555_ );
or   ( new_n52574_, new_n52155_, new_n7734_ );
or   ( new_n52575_, new_n52417_, new_n7732_ );
and  ( new_n52576_, new_n52575_, new_n52574_ );
or   ( new_n52577_, new_n52158_, new_n4711_ );
or   ( new_n52578_, new_n52412_, new_n4709_ );
and  ( new_n52579_, new_n52578_, new_n52577_ );
nor  ( new_n52580_, new_n52579_, new_n52576_ );
and  ( new_n52581_, new_n52441_, new_n6910_ );
and  ( new_n52582_, new_n52164_, new_n6908_ );
nor  ( new_n52583_, new_n52582_, new_n52581_ );
and  ( new_n52584_, new_n52579_, new_n52576_ );
nor  ( new_n52585_, new_n52584_, new_n52583_ );
nor  ( new_n52586_, new_n52585_, new_n52580_ );
nor  ( new_n52587_, new_n52586_, new_n52573_ );
nor  ( new_n52588_, new_n52587_, new_n52572_ );
nor  ( new_n52589_, new_n52588_, new_n52541_ );
nor  ( new_n52590_, new_n52589_, new_n52540_ );
not  ( new_n52591_, new_n52590_ );
xor  ( new_n52592_, new_n52114_, new_n52113_ );
and  ( new_n52593_, new_n52592_, new_n52591_ );
xor  ( new_n52594_, new_n52592_, new_n52591_ );
not  ( new_n52595_, new_n52594_ );
xnor ( new_n52596_, new_n52169_, new_n52153_ );
nor  ( new_n52597_, new_n51860_, new_n6175_ );
xor  ( new_n52598_, new_n43985_, RIbb2e080_47 );
and  ( new_n52599_, new_n52598_, new_n5917_ );
or   ( new_n52600_, new_n52599_, new_n52597_ );
xor  ( new_n52601_, new_n51768_, new_n51761_ );
and  ( new_n52602_, new_n52601_, new_n52600_ );
nor  ( new_n52603_, new_n51884_, new_n2809_ );
xor  ( new_n52604_, new_n45584_, RIbb2e800_31 );
and  ( new_n52605_, new_n52604_, new_n2615_ );
nor  ( new_n52606_, new_n52605_, new_n52603_ );
not  ( new_n52607_, new_n52606_ );
xor  ( new_n52608_, new_n52601_, new_n52600_ );
and  ( new_n52609_, new_n52608_, new_n52607_ );
nor  ( new_n52610_, new_n52609_, new_n52602_ );
xor  ( new_n52611_, new_n51972_, new_n51971_ );
xnor ( new_n52612_, new_n51792_, new_n51788_ );
xor  ( new_n52613_, new_n52612_, new_n51797_ );
xor  ( new_n52614_, new_n52613_, new_n52611_ );
xor  ( new_n52615_, new_n52614_, new_n52610_ );
or   ( new_n52616_, new_n52615_, new_n52596_ );
nand ( new_n52617_, new_n52615_, new_n52596_ );
xnor ( new_n52618_, new_n52103_, new_n52099_ );
xor  ( new_n52619_, new_n52618_, new_n52109_ );
xnor ( new_n52620_, new_n52080_, new_n52076_ );
xor  ( new_n52621_, new_n52620_, new_n52086_ );
nor  ( new_n52622_, new_n52621_, new_n52619_ );
and  ( new_n52623_, new_n52621_, new_n52619_ );
xor  ( new_n52624_, new_n52608_, new_n52607_ );
nor  ( new_n52625_, new_n52624_, new_n52623_ );
nor  ( new_n52626_, new_n52625_, new_n52622_ );
nand ( new_n52627_, new_n52626_, new_n52617_ );
and  ( new_n52628_, new_n52627_, new_n52616_ );
nor  ( new_n52629_, new_n52628_, new_n52595_ );
or   ( new_n52630_, new_n52629_, new_n52593_ );
and  ( new_n52631_, new_n52257_, new_n52242_ );
and  ( new_n52632_, new_n52260_, new_n52258_ );
or   ( new_n52633_, new_n52632_, new_n52631_ );
xnor ( new_n52634_, new_n51629_, new_n51627_ );
xor  ( new_n52635_, new_n52634_, new_n51631_ );
xor  ( new_n52636_, new_n51800_, new_n51784_ );
xor  ( new_n52637_, new_n51990_, new_n51974_ );
xor  ( new_n52638_, new_n52637_, new_n51993_ );
nand ( new_n52639_, new_n52638_, new_n52636_ );
nor  ( new_n52640_, new_n52638_, new_n52636_ );
and  ( new_n52641_, new_n52613_, new_n52611_ );
nor  ( new_n52642_, new_n52613_, new_n52611_ );
nor  ( new_n52643_, new_n52642_, new_n52610_ );
nor  ( new_n52644_, new_n52643_, new_n52641_ );
or   ( new_n52645_, new_n52644_, new_n52640_ );
and  ( new_n52646_, new_n52645_, new_n52639_ );
xor  ( new_n52647_, new_n52646_, new_n52635_ );
xor  ( new_n52648_, new_n52647_, new_n52633_ );
nand ( new_n52649_, new_n52648_, new_n52630_ );
not  ( new_n52650_, new_n52034_ );
or   ( new_n52651_, new_n52650_, new_n44007_ );
or   ( new_n52652_, new_n51762_, new_n302_ );
and  ( new_n52653_, new_n52652_, new_n52651_ );
xor  ( new_n52654_, new_n52280_, new_n43945_ );
not  ( new_n52655_, new_n52654_ );
or   ( new_n52656_, new_n52655_, new_n43983_ );
nor  ( new_n52657_, new_n51758_, new_n43880_ );
or   ( new_n52658_, new_n51759_, new_n43977_ );
or   ( new_n52659_, new_n52658_, new_n52657_ );
and  ( new_n52660_, new_n52659_, new_n52656_ );
or   ( new_n52661_, new_n52660_, new_n52653_ );
nor  ( new_n52662_, new_n52285_, new_n340_ );
xor  ( new_n52663_, new_n50115_, new_n329_ );
nor  ( new_n52664_, new_n52663_, new_n337_ );
or   ( new_n52665_, new_n52664_, new_n52662_ );
xor  ( new_n52666_, new_n52660_, new_n52653_ );
nand ( new_n52667_, new_n52666_, new_n52665_ );
and  ( new_n52668_, new_n52667_, new_n52661_ );
nand ( new_n52669_, new_n52598_, new_n5915_ );
or   ( new_n52670_, new_n52399_, new_n6173_ );
and  ( new_n52671_, new_n52670_, new_n52669_ );
nor  ( new_n52672_, new_n52671_, new_n52668_ );
and  ( new_n52673_, new_n52405_, new_n2615_ );
and  ( new_n52674_, new_n52604_, new_n2613_ );
nor  ( new_n52675_, new_n52674_, new_n52673_ );
not  ( new_n52676_, new_n52675_ );
xor  ( new_n52677_, new_n52671_, new_n52668_ );
and  ( new_n52678_, new_n52677_, new_n52676_ );
or   ( new_n52679_, new_n52678_, new_n52672_ );
xor  ( new_n52680_, new_n52147_, new_n52146_ );
nand ( new_n52681_, new_n52680_, new_n52679_ );
xor  ( new_n52682_, new_n52680_, new_n52679_ );
xnor ( new_n52683_, new_n52179_, new_n52175_ );
xor  ( new_n52684_, new_n52683_, new_n52185_ );
nand ( new_n52685_, new_n52684_, new_n52682_ );
and  ( new_n52686_, new_n52685_, new_n52681_ );
xor  ( new_n52687_, new_n52219_, new_n52218_ );
xnor ( new_n52688_, new_n52195_, new_n52191_ );
xor  ( new_n52689_, new_n52688_, new_n52200_ );
nand ( new_n52690_, new_n52689_, new_n52687_ );
or   ( new_n52691_, new_n52689_, new_n52687_ );
xor  ( new_n52692_, new_n52161_, new_n52157_ );
xnor ( new_n52693_, new_n52692_, new_n52166_ );
nand ( new_n52694_, new_n52693_, new_n52691_ );
and  ( new_n52695_, new_n52694_, new_n52690_ );
nor  ( new_n52696_, new_n52695_, new_n52686_ );
nand ( new_n52697_, new_n52695_, new_n52686_ );
xor  ( new_n52698_, new_n52203_, new_n52187_ );
xnor ( new_n52699_, new_n52698_, new_n52221_ );
and  ( new_n52700_, new_n52699_, new_n52697_ );
or   ( new_n52701_, new_n52700_, new_n52696_ );
xnor ( new_n52702_, new_n52638_, new_n52636_ );
xor  ( new_n52703_, new_n52702_, new_n52644_ );
and  ( new_n52704_, new_n52703_, new_n52701_ );
xor  ( new_n52705_, new_n52703_, new_n52701_ );
xor  ( new_n52706_, new_n52235_, new_n52234_ );
and  ( new_n52707_, new_n52706_, new_n52705_ );
or   ( new_n52708_, new_n52707_, new_n52704_ );
xor  ( new_n52709_, new_n52648_, new_n52630_ );
nand ( new_n52710_, new_n52709_, new_n52708_ );
and  ( new_n52711_, new_n52710_, new_n52649_ );
xor  ( new_n52712_, new_n52711_, new_n52504_ );
nand ( new_n52713_, new_n52239_, new_n52238_ );
nand ( new_n52714_, new_n52240_, new_n52237_ );
and  ( new_n52715_, new_n52714_, new_n52713_ );
nor  ( new_n52716_, new_n52646_, new_n52635_ );
and  ( new_n52717_, new_n52647_, new_n52633_ );
or   ( new_n52718_, new_n52717_, new_n52716_ );
xor  ( new_n52719_, new_n51940_, new_n51898_ );
xor  ( new_n52720_, new_n52719_, new_n52718_ );
xor  ( new_n52721_, new_n52720_, new_n52715_ );
xor  ( new_n52722_, new_n52721_, new_n52712_ );
nand ( new_n52723_, new_n52500_, new_n52498_ );
nand ( new_n52724_, new_n52501_, new_n52494_ );
and  ( new_n52725_, new_n52724_, new_n52723_ );
xnor ( new_n52726_, new_n52007_, new_n52005_ );
xor  ( new_n52727_, new_n52025_, new_n52023_ );
xor  ( new_n52728_, new_n52727_, new_n52119_ );
xor  ( new_n52729_, new_n52728_, new_n52726_ );
xor  ( new_n52730_, new_n52729_, new_n52725_ );
or   ( new_n52731_, new_n52730_, new_n52722_ );
and  ( new_n52732_, new_n52730_, new_n52722_ );
xor  ( new_n52733_, new_n52628_, new_n52595_ );
not  ( new_n52734_, new_n52733_ );
xor  ( new_n52735_, new_n52358_, new_n52357_ );
xor  ( new_n52736_, new_n52588_, new_n52541_ );
nand ( new_n52737_, new_n52736_, new_n52735_ );
nor  ( new_n52738_, new_n52736_, new_n52735_ );
xor  ( new_n52739_, new_n51142_, new_n275_ );
or   ( new_n52740_, new_n52739_, new_n283_ );
or   ( new_n52741_, new_n52268_, new_n286_ );
and  ( new_n52742_, new_n52741_, new_n52740_ );
or   ( new_n52743_, new_n52264_, new_n320_ );
xor  ( new_n52744_, new_n50788_, new_n309_ );
or   ( new_n52745_, new_n52744_, new_n317_ );
and  ( new_n52746_, new_n52745_, new_n52743_ );
or   ( new_n52747_, new_n52746_, new_n52742_ );
and  ( new_n52748_, new_n52522_, new_n371_ );
xor  ( new_n52749_, new_n49488_, RIbb2f160_11 );
and  ( new_n52750_, new_n52749_, new_n373_ );
or   ( new_n52751_, new_n52750_, new_n52748_ );
xor  ( new_n52752_, new_n52746_, new_n52742_ );
nand ( new_n52753_, new_n52752_, new_n52751_ );
and  ( new_n52754_, new_n52753_, new_n52747_ );
or   ( new_n52755_, new_n52510_, new_n2124_ );
xor  ( new_n52756_, new_n46427_, new_n1840_ );
or   ( new_n52757_, new_n52756_, new_n2122_ );
and  ( new_n52758_, new_n52757_, new_n52755_ );
or   ( new_n52759_, new_n52308_, new_n1846_ );
xor  ( new_n52760_, new_n46789_, new_n1583_ );
or   ( new_n52761_, new_n52760_, new_n1844_ );
and  ( new_n52762_, new_n52761_, new_n52759_ );
or   ( new_n52763_, new_n52762_, new_n52758_ );
and  ( new_n52764_, new_n52762_, new_n52758_ );
xor  ( new_n52765_, new_n46958_, RIbb2ebc0_23 );
nand ( new_n52766_, new_n52765_, new_n1476_ );
or   ( new_n52767_, new_n52303_, new_n1595_ );
and  ( new_n52768_, new_n52767_, new_n52766_ );
or   ( new_n52769_, new_n52768_, new_n52764_ );
and  ( new_n52770_, new_n52769_, new_n52763_ );
nor  ( new_n52771_, new_n52770_, new_n52754_ );
or   ( new_n52772_, new_n52317_, new_n1366_ );
xor  ( new_n52773_, new_n47046_, new_n1126_ );
or   ( new_n52774_, new_n52773_, new_n1364_ );
and  ( new_n52775_, new_n52774_, new_n52772_ );
nand ( new_n52776_, new_n52327_, new_n820_ );
xor  ( new_n52777_, new_n48291_, RIbb2ee90_17 );
nand ( new_n52778_, new_n52777_, new_n822_ );
and  ( new_n52779_, new_n52778_, new_n52776_ );
nor  ( new_n52780_, new_n52779_, new_n52775_ );
and  ( new_n52781_, new_n52779_, new_n52775_ );
and  ( new_n52782_, new_n52322_, new_n1040_ );
xor  ( new_n52783_, new_n47640_, new_n893_ );
nor  ( new_n52784_, new_n52783_, new_n1135_ );
nor  ( new_n52785_, new_n52784_, new_n52782_ );
nor  ( new_n52786_, new_n52785_, new_n52781_ );
nor  ( new_n52787_, new_n52786_, new_n52780_ );
not  ( new_n52788_, new_n52787_ );
xor  ( new_n52789_, new_n52770_, new_n52754_ );
and  ( new_n52790_, new_n52789_, new_n52788_ );
or   ( new_n52791_, new_n52790_, new_n52771_ );
xnor ( new_n52792_, new_n52289_, new_n52277_ );
xor  ( new_n52793_, new_n52792_, new_n52313_ );
and  ( new_n52794_, new_n52793_, new_n52791_ );
nor  ( new_n52795_, new_n52793_, new_n52791_ );
not  ( new_n52796_, new_n52795_ );
xor  ( new_n52797_, new_n52355_, new_n52337_ );
and  ( new_n52798_, new_n52797_, new_n52796_ );
nor  ( new_n52799_, new_n52798_, new_n52794_ );
or   ( new_n52800_, new_n52799_, new_n52738_ );
and  ( new_n52801_, new_n52800_, new_n52737_ );
nor  ( new_n52802_, new_n52801_, new_n52734_ );
xor  ( new_n52803_, new_n52801_, new_n52734_ );
xor  ( new_n52804_, new_n52706_, new_n52705_ );
and  ( new_n52805_, new_n52804_, new_n52803_ );
nor  ( new_n52806_, new_n52805_, new_n52802_ );
not  ( new_n52807_, new_n52806_ );
xor  ( new_n52808_, new_n52709_, new_n52708_ );
and  ( new_n52809_, new_n52808_, new_n52807_ );
xor  ( new_n52810_, new_n52808_, new_n52807_ );
xor  ( new_n52811_, new_n52502_, new_n52493_ );
and  ( new_n52812_, new_n52811_, new_n52810_ );
nor  ( new_n52813_, new_n52812_, new_n52809_ );
or   ( new_n52814_, new_n52813_, new_n52732_ );
and  ( new_n52815_, new_n52814_, new_n52731_ );
xor  ( new_n52816_, new_n52011_, new_n52010_ );
not  ( new_n52817_, new_n52816_ );
nand ( new_n52818_, new_n52719_, new_n52718_ );
nor  ( new_n52819_, new_n52719_, new_n52718_ );
or   ( new_n52820_, new_n52819_, new_n52715_ );
and  ( new_n52821_, new_n52820_, new_n52818_ );
xor  ( new_n52822_, new_n52821_, new_n52817_ );
or   ( new_n52823_, new_n52728_, new_n52726_ );
and  ( new_n52824_, new_n52728_, new_n52726_ );
or   ( new_n52825_, new_n52824_, new_n52725_ );
nand ( new_n52826_, new_n52825_, new_n52823_ );
xnor ( new_n52827_, new_n52826_, new_n52822_ );
xor  ( new_n52828_, new_n52021_, new_n52019_ );
xor  ( new_n52829_, new_n52828_, new_n52122_ );
xor  ( new_n52830_, new_n52829_, new_n52827_ );
or   ( new_n52831_, new_n52711_, new_n52504_ );
and  ( new_n52832_, new_n52711_, new_n52504_ );
or   ( new_n52833_, new_n52721_, new_n52832_ );
and  ( new_n52834_, new_n52833_, new_n52831_ );
xor  ( new_n52835_, new_n52834_, new_n52830_ );
nor  ( new_n52836_, new_n52835_, new_n52815_ );
xnor ( new_n52837_, new_n52811_, new_n52810_ );
xor  ( new_n52838_, new_n52684_, new_n52682_ );
xor  ( new_n52839_, new_n52689_, new_n52687_ );
xor  ( new_n52840_, new_n52839_, new_n52693_ );
nand ( new_n52841_, new_n52840_, new_n52838_ );
xor  ( new_n52842_, new_n52666_, new_n52665_ );
xor  ( new_n52843_, new_n52752_, new_n52751_ );
nand ( new_n52844_, new_n52843_, new_n52842_ );
or   ( new_n52845_, new_n52477_, new_n526_ );
xor  ( new_n52846_, new_n49427_, new_n400_ );
or   ( new_n52847_, new_n52846_, new_n524_ );
and  ( new_n52848_, new_n52847_, new_n52845_ );
nor  ( new_n52849_, RIbb2d900_63, RIbb2d978_62 );
or   ( new_n52850_, new_n52849_, new_n9421_ );
xor  ( new_n52851_, new_n43793_, RIbb2d9f0_61 );
or   ( new_n52852_, new_n52851_, new_n10059_ );
and  ( new_n52853_, new_n52852_, new_n52850_ );
nor  ( new_n52854_, new_n52853_, new_n52848_ );
xor  ( new_n52855_, new_n48908_, new_n520_ );
nor  ( new_n52856_, new_n52855_, new_n755_ );
and  ( new_n52857_, new_n52471_, new_n660_ );
or   ( new_n52858_, new_n52857_, new_n52856_ );
xor  ( new_n52859_, new_n52853_, new_n52848_ );
and  ( new_n52860_, new_n52859_, new_n52858_ );
or   ( new_n52861_, new_n52860_, new_n52854_ );
xor  ( new_n52862_, new_n52843_, new_n52842_ );
nand ( new_n52863_, new_n52862_, new_n52861_ );
and  ( new_n52864_, new_n52863_, new_n52844_ );
xor  ( new_n52865_, new_n50894_, new_n309_ );
or   ( new_n52866_, new_n52865_, new_n317_ );
or   ( new_n52867_, new_n52744_, new_n320_ );
and  ( new_n52868_, new_n52867_, new_n52866_ );
or   ( new_n52869_, new_n52756_, new_n2124_ );
xor  ( new_n52870_, new_n46619_, new_n1840_ );
or   ( new_n52871_, new_n52870_, new_n2122_ );
and  ( new_n52872_, new_n52871_, new_n52869_ );
or   ( new_n52873_, new_n52872_, new_n52868_ );
xor  ( new_n52874_, new_n46962_, new_n1583_ );
nor  ( new_n52875_, new_n52874_, new_n1844_ );
nor  ( new_n52876_, new_n52760_, new_n1846_ );
or   ( new_n52877_, new_n52876_, new_n52875_ );
xor  ( new_n52878_, new_n52872_, new_n52868_ );
nand ( new_n52879_, new_n52878_, new_n52877_ );
and  ( new_n52880_, new_n52879_, new_n52873_ );
or   ( new_n52881_, new_n52783_, new_n1137_ );
xor  ( new_n52882_, new_n48039_, new_n893_ );
or   ( new_n52883_, new_n52882_, new_n1135_ );
and  ( new_n52884_, new_n52883_, new_n52881_ );
xor  ( new_n52885_, new_n47296_, RIbb2ecb0_21 );
nand ( new_n52886_, new_n52885_, new_n1253_ );
or   ( new_n52887_, new_n52773_, new_n1366_ );
and  ( new_n52888_, new_n52887_, new_n52886_ );
or   ( new_n52889_, new_n52888_, new_n52884_ );
and  ( new_n52890_, new_n52777_, new_n820_ );
xor  ( new_n52891_, new_n48518_, RIbb2ee90_17 );
and  ( new_n52892_, new_n52891_, new_n822_ );
nor  ( new_n52893_, new_n52892_, new_n52890_ );
and  ( new_n52894_, new_n52888_, new_n52884_ );
or   ( new_n52895_, new_n52894_, new_n52893_ );
and  ( new_n52896_, new_n52895_, new_n52889_ );
or   ( new_n52897_, new_n52896_, new_n52880_ );
and  ( new_n52898_, new_n52293_, new_n43879_ );
or   ( new_n52899_, new_n52294_, new_n43977_ );
or   ( new_n52900_, new_n52899_, new_n52898_ );
xor  ( new_n52901_, RIbb33210_189, new_n9679_ );
xor  ( new_n52902_, new_n52901_, new_n43528_ );
xor  ( new_n52903_, new_n52902_, new_n43945_ );
or   ( new_n52904_, new_n52903_, new_n43983_ );
and  ( new_n52905_, new_n52904_, new_n52900_ );
and  ( new_n52906_, new_n52905_, RIbb2d900_63 );
xor  ( new_n52907_, RIbb33288_190, new_n10220_ );
xor  ( new_n52908_, new_n52907_, new_n43526_ );
or   ( new_n52909_, new_n52908_, new_n43879_ );
or   ( new_n52910_, new_n52650_, new_n302_ );
or   ( new_n52911_, new_n52654_, new_n44007_ );
and  ( new_n52912_, new_n52911_, new_n52910_ );
or   ( new_n52913_, new_n52912_, new_n52909_ );
xor  ( new_n52914_, new_n51446_, RIbb2f430_5 );
and  ( new_n52915_, new_n52914_, new_n280_ );
xor  ( new_n52916_, new_n51477_, RIbb2f430_5 );
and  ( new_n52917_, new_n52916_, new_n282_ );
or   ( new_n52918_, new_n52917_, new_n52915_ );
xor  ( new_n52919_, new_n52912_, new_n52909_ );
nand ( new_n52920_, new_n52919_, new_n52918_ );
and  ( new_n52921_, new_n52920_, new_n52913_ );
nor  ( new_n52922_, new_n52921_, new_n52906_ );
xor  ( new_n52923_, new_n47303_, new_n1355_ );
nor  ( new_n52924_, new_n52923_, new_n1593_ );
and  ( new_n52925_, new_n52765_, new_n1474_ );
nor  ( new_n52926_, new_n52925_, new_n52924_ );
and  ( new_n52927_, new_n52921_, new_n52906_ );
nor  ( new_n52928_, new_n52927_, new_n52926_ );
nor  ( new_n52929_, new_n52928_, new_n52922_ );
and  ( new_n52930_, new_n52896_, new_n52880_ );
or   ( new_n52931_, new_n52930_, new_n52929_ );
and  ( new_n52932_, new_n52931_, new_n52897_ );
nor  ( new_n52933_, new_n52932_, new_n52864_ );
xor  ( new_n52934_, new_n43937_, RIbb2ddb0_53 );
nand ( new_n52935_, new_n52934_, new_n7489_ );
or   ( new_n52936_, new_n52419_, new_n7734_ );
and  ( new_n52937_, new_n52936_, new_n52935_ );
nand ( new_n52938_, new_n52425_, new_n4958_ );
xor  ( new_n52939_, new_n44506_, new_n4705_ );
or   ( new_n52940_, new_n52939_, new_n5207_ );
and  ( new_n52941_, new_n52940_, new_n52938_ );
or   ( new_n52942_, new_n52941_, new_n52937_ );
xor  ( new_n52943_, new_n44681_, RIbb2e350_41 );
and  ( new_n52944_, new_n52943_, new_n4543_ );
and  ( new_n52945_, new_n52414_, new_n4541_ );
or   ( new_n52946_, new_n52945_, new_n52944_ );
xor  ( new_n52947_, new_n52941_, new_n52937_ );
nand ( new_n52948_, new_n52947_, new_n52946_ );
and  ( new_n52949_, new_n52948_, new_n52942_ );
xor  ( new_n52950_, new_n44183_, new_n5594_ );
or   ( new_n52951_, new_n52950_, new_n6173_ );
or   ( new_n52952_, new_n52397_, new_n6175_ );
and  ( new_n52953_, new_n52952_, new_n52951_ );
nand ( new_n52954_, new_n52403_, new_n2613_ );
xor  ( new_n52955_, new_n45928_, new_n2421_ );
or   ( new_n52956_, new_n52955_, new_n2807_ );
and  ( new_n52957_, new_n52956_, new_n52954_ );
or   ( new_n52958_, new_n52957_, new_n52953_ );
nor  ( new_n52959_, new_n52394_, new_n2427_ );
xor  ( new_n52960_, new_n46137_, RIbb2e8f0_29 );
and  ( new_n52961_, new_n52960_, new_n2244_ );
nor  ( new_n52962_, new_n52961_, new_n52959_ );
and  ( new_n52963_, new_n52957_, new_n52953_ );
or   ( new_n52964_, new_n52963_, new_n52962_ );
and  ( new_n52965_, new_n52964_, new_n52958_ );
nor  ( new_n52966_, new_n52965_, new_n52949_ );
nand ( new_n52967_, new_n52965_, new_n52949_ );
or   ( new_n52968_, new_n52379_, new_n9424_ );
xor  ( new_n52969_, new_n43898_, new_n8870_ );
or   ( new_n52970_, new_n52969_, new_n9422_ );
and  ( new_n52971_, new_n52970_, new_n52968_ );
xor  ( new_n52972_, new_n43884_, new_n7722_ );
or   ( new_n52973_, new_n52972_, new_n8264_ );
or   ( new_n52974_, new_n52374_, new_n8266_ );
and  ( new_n52975_, new_n52974_, new_n52973_ );
nor  ( new_n52976_, new_n52975_, new_n52971_ );
xor  ( new_n52977_, new_n44319_, RIbb2e170_45 );
and  ( new_n52978_, new_n52977_, new_n5373_ );
and  ( new_n52979_, new_n52386_, new_n5371_ );
or   ( new_n52980_, new_n52979_, new_n52978_ );
xor  ( new_n52981_, new_n52975_, new_n52971_ );
and  ( new_n52982_, new_n52981_, new_n52980_ );
or   ( new_n52983_, new_n52982_, new_n52976_ );
and  ( new_n52984_, new_n52983_, new_n52967_ );
or   ( new_n52985_, new_n52984_, new_n52966_ );
xor  ( new_n52986_, new_n52932_, new_n52864_ );
and  ( new_n52987_, new_n52986_, new_n52985_ );
nor  ( new_n52988_, new_n52987_, new_n52933_ );
not  ( new_n52989_, new_n52988_ );
xor  ( new_n52990_, new_n52840_, new_n52838_ );
nand ( new_n52991_, new_n52990_, new_n52989_ );
and  ( new_n52992_, new_n52991_, new_n52841_ );
xnor ( new_n52993_, new_n52695_, new_n52686_ );
xor  ( new_n52994_, new_n52993_, new_n52699_ );
nor  ( new_n52995_, new_n52994_, new_n52992_ );
xor  ( new_n52996_, new_n52994_, new_n52992_ );
xor  ( new_n52997_, new_n52487_, new_n52373_ );
and  ( new_n52998_, new_n52997_, new_n52996_ );
or   ( new_n52999_, new_n52998_, new_n52995_ );
xor  ( new_n53000_, new_n52532_, new_n52531_ );
xor  ( new_n53001_, new_n52569_, new_n52568_ );
and  ( new_n53002_, new_n53001_, new_n53000_ );
xor  ( new_n53003_, new_n53001_, new_n53000_ );
xnor ( new_n53004_, new_n52512_, new_n52508_ );
xor  ( new_n53005_, new_n53004_, new_n52516_ );
and  ( new_n53006_, new_n53005_, new_n53003_ );
nor  ( new_n53007_, new_n53006_, new_n53002_ );
xnor ( new_n53008_, new_n52311_, new_n52310_ );
or   ( new_n53009_, new_n52557_, new_n3463_ );
xor  ( new_n53010_, new_n45204_, new_n3113_ );
or   ( new_n53011_, new_n53010_, new_n3461_ );
and  ( new_n53012_, new_n53011_, new_n53009_ );
xor  ( new_n53013_, new_n44974_, new_n3457_ );
or   ( new_n53014_, new_n53013_, new_n3896_ );
or   ( new_n53015_, new_n52546_, new_n3898_ );
and  ( new_n53016_, new_n53015_, new_n53014_ );
or   ( new_n53017_, new_n53016_, new_n53012_ );
nor  ( new_n53018_, new_n52560_, new_n6647_ );
xor  ( new_n53019_, new_n43985_, RIbb2df90_49 );
and  ( new_n53020_, new_n53019_, new_n6510_ );
nor  ( new_n53021_, new_n53020_, new_n53018_ );
and  ( new_n53022_, new_n53016_, new_n53012_ );
or   ( new_n53023_, new_n53022_, new_n53021_ );
and  ( new_n53024_, new_n53023_, new_n53017_ );
nand ( new_n53025_, new_n53024_, new_n53008_ );
xor  ( new_n53026_, new_n52677_, new_n52676_ );
nor  ( new_n53027_, new_n53024_, new_n53008_ );
or   ( new_n53028_, new_n53027_, new_n53026_ );
nand ( new_n53029_, new_n53028_, new_n53025_ );
nor  ( new_n53030_, new_n53029_, new_n53007_ );
xnor ( new_n53031_, new_n53029_, new_n53007_ );
xnor ( new_n53032_, new_n52621_, new_n52619_ );
xor  ( new_n53033_, new_n53032_, new_n52624_ );
nor  ( new_n53034_, new_n53033_, new_n53031_ );
or   ( new_n53035_, new_n53034_, new_n53030_ );
xor  ( new_n53036_, new_n52615_, new_n52596_ );
xor  ( new_n53037_, new_n53036_, new_n52626_ );
or   ( new_n53038_, new_n53037_, new_n53035_ );
nand ( new_n53039_, new_n53037_, new_n53035_ );
or   ( new_n53040_, new_n52902_, new_n43879_ );
xor  ( new_n53041_, new_n52293_, new_n43945_ );
or   ( new_n53042_, new_n53041_, new_n43983_ );
nor  ( new_n53043_, new_n52280_, new_n43880_ );
or   ( new_n53044_, new_n52281_, new_n43977_ );
or   ( new_n53045_, new_n53044_, new_n53043_ );
and  ( new_n53046_, new_n53045_, new_n53042_ );
or   ( new_n53047_, new_n53046_, new_n53040_ );
xor  ( new_n53048_, new_n53046_, new_n53040_ );
nand ( new_n53049_, new_n53048_, new_n52653_ );
and  ( new_n53050_, new_n53049_, new_n53047_ );
nand ( new_n53051_, new_n52749_, new_n371_ );
xor  ( new_n53052_, new_n49758_, new_n325_ );
or   ( new_n53053_, new_n53052_, new_n409_ );
and  ( new_n53054_, new_n53053_, new_n53051_ );
or   ( new_n53055_, new_n52739_, new_n286_ );
nand ( new_n53056_, new_n52914_, new_n282_ );
and  ( new_n53057_, new_n53056_, new_n53055_ );
nor  ( new_n53058_, new_n53057_, new_n53054_ );
nor  ( new_n53059_, new_n52663_, new_n340_ );
xor  ( new_n53060_, new_n50487_, new_n329_ );
nor  ( new_n53061_, new_n53060_, new_n337_ );
nor  ( new_n53062_, new_n53061_, new_n53059_ );
and  ( new_n53063_, new_n53057_, new_n53054_ );
nor  ( new_n53064_, new_n53063_, new_n53062_ );
nor  ( new_n53065_, new_n53064_, new_n53058_ );
nor  ( new_n53066_, new_n53065_, new_n53050_ );
xor  ( new_n53067_, new_n45584_, RIbb2e710_33 );
and  ( new_n53068_, new_n53067_, new_n2930_ );
nor  ( new_n53069_, new_n52566_, new_n3119_ );
nor  ( new_n53070_, new_n53069_, new_n53068_ );
not  ( new_n53071_, new_n53070_ );
xor  ( new_n53072_, new_n53065_, new_n53050_ );
and  ( new_n53073_, new_n53072_, new_n53071_ );
nor  ( new_n53074_, new_n53073_, new_n53066_ );
not  ( new_n53075_, new_n53074_ );
xnor ( new_n53076_, new_n52548_, new_n52544_ );
nand ( new_n53077_, new_n53076_, new_n52552_ );
not  ( new_n53078_, new_n52554_ );
or   ( new_n53079_, new_n53078_, new_n52549_ );
and  ( new_n53080_, new_n53079_, new_n53077_ );
and  ( new_n53081_, new_n53080_, new_n53075_ );
xor  ( new_n53082_, new_n53080_, new_n53075_ );
xnor ( new_n53083_, new_n52579_, new_n52576_ );
xor  ( new_n53084_, new_n53083_, new_n52583_ );
and  ( new_n53085_, new_n53084_, new_n53082_ );
or   ( new_n53086_, new_n53085_, new_n53081_ );
xnor ( new_n53087_, new_n52571_, new_n52555_ );
nand ( new_n53088_, new_n53087_, new_n52586_ );
not  ( new_n53089_, new_n52587_ );
or   ( new_n53090_, new_n53089_, new_n52572_ );
and  ( new_n53091_, new_n53090_, new_n53088_ );
and  ( new_n53092_, new_n53091_, new_n53086_ );
nor  ( new_n53093_, new_n53091_, new_n53086_ );
not  ( new_n53094_, new_n53093_ );
xor  ( new_n53095_, new_n52536_, new_n52535_ );
and  ( new_n53096_, new_n53095_, new_n53094_ );
nor  ( new_n53097_, new_n53096_, new_n53092_ );
nand ( new_n53098_, new_n53097_, new_n53039_ );
and  ( new_n53099_, new_n53098_, new_n53038_ );
nand ( new_n53100_, new_n53099_, new_n52999_ );
nor  ( new_n53101_, new_n53099_, new_n52999_ );
xor  ( new_n53102_, new_n52366_, new_n52261_ );
xor  ( new_n53103_, new_n53102_, new_n52489_ );
or   ( new_n53104_, new_n53103_, new_n53101_ );
and  ( new_n53105_, new_n53104_, new_n53100_ );
nor  ( new_n53106_, new_n53105_, new_n52837_ );
nand ( new_n53107_, new_n53105_, new_n52837_ );
xnor ( new_n53108_, new_n52804_, new_n52803_ );
xor  ( new_n53109_, new_n52997_, new_n52996_ );
xnor ( new_n53110_, new_n52462_, new_n52433_ );
xor  ( new_n53111_, new_n53110_, new_n52485_ );
xor  ( new_n53112_, new_n53091_, new_n53086_ );
xor  ( new_n53113_, new_n53112_, new_n53095_ );
or   ( new_n53114_, new_n53113_, new_n53111_ );
and  ( new_n53115_, new_n53113_, new_n53111_ );
xor  ( new_n53116_, new_n53033_, new_n53031_ );
or   ( new_n53117_, new_n53116_, new_n53115_ );
and  ( new_n53118_, new_n53117_, new_n53114_ );
nand ( new_n53119_, new_n53118_, new_n53109_ );
nor  ( new_n53120_, new_n53118_, new_n53109_ );
xor  ( new_n53121_, new_n53084_, new_n53082_ );
xor  ( new_n53122_, new_n53005_, new_n53003_ );
nand ( new_n53123_, new_n53122_, new_n53121_ );
xor  ( new_n53124_, new_n53122_, new_n53121_ );
xor  ( new_n53125_, new_n52986_, new_n52985_ );
nand ( new_n53126_, new_n53125_, new_n53124_ );
and  ( new_n53127_, new_n53126_, new_n53123_ );
xor  ( new_n53128_, new_n52450_, new_n52449_ );
xnor ( new_n53129_, new_n52401_, new_n52396_ );
xor  ( new_n53130_, new_n53129_, new_n52407_ );
nor  ( new_n53131_, new_n53130_, new_n53128_ );
and  ( new_n53132_, new_n53130_, new_n53128_ );
xor  ( new_n53133_, new_n53072_, new_n53071_ );
nor  ( new_n53134_, new_n53133_, new_n53132_ );
or   ( new_n53135_, new_n53134_, new_n53131_ );
xnor ( new_n53136_, new_n53024_, new_n53008_ );
xor  ( new_n53137_, new_n53136_, new_n53026_ );
or   ( new_n53138_, new_n53137_, new_n53135_ );
and  ( new_n53139_, new_n53137_, new_n53135_ );
nor  ( new_n53140_, new_n53052_, new_n411_ );
xor  ( new_n53141_, new_n50115_, new_n325_ );
nor  ( new_n53142_, new_n53141_, new_n409_ );
nor  ( new_n53143_, new_n53142_, new_n53140_ );
or   ( new_n53144_, new_n52865_, new_n320_ );
xor  ( new_n53145_, new_n51142_, new_n309_ );
or   ( new_n53146_, new_n53145_, new_n317_ );
and  ( new_n53147_, new_n53146_, new_n53144_ );
nor  ( new_n53148_, new_n53147_, new_n53143_ );
xor  ( new_n53149_, new_n53048_, new_n52653_ );
and  ( new_n53150_, new_n53149_, new_n53148_ );
and  ( new_n53151_, new_n53067_, new_n2928_ );
xor  ( new_n53152_, new_n45738_, RIbb2e710_33 );
and  ( new_n53153_, new_n53152_, new_n2930_ );
nor  ( new_n53154_, new_n53153_, new_n53151_ );
not  ( new_n53155_, new_n53154_ );
xor  ( new_n53156_, new_n53149_, new_n53148_ );
and  ( new_n53157_, new_n53156_, new_n53155_ );
or   ( new_n53158_, new_n53157_, new_n53150_ );
xnor ( new_n53159_, new_n52382_, new_n52378_ );
nand ( new_n53160_, new_n53159_, new_n52388_ );
not  ( new_n53161_, new_n52390_ );
or   ( new_n53162_, new_n53161_, new_n52383_ );
and  ( new_n53163_, new_n53162_, new_n53160_ );
nand ( new_n53164_, new_n53163_, new_n53158_ );
xor  ( new_n53165_, new_n53163_, new_n53158_ );
xnor ( new_n53166_, new_n52421_, new_n52416_ );
nand ( new_n53167_, new_n53166_, new_n52427_ );
not  ( new_n53168_, new_n52429_ );
or   ( new_n53169_, new_n53168_, new_n52422_ );
and  ( new_n53170_, new_n53169_, new_n53167_ );
nand ( new_n53171_, new_n53170_, new_n53165_ );
and  ( new_n53172_, new_n53171_, new_n53164_ );
or   ( new_n53173_, new_n53172_, new_n53139_ );
and  ( new_n53174_, new_n53173_, new_n53138_ );
nor  ( new_n53175_, new_n53174_, new_n53127_ );
xor  ( new_n53176_, new_n52990_, new_n52989_ );
xor  ( new_n53177_, new_n53174_, new_n53127_ );
and  ( new_n53178_, new_n53177_, new_n53176_ );
nor  ( new_n53179_, new_n53178_, new_n53175_ );
or   ( new_n53180_, new_n53179_, new_n53120_ );
and  ( new_n53181_, new_n53180_, new_n53119_ );
nor  ( new_n53182_, new_n53181_, new_n53108_ );
nand ( new_n53183_, new_n53181_, new_n53108_ );
xor  ( new_n53184_, new_n52789_, new_n52788_ );
xor  ( new_n53185_, new_n52467_, new_n52465_ );
xnor ( new_n53186_, new_n53185_, new_n52483_ );
and  ( new_n53187_, new_n53186_, new_n53184_ );
xnor ( new_n53188_, new_n53186_, new_n53184_ );
xor  ( new_n53189_, new_n52779_, new_n52775_ );
xor  ( new_n53190_, new_n53189_, new_n52785_ );
or   ( new_n53191_, new_n53010_, new_n3463_ );
xor  ( new_n53192_, new_n45403_, new_n3113_ );
or   ( new_n53193_, new_n53192_, new_n3461_ );
and  ( new_n53194_, new_n53193_, new_n53191_ );
or   ( new_n53195_, new_n53013_, new_n3898_ );
xor  ( new_n53196_, new_n45119_, new_n3457_ );
or   ( new_n53197_, new_n53196_, new_n3896_ );
and  ( new_n53198_, new_n53197_, new_n53195_ );
or   ( new_n53199_, new_n53198_, new_n53194_ );
xor  ( new_n53200_, new_n43812_, RIbb2df90_49 );
and  ( new_n53201_, new_n53200_, new_n6510_ );
and  ( new_n53202_, new_n53019_, new_n6508_ );
nor  ( new_n53203_, new_n53202_, new_n53201_ );
and  ( new_n53204_, new_n53198_, new_n53194_ );
or   ( new_n53205_, new_n53204_, new_n53203_ );
and  ( new_n53206_, new_n53205_, new_n53199_ );
or   ( new_n53207_, new_n53206_, new_n53190_ );
nand ( new_n53208_, new_n53206_, new_n53190_ );
xor  ( new_n53209_, new_n52481_, new_n52480_ );
nand ( new_n53210_, new_n53209_, new_n53208_ );
and  ( new_n53211_, new_n53210_, new_n53207_ );
nor  ( new_n53212_, new_n53211_, new_n53188_ );
or   ( new_n53213_, new_n53212_, new_n53187_ );
xor  ( new_n53214_, new_n52793_, new_n52791_ );
xor  ( new_n53215_, new_n53214_, new_n52797_ );
and  ( new_n53216_, new_n53215_, new_n53213_ );
or   ( new_n53217_, new_n53215_, new_n53213_ );
xnor ( new_n53218_, new_n52431_, new_n52430_ );
xor  ( new_n53219_, new_n52762_, new_n52758_ );
xor  ( new_n53220_, new_n53219_, new_n52768_ );
or   ( new_n53221_, new_n52439_, new_n7186_ );
xor  ( new_n53222_, new_n43952_, new_n6635_ );
or   ( new_n53223_, new_n53222_, new_n7184_ );
and  ( new_n53224_, new_n53223_, new_n53221_ );
or   ( new_n53225_, new_n52434_, new_n8876_ );
xor  ( new_n53226_, new_n43799_, new_n8254_ );
or   ( new_n53227_, new_n53226_, new_n8874_ );
and  ( new_n53228_, new_n53227_, new_n53225_ );
or   ( new_n53229_, new_n53228_, new_n53224_ );
and  ( new_n53230_, new_n52447_, new_n4032_ );
xor  ( new_n53231_, new_n44877_, RIbb2e440_39 );
and  ( new_n53232_, new_n53231_, new_n4034_ );
nor  ( new_n53233_, new_n53232_, new_n53230_ );
and  ( new_n53234_, new_n53228_, new_n53224_ );
or   ( new_n53235_, new_n53234_, new_n53233_ );
and  ( new_n53236_, new_n53235_, new_n53229_ );
or   ( new_n53237_, new_n53236_, new_n53220_ );
nand ( new_n53238_, new_n53236_, new_n53220_ );
xor  ( new_n53239_, new_n53016_, new_n53012_ );
xnor ( new_n53240_, new_n53239_, new_n53021_ );
nand ( new_n53241_, new_n53240_, new_n53238_ );
and  ( new_n53242_, new_n53241_, new_n53237_ );
nor  ( new_n53243_, new_n53242_, new_n53218_ );
nand ( new_n53244_, new_n53242_, new_n53218_ );
xor  ( new_n53245_, new_n52453_, new_n52452_ );
xor  ( new_n53246_, new_n53245_, new_n52460_ );
and  ( new_n53247_, new_n53246_, new_n53244_ );
or   ( new_n53248_, new_n53247_, new_n53243_ );
and  ( new_n53249_, new_n53248_, new_n53217_ );
or   ( new_n53250_, new_n53249_, new_n53216_ );
xnor ( new_n53251_, new_n52736_, new_n52735_ );
xor  ( new_n53252_, new_n53251_, new_n52799_ );
or   ( new_n53253_, new_n53252_, new_n53250_ );
xor  ( new_n53254_, new_n53252_, new_n53250_ );
xor  ( new_n53255_, new_n53037_, new_n53035_ );
xor  ( new_n53256_, new_n53255_, new_n53097_ );
nand ( new_n53257_, new_n53256_, new_n53254_ );
and  ( new_n53258_, new_n53257_, new_n53253_ );
and  ( new_n53259_, new_n53258_, new_n53183_ );
or   ( new_n53260_, new_n53259_, new_n53182_ );
and  ( new_n53261_, new_n53260_, new_n53107_ );
or   ( new_n53262_, new_n53261_, new_n53106_ );
xnor ( new_n53263_, new_n52730_, new_n52722_ );
xor  ( new_n53264_, new_n53263_, new_n52813_ );
and  ( new_n53265_, new_n53264_, new_n53262_ );
nor  ( new_n53266_, new_n53264_, new_n53262_ );
not  ( new_n53267_, new_n53266_ );
xor  ( new_n53268_, new_n53099_, new_n52999_ );
xor  ( new_n53269_, new_n53268_, new_n53103_ );
xnor ( new_n53270_, new_n52921_, new_n52906_ );
xor  ( new_n53271_, new_n53270_, new_n52926_ );
xor  ( new_n53272_, new_n52859_, new_n52858_ );
and  ( new_n53273_, new_n53272_, new_n53271_ );
xnor ( new_n53274_, new_n52888_, new_n52884_ );
xor  ( new_n53275_, new_n53274_, new_n52893_ );
xor  ( new_n53276_, new_n53272_, new_n53271_ );
and  ( new_n53277_, new_n53276_, new_n53275_ );
nor  ( new_n53278_, new_n53277_, new_n53273_ );
not  ( new_n53279_, new_n53278_ );
xor  ( new_n53280_, new_n52862_, new_n52861_ );
and  ( new_n53281_, new_n53280_, new_n53279_ );
xor  ( new_n53282_, new_n53280_, new_n53279_ );
xnor ( new_n53283_, new_n52896_, new_n52880_ );
xor  ( new_n53284_, new_n53283_, new_n52929_ );
and  ( new_n53285_, new_n53284_, new_n53282_ );
or   ( new_n53286_, new_n53285_, new_n53281_ );
xor  ( new_n53287_, new_n53211_, new_n53188_ );
and  ( new_n53288_, new_n53287_, new_n53286_ );
or   ( new_n53289_, new_n53060_, new_n340_ );
xor  ( new_n53290_, new_n50788_, new_n329_ );
or   ( new_n53291_, new_n53290_, new_n337_ );
and  ( new_n53292_, new_n53291_, new_n53289_ );
or   ( new_n53293_, new_n52846_, new_n526_ );
xor  ( new_n53294_, new_n49488_, new_n400_ );
or   ( new_n53295_, new_n53294_, new_n524_ );
and  ( new_n53296_, new_n53295_, new_n53293_ );
or   ( new_n53297_, new_n53296_, new_n53292_ );
xor  ( new_n53298_, new_n46789_, new_n1840_ );
nor  ( new_n53299_, new_n53298_, new_n2122_ );
nor  ( new_n53300_, new_n52870_, new_n2124_ );
or   ( new_n53301_, new_n53300_, new_n53299_ );
xor  ( new_n53302_, new_n53296_, new_n53292_ );
nand ( new_n53303_, new_n53302_, new_n53301_ );
and  ( new_n53304_, new_n53303_, new_n53297_ );
xor  ( new_n53305_, RIbb33300_191, new_n10541_ );
xor  ( new_n53306_, new_n53305_, new_n43019_ );
or   ( new_n53307_, new_n53306_, new_n43879_ );
xor  ( new_n53308_, new_n52908_, new_n43945_ );
or   ( new_n53309_, new_n53308_, new_n43983_ );
xor  ( new_n53310_, new_n52902_, new_n43880_ );
or   ( new_n53311_, new_n53310_, new_n43977_ );
and  ( new_n53312_, new_n53311_, new_n53309_ );
or   ( new_n53313_, new_n53312_, new_n53307_ );
and  ( new_n53314_, new_n52655_, new_n295_ );
and  ( new_n53315_, new_n53041_, new_n43949_ );
or   ( new_n53316_, new_n53315_, new_n53314_ );
xor  ( new_n53317_, new_n53312_, new_n53307_ );
nand ( new_n53318_, new_n53317_, new_n53316_ );
and  ( new_n53319_, new_n53318_, new_n53313_ );
xor  ( new_n53320_, new_n52905_, RIbb2d900_63 );
or   ( new_n53321_, new_n53320_, new_n53319_ );
and  ( new_n53322_, new_n52960_, new_n2242_ );
xor  ( new_n53323_, new_n46427_, RIbb2e8f0_29 );
and  ( new_n53324_, new_n53323_, new_n2244_ );
or   ( new_n53325_, new_n53324_, new_n53322_ );
xor  ( new_n53326_, new_n53320_, new_n53319_ );
nand ( new_n53327_, new_n53326_, new_n53325_ );
and  ( new_n53328_, new_n53327_, new_n53321_ );
or   ( new_n53329_, new_n53328_, new_n53304_ );
or   ( new_n53330_, new_n52923_, new_n1595_ );
xor  ( new_n53331_, new_n47046_, new_n1355_ );
or   ( new_n53332_, new_n53331_, new_n1593_ );
and  ( new_n53333_, new_n53332_, new_n53330_ );
or   ( new_n53334_, new_n52874_, new_n1846_ );
xor  ( new_n53335_, new_n46958_, RIbb2ead0_25 );
nand ( new_n53336_, new_n53335_, new_n1741_ );
and  ( new_n53337_, new_n53336_, new_n53334_ );
nor  ( new_n53338_, new_n53337_, new_n53333_ );
and  ( new_n53339_, new_n52885_, new_n1251_ );
xor  ( new_n53340_, new_n47640_, new_n1126_ );
nor  ( new_n53341_, new_n53340_, new_n1364_ );
nor  ( new_n53342_, new_n53341_, new_n53339_ );
and  ( new_n53343_, new_n53337_, new_n53333_ );
nor  ( new_n53344_, new_n53343_, new_n53342_ );
nor  ( new_n53345_, new_n53344_, new_n53338_ );
not  ( new_n53346_, new_n53345_ );
xor  ( new_n53347_, new_n53328_, new_n53304_ );
nand ( new_n53348_, new_n53347_, new_n53346_ );
and  ( new_n53349_, new_n53348_, new_n53329_ );
xor  ( new_n53350_, new_n48291_, RIbb2eda0_19 );
nand ( new_n53351_, new_n53350_, new_n1042_ );
or   ( new_n53352_, new_n52882_, new_n1137_ );
and  ( new_n53353_, new_n53352_, new_n53351_ );
xor  ( new_n53354_, new_n48756_, RIbb2ee90_17 );
nand ( new_n53355_, new_n53354_, new_n822_ );
nand ( new_n53356_, new_n52891_, new_n820_ );
and  ( new_n53357_, new_n53356_, new_n53355_ );
nor  ( new_n53358_, new_n53357_, new_n53353_ );
xor  ( new_n53359_, new_n49265_, new_n520_ );
nor  ( new_n53360_, new_n53359_, new_n755_ );
nor  ( new_n53361_, new_n52855_, new_n757_ );
nor  ( new_n53362_, new_n53361_, new_n53360_ );
and  ( new_n53363_, new_n53357_, new_n53353_ );
nor  ( new_n53364_, new_n53363_, new_n53362_ );
nor  ( new_n53365_, new_n53364_, new_n53358_ );
xnor ( new_n53366_, new_n53057_, new_n53054_ );
nand ( new_n53367_, new_n53366_, new_n53062_ );
not  ( new_n53368_, new_n53064_ );
or   ( new_n53369_, new_n53368_, new_n53058_ );
nand ( new_n53370_, new_n53369_, new_n53367_ );
or   ( new_n53371_, new_n53370_, new_n53365_ );
xnor ( new_n53372_, new_n53370_, new_n53365_ );
xor  ( new_n53373_, new_n46037_, new_n2421_ );
or   ( new_n53374_, new_n53373_, new_n2807_ );
or   ( new_n53375_, new_n52955_, new_n2809_ );
and  ( new_n53376_, new_n53375_, new_n53374_ );
xor  ( new_n53377_, new_n43914_, RIbb2df90_49 );
nand ( new_n53378_, new_n53377_, new_n6510_ );
nand ( new_n53379_, new_n53200_, new_n6508_ );
and  ( new_n53380_, new_n53379_, new_n53378_ );
nor  ( new_n53381_, new_n53380_, new_n53376_ );
xor  ( new_n53382_, new_n45597_, RIbb2e710_33 );
and  ( new_n53383_, new_n53382_, new_n2930_ );
and  ( new_n53384_, new_n53152_, new_n2928_ );
nor  ( new_n53385_, new_n53384_, new_n53383_ );
and  ( new_n53386_, new_n53380_, new_n53376_ );
nor  ( new_n53387_, new_n53386_, new_n53385_ );
nor  ( new_n53388_, new_n53387_, new_n53381_ );
or   ( new_n53389_, new_n53388_, new_n53372_ );
and  ( new_n53390_, new_n53389_, new_n53371_ );
nor  ( new_n53391_, new_n53390_, new_n53349_ );
xor  ( new_n53392_, new_n43985_, new_n6635_ );
or   ( new_n53393_, new_n53392_, new_n7184_ );
or   ( new_n53394_, new_n53222_, new_n7186_ );
and  ( new_n53395_, new_n53394_, new_n53393_ );
nand ( new_n53396_, new_n53231_, new_n4032_ );
xor  ( new_n53397_, new_n44974_, new_n3892_ );
or   ( new_n53398_, new_n53397_, new_n4302_ );
and  ( new_n53399_, new_n53398_, new_n53396_ );
or   ( new_n53400_, new_n53399_, new_n53395_ );
xor  ( new_n53401_, new_n45204_, RIbb2e530_37 );
and  ( new_n53402_, new_n53401_, new_n3733_ );
nor  ( new_n53403_, new_n53196_, new_n3898_ );
or   ( new_n53404_, new_n53403_, new_n53402_ );
xor  ( new_n53405_, new_n53399_, new_n53395_ );
nand ( new_n53406_, new_n53405_, new_n53404_ );
and  ( new_n53407_, new_n53406_, new_n53400_ );
xor  ( new_n53408_, new_n44785_, RIbb2e350_41 );
nand ( new_n53409_, new_n53408_, new_n4543_ );
nand ( new_n53410_, new_n52943_, new_n4541_ );
and  ( new_n53411_, new_n53410_, new_n53409_ );
xor  ( new_n53412_, new_n43894_, new_n8870_ );
or   ( new_n53413_, new_n53412_, new_n9422_ );
or   ( new_n53414_, new_n52969_, new_n9424_ );
and  ( new_n53415_, new_n53414_, new_n53413_ );
or   ( new_n53416_, new_n53415_, new_n53411_ );
xor  ( new_n53417_, new_n43956_, new_n7174_ );
nor  ( new_n53418_, new_n53417_, new_n7732_ );
and  ( new_n53419_, new_n52934_, new_n7487_ );
nor  ( new_n53420_, new_n53419_, new_n53418_ );
and  ( new_n53421_, new_n53415_, new_n53411_ );
or   ( new_n53422_, new_n53421_, new_n53420_ );
and  ( new_n53423_, new_n53422_, new_n53416_ );
nor  ( new_n53424_, new_n53423_, new_n53407_ );
xor  ( new_n53425_, new_n43787_, RIbb2d9f0_61 );
nand ( new_n53426_, new_n53425_, new_n9740_ );
or   ( new_n53427_, new_n52851_, new_n10061_ );
and  ( new_n53428_, new_n53427_, new_n53426_ );
or   ( new_n53429_, new_n52950_, new_n6175_ );
xor  ( new_n53430_, new_n44218_, new_n5594_ );
or   ( new_n53431_, new_n53430_, new_n6173_ );
and  ( new_n53432_, new_n53431_, new_n53429_ );
nor  ( new_n53433_, new_n53432_, new_n53428_ );
xor  ( new_n53434_, new_n43803_, RIbb2dbd0_57 );
and  ( new_n53435_, new_n53434_, new_n8651_ );
nor  ( new_n53436_, new_n53226_, new_n8876_ );
or   ( new_n53437_, new_n53436_, new_n53435_ );
xor  ( new_n53438_, new_n53432_, new_n53428_ );
and  ( new_n53439_, new_n53438_, new_n53437_ );
or   ( new_n53440_, new_n53439_, new_n53433_ );
xor  ( new_n53441_, new_n53423_, new_n53407_ );
and  ( new_n53442_, new_n53441_, new_n53440_ );
or   ( new_n53443_, new_n53442_, new_n53424_ );
xor  ( new_n53444_, new_n53390_, new_n53349_ );
and  ( new_n53445_, new_n53444_, new_n53443_ );
or   ( new_n53446_, new_n53445_, new_n53391_ );
xor  ( new_n53447_, new_n53287_, new_n53286_ );
and  ( new_n53448_, new_n53447_, new_n53446_ );
or   ( new_n53449_, new_n53448_, new_n53288_ );
xor  ( new_n53450_, new_n53215_, new_n53213_ );
xor  ( new_n53451_, new_n53450_, new_n53248_ );
nand ( new_n53452_, new_n53451_, new_n53449_ );
xor  ( new_n53453_, new_n51758_, new_n275_ );
or   ( new_n53454_, new_n53453_, new_n283_ );
nand ( new_n53455_, new_n52916_, new_n280_ );
and  ( new_n53456_, new_n53455_, new_n53454_ );
or   ( new_n53457_, new_n53294_, new_n526_ );
xor  ( new_n53458_, new_n49758_, new_n400_ );
or   ( new_n53459_, new_n53458_, new_n524_ );
and  ( new_n53460_, new_n53459_, new_n53457_ );
nor  ( new_n53461_, new_n53460_, new_n53456_ );
nor  ( new_n53462_, new_n53145_, new_n320_ );
xor  ( new_n53463_, new_n51446_, RIbb2f340_7 );
and  ( new_n53464_, new_n53463_, new_n316_ );
nor  ( new_n53465_, new_n53464_, new_n53462_ );
not  ( new_n53466_, new_n53465_ );
xor  ( new_n53467_, new_n53460_, new_n53456_ );
and  ( new_n53468_, new_n53467_, new_n53466_ );
or   ( new_n53469_, new_n53468_, new_n53461_ );
xor  ( new_n53470_, new_n52919_, new_n52918_ );
and  ( new_n53471_, new_n53470_, new_n53469_ );
nor  ( new_n53472_, new_n53192_, new_n3463_ );
xor  ( new_n53473_, new_n45584_, RIbb2e620_35 );
and  ( new_n53474_, new_n53473_, new_n3293_ );
nor  ( new_n53475_, new_n53474_, new_n53472_ );
not  ( new_n53476_, new_n53475_ );
xor  ( new_n53477_, new_n53470_, new_n53469_ );
and  ( new_n53478_, new_n53477_, new_n53476_ );
or   ( new_n53479_, new_n53478_, new_n53471_ );
xor  ( new_n53480_, new_n52981_, new_n52980_ );
and  ( new_n53481_, new_n53480_, new_n53479_ );
xor  ( new_n53482_, new_n52957_, new_n52953_ );
xnor ( new_n53483_, new_n53482_, new_n52962_ );
xor  ( new_n53484_, new_n53480_, new_n53479_ );
and  ( new_n53485_, new_n53484_, new_n53483_ );
nor  ( new_n53486_, new_n53485_, new_n53481_ );
not  ( new_n53487_, new_n53486_ );
xor  ( new_n53488_, new_n52947_, new_n52946_ );
xnor ( new_n53489_, new_n53228_, new_n53224_ );
xor  ( new_n53490_, new_n53489_, new_n53233_ );
or   ( new_n53491_, new_n53490_, new_n53488_ );
and  ( new_n53492_, new_n53490_, new_n53488_ );
xor  ( new_n53493_, new_n53156_, new_n53155_ );
or   ( new_n53494_, new_n53493_, new_n53492_ );
and  ( new_n53495_, new_n53494_, new_n53491_ );
and  ( new_n53496_, new_n53495_, new_n53487_ );
xor  ( new_n53497_, new_n53495_, new_n53487_ );
xor  ( new_n53498_, new_n53236_, new_n53220_ );
xor  ( new_n53499_, new_n53498_, new_n53240_ );
and  ( new_n53500_, new_n53499_, new_n53497_ );
nor  ( new_n53501_, new_n53500_, new_n53496_ );
not  ( new_n53502_, new_n53501_ );
xor  ( new_n53503_, new_n43888_, new_n7722_ );
or   ( new_n53504_, new_n53503_, new_n8264_ );
or   ( new_n53505_, new_n52972_, new_n8266_ );
and  ( new_n53506_, new_n53505_, new_n53504_ );
xor  ( new_n53507_, new_n44600_, RIbb2e260_43 );
nand ( new_n53508_, new_n53507_, new_n4960_ );
or   ( new_n53509_, new_n52939_, new_n5209_ );
and  ( new_n53510_, new_n53509_, new_n53508_ );
nor  ( new_n53511_, new_n53510_, new_n53506_ );
and  ( new_n53512_, new_n52977_, new_n5371_ );
xor  ( new_n53513_, new_n44407_, RIbb2e170_45 );
and  ( new_n53514_, new_n53513_, new_n5373_ );
or   ( new_n53515_, new_n53514_, new_n53512_ );
nand ( new_n53516_, new_n53510_, new_n53506_ );
and  ( new_n53517_, new_n53516_, new_n53515_ );
or   ( new_n53518_, new_n53517_, new_n53511_ );
xor  ( new_n53519_, new_n52878_, new_n52877_ );
and  ( new_n53520_, new_n53519_, new_n53518_ );
xor  ( new_n53521_, new_n53519_, new_n53518_ );
xnor ( new_n53522_, new_n53198_, new_n53194_ );
xor  ( new_n53523_, new_n53522_, new_n53203_ );
and  ( new_n53524_, new_n53523_, new_n53521_ );
or   ( new_n53525_, new_n53524_, new_n53520_ );
xor  ( new_n53526_, new_n52965_, new_n52949_ );
xor  ( new_n53527_, new_n53526_, new_n52983_ );
or   ( new_n53528_, new_n53527_, new_n53525_ );
and  ( new_n53529_, new_n53527_, new_n53525_ );
xor  ( new_n53530_, new_n53206_, new_n53190_ );
xor  ( new_n53531_, new_n53530_, new_n53209_ );
or   ( new_n53532_, new_n53531_, new_n53529_ );
and  ( new_n53533_, new_n53532_, new_n53528_ );
and  ( new_n53534_, new_n53533_, new_n53502_ );
xor  ( new_n53535_, new_n53533_, new_n53502_ );
xor  ( new_n53536_, new_n53242_, new_n53218_ );
xor  ( new_n53537_, new_n53536_, new_n53246_ );
and  ( new_n53538_, new_n53537_, new_n53535_ );
or   ( new_n53539_, new_n53538_, new_n53534_ );
xor  ( new_n53540_, new_n53451_, new_n53449_ );
nand ( new_n53541_, new_n53540_, new_n53539_ );
and  ( new_n53542_, new_n53541_, new_n53452_ );
xor  ( new_n53543_, new_n53256_, new_n53254_ );
nand ( new_n53544_, new_n53543_, new_n53542_ );
nor  ( new_n53545_, new_n53543_, new_n53542_ );
xor  ( new_n53546_, new_n53118_, new_n53109_ );
xnor ( new_n53547_, new_n53546_, new_n53179_ );
or   ( new_n53548_, new_n53547_, new_n53545_ );
nand ( new_n53549_, new_n53548_, new_n53544_ );
and  ( new_n53550_, new_n53549_, new_n53269_ );
xnor ( new_n53551_, new_n53549_, new_n53269_ );
xor  ( new_n53552_, new_n53181_, new_n53108_ );
xor  ( new_n53553_, new_n53552_, new_n53258_ );
nor  ( new_n53554_, new_n53553_, new_n53551_ );
nor  ( new_n53555_, new_n53554_, new_n53550_ );
xor  ( new_n53556_, new_n53105_, new_n52837_ );
xor  ( new_n53557_, new_n53556_, new_n53260_ );
nor  ( new_n53558_, new_n53557_, new_n53555_ );
and  ( new_n53559_, new_n53557_, new_n53555_ );
xor  ( new_n53560_, new_n53177_, new_n53176_ );
xor  ( new_n53561_, new_n53113_, new_n53111_ );
xor  ( new_n53562_, new_n53561_, new_n53116_ );
and  ( new_n53563_, new_n53562_, new_n53560_ );
xnor ( new_n53564_, new_n53562_, new_n53560_ );
xnor ( new_n53565_, new_n53125_, new_n53124_ );
xor  ( new_n53566_, new_n53137_, new_n53135_ );
xor  ( new_n53567_, new_n53566_, new_n53172_ );
or   ( new_n53568_, new_n53567_, new_n53565_ );
and  ( new_n53569_, new_n53567_, new_n53565_ );
xor  ( new_n53570_, new_n53170_, new_n53165_ );
xor  ( new_n53571_, new_n53130_, new_n53128_ );
xor  ( new_n53572_, new_n53571_, new_n53133_ );
nand ( new_n53573_, new_n53572_, new_n53570_ );
xor  ( new_n53574_, new_n53347_, new_n53346_ );
xor  ( new_n53575_, new_n53388_, new_n53372_ );
and  ( new_n53576_, new_n53575_, new_n53574_ );
xnor ( new_n53577_, new_n53575_, new_n53574_ );
or   ( new_n53578_, new_n53503_, new_n8266_ );
xor  ( new_n53579_, new_n43937_, RIbb2dcc0_55 );
nand ( new_n53580_, new_n53579_, new_n8042_ );
and  ( new_n53581_, new_n53580_, new_n53578_ );
nand ( new_n53582_, new_n53513_, new_n5371_ );
xor  ( new_n53583_, new_n44506_, new_n5203_ );
or   ( new_n53584_, new_n53583_, new_n5604_ );
and  ( new_n53585_, new_n53584_, new_n53582_ );
or   ( new_n53586_, new_n53585_, new_n53581_ );
and  ( new_n53587_, new_n53507_, new_n4958_ );
xor  ( new_n53588_, new_n44681_, RIbb2e260_43 );
and  ( new_n53589_, new_n53588_, new_n4960_ );
or   ( new_n53590_, new_n53589_, new_n53587_ );
xor  ( new_n53591_, new_n53585_, new_n53581_ );
nand ( new_n53592_, new_n53591_, new_n53590_ );
and  ( new_n53593_, new_n53592_, new_n53586_ );
xor  ( new_n53594_, new_n43952_, new_n7174_ );
or   ( new_n53595_, new_n53594_, new_n7732_ );
or   ( new_n53596_, new_n53417_, new_n7734_ );
and  ( new_n53597_, new_n53596_, new_n53595_ );
xor  ( new_n53598_, new_n43799_, new_n8870_ );
or   ( new_n53599_, new_n53598_, new_n9422_ );
or   ( new_n53600_, new_n53412_, new_n9424_ );
and  ( new_n53601_, new_n53600_, new_n53599_ );
nor  ( new_n53602_, new_n53601_, new_n53597_ );
and  ( new_n53603_, new_n53601_, new_n53597_ );
and  ( new_n53604_, new_n53408_, new_n4541_ );
xor  ( new_n53605_, new_n44877_, RIbb2e350_41 );
and  ( new_n53606_, new_n53605_, new_n4543_ );
nor  ( new_n53607_, new_n53606_, new_n53604_ );
nor  ( new_n53608_, new_n53607_, new_n53603_ );
nor  ( new_n53609_, new_n53608_, new_n53602_ );
or   ( new_n53610_, new_n53609_, new_n53593_ );
or   ( new_n53611_, new_n53373_, new_n2809_ );
xor  ( new_n53612_, new_n46137_, RIbb2e800_31 );
nand ( new_n53613_, new_n53612_, new_n2615_ );
and  ( new_n53614_, new_n53613_, new_n53611_ );
nand ( new_n53615_, new_n53382_, new_n2928_ );
xor  ( new_n53616_, new_n45928_, new_n2797_ );
or   ( new_n53617_, new_n53616_, new_n3117_ );
and  ( new_n53618_, new_n53617_, new_n53615_ );
nor  ( new_n53619_, new_n53618_, new_n53614_ );
and  ( new_n53620_, new_n53377_, new_n6508_ );
xor  ( new_n53621_, new_n44183_, RIbb2df90_49 );
and  ( new_n53622_, new_n53621_, new_n6510_ );
or   ( new_n53623_, new_n53622_, new_n53620_ );
xor  ( new_n53624_, new_n53618_, new_n53614_ );
and  ( new_n53625_, new_n53624_, new_n53623_ );
nor  ( new_n53626_, new_n53625_, new_n53619_ );
and  ( new_n53627_, new_n53609_, new_n53593_ );
or   ( new_n53628_, new_n53627_, new_n53626_ );
and  ( new_n53629_, new_n53628_, new_n53610_ );
nor  ( new_n53630_, new_n53629_, new_n53577_ );
or   ( new_n53631_, new_n53630_, new_n53576_ );
xor  ( new_n53632_, new_n53572_, new_n53570_ );
nand ( new_n53633_, new_n53632_, new_n53631_ );
and  ( new_n53634_, new_n53633_, new_n53573_ );
or   ( new_n53635_, new_n53634_, new_n53569_ );
and  ( new_n53636_, new_n53635_, new_n53568_ );
nor  ( new_n53637_, new_n53636_, new_n53564_ );
nor  ( new_n53638_, new_n53637_, new_n53563_ );
xnor ( new_n53639_, new_n53284_, new_n53282_ );
xor  ( new_n53640_, new_n53147_, new_n53143_ );
not  ( new_n53641_, new_n53640_ );
xor  ( new_n53642_, new_n49427_, RIbb2ef80_15 );
and  ( new_n53643_, new_n53642_, new_n662_ );
nor  ( new_n53644_, new_n53359_, new_n757_ );
or   ( new_n53645_, new_n53644_, new_n53643_ );
or   ( new_n53646_, new_n43793_, RIbb2d888_64 );
and  ( new_n53647_, new_n53646_, RIbb2d900_63 );
nand ( new_n53648_, new_n53647_, new_n53645_ );
nor  ( new_n53649_, new_n53647_, new_n53645_ );
xor  ( new_n53650_, new_n48908_, new_n745_ );
nor  ( new_n53651_, new_n53650_, new_n897_ );
and  ( new_n53652_, new_n53354_, new_n820_ );
nor  ( new_n53653_, new_n53652_, new_n53651_ );
or   ( new_n53654_, new_n53653_, new_n53649_ );
and  ( new_n53655_, new_n53654_, new_n53648_ );
nor  ( new_n53656_, new_n53655_, new_n53641_ );
xor  ( new_n53657_, new_n53655_, new_n53641_ );
xor  ( new_n53658_, new_n53302_, new_n53301_ );
and  ( new_n53659_, new_n53658_, new_n53657_ );
nor  ( new_n53660_, new_n53659_, new_n53656_ );
or   ( new_n53661_, new_n53290_, new_n340_ );
xor  ( new_n53662_, new_n50894_, new_n329_ );
or   ( new_n53663_, new_n53662_, new_n337_ );
and  ( new_n53664_, new_n53663_, new_n53661_ );
or   ( new_n53665_, new_n53141_, new_n411_ );
xor  ( new_n53666_, new_n50487_, new_n325_ );
or   ( new_n53667_, new_n53666_, new_n409_ );
and  ( new_n53668_, new_n53667_, new_n53665_ );
or   ( new_n53669_, new_n53668_, new_n53664_ );
xor  ( new_n53670_, new_n46962_, new_n1840_ );
nor  ( new_n53671_, new_n53670_, new_n2122_ );
nor  ( new_n53672_, new_n53298_, new_n2124_ );
or   ( new_n53673_, new_n53672_, new_n53671_ );
xor  ( new_n53674_, new_n53668_, new_n53664_ );
nand ( new_n53675_, new_n53674_, new_n53673_ );
and  ( new_n53676_, new_n53675_, new_n53669_ );
xor  ( new_n53677_, new_n48039_, new_n1126_ );
or   ( new_n53678_, new_n53677_, new_n1364_ );
or   ( new_n53679_, new_n53340_, new_n1366_ );
and  ( new_n53680_, new_n53679_, new_n53678_ );
or   ( new_n53681_, new_n53331_, new_n1595_ );
xor  ( new_n53682_, new_n47296_, new_n1355_ );
or   ( new_n53683_, new_n53682_, new_n1593_ );
and  ( new_n53684_, new_n53683_, new_n53681_ );
nor  ( new_n53685_, new_n53684_, new_n53680_ );
and  ( new_n53686_, new_n53350_, new_n1040_ );
xor  ( new_n53687_, new_n48518_, RIbb2eda0_19 );
and  ( new_n53688_, new_n53687_, new_n1042_ );
nor  ( new_n53689_, new_n53688_, new_n53686_ );
and  ( new_n53690_, new_n53684_, new_n53680_ );
nor  ( new_n53691_, new_n53690_, new_n53689_ );
nor  ( new_n53692_, new_n53691_, new_n53685_ );
or   ( new_n53693_, new_n53692_, new_n53676_ );
xor  ( new_n53694_, RIbb33378_192, RIbb31578_128 );
not  ( new_n53695_, new_n53694_ );
or   ( new_n53696_, new_n53695_, new_n43879_ );
xor  ( new_n53697_, new_n53306_, new_n43945_ );
or   ( new_n53698_, new_n53697_, new_n43983_ );
xor  ( new_n53699_, new_n52908_, new_n43880_ );
or   ( new_n53700_, new_n53699_, new_n43977_ );
and  ( new_n53701_, new_n53700_, new_n53698_ );
or   ( new_n53702_, new_n53701_, new_n53696_ );
and  ( new_n53703_, new_n53463_, new_n314_ );
xor  ( new_n53704_, new_n51477_, RIbb2f340_7 );
and  ( new_n53705_, new_n53704_, new_n316_ );
or   ( new_n53706_, new_n53705_, new_n53703_ );
xor  ( new_n53707_, new_n53701_, new_n53696_ );
nand ( new_n53708_, new_n53707_, new_n53706_ );
and  ( new_n53709_, new_n53708_, new_n53702_ );
nand ( new_n53710_, new_n53323_, new_n2242_ );
xor  ( new_n53711_, new_n46619_, new_n2118_ );
or   ( new_n53712_, new_n53711_, new_n2425_ );
and  ( new_n53713_, new_n53712_, new_n53710_ );
or   ( new_n53714_, new_n53713_, new_n53709_ );
xor  ( new_n53715_, new_n47303_, new_n1583_ );
nor  ( new_n53716_, new_n53715_, new_n1844_ );
and  ( new_n53717_, new_n53335_, new_n1739_ );
or   ( new_n53718_, new_n53717_, new_n53716_ );
xor  ( new_n53719_, new_n53713_, new_n53709_ );
nand ( new_n53720_, new_n53719_, new_n53718_ );
and  ( new_n53721_, new_n53720_, new_n53714_ );
and  ( new_n53722_, new_n53692_, new_n53676_ );
or   ( new_n53723_, new_n53722_, new_n53721_ );
and  ( new_n53724_, new_n53723_, new_n53693_ );
or   ( new_n53725_, new_n53724_, new_n53660_ );
and  ( new_n53726_, new_n53724_, new_n53660_ );
xnor ( new_n53727_, new_n53357_, new_n53353_ );
xor  ( new_n53728_, new_n53727_, new_n53362_ );
xnor ( new_n53729_, new_n53337_, new_n53333_ );
nand ( new_n53730_, new_n53729_, new_n53342_ );
not  ( new_n53731_, new_n53344_ );
or   ( new_n53732_, new_n53731_, new_n53338_ );
and  ( new_n53733_, new_n53732_, new_n53730_ );
nand ( new_n53734_, new_n53733_, new_n53728_ );
nor  ( new_n53735_, new_n53733_, new_n53728_ );
xor  ( new_n53736_, new_n45119_, new_n3892_ );
or   ( new_n53737_, new_n53736_, new_n4302_ );
or   ( new_n53738_, new_n53397_, new_n4304_ );
and  ( new_n53739_, new_n53738_, new_n53737_ );
xor  ( new_n53740_, new_n43812_, new_n6635_ );
or   ( new_n53741_, new_n53740_, new_n7184_ );
or   ( new_n53742_, new_n53392_, new_n7186_ );
and  ( new_n53743_, new_n53742_, new_n53741_ );
or   ( new_n53744_, new_n53743_, new_n53739_ );
and  ( new_n53745_, new_n53401_, new_n3731_ );
xor  ( new_n53746_, new_n45403_, new_n3457_ );
nor  ( new_n53747_, new_n53746_, new_n3896_ );
nor  ( new_n53748_, new_n53747_, new_n53745_ );
and  ( new_n53749_, new_n53743_, new_n53739_ );
or   ( new_n53750_, new_n53749_, new_n53748_ );
and  ( new_n53751_, new_n53750_, new_n53744_ );
or   ( new_n53752_, new_n53751_, new_n53735_ );
and  ( new_n53753_, new_n53752_, new_n53734_ );
or   ( new_n53754_, new_n53753_, new_n53726_ );
and  ( new_n53755_, new_n53754_, new_n53725_ );
nor  ( new_n53756_, new_n53755_, new_n53639_ );
xor  ( new_n53757_, new_n53755_, new_n53639_ );
xor  ( new_n53758_, new_n53444_, new_n53443_ );
and  ( new_n53759_, new_n53758_, new_n53757_ );
or   ( new_n53760_, new_n53759_, new_n53756_ );
xor  ( new_n53761_, new_n53447_, new_n53446_ );
and  ( new_n53762_, new_n53761_, new_n53760_ );
xor  ( new_n53763_, new_n52280_, new_n275_ );
or   ( new_n53764_, new_n53763_, new_n283_ );
or   ( new_n53765_, new_n53453_, new_n286_ );
and  ( new_n53766_, new_n53765_, new_n53764_ );
not  ( new_n53767_, new_n52903_ );
or   ( new_n53768_, new_n53767_, new_n44007_ );
nand ( new_n53769_, new_n53041_, new_n295_ );
and  ( new_n53770_, new_n53769_, new_n53768_ );
nor  ( new_n53771_, new_n53770_, new_n53766_ );
and  ( new_n53772_, new_n53704_, new_n314_ );
xor  ( new_n53773_, new_n51758_, new_n309_ );
nor  ( new_n53774_, new_n53773_, new_n317_ );
nor  ( new_n53775_, new_n53774_, new_n53772_ );
not  ( new_n53776_, new_n53775_ );
and  ( new_n53777_, new_n53695_, new_n43945_ );
or   ( new_n53778_, new_n53777_, new_n43976_ );
or   ( new_n53779_, new_n53695_, new_n43945_ );
and  ( new_n53780_, new_n53779_, new_n43880_ );
and  ( new_n53781_, new_n53780_, new_n53778_ );
and  ( new_n53782_, new_n53781_, new_n53776_ );
xor  ( new_n53783_, new_n53770_, new_n53766_ );
and  ( new_n53784_, new_n53783_, new_n53782_ );
or   ( new_n53785_, new_n53784_, new_n53771_ );
xor  ( new_n53786_, new_n53317_, new_n53316_ );
and  ( new_n53787_, new_n53786_, new_n53785_ );
xor  ( new_n53788_, new_n45738_, RIbb2e620_35 );
and  ( new_n53789_, new_n53788_, new_n3293_ );
and  ( new_n53790_, new_n53473_, new_n3291_ );
or   ( new_n53791_, new_n53790_, new_n53789_ );
xor  ( new_n53792_, new_n53786_, new_n53785_ );
and  ( new_n53793_, new_n53792_, new_n53791_ );
nor  ( new_n53794_, new_n53793_, new_n53787_ );
xnor ( new_n53795_, new_n53326_, new_n53325_ );
nor  ( new_n53796_, new_n53795_, new_n53794_ );
xnor ( new_n53797_, new_n53795_, new_n53794_ );
or   ( new_n53798_, new_n53430_, new_n6175_ );
xor  ( new_n53799_, new_n44319_, RIbb2e080_47 );
nand ( new_n53800_, new_n53799_, new_n5917_ );
and  ( new_n53801_, new_n53800_, new_n53798_ );
nand ( new_n53802_, new_n53434_, new_n8649_ );
xor  ( new_n53803_, new_n43884_, RIbb2dbd0_57 );
nand ( new_n53804_, new_n53803_, new_n8651_ );
and  ( new_n53805_, new_n53804_, new_n53802_ );
or   ( new_n53806_, new_n53805_, new_n53801_ );
and  ( new_n53807_, new_n53425_, new_n9738_ );
xor  ( new_n53808_, new_n43898_, new_n9418_ );
nor  ( new_n53809_, new_n53808_, new_n10059_ );
nor  ( new_n53810_, new_n53809_, new_n53807_ );
and  ( new_n53811_, new_n53805_, new_n53801_ );
or   ( new_n53812_, new_n53811_, new_n53810_ );
and  ( new_n53813_, new_n53812_, new_n53806_ );
nor  ( new_n53814_, new_n53813_, new_n53797_ );
nor  ( new_n53815_, new_n53814_, new_n53796_ );
not  ( new_n53816_, new_n53815_ );
xor  ( new_n53817_, new_n53276_, new_n53275_ );
and  ( new_n53818_, new_n53817_, new_n53816_ );
xor  ( new_n53819_, new_n53817_, new_n53816_ );
xor  ( new_n53820_, new_n53441_, new_n53440_ );
and  ( new_n53821_, new_n53820_, new_n53819_ );
nor  ( new_n53822_, new_n53821_, new_n53818_ );
xor  ( new_n53823_, new_n53510_, new_n53506_ );
xor  ( new_n53824_, new_n53823_, new_n53515_ );
xnor ( new_n53825_, new_n53415_, new_n53411_ );
xor  ( new_n53826_, new_n53825_, new_n53420_ );
or   ( new_n53827_, new_n53826_, new_n53824_ );
and  ( new_n53828_, new_n53826_, new_n53824_ );
xor  ( new_n53829_, new_n53405_, new_n53404_ );
or   ( new_n53830_, new_n53829_, new_n53828_ );
and  ( new_n53831_, new_n53830_, new_n53827_ );
xor  ( new_n53832_, new_n53438_, new_n53437_ );
xnor ( new_n53833_, new_n53380_, new_n53376_ );
nand ( new_n53834_, new_n53833_, new_n53385_ );
not  ( new_n53835_, new_n53387_ );
or   ( new_n53836_, new_n53835_, new_n53381_ );
and  ( new_n53837_, new_n53836_, new_n53834_ );
or   ( new_n53838_, new_n53837_, new_n53832_ );
and  ( new_n53839_, new_n53837_, new_n53832_ );
xor  ( new_n53840_, new_n53477_, new_n53476_ );
or   ( new_n53841_, new_n53840_, new_n53839_ );
and  ( new_n53842_, new_n53841_, new_n53838_ );
nand ( new_n53843_, new_n53842_, new_n53831_ );
xor  ( new_n53844_, new_n53523_, new_n53521_ );
xor  ( new_n53845_, new_n53842_, new_n53831_ );
nand ( new_n53846_, new_n53845_, new_n53844_ );
and  ( new_n53847_, new_n53846_, new_n53843_ );
nor  ( new_n53848_, new_n53847_, new_n53822_ );
xor  ( new_n53849_, new_n53847_, new_n53822_ );
not  ( new_n53850_, new_n53849_ );
xnor ( new_n53851_, new_n53527_, new_n53525_ );
xor  ( new_n53852_, new_n53851_, new_n53531_ );
nor  ( new_n53853_, new_n53852_, new_n53850_ );
nor  ( new_n53854_, new_n53853_, new_n53848_ );
xnor ( new_n53855_, new_n53761_, new_n53760_ );
nor  ( new_n53856_, new_n53855_, new_n53854_ );
nor  ( new_n53857_, new_n53856_, new_n53762_ );
xnor ( new_n53858_, new_n53540_, new_n53539_ );
or   ( new_n53859_, new_n53858_, new_n53857_ );
xnor ( new_n53860_, new_n53858_, new_n53857_ );
xnor ( new_n53861_, new_n53537_, new_n53535_ );
xor  ( new_n53862_, new_n53567_, new_n53565_ );
xor  ( new_n53863_, new_n53862_, new_n53634_ );
or   ( new_n53864_, new_n53863_, new_n53861_ );
and  ( new_n53865_, new_n53863_, new_n53861_ );
xnor ( new_n53866_, new_n53499_, new_n53497_ );
xnor ( new_n53867_, new_n53484_, new_n53483_ );
xnor ( new_n53868_, new_n53490_, new_n53488_ );
xor  ( new_n53869_, new_n53868_, new_n53493_ );
or   ( new_n53870_, new_n53869_, new_n53867_ );
and  ( new_n53871_, new_n53869_, new_n53867_ );
xnor ( new_n53872_, new_n53658_, new_n53657_ );
nand ( new_n53873_, new_n53621_, new_n6508_ );
xor  ( new_n53874_, new_n44218_, new_n6163_ );
or   ( new_n53875_, new_n53874_, new_n6645_ );
and  ( new_n53876_, new_n53875_, new_n53873_ );
and  ( new_n53877_, new_n43793_, new_n10052_ );
nor  ( new_n53878_, new_n43793_, new_n10052_ );
or   ( new_n53879_, new_n53878_, new_n21077_ );
or   ( new_n53880_, new_n53879_, new_n53877_ );
or   ( new_n53881_, new_n43787_, new_n10052_ );
or   ( new_n53882_, new_n53881_, RIbb2d888_64 );
and  ( new_n53883_, new_n53882_, new_n53880_ );
nor  ( new_n53884_, new_n53883_, new_n53876_ );
and  ( new_n53885_, new_n53799_, new_n5915_ );
xor  ( new_n53886_, new_n44407_, RIbb2e080_47 );
and  ( new_n53887_, new_n53886_, new_n5917_ );
or   ( new_n53888_, new_n53887_, new_n53885_ );
xor  ( new_n53889_, new_n53883_, new_n53876_ );
and  ( new_n53890_, new_n53889_, new_n53888_ );
nor  ( new_n53891_, new_n53890_, new_n53884_ );
not  ( new_n53892_, new_n53891_ );
or   ( new_n53893_, new_n53650_, new_n899_ );
xor  ( new_n53894_, new_n49265_, new_n745_ );
or   ( new_n53895_, new_n53894_, new_n897_ );
and  ( new_n53896_, new_n53895_, new_n53893_ );
xor  ( new_n53897_, new_n46037_, new_n2797_ );
or   ( new_n53898_, new_n53897_, new_n3117_ );
or   ( new_n53899_, new_n53616_, new_n3119_ );
and  ( new_n53900_, new_n53899_, new_n53898_ );
nor  ( new_n53901_, new_n53900_, new_n53896_ );
and  ( new_n53902_, new_n53900_, new_n53896_ );
and  ( new_n53903_, new_n53803_, new_n8649_ );
xor  ( new_n53904_, new_n43888_, RIbb2dbd0_57 );
and  ( new_n53905_, new_n53904_, new_n8651_ );
nor  ( new_n53906_, new_n53905_, new_n53903_ );
nor  ( new_n53907_, new_n53906_, new_n53902_ );
nor  ( new_n53908_, new_n53907_, new_n53901_ );
not  ( new_n53909_, new_n53908_ );
and  ( new_n53910_, new_n53909_, new_n53892_ );
and  ( new_n53911_, new_n53908_, new_n53891_ );
or   ( new_n53912_, new_n53598_, new_n9424_ );
xor  ( new_n53913_, new_n43803_, new_n8870_ );
or   ( new_n53914_, new_n53913_, new_n9422_ );
and  ( new_n53915_, new_n53914_, new_n53912_ );
xor  ( new_n53916_, new_n44974_, new_n4292_ );
or   ( new_n53917_, new_n53916_, new_n4709_ );
nand ( new_n53918_, new_n53605_, new_n4541_ );
and  ( new_n53919_, new_n53918_, new_n53917_ );
nor  ( new_n53920_, new_n53919_, new_n53915_ );
and  ( new_n53921_, new_n53588_, new_n4958_ );
xor  ( new_n53922_, new_n44785_, RIbb2e260_43 );
and  ( new_n53923_, new_n53922_, new_n4960_ );
nor  ( new_n53924_, new_n53923_, new_n53921_ );
and  ( new_n53925_, new_n53919_, new_n53915_ );
nor  ( new_n53926_, new_n53925_, new_n53924_ );
nor  ( new_n53927_, new_n53926_, new_n53920_ );
nor  ( new_n53928_, new_n53927_, new_n53911_ );
nor  ( new_n53929_, new_n53928_, new_n53910_ );
or   ( new_n53930_, new_n53929_, new_n53872_ );
nor  ( new_n53931_, new_n53594_, new_n7734_ );
xor  ( new_n53932_, new_n43985_, RIbb2ddb0_53 );
and  ( new_n53933_, new_n53932_, new_n7489_ );
or   ( new_n53934_, new_n53933_, new_n53931_ );
xor  ( new_n53935_, new_n53707_, new_n53706_ );
and  ( new_n53936_, new_n53935_, new_n53934_ );
nor  ( new_n53937_, new_n53736_, new_n4304_ );
xor  ( new_n53938_, new_n45204_, RIbb2e440_39 );
and  ( new_n53939_, new_n53938_, new_n4034_ );
or   ( new_n53940_, new_n53939_, new_n53937_ );
xor  ( new_n53941_, new_n53935_, new_n53934_ );
and  ( new_n53942_, new_n53941_, new_n53940_ );
nor  ( new_n53943_, new_n53942_, new_n53936_ );
or   ( new_n53944_, new_n53746_, new_n3898_ );
xor  ( new_n53945_, new_n45584_, RIbb2e530_37 );
nand ( new_n53946_, new_n53945_, new_n3733_ );
and  ( new_n53947_, new_n53946_, new_n53944_ );
or   ( new_n53948_, new_n53740_, new_n7186_ );
xor  ( new_n53949_, new_n43914_, new_n6635_ );
or   ( new_n53950_, new_n53949_, new_n7184_ );
and  ( new_n53951_, new_n53950_, new_n53948_ );
or   ( new_n53952_, new_n53951_, new_n53947_ );
xor  ( new_n53953_, new_n45597_, RIbb2e620_35 );
and  ( new_n53954_, new_n53953_, new_n3293_ );
and  ( new_n53955_, new_n53788_, new_n3291_ );
or   ( new_n53956_, new_n53955_, new_n53954_ );
xor  ( new_n53957_, new_n53951_, new_n53947_ );
nand ( new_n53958_, new_n53957_, new_n53956_ );
and  ( new_n53959_, new_n53958_, new_n53952_ );
nor  ( new_n53960_, new_n53959_, new_n53943_ );
xor  ( new_n53961_, new_n53959_, new_n53943_ );
xnor ( new_n53962_, new_n53647_, new_n53645_ );
xor  ( new_n53963_, new_n53962_, new_n53653_ );
and  ( new_n53964_, new_n53963_, new_n53961_ );
nor  ( new_n53965_, new_n53964_, new_n53960_ );
not  ( new_n53966_, new_n53965_ );
xor  ( new_n53967_, new_n53929_, new_n53872_ );
nand ( new_n53968_, new_n53967_, new_n53966_ );
and  ( new_n53969_, new_n53968_, new_n53930_ );
or   ( new_n53970_, new_n53969_, new_n53871_ );
and  ( new_n53971_, new_n53970_, new_n53870_ );
or   ( new_n53972_, new_n53971_, new_n53866_ );
xor  ( new_n53973_, new_n53971_, new_n53866_ );
xor  ( new_n53974_, new_n53632_, new_n53631_ );
nand ( new_n53975_, new_n53974_, new_n53973_ );
and  ( new_n53976_, new_n53975_, new_n53972_ );
or   ( new_n53977_, new_n53976_, new_n53865_ );
and  ( new_n53978_, new_n53977_, new_n53864_ );
or   ( new_n53979_, new_n53978_, new_n53860_ );
and  ( new_n53980_, new_n53979_, new_n53859_ );
or   ( new_n53981_, new_n53980_, new_n53638_ );
xnor ( new_n53982_, new_n53980_, new_n53638_ );
xnor ( new_n53983_, new_n53543_, new_n53542_ );
xor  ( new_n53984_, new_n53983_, new_n53547_ );
or   ( new_n53985_, new_n53984_, new_n53982_ );
and  ( new_n53986_, new_n53985_, new_n53981_ );
xor  ( new_n53987_, new_n53553_, new_n53551_ );
and  ( new_n53988_, new_n53987_, new_n53986_ );
nor  ( new_n53989_, new_n53987_, new_n53986_ );
xnor ( new_n53990_, new_n53855_, new_n53854_ );
xor  ( new_n53991_, new_n53467_, new_n53466_ );
xor  ( new_n53992_, new_n53674_, new_n53673_ );
and  ( new_n53993_, new_n53992_, new_n53991_ );
xor  ( new_n53994_, new_n53992_, new_n53991_ );
not  ( new_n53995_, new_n53994_ );
xor  ( new_n53996_, new_n48291_, RIbb2ecb0_21 );
nand ( new_n53997_, new_n53996_, new_n1253_ );
or   ( new_n53998_, new_n53677_, new_n1366_ );
and  ( new_n53999_, new_n53998_, new_n53997_ );
nand ( new_n54000_, new_n53687_, new_n1040_ );
xor  ( new_n54001_, new_n48756_, RIbb2eda0_19 );
nand ( new_n54002_, new_n54001_, new_n1042_ );
and  ( new_n54003_, new_n54002_, new_n54000_ );
nor  ( new_n54004_, new_n54003_, new_n53999_ );
and  ( new_n54005_, new_n53612_, new_n2613_ );
xor  ( new_n54006_, new_n46427_, RIbb2e800_31 );
and  ( new_n54007_, new_n54006_, new_n2615_ );
nor  ( new_n54008_, new_n54007_, new_n54005_ );
and  ( new_n54009_, new_n54003_, new_n53999_ );
nor  ( new_n54010_, new_n54009_, new_n54008_ );
nor  ( new_n54011_, new_n54010_, new_n54004_ );
nor  ( new_n54012_, new_n54011_, new_n53995_ );
nor  ( new_n54013_, new_n54012_, new_n53993_ );
nor  ( new_n54014_, new_n53662_, new_n340_ );
xor  ( new_n54015_, new_n51142_, new_n329_ );
nor  ( new_n54016_, new_n54015_, new_n337_ );
nor  ( new_n54017_, new_n54016_, new_n54014_ );
or   ( new_n54018_, new_n53666_, new_n411_ );
xor  ( new_n54019_, new_n50788_, new_n325_ );
or   ( new_n54020_, new_n54019_, new_n409_ );
and  ( new_n54021_, new_n54020_, new_n54018_ );
nor  ( new_n54022_, new_n54021_, new_n54017_ );
and  ( new_n54023_, new_n53642_, new_n660_ );
xor  ( new_n54024_, new_n49488_, RIbb2ef80_15 );
and  ( new_n54025_, new_n54024_, new_n662_ );
nor  ( new_n54026_, new_n54025_, new_n54023_ );
and  ( new_n54027_, new_n54021_, new_n54017_ );
nor  ( new_n54028_, new_n54027_, new_n54026_ );
nor  ( new_n54029_, new_n54028_, new_n54022_ );
or   ( new_n54030_, new_n53458_, new_n526_ );
xor  ( new_n54031_, new_n50115_, new_n400_ );
or   ( new_n54032_, new_n54031_, new_n524_ );
and  ( new_n54033_, new_n54032_, new_n54030_ );
or   ( new_n54034_, new_n53711_, new_n2427_ );
xor  ( new_n54035_, new_n46789_, new_n2118_ );
or   ( new_n54036_, new_n54035_, new_n2425_ );
and  ( new_n54037_, new_n54036_, new_n54034_ );
or   ( new_n54038_, new_n54037_, new_n54033_ );
xor  ( new_n54039_, new_n46958_, RIbb2e9e0_27 );
and  ( new_n54040_, new_n54039_, new_n2002_ );
nor  ( new_n54041_, new_n53670_, new_n2124_ );
or   ( new_n54042_, new_n54041_, new_n54040_ );
xor  ( new_n54043_, new_n54037_, new_n54033_ );
nand ( new_n54044_, new_n54043_, new_n54042_ );
and  ( new_n54045_, new_n54044_, new_n54038_ );
or   ( new_n54046_, new_n54045_, new_n54029_ );
xnor ( new_n54047_, new_n54045_, new_n54029_ );
nor  ( new_n54048_, new_n53715_, new_n1846_ );
xor  ( new_n54049_, new_n47046_, new_n1583_ );
nor  ( new_n54050_, new_n54049_, new_n1844_ );
nor  ( new_n54051_, new_n54050_, new_n54048_ );
or   ( new_n54052_, new_n53682_, new_n1595_ );
xor  ( new_n54053_, new_n47640_, new_n1355_ );
or   ( new_n54054_, new_n54053_, new_n1593_ );
and  ( new_n54055_, new_n54054_, new_n54052_ );
nor  ( new_n54056_, new_n54055_, new_n54051_ );
and  ( new_n54057_, new_n54055_, new_n54051_ );
not  ( new_n54058_, new_n53308_ );
or   ( new_n54059_, new_n54058_, new_n44007_ );
or   ( new_n54060_, new_n53767_, new_n302_ );
and  ( new_n54061_, new_n54060_, new_n54059_ );
xor  ( new_n54062_, new_n53694_, new_n43950_ );
or   ( new_n54063_, new_n54062_, new_n43983_ );
xor  ( new_n54064_, new_n53306_, new_n43880_ );
or   ( new_n54065_, new_n54064_, new_n43977_ );
and  ( new_n54066_, new_n54065_, new_n54063_ );
nor  ( new_n54067_, new_n54066_, new_n54061_ );
nor  ( new_n54068_, new_n53763_, new_n286_ );
xor  ( new_n54069_, new_n52293_, RIbb2f430_5 );
nor  ( new_n54070_, new_n54069_, new_n283_ );
nor  ( new_n54071_, new_n54070_, new_n54068_ );
xnor ( new_n54072_, new_n54066_, new_n54061_ );
nor  ( new_n54073_, new_n54072_, new_n54071_ );
nor  ( new_n54074_, new_n54073_, new_n54067_ );
nor  ( new_n54075_, new_n54074_, new_n54057_ );
nor  ( new_n54076_, new_n54075_, new_n54056_ );
or   ( new_n54077_, new_n54076_, new_n54047_ );
and  ( new_n54078_, new_n54077_, new_n54046_ );
nor  ( new_n54079_, new_n54078_, new_n54013_ );
xor  ( new_n54080_, new_n54078_, new_n54013_ );
xor  ( new_n54081_, new_n53719_, new_n53718_ );
xnor ( new_n54082_, new_n53684_, new_n53680_ );
nand ( new_n54083_, new_n54082_, new_n53689_ );
not  ( new_n54084_, new_n53691_ );
or   ( new_n54085_, new_n54084_, new_n53685_ );
and  ( new_n54086_, new_n54085_, new_n54083_ );
or   ( new_n54087_, new_n54086_, new_n54081_ );
and  ( new_n54088_, new_n54086_, new_n54081_ );
or   ( new_n54089_, new_n53583_, new_n5606_ );
xor  ( new_n54090_, new_n44600_, RIbb2e170_45 );
nand ( new_n54091_, new_n54090_, new_n5373_ );
and  ( new_n54092_, new_n54091_, new_n54089_ );
xor  ( new_n54093_, new_n43894_, new_n9418_ );
or   ( new_n54094_, new_n54093_, new_n10059_ );
or   ( new_n54095_, new_n53808_, new_n10061_ );
and  ( new_n54096_, new_n54095_, new_n54094_ );
nor  ( new_n54097_, new_n54096_, new_n54092_ );
xor  ( new_n54098_, new_n43956_, new_n7722_ );
nor  ( new_n54099_, new_n54098_, new_n8264_ );
and  ( new_n54100_, new_n53579_, new_n8040_ );
or   ( new_n54101_, new_n54100_, new_n54099_ );
xor  ( new_n54102_, new_n54096_, new_n54092_ );
and  ( new_n54103_, new_n54102_, new_n54101_ );
or   ( new_n54104_, new_n54103_, new_n54097_ );
or   ( new_n54105_, new_n54104_, new_n54088_ );
and  ( new_n54106_, new_n54105_, new_n54087_ );
and  ( new_n54107_, new_n54106_, new_n54080_ );
or   ( new_n54108_, new_n54107_, new_n54079_ );
xnor ( new_n54109_, new_n53753_, new_n53660_ );
xor  ( new_n54110_, new_n54109_, new_n53724_ );
and  ( new_n54111_, new_n54110_, new_n54108_ );
xor  ( new_n54112_, new_n53692_, new_n53676_ );
xor  ( new_n54113_, new_n54112_, new_n53721_ );
xor  ( new_n54114_, new_n53733_, new_n53728_ );
xor  ( new_n54115_, new_n54114_, new_n53751_ );
nor  ( new_n54116_, new_n54115_, new_n54113_ );
xor  ( new_n54117_, new_n53609_, new_n53593_ );
xnor ( new_n54118_, new_n54117_, new_n53626_ );
xor  ( new_n54119_, new_n54115_, new_n54113_ );
and  ( new_n54120_, new_n54119_, new_n54118_ );
nor  ( new_n54121_, new_n54120_, new_n54116_ );
nor  ( new_n54122_, new_n54110_, new_n54108_ );
nor  ( new_n54123_, new_n54122_, new_n54121_ );
or   ( new_n54124_, new_n54123_, new_n54111_ );
xor  ( new_n54125_, new_n53758_, new_n53757_ );
nand ( new_n54126_, new_n54125_, new_n54124_ );
or   ( new_n54127_, new_n54125_, new_n54124_ );
xor  ( new_n54128_, new_n53852_, new_n53850_ );
nand ( new_n54129_, new_n54128_, new_n54127_ );
and  ( new_n54130_, new_n54129_, new_n54126_ );
nor  ( new_n54131_, new_n54130_, new_n53990_ );
xor  ( new_n54132_, new_n53629_, new_n53577_ );
xnor ( new_n54133_, new_n53743_, new_n53739_ );
xor  ( new_n54134_, new_n54133_, new_n53748_ );
xnor ( new_n54135_, new_n53601_, new_n53597_ );
nand ( new_n54136_, new_n54135_, new_n53607_ );
not  ( new_n54137_, new_n53608_ );
or   ( new_n54138_, new_n54137_, new_n53602_ );
and  ( new_n54139_, new_n54138_, new_n54136_ );
or   ( new_n54140_, new_n54139_, new_n54134_ );
and  ( new_n54141_, new_n54139_, new_n54134_ );
xor  ( new_n54142_, new_n53591_, new_n53590_ );
or   ( new_n54143_, new_n54142_, new_n54141_ );
and  ( new_n54144_, new_n54143_, new_n54140_ );
xor  ( new_n54145_, new_n53813_, new_n53797_ );
or   ( new_n54146_, new_n54145_, new_n54144_ );
xor  ( new_n54147_, new_n53624_, new_n53623_ );
xnor ( new_n54148_, new_n53805_, new_n53801_ );
xor  ( new_n54149_, new_n54148_, new_n53810_ );
or   ( new_n54150_, new_n54149_, new_n54147_ );
and  ( new_n54151_, new_n54149_, new_n54147_ );
xor  ( new_n54152_, new_n53792_, new_n53791_ );
or   ( new_n54153_, new_n54152_, new_n54151_ );
and  ( new_n54154_, new_n54153_, new_n54150_ );
and  ( new_n54155_, new_n54145_, new_n54144_ );
or   ( new_n54156_, new_n54155_, new_n54154_ );
and  ( new_n54157_, new_n54156_, new_n54146_ );
nand ( new_n54158_, new_n54157_, new_n54132_ );
xor  ( new_n54159_, new_n53845_, new_n53844_ );
xor  ( new_n54160_, new_n54157_, new_n54132_ );
nand ( new_n54161_, new_n54160_, new_n54159_ );
and  ( new_n54162_, new_n54161_, new_n54158_ );
xor  ( new_n54163_, new_n53820_, new_n53819_ );
xor  ( new_n54164_, new_n54011_, new_n53995_ );
xor  ( new_n54165_, new_n54043_, new_n54042_ );
xnor ( new_n54166_, new_n54003_, new_n53999_ );
nand ( new_n54167_, new_n54166_, new_n54008_ );
not  ( new_n54168_, new_n54010_ );
or   ( new_n54169_, new_n54168_, new_n54004_ );
and  ( new_n54170_, new_n54169_, new_n54167_ );
nand ( new_n54171_, new_n54170_, new_n54165_ );
nor  ( new_n54172_, new_n54170_, new_n54165_ );
or   ( new_n54173_, new_n54098_, new_n8266_ );
xor  ( new_n54174_, new_n43952_, new_n7722_ );
or   ( new_n54175_, new_n54174_, new_n8264_ );
and  ( new_n54176_, new_n54175_, new_n54173_ );
xor  ( new_n54177_, new_n44877_, RIbb2e260_43 );
nand ( new_n54178_, new_n54177_, new_n4960_ );
nand ( new_n54179_, new_n53922_, new_n4958_ );
and  ( new_n54180_, new_n54179_, new_n54178_ );
nor  ( new_n54181_, new_n54180_, new_n54176_ );
and  ( new_n54182_, new_n54090_, new_n5371_ );
xor  ( new_n54183_, new_n44681_, RIbb2e170_45 );
and  ( new_n54184_, new_n54183_, new_n5373_ );
or   ( new_n54185_, new_n54184_, new_n54182_ );
xor  ( new_n54186_, new_n54180_, new_n54176_ );
and  ( new_n54187_, new_n54186_, new_n54185_ );
nor  ( new_n54188_, new_n54187_, new_n54181_ );
or   ( new_n54189_, new_n54188_, new_n54172_ );
nand ( new_n54190_, new_n54189_, new_n54171_ );
and  ( new_n54191_, new_n54190_, new_n54164_ );
xnor ( new_n54192_, new_n54190_, new_n54164_ );
xnor ( new_n54193_, new_n54021_, new_n54017_ );
and  ( new_n54194_, new_n54193_, new_n54026_ );
not  ( new_n54195_, new_n54022_ );
and  ( new_n54196_, new_n54028_, new_n54195_ );
or   ( new_n54197_, new_n54196_, new_n54194_ );
xor  ( new_n54198_, new_n44319_, RIbb2df90_49 );
nand ( new_n54199_, new_n54198_, new_n6510_ );
or   ( new_n54200_, new_n53874_, new_n6647_ );
and  ( new_n54201_, new_n54200_, new_n54199_ );
or   ( new_n54202_, new_n53897_, new_n3119_ );
xor  ( new_n54203_, new_n46137_, RIbb2e710_33 );
nand ( new_n54204_, new_n54203_, new_n2930_ );
and  ( new_n54205_, new_n54204_, new_n54202_ );
nor  ( new_n54206_, new_n54205_, new_n54201_ );
and  ( new_n54207_, new_n54205_, new_n54201_ );
xor  ( new_n54208_, new_n43937_, RIbb2dbd0_57 );
and  ( new_n54209_, new_n54208_, new_n8651_ );
and  ( new_n54210_, new_n53904_, new_n8649_ );
nor  ( new_n54211_, new_n54210_, new_n54209_ );
nor  ( new_n54212_, new_n54211_, new_n54207_ );
nor  ( new_n54213_, new_n54212_, new_n54206_ );
or   ( new_n54214_, new_n54213_, new_n54197_ );
nand ( new_n54215_, new_n54213_, new_n54197_ );
xor  ( new_n54216_, new_n54055_, new_n54051_ );
not  ( new_n54217_, new_n54216_ );
and  ( new_n54218_, new_n54217_, new_n54074_ );
not  ( new_n54219_, new_n54056_ );
and  ( new_n54220_, new_n54075_, new_n54219_ );
nor  ( new_n54221_, new_n54220_, new_n54218_ );
nand ( new_n54222_, new_n54221_, new_n54215_ );
and  ( new_n54223_, new_n54222_, new_n54214_ );
nor  ( new_n54224_, new_n54223_, new_n54192_ );
or   ( new_n54225_, new_n54224_, new_n54191_ );
xor  ( new_n54226_, new_n53826_, new_n53824_ );
xor  ( new_n54227_, new_n54226_, new_n53829_ );
nand ( new_n54228_, new_n54227_, new_n54225_ );
nor  ( new_n54229_, new_n54227_, new_n54225_ );
xor  ( new_n54230_, new_n53837_, new_n53832_ );
xnor ( new_n54231_, new_n54230_, new_n53840_ );
or   ( new_n54232_, new_n54231_, new_n54229_ );
nand ( new_n54233_, new_n54232_, new_n54228_ );
nand ( new_n54234_, new_n54233_, new_n54163_ );
xnor ( new_n54235_, new_n54233_, new_n54163_ );
xor  ( new_n54236_, new_n53869_, new_n53867_ );
xor  ( new_n54237_, new_n54236_, new_n53969_ );
or   ( new_n54238_, new_n54237_, new_n54235_ );
and  ( new_n54239_, new_n54238_, new_n54234_ );
nor  ( new_n54240_, new_n54239_, new_n54162_ );
xor  ( new_n54241_, new_n54239_, new_n54162_ );
xor  ( new_n54242_, new_n53974_, new_n53973_ );
and  ( new_n54243_, new_n54242_, new_n54241_ );
nor  ( new_n54244_, new_n54243_, new_n54240_ );
xnor ( new_n54245_, new_n54130_, new_n53990_ );
nor  ( new_n54246_, new_n54245_, new_n54244_ );
nor  ( new_n54247_, new_n54246_, new_n54131_ );
not  ( new_n54248_, new_n54247_ );
xor  ( new_n54249_, new_n53636_, new_n53564_ );
and  ( new_n54250_, new_n54249_, new_n54248_ );
xor  ( new_n54251_, new_n54249_, new_n54248_ );
xor  ( new_n54252_, new_n53978_, new_n53860_ );
and  ( new_n54253_, new_n54252_, new_n54251_ );
or   ( new_n54254_, new_n54253_, new_n54250_ );
xor  ( new_n54255_, new_n53984_, new_n53982_ );
nor  ( new_n54256_, new_n54255_, new_n54254_ );
and  ( new_n54257_, new_n54255_, new_n54254_ );
xor  ( new_n54258_, new_n54252_, new_n54251_ );
xnor ( new_n54259_, new_n54245_, new_n54244_ );
xor  ( new_n54260_, new_n53863_, new_n53861_ );
xor  ( new_n54261_, new_n54260_, new_n53976_ );
nor  ( new_n54262_, new_n54261_, new_n54259_ );
xor  ( new_n54263_, new_n54110_, new_n54108_ );
xor  ( new_n54264_, new_n54263_, new_n54121_ );
xor  ( new_n54265_, new_n54106_, new_n54080_ );
xor  ( new_n54266_, new_n54086_, new_n54081_ );
xor  ( new_n54267_, new_n54266_, new_n54104_ );
xnor ( new_n54268_, new_n53900_, new_n53896_ );
nand ( new_n54269_, new_n54268_, new_n53906_ );
not  ( new_n54270_, new_n53907_ );
or   ( new_n54271_, new_n54270_, new_n53901_ );
and  ( new_n54272_, new_n54271_, new_n54269_ );
xor  ( new_n54273_, new_n53889_, new_n53888_ );
or   ( new_n54274_, new_n54273_, new_n54272_ );
and  ( new_n54275_, new_n54273_, new_n54272_ );
xnor ( new_n54276_, new_n53919_, new_n53915_ );
xor  ( new_n54277_, new_n54276_, new_n53924_ );
or   ( new_n54278_, new_n54277_, new_n54275_ );
and  ( new_n54279_, new_n54278_, new_n54274_ );
nor  ( new_n54280_, new_n54279_, new_n54267_ );
and  ( new_n54281_, new_n54279_, new_n54267_ );
xor  ( new_n54282_, new_n53957_, new_n53956_ );
xor  ( new_n54283_, new_n54102_, new_n54101_ );
nor  ( new_n54284_, new_n54283_, new_n54282_ );
and  ( new_n54285_, new_n54283_, new_n54282_ );
xnor ( new_n54286_, new_n54072_, new_n54071_ );
nand ( new_n54287_, new_n53953_, new_n3291_ );
xor  ( new_n54288_, new_n45928_, new_n3113_ );
or   ( new_n54289_, new_n54288_, new_n3461_ );
and  ( new_n54290_, new_n54289_, new_n54287_ );
and  ( new_n54291_, new_n54290_, new_n54286_ );
xor  ( new_n54292_, new_n50788_, new_n400_ );
or   ( new_n54293_, new_n54292_, new_n524_ );
xor  ( new_n54294_, new_n50487_, new_n400_ );
or   ( new_n54295_, new_n54294_, new_n526_ );
and  ( new_n54296_, new_n54295_, new_n54293_ );
xor  ( new_n54297_, new_n51142_, new_n325_ );
or   ( new_n54298_, new_n54297_, new_n409_ );
xor  ( new_n54299_, new_n50894_, new_n325_ );
or   ( new_n54300_, new_n54299_, new_n411_ );
and  ( new_n54301_, new_n54300_, new_n54298_ );
nor  ( new_n54302_, new_n54301_, new_n54296_ );
xor  ( new_n54303_, new_n50115_, new_n520_ );
nor  ( new_n54304_, new_n54303_, new_n755_ );
xor  ( new_n54305_, new_n49758_, new_n520_ );
nor  ( new_n54306_, new_n54305_, new_n757_ );
nor  ( new_n54307_, new_n54306_, new_n54304_ );
and  ( new_n54308_, new_n54301_, new_n54296_ );
nor  ( new_n54309_, new_n54308_, new_n54307_ );
nor  ( new_n54310_, new_n54309_, new_n54302_ );
nor  ( new_n54311_, new_n54290_, new_n54286_ );
not  ( new_n54312_, new_n54311_ );
and  ( new_n54313_, new_n54312_, new_n54310_ );
nor  ( new_n54314_, new_n54313_, new_n54291_ );
nor  ( new_n54315_, new_n54314_, new_n54285_ );
nor  ( new_n54316_, new_n54315_, new_n54284_ );
nor  ( new_n54317_, new_n54316_, new_n54281_ );
nor  ( new_n54318_, new_n54317_, new_n54280_ );
and  ( new_n54319_, new_n54318_, new_n54265_ );
nor  ( new_n54320_, new_n54318_, new_n54265_ );
xnor ( new_n54321_, new_n53783_, new_n53782_ );
or   ( new_n54322_, new_n54015_, new_n340_ );
xor  ( new_n54323_, new_n51446_, RIbb2f250_9 );
nand ( new_n54324_, new_n54323_, new_n336_ );
and  ( new_n54325_, new_n54324_, new_n54322_ );
or   ( new_n54326_, new_n54019_, new_n411_ );
or   ( new_n54327_, new_n54299_, new_n409_ );
and  ( new_n54328_, new_n54327_, new_n54326_ );
or   ( new_n54329_, new_n54328_, new_n54325_ );
nand ( new_n54330_, new_n54328_, new_n54325_ );
xor  ( new_n54331_, new_n53781_, new_n53776_ );
nand ( new_n54332_, new_n54331_, new_n54330_ );
and  ( new_n54333_, new_n54332_, new_n54329_ );
or   ( new_n54334_, new_n54333_, new_n54321_ );
or   ( new_n54335_, new_n54294_, new_n524_ );
or   ( new_n54336_, new_n54031_, new_n526_ );
and  ( new_n54337_, new_n54336_, new_n54335_ );
or   ( new_n54338_, new_n54305_, new_n755_ );
nand ( new_n54339_, new_n54024_, new_n660_ );
and  ( new_n54340_, new_n54339_, new_n54338_ );
nor  ( new_n54341_, new_n54340_, new_n54337_ );
xor  ( new_n54342_, new_n46962_, new_n2118_ );
nor  ( new_n54343_, new_n54342_, new_n2425_ );
nor  ( new_n54344_, new_n54035_, new_n2427_ );
or   ( new_n54345_, new_n54344_, new_n54343_ );
xor  ( new_n54346_, new_n54340_, new_n54337_ );
and  ( new_n54347_, new_n54346_, new_n54345_ );
or   ( new_n54348_, new_n54347_, new_n54341_ );
xor  ( new_n54349_, new_n54333_, new_n54321_ );
nand ( new_n54350_, new_n54349_, new_n54348_ );
and  ( new_n54351_, new_n54350_, new_n54334_ );
or   ( new_n54352_, new_n53913_, new_n9424_ );
xor  ( new_n54353_, new_n43884_, RIbb2dae0_59 );
nand ( new_n54354_, new_n54353_, new_n9187_ );
and  ( new_n54355_, new_n54354_, new_n54352_ );
or   ( new_n54356_, new_n53916_, new_n4711_ );
xor  ( new_n54357_, new_n45119_, new_n4292_ );
or   ( new_n54358_, new_n54357_, new_n4709_ );
and  ( new_n54359_, new_n54358_, new_n54356_ );
or   ( new_n54360_, new_n54359_, new_n54355_ );
xor  ( new_n54361_, new_n43812_, RIbb2ddb0_53 );
and  ( new_n54362_, new_n54361_, new_n7489_ );
and  ( new_n54363_, new_n53932_, new_n7487_ );
nor  ( new_n54364_, new_n54363_, new_n54362_ );
not  ( new_n54365_, new_n54364_ );
xor  ( new_n54366_, new_n54359_, new_n54355_ );
nand ( new_n54367_, new_n54366_, new_n54365_ );
and  ( new_n54368_, new_n54367_, new_n54360_ );
nand ( new_n54369_, new_n53886_, new_n5915_ );
xor  ( new_n54370_, new_n44506_, new_n5594_ );
or   ( new_n54371_, new_n54370_, new_n6173_ );
and  ( new_n54372_, new_n54371_, new_n54369_ );
or   ( new_n54373_, new_n54093_, new_n10061_ );
xor  ( new_n54374_, new_n43799_, new_n9418_ );
or   ( new_n54375_, new_n54374_, new_n10059_ );
and  ( new_n54376_, new_n54375_, new_n54373_ );
or   ( new_n54377_, new_n54376_, new_n54372_ );
and  ( new_n54378_, new_n54376_, new_n54372_ );
xor  ( new_n54379_, new_n43787_, new_n10052_ );
nor  ( new_n54380_, new_n54379_, new_n21077_ );
nor  ( new_n54381_, new_n43898_, new_n10052_ );
and  ( new_n54382_, new_n54381_, new_n21077_ );
nor  ( new_n54383_, new_n54382_, new_n54380_ );
or   ( new_n54384_, new_n54383_, new_n54378_ );
and  ( new_n54385_, new_n54384_, new_n54377_ );
or   ( new_n54386_, new_n54385_, new_n54368_ );
and  ( new_n54387_, new_n54385_, new_n54368_ );
xor  ( new_n54388_, new_n44183_, RIbb2dea0_51 );
nand ( new_n54389_, new_n54388_, new_n6910_ );
or   ( new_n54390_, new_n53949_, new_n7186_ );
and  ( new_n54391_, new_n54390_, new_n54389_ );
nand ( new_n54392_, new_n53938_, new_n4032_ );
xor  ( new_n54393_, new_n45403_, new_n3892_ );
or   ( new_n54394_, new_n54393_, new_n4302_ );
and  ( new_n54395_, new_n54394_, new_n54392_ );
nor  ( new_n54396_, new_n54395_, new_n54391_ );
and  ( new_n54397_, new_n53945_, new_n3731_ );
xor  ( new_n54398_, new_n45738_, RIbb2e530_37 );
and  ( new_n54399_, new_n54398_, new_n3733_ );
nor  ( new_n54400_, new_n54399_, new_n54397_ );
and  ( new_n54401_, new_n54395_, new_n54391_ );
nor  ( new_n54402_, new_n54401_, new_n54400_ );
nor  ( new_n54403_, new_n54402_, new_n54396_ );
or   ( new_n54404_, new_n54403_, new_n54387_ );
and  ( new_n54405_, new_n54404_, new_n54386_ );
nor  ( new_n54406_, new_n54405_, new_n54351_ );
nor  ( new_n54407_, new_n54053_, new_n1595_ );
xor  ( new_n54408_, new_n48039_, RIbb2ebc0_23 );
and  ( new_n54409_, new_n54408_, new_n1476_ );
nor  ( new_n54410_, new_n54409_, new_n54407_ );
xor  ( new_n54411_, new_n47296_, new_n1583_ );
or   ( new_n54412_, new_n54411_, new_n1844_ );
or   ( new_n54413_, new_n54049_, new_n1846_ );
and  ( new_n54414_, new_n54413_, new_n54412_ );
nor  ( new_n54415_, new_n54414_, new_n54410_ );
and  ( new_n54416_, new_n53996_, new_n1251_ );
xor  ( new_n54417_, new_n48518_, RIbb2ecb0_21 );
and  ( new_n54418_, new_n54417_, new_n1253_ );
nor  ( new_n54419_, new_n54418_, new_n54416_ );
and  ( new_n54420_, new_n54414_, new_n54410_ );
nor  ( new_n54421_, new_n54420_, new_n54419_ );
nor  ( new_n54422_, new_n54421_, new_n54415_ );
nor  ( new_n54423_, new_n54069_, new_n286_ );
xor  ( new_n54424_, new_n52902_, RIbb2f430_5 );
nor  ( new_n54425_, new_n54424_, new_n283_ );
or   ( new_n54426_, new_n54425_, new_n54423_ );
and  ( new_n54427_, new_n53694_, new_n43978_ );
nand ( new_n54428_, new_n54427_, new_n54426_ );
nor  ( new_n54429_, new_n54424_, new_n286_ );
xor  ( new_n54430_, new_n52908_, RIbb2f430_5 );
nor  ( new_n54431_, new_n54430_, new_n283_ );
or   ( new_n54432_, new_n54431_, new_n54429_ );
or   ( new_n54433_, new_n53695_, new_n43947_ );
and  ( new_n54434_, new_n54433_, new_n291_ );
and  ( new_n54435_, new_n54434_, new_n43950_ );
and  ( new_n54436_, new_n54435_, new_n54432_ );
xor  ( new_n54437_, new_n54427_, new_n54426_ );
nand ( new_n54438_, new_n54437_, new_n54436_ );
and  ( new_n54439_, new_n54438_, new_n54428_ );
xor  ( new_n54440_, new_n52280_, new_n309_ );
or   ( new_n54441_, new_n54440_, new_n317_ );
or   ( new_n54442_, new_n53773_, new_n320_ );
and  ( new_n54443_, new_n54442_, new_n54441_ );
not  ( new_n54444_, new_n53697_ );
or   ( new_n54445_, new_n54444_, new_n44007_ );
or   ( new_n54446_, new_n54058_, new_n302_ );
and  ( new_n54447_, new_n54446_, new_n54445_ );
or   ( new_n54448_, new_n54447_, new_n54443_ );
and  ( new_n54449_, new_n54323_, new_n334_ );
xor  ( new_n54450_, new_n51477_, RIbb2f250_9 );
and  ( new_n54451_, new_n54450_, new_n336_ );
or   ( new_n54452_, new_n54451_, new_n54449_ );
xor  ( new_n54453_, new_n54447_, new_n54443_ );
nand ( new_n54454_, new_n54453_, new_n54452_ );
and  ( new_n54455_, new_n54454_, new_n54448_ );
or   ( new_n54456_, new_n54455_, new_n54439_ );
xor  ( new_n54457_, new_n47303_, new_n1840_ );
nor  ( new_n54458_, new_n54457_, new_n2122_ );
and  ( new_n54459_, new_n54039_, new_n2000_ );
nor  ( new_n54460_, new_n54459_, new_n54458_ );
not  ( new_n54461_, new_n54460_ );
xor  ( new_n54462_, new_n54455_, new_n54439_ );
nand ( new_n54463_, new_n54462_, new_n54461_ );
and  ( new_n54464_, new_n54463_, new_n54456_ );
nor  ( new_n54465_, new_n54464_, new_n54422_ );
xor  ( new_n54466_, new_n54464_, new_n54422_ );
not  ( new_n54467_, new_n54466_ );
xor  ( new_n54468_, new_n48908_, new_n893_ );
nor  ( new_n54469_, new_n54468_, new_n1135_ );
and  ( new_n54470_, new_n54001_, new_n1040_ );
nor  ( new_n54471_, new_n54470_, new_n54469_ );
nand ( new_n54472_, new_n54006_, new_n2613_ );
xor  ( new_n54473_, new_n46619_, new_n2421_ );
or   ( new_n54474_, new_n54473_, new_n2807_ );
and  ( new_n54475_, new_n54474_, new_n54472_ );
nor  ( new_n54476_, new_n54475_, new_n54471_ );
and  ( new_n54477_, new_n54475_, new_n54471_ );
nor  ( new_n54478_, new_n53894_, new_n899_ );
xor  ( new_n54479_, new_n49427_, RIbb2ee90_17 );
and  ( new_n54480_, new_n54479_, new_n822_ );
nor  ( new_n54481_, new_n54480_, new_n54478_ );
nor  ( new_n54482_, new_n54481_, new_n54477_ );
nor  ( new_n54483_, new_n54482_, new_n54476_ );
nor  ( new_n54484_, new_n54483_, new_n54467_ );
or   ( new_n54485_, new_n54484_, new_n54465_ );
xor  ( new_n54486_, new_n54405_, new_n54351_ );
and  ( new_n54487_, new_n54486_, new_n54485_ );
nor  ( new_n54488_, new_n54487_, new_n54406_ );
nor  ( new_n54489_, new_n54488_, new_n54320_ );
nor  ( new_n54490_, new_n54489_, new_n54319_ );
nor  ( new_n54491_, new_n54490_, new_n54264_ );
xor  ( new_n54492_, new_n54490_, new_n54264_ );
xor  ( new_n54493_, new_n54160_, new_n54159_ );
and  ( new_n54494_, new_n54493_, new_n54492_ );
or   ( new_n54495_, new_n54494_, new_n54491_ );
xor  ( new_n54496_, new_n54125_, new_n54124_ );
xor  ( new_n54497_, new_n54496_, new_n54128_ );
and  ( new_n54498_, new_n54497_, new_n54495_ );
xor  ( new_n54499_, new_n54242_, new_n54241_ );
xor  ( new_n54500_, new_n54497_, new_n54495_ );
and  ( new_n54501_, new_n54500_, new_n54499_ );
nor  ( new_n54502_, new_n54501_, new_n54498_ );
and  ( new_n54503_, new_n54261_, new_n54259_ );
nor  ( new_n54504_, new_n54503_, new_n54502_ );
nor  ( new_n54505_, new_n54504_, new_n54262_ );
not  ( new_n54506_, new_n54505_ );
and  ( new_n54507_, new_n54506_, new_n54258_ );
xor  ( new_n54508_, new_n54483_, new_n54467_ );
not  ( new_n54509_, new_n54508_ );
xnor ( new_n54510_, new_n54475_, new_n54471_ );
and  ( new_n54511_, new_n54510_, new_n54481_ );
not  ( new_n54512_, new_n54476_ );
and  ( new_n54513_, new_n54482_, new_n54512_ );
or   ( new_n54514_, new_n54513_, new_n54511_ );
xor  ( new_n54515_, new_n44974_, RIbb2e260_43 );
and  ( new_n54516_, new_n54515_, new_n4960_ );
and  ( new_n54517_, new_n54177_, new_n4958_ );
nor  ( new_n54518_, new_n54517_, new_n54516_ );
or   ( new_n54519_, new_n54357_, new_n4711_ );
xor  ( new_n54520_, new_n45204_, new_n4292_ );
or   ( new_n54521_, new_n54520_, new_n4709_ );
and  ( new_n54522_, new_n54521_, new_n54519_ );
nor  ( new_n54523_, new_n54522_, new_n54518_ );
and  ( new_n54524_, new_n54522_, new_n54518_ );
xor  ( new_n54525_, new_n43888_, RIbb2dae0_59 );
and  ( new_n54526_, new_n54525_, new_n9187_ );
and  ( new_n54527_, new_n54353_, new_n9185_ );
nor  ( new_n54528_, new_n54527_, new_n54526_ );
nor  ( new_n54529_, new_n54528_, new_n54524_ );
nor  ( new_n54530_, new_n54529_, new_n54523_ );
or   ( new_n54531_, new_n54530_, new_n54514_ );
and  ( new_n54532_, new_n54530_, new_n54514_ );
and  ( new_n54533_, new_n54388_, new_n6908_ );
xor  ( new_n54534_, new_n44218_, RIbb2dea0_51 );
and  ( new_n54535_, new_n54534_, new_n6910_ );
or   ( new_n54536_, new_n54535_, new_n54533_ );
xor  ( new_n54537_, new_n54453_, new_n54452_ );
and  ( new_n54538_, new_n54537_, new_n54536_ );
and  ( new_n54539_, new_n54398_, new_n3731_ );
xor  ( new_n54540_, new_n45597_, RIbb2e530_37 );
and  ( new_n54541_, new_n54540_, new_n3733_ );
or   ( new_n54542_, new_n54541_, new_n54539_ );
xor  ( new_n54543_, new_n54537_, new_n54536_ );
and  ( new_n54544_, new_n54543_, new_n54542_ );
nor  ( new_n54545_, new_n54544_, new_n54538_ );
or   ( new_n54546_, new_n54545_, new_n54532_ );
and  ( new_n54547_, new_n54546_, new_n54531_ );
nor  ( new_n54548_, new_n54547_, new_n54509_ );
xor  ( new_n54549_, new_n54547_, new_n54509_ );
xor  ( new_n54550_, new_n44600_, RIbb2e080_47 );
nand ( new_n54551_, new_n54550_, new_n5917_ );
or   ( new_n54552_, new_n54370_, new_n6175_ );
and  ( new_n54553_, new_n54552_, new_n54551_ );
or   ( new_n54554_, new_n54374_, new_n10061_ );
xor  ( new_n54555_, new_n43803_, RIbb2d9f0_61 );
nand ( new_n54556_, new_n54555_, new_n9740_ );
and  ( new_n54557_, new_n54556_, new_n54554_ );
nor  ( new_n54558_, new_n54557_, new_n54553_ );
and  ( new_n54559_, new_n54208_, new_n8649_ );
xor  ( new_n54560_, new_n43956_, new_n8254_ );
nor  ( new_n54561_, new_n54560_, new_n8874_ );
nor  ( new_n54562_, new_n54561_, new_n54559_ );
and  ( new_n54563_, new_n54557_, new_n54553_ );
nor  ( new_n54564_, new_n54563_, new_n54562_ );
nor  ( new_n54565_, new_n54564_, new_n54558_ );
xor  ( new_n54566_, new_n43985_, new_n7722_ );
or   ( new_n54567_, new_n54566_, new_n8264_ );
or   ( new_n54568_, new_n54174_, new_n8266_ );
and  ( new_n54569_, new_n54568_, new_n54567_ );
xor  ( new_n54570_, new_n44785_, new_n5203_ );
or   ( new_n54571_, new_n54570_, new_n5604_ );
nand ( new_n54572_, new_n54183_, new_n5371_ );
and  ( new_n54573_, new_n54572_, new_n54571_ );
or   ( new_n54574_, new_n54573_, new_n54569_ );
and  ( new_n54575_, new_n54573_, new_n54569_ );
xor  ( new_n54576_, new_n43898_, new_n10052_ );
nor  ( new_n54577_, new_n54576_, new_n21077_ );
and  ( new_n54578_, new_n44104_, RIbb2d900_63 );
and  ( new_n54579_, new_n54578_, new_n21077_ );
nor  ( new_n54580_, new_n54579_, new_n54577_ );
or   ( new_n54581_, new_n54580_, new_n54575_ );
and  ( new_n54582_, new_n54581_, new_n54574_ );
or   ( new_n54583_, new_n54582_, new_n54565_ );
and  ( new_n54584_, new_n54582_, new_n54565_ );
or   ( new_n54585_, new_n54288_, new_n3463_ );
xor  ( new_n54586_, new_n46037_, new_n3113_ );
or   ( new_n54587_, new_n54586_, new_n3461_ );
and  ( new_n54588_, new_n54587_, new_n54585_ );
xor  ( new_n54589_, new_n45584_, RIbb2e440_39 );
nand ( new_n54590_, new_n54589_, new_n4034_ );
or   ( new_n54591_, new_n54393_, new_n4304_ );
and  ( new_n54592_, new_n54591_, new_n54590_ );
nor  ( new_n54593_, new_n54592_, new_n54588_ );
and  ( new_n54594_, new_n54361_, new_n7487_ );
xor  ( new_n54595_, new_n43914_, RIbb2ddb0_53 );
and  ( new_n54596_, new_n54595_, new_n7489_ );
nor  ( new_n54597_, new_n54596_, new_n54594_ );
and  ( new_n54598_, new_n54592_, new_n54588_ );
nor  ( new_n54599_, new_n54598_, new_n54597_ );
nor  ( new_n54600_, new_n54599_, new_n54593_ );
or   ( new_n54601_, new_n54600_, new_n54584_ );
nand ( new_n54602_, new_n54601_, new_n54583_ );
and  ( new_n54603_, new_n54602_, new_n54549_ );
nor  ( new_n54604_, new_n54603_, new_n54548_ );
not  ( new_n54605_, new_n54604_ );
xor  ( new_n54606_, new_n54486_, new_n54485_ );
and  ( new_n54607_, new_n54606_, new_n54605_ );
xor  ( new_n54608_, new_n54606_, new_n54605_ );
xor  ( new_n54609_, new_n54223_, new_n54192_ );
and  ( new_n54610_, new_n54609_, new_n54608_ );
or   ( new_n54611_, new_n54610_, new_n54607_ );
xnor ( new_n54612_, new_n54318_, new_n54265_ );
nand ( new_n54613_, new_n54612_, new_n54488_ );
or   ( new_n54614_, new_n54488_, new_n54320_ );
or   ( new_n54615_, new_n54614_, new_n54319_ );
and  ( new_n54616_, new_n54615_, new_n54613_ );
and  ( new_n54617_, new_n54616_, new_n54611_ );
nor  ( new_n54618_, new_n54616_, new_n54611_ );
not  ( new_n54619_, new_n54618_ );
xor  ( new_n54620_, new_n53967_, new_n53966_ );
not  ( new_n54621_, new_n54620_ );
xor  ( new_n54622_, new_n54076_, new_n54047_ );
xor  ( new_n54623_, new_n53908_, new_n53892_ );
nand ( new_n54624_, new_n54623_, new_n53927_ );
or   ( new_n54625_, new_n53927_, new_n53911_ );
or   ( new_n54626_, new_n54625_, new_n53910_ );
and  ( new_n54627_, new_n54626_, new_n54624_ );
nand ( new_n54628_, new_n54627_, new_n54622_ );
or   ( new_n54629_, new_n54627_, new_n54622_ );
xor  ( new_n54630_, new_n53963_, new_n53961_ );
nand ( new_n54631_, new_n54630_, new_n54629_ );
and  ( new_n54632_, new_n54631_, new_n54628_ );
xor  ( new_n54633_, new_n54632_, new_n54621_ );
not  ( new_n54634_, new_n54633_ );
xor  ( new_n54635_, new_n54149_, new_n54147_ );
xor  ( new_n54636_, new_n54635_, new_n54152_ );
xor  ( new_n54637_, new_n54139_, new_n54134_ );
xor  ( new_n54638_, new_n54637_, new_n54142_ );
nand ( new_n54639_, new_n54638_, new_n54636_ );
nor  ( new_n54640_, new_n54638_, new_n54636_ );
xor  ( new_n54641_, new_n54349_, new_n54348_ );
xor  ( new_n54642_, new_n53941_, new_n53940_ );
and  ( new_n54643_, new_n54642_, new_n54641_ );
nor  ( new_n54644_, new_n54642_, new_n54641_ );
or   ( new_n54645_, new_n54468_, new_n1137_ );
xor  ( new_n54646_, new_n49265_, new_n893_ );
or   ( new_n54647_, new_n54646_, new_n1135_ );
and  ( new_n54648_, new_n54647_, new_n54645_ );
xor  ( new_n54649_, new_n48291_, RIbb2ebc0_23 );
nand ( new_n54650_, new_n54649_, new_n1476_ );
nand ( new_n54651_, new_n54408_, new_n1474_ );
and  ( new_n54652_, new_n54651_, new_n54650_ );
or   ( new_n54653_, new_n54652_, new_n54648_ );
and  ( new_n54654_, new_n54417_, new_n1251_ );
xor  ( new_n54655_, new_n48756_, RIbb2ecb0_21 );
and  ( new_n54656_, new_n54655_, new_n1253_ );
or   ( new_n54657_, new_n54656_, new_n54654_ );
xor  ( new_n54658_, new_n54652_, new_n54648_ );
nand ( new_n54659_, new_n54658_, new_n54657_ );
and  ( new_n54660_, new_n54659_, new_n54653_ );
or   ( new_n54661_, new_n54440_, new_n320_ );
xor  ( new_n54662_, new_n52293_, RIbb2f340_7 );
or   ( new_n54663_, new_n54662_, new_n317_ );
and  ( new_n54664_, new_n54663_, new_n54661_ );
or   ( new_n54665_, new_n54444_, new_n302_ );
nand ( new_n54666_, new_n54062_, new_n43949_ );
and  ( new_n54667_, new_n54666_, new_n54665_ );
or   ( new_n54668_, new_n54667_, new_n54664_ );
and  ( new_n54669_, new_n54450_, new_n334_ );
xor  ( new_n54670_, new_n51758_, new_n329_ );
nor  ( new_n54671_, new_n54670_, new_n337_ );
or   ( new_n54672_, new_n54671_, new_n54669_ );
xor  ( new_n54673_, new_n54667_, new_n54664_ );
nand ( new_n54674_, new_n54673_, new_n54672_ );
and  ( new_n54675_, new_n54674_, new_n54668_ );
or   ( new_n54676_, new_n54411_, new_n1846_ );
xor  ( new_n54677_, new_n47640_, new_n1583_ );
or   ( new_n54678_, new_n54677_, new_n1844_ );
and  ( new_n54679_, new_n54678_, new_n54676_ );
or   ( new_n54680_, new_n54679_, new_n54675_ );
nor  ( new_n54681_, new_n54457_, new_n2124_ );
xor  ( new_n54682_, new_n47046_, new_n1840_ );
nor  ( new_n54683_, new_n54682_, new_n2122_ );
or   ( new_n54684_, new_n54683_, new_n54681_ );
xor  ( new_n54685_, new_n54679_, new_n54675_ );
nand ( new_n54686_, new_n54685_, new_n54684_ );
and  ( new_n54687_, new_n54686_, new_n54680_ );
nor  ( new_n54688_, new_n54687_, new_n54660_ );
and  ( new_n54689_, new_n54687_, new_n54660_ );
xor  ( new_n54690_, new_n46958_, RIbb2e8f0_29 );
nand ( new_n54691_, new_n54690_, new_n2244_ );
or   ( new_n54692_, new_n54342_, new_n2427_ );
and  ( new_n54693_, new_n54692_, new_n54691_ );
xor  ( new_n54694_, new_n46789_, new_n2421_ );
or   ( new_n54695_, new_n54694_, new_n2807_ );
or   ( new_n54696_, new_n54473_, new_n2809_ );
and  ( new_n54697_, new_n54696_, new_n54695_ );
nor  ( new_n54698_, new_n54697_, new_n54693_ );
and  ( new_n54699_, new_n54479_, new_n820_ );
xor  ( new_n54700_, new_n49488_, RIbb2ee90_17 );
and  ( new_n54701_, new_n54700_, new_n822_ );
nor  ( new_n54702_, new_n54701_, new_n54699_ );
and  ( new_n54703_, new_n54697_, new_n54693_ );
nor  ( new_n54704_, new_n54703_, new_n54702_ );
nor  ( new_n54705_, new_n54704_, new_n54698_ );
nor  ( new_n54706_, new_n54705_, new_n54689_ );
nor  ( new_n54707_, new_n54706_, new_n54688_ );
nor  ( new_n54708_, new_n54707_, new_n54644_ );
nor  ( new_n54709_, new_n54708_, new_n54643_ );
or   ( new_n54710_, new_n54709_, new_n54640_ );
and  ( new_n54711_, new_n54710_, new_n54639_ );
xor  ( new_n54712_, new_n54711_, new_n54634_ );
and  ( new_n54713_, new_n54712_, new_n54619_ );
nor  ( new_n54714_, new_n54713_, new_n54617_ );
xor  ( new_n54715_, new_n54346_, new_n54345_ );
xor  ( new_n54716_, new_n54328_, new_n54325_ );
xor  ( new_n54717_, new_n54716_, new_n54331_ );
and  ( new_n54718_, new_n54717_, new_n54715_ );
and  ( new_n54719_, new_n54203_, new_n2928_ );
xor  ( new_n54720_, new_n46427_, RIbb2e710_33 );
and  ( new_n54721_, new_n54720_, new_n2930_ );
or   ( new_n54722_, new_n54721_, new_n54719_ );
xor  ( new_n54723_, new_n54437_, new_n54436_ );
and  ( new_n54724_, new_n54723_, new_n54722_ );
xor  ( new_n54725_, new_n44407_, RIbb2df90_49 );
and  ( new_n54726_, new_n54725_, new_n6510_ );
and  ( new_n54727_, new_n54198_, new_n6508_ );
or   ( new_n54728_, new_n54727_, new_n54726_ );
xor  ( new_n54729_, new_n54723_, new_n54722_ );
and  ( new_n54730_, new_n54729_, new_n54728_ );
or   ( new_n54731_, new_n54730_, new_n54724_ );
xor  ( new_n54732_, new_n54717_, new_n54715_ );
and  ( new_n54733_, new_n54732_, new_n54731_ );
nor  ( new_n54734_, new_n54733_, new_n54718_ );
xnor ( new_n54735_, new_n54385_, new_n54368_ );
xnor ( new_n54736_, new_n54735_, new_n54403_ );
nor  ( new_n54737_, new_n54736_, new_n54734_ );
xnor ( new_n54738_, new_n54736_, new_n54734_ );
xnor ( new_n54739_, new_n54205_, new_n54201_ );
nand ( new_n54740_, new_n54739_, new_n54211_ );
not  ( new_n54741_, new_n54212_ );
or   ( new_n54742_, new_n54741_, new_n54206_ );
and  ( new_n54743_, new_n54742_, new_n54740_ );
xnor ( new_n54744_, new_n54395_, new_n54391_ );
xor  ( new_n54745_, new_n54744_, new_n54400_ );
nand ( new_n54746_, new_n54745_, new_n54743_ );
or   ( new_n54747_, new_n54745_, new_n54743_ );
xor  ( new_n54748_, new_n54376_, new_n54372_ );
xnor ( new_n54749_, new_n54748_, new_n54383_ );
nand ( new_n54750_, new_n54749_, new_n54747_ );
and  ( new_n54751_, new_n54750_, new_n54746_ );
nor  ( new_n54752_, new_n54751_, new_n54738_ );
or   ( new_n54753_, new_n54752_, new_n54737_ );
xor  ( new_n54754_, new_n54279_, new_n54267_ );
xor  ( new_n54755_, new_n54754_, new_n54316_ );
nand ( new_n54756_, new_n54755_, new_n54753_ );
nor  ( new_n54757_, new_n54755_, new_n54753_ );
xnor ( new_n54758_, new_n54170_, new_n54165_ );
xor  ( new_n54759_, new_n54758_, new_n54188_ );
xor  ( new_n54760_, new_n54213_, new_n54197_ );
xor  ( new_n54761_, new_n54760_, new_n54221_ );
and  ( new_n54762_, new_n54761_, new_n54759_ );
nor  ( new_n54763_, new_n54761_, new_n54759_ );
xnor ( new_n54764_, new_n54414_, new_n54410_ );
and  ( new_n54765_, new_n54764_, new_n54419_ );
not  ( new_n54766_, new_n54415_ );
and  ( new_n54767_, new_n54421_, new_n54766_ );
or   ( new_n54768_, new_n54767_, new_n54765_ );
xor  ( new_n54769_, new_n54290_, new_n54286_ );
xor  ( new_n54770_, new_n54769_, new_n54310_ );
nor  ( new_n54771_, new_n54770_, new_n54768_ );
and  ( new_n54772_, new_n54770_, new_n54768_ );
not  ( new_n54773_, new_n54772_ );
xor  ( new_n54774_, new_n54462_, new_n54461_ );
and  ( new_n54775_, new_n54774_, new_n54773_ );
nor  ( new_n54776_, new_n54775_, new_n54771_ );
nor  ( new_n54777_, new_n54776_, new_n54763_ );
nor  ( new_n54778_, new_n54777_, new_n54762_ );
or   ( new_n54779_, new_n54778_, new_n54757_ );
and  ( new_n54780_, new_n54779_, new_n54756_ );
xor  ( new_n54781_, new_n54283_, new_n54282_ );
xor  ( new_n54782_, new_n54781_, new_n54314_ );
xor  ( new_n54783_, new_n54273_, new_n54272_ );
xor  ( new_n54784_, new_n54783_, new_n54277_ );
and  ( new_n54785_, new_n54784_, new_n54782_ );
or   ( new_n54786_, new_n54784_, new_n54782_ );
xor  ( new_n54787_, new_n54366_, new_n54365_ );
or   ( new_n54788_, new_n54297_, new_n411_ );
xor  ( new_n54789_, new_n51446_, RIbb2f160_11 );
nand ( new_n54790_, new_n54789_, new_n373_ );
and  ( new_n54791_, new_n54790_, new_n54788_ );
or   ( new_n54792_, new_n54303_, new_n757_ );
xor  ( new_n54793_, new_n50487_, new_n520_ );
or   ( new_n54794_, new_n54793_, new_n755_ );
and  ( new_n54795_, new_n54794_, new_n54792_ );
nor  ( new_n54796_, new_n54795_, new_n54791_ );
xor  ( new_n54797_, new_n49758_, new_n745_ );
nor  ( new_n54798_, new_n54797_, new_n897_ );
and  ( new_n54799_, new_n54700_, new_n820_ );
or   ( new_n54800_, new_n54799_, new_n54798_ );
xor  ( new_n54801_, new_n54795_, new_n54791_ );
and  ( new_n54802_, new_n54801_, new_n54800_ );
nor  ( new_n54803_, new_n54802_, new_n54796_ );
nor  ( new_n54804_, new_n54430_, new_n286_ );
xor  ( new_n54805_, new_n53306_, RIbb2f430_5 );
nor  ( new_n54806_, new_n54805_, new_n283_ );
or   ( new_n54807_, new_n54806_, new_n54804_ );
and  ( new_n54808_, new_n53694_, new_n295_ );
and  ( new_n54809_, new_n54808_, new_n54807_ );
xor  ( new_n54810_, new_n52902_, RIbb2f340_7 );
nor  ( new_n54811_, new_n54810_, new_n317_ );
nor  ( new_n54812_, new_n54662_, new_n320_ );
or   ( new_n54813_, new_n54812_, new_n54811_ );
xor  ( new_n54814_, new_n54808_, new_n54807_ );
and  ( new_n54815_, new_n54814_, new_n54813_ );
or   ( new_n54816_, new_n54815_, new_n54809_ );
xor  ( new_n54817_, new_n54435_, new_n54432_ );
and  ( new_n54818_, new_n54817_, new_n54816_ );
xor  ( new_n54819_, new_n50894_, new_n400_ );
nor  ( new_n54820_, new_n54819_, new_n524_ );
nor  ( new_n54821_, new_n54292_, new_n526_ );
or   ( new_n54822_, new_n54821_, new_n54820_ );
xor  ( new_n54823_, new_n54817_, new_n54816_ );
and  ( new_n54824_, new_n54823_, new_n54822_ );
or   ( new_n54825_, new_n54824_, new_n54818_ );
xnor ( new_n54826_, new_n54301_, new_n54296_ );
nand ( new_n54827_, new_n54826_, new_n54307_ );
not  ( new_n54828_, new_n54309_ );
or   ( new_n54829_, new_n54828_, new_n54302_ );
and  ( new_n54830_, new_n54829_, new_n54827_ );
nand ( new_n54831_, new_n54830_, new_n54825_ );
nand ( new_n54832_, new_n54831_, new_n54803_ );
or   ( new_n54833_, new_n54830_, new_n54825_ );
and  ( new_n54834_, new_n54833_, new_n54832_ );
and  ( new_n54835_, new_n54834_, new_n54787_ );
xor  ( new_n54836_, new_n54834_, new_n54787_ );
xor  ( new_n54837_, new_n54186_, new_n54185_ );
and  ( new_n54838_, new_n54837_, new_n54836_ );
or   ( new_n54839_, new_n54838_, new_n54835_ );
and  ( new_n54840_, new_n54839_, new_n54786_ );
or   ( new_n54841_, new_n54840_, new_n54785_ );
xor  ( new_n54842_, new_n54627_, new_n54622_ );
xor  ( new_n54843_, new_n54842_, new_n54630_ );
nand ( new_n54844_, new_n54843_, new_n54841_ );
or   ( new_n54845_, new_n54843_, new_n54841_ );
xor  ( new_n54846_, new_n54638_, new_n54636_ );
xnor ( new_n54847_, new_n54846_, new_n54709_ );
nand ( new_n54848_, new_n54847_, new_n54845_ );
and  ( new_n54849_, new_n54848_, new_n54844_ );
or   ( new_n54850_, new_n54849_, new_n54780_ );
and  ( new_n54851_, new_n54849_, new_n54780_ );
xor  ( new_n54852_, new_n54119_, new_n54118_ );
xor  ( new_n54853_, new_n54145_, new_n54144_ );
xor  ( new_n54854_, new_n54853_, new_n54154_ );
xor  ( new_n54855_, new_n54854_, new_n54852_ );
xnor ( new_n54856_, new_n54227_, new_n54225_ );
xor  ( new_n54857_, new_n54856_, new_n54231_ );
xnor ( new_n54858_, new_n54857_, new_n54855_ );
or   ( new_n54859_, new_n54858_, new_n54851_ );
and  ( new_n54860_, new_n54859_, new_n54850_ );
xor  ( new_n54861_, new_n54860_, new_n54714_ );
xor  ( new_n54862_, new_n54493_, new_n54492_ );
xor  ( new_n54863_, new_n54862_, new_n54861_ );
xor  ( new_n54864_, new_n54732_, new_n54731_ );
xor  ( new_n54865_, new_n48039_, new_n1583_ );
or   ( new_n54866_, new_n54865_, new_n1844_ );
or   ( new_n54867_, new_n54677_, new_n1846_ );
and  ( new_n54868_, new_n54867_, new_n54866_ );
or   ( new_n54869_, new_n54682_, new_n2124_ );
xor  ( new_n54870_, new_n47296_, RIbb2e9e0_27 );
nand ( new_n54871_, new_n54870_, new_n2002_ );
and  ( new_n54872_, new_n54871_, new_n54869_ );
or   ( new_n54873_, new_n54872_, new_n54868_ );
and  ( new_n54874_, new_n54649_, new_n1474_ );
xor  ( new_n54875_, new_n48518_, RIbb2ebc0_23 );
and  ( new_n54876_, new_n54875_, new_n1476_ );
or   ( new_n54877_, new_n54876_, new_n54874_ );
xor  ( new_n54878_, new_n54872_, new_n54868_ );
nand ( new_n54879_, new_n54878_, new_n54877_ );
and  ( new_n54880_, new_n54879_, new_n54873_ );
nand ( new_n54881_, new_n54655_, new_n1251_ );
xor  ( new_n54882_, new_n48908_, new_n1126_ );
or   ( new_n54883_, new_n54882_, new_n1364_ );
and  ( new_n54884_, new_n54883_, new_n54881_ );
xor  ( new_n54885_, new_n46619_, new_n2797_ );
or   ( new_n54886_, new_n54885_, new_n3117_ );
nand ( new_n54887_, new_n54720_, new_n2928_ );
and  ( new_n54888_, new_n54887_, new_n54886_ );
nor  ( new_n54889_, new_n54888_, new_n54884_ );
and  ( new_n54890_, new_n54888_, new_n54884_ );
nor  ( new_n54891_, new_n54646_, new_n1137_ );
xor  ( new_n54892_, new_n49427_, RIbb2eda0_19 );
and  ( new_n54893_, new_n54892_, new_n1042_ );
nor  ( new_n54894_, new_n54893_, new_n54891_ );
nor  ( new_n54895_, new_n54894_, new_n54890_ );
nor  ( new_n54896_, new_n54895_, new_n54889_ );
nand ( new_n54897_, new_n54896_, new_n54880_ );
nor  ( new_n54898_, new_n54896_, new_n54880_ );
xor  ( new_n54899_, new_n46962_, new_n2421_ );
nor  ( new_n54900_, new_n54899_, new_n2807_ );
nor  ( new_n54901_, new_n54694_, new_n2809_ );
or   ( new_n54902_, new_n54901_, new_n54900_ );
or   ( new_n54903_, RIbb2f3b8_6, RIbb2f340_7 );
and  ( new_n54904_, new_n53694_, new_n54903_ );
or   ( new_n54905_, new_n54904_, new_n278_ );
or   ( new_n54906_, new_n54805_, new_n286_ );
nor  ( new_n54907_, RIbb2f3b8_6, new_n275_ );
and  ( new_n54908_, new_n53694_, RIbb2f340_7 );
nor  ( new_n54909_, new_n54908_, new_n54907_ );
and  ( new_n54910_, RIbb2f3b8_6, new_n275_ );
nor  ( new_n54911_, new_n53694_, RIbb2f340_7 );
nor  ( new_n54912_, new_n54911_, new_n54910_ );
or   ( new_n54913_, new_n54912_, new_n54909_ );
and  ( new_n54914_, new_n54913_, new_n54906_ );
or   ( new_n54915_, new_n54914_, new_n54905_ );
xor  ( new_n54916_, new_n52280_, new_n329_ );
or   ( new_n54917_, new_n54916_, new_n337_ );
or   ( new_n54918_, new_n54670_, new_n340_ );
and  ( new_n54919_, new_n54918_, new_n54917_ );
nand ( new_n54920_, new_n54919_, new_n54915_ );
or   ( new_n54921_, new_n54919_, new_n54915_ );
and  ( new_n54922_, new_n54789_, new_n371_ );
xor  ( new_n54923_, new_n51477_, RIbb2f160_11 );
and  ( new_n54924_, new_n54923_, new_n373_ );
nor  ( new_n54925_, new_n54924_, new_n54922_ );
nand ( new_n54926_, new_n54925_, new_n54921_ );
and  ( new_n54927_, new_n54926_, new_n54920_ );
nor  ( new_n54928_, new_n54927_, new_n54902_ );
xor  ( new_n54929_, new_n47303_, new_n2118_ );
nor  ( new_n54930_, new_n54929_, new_n2425_ );
and  ( new_n54931_, new_n54690_, new_n2242_ );
nor  ( new_n54932_, new_n54931_, new_n54930_ );
xor  ( new_n54933_, new_n54927_, new_n54902_ );
and  ( new_n54934_, new_n54933_, new_n54932_ );
nor  ( new_n54935_, new_n54934_, new_n54928_ );
or   ( new_n54936_, new_n54935_, new_n54898_ );
and  ( new_n54937_, new_n54936_, new_n54897_ );
and  ( new_n54938_, new_n54937_, new_n54864_ );
nand ( new_n54939_, new_n54540_, new_n3731_ );
xor  ( new_n54940_, new_n45928_, new_n3457_ );
or   ( new_n54941_, new_n54940_, new_n3896_ );
and  ( new_n54942_, new_n54941_, new_n54939_ );
xor  ( new_n54943_, new_n44319_, new_n6635_ );
or   ( new_n54944_, new_n54943_, new_n7184_ );
nand ( new_n54945_, new_n54534_, new_n6908_ );
and  ( new_n54946_, new_n54945_, new_n54944_ );
nor  ( new_n54947_, new_n54946_, new_n54942_ );
and  ( new_n54948_, new_n54589_, new_n4032_ );
xor  ( new_n54949_, new_n45738_, RIbb2e440_39 );
and  ( new_n54950_, new_n54949_, new_n4034_ );
or   ( new_n54951_, new_n54950_, new_n54948_ );
xor  ( new_n54952_, new_n54946_, new_n54942_ );
and  ( new_n54953_, new_n54952_, new_n54951_ );
nor  ( new_n54954_, new_n54953_, new_n54947_ );
not  ( new_n54955_, new_n54954_ );
xor  ( new_n54956_, new_n54658_, new_n54657_ );
and  ( new_n54957_, new_n54956_, new_n54955_ );
xor  ( new_n54958_, new_n54956_, new_n54955_ );
xor  ( new_n54959_, new_n54729_, new_n54728_ );
and  ( new_n54960_, new_n54959_, new_n54958_ );
nor  ( new_n54961_, new_n54960_, new_n54957_ );
xnor ( new_n54962_, new_n54937_, new_n54864_ );
nor  ( new_n54963_, new_n54962_, new_n54961_ );
or   ( new_n54964_, new_n54963_, new_n54938_ );
xnor ( new_n54965_, new_n54642_, new_n54641_ );
xor  ( new_n54966_, new_n54965_, new_n54707_ );
nand ( new_n54967_, new_n54966_, new_n54964_ );
nor  ( new_n54968_, new_n54966_, new_n54964_ );
or   ( new_n54969_, new_n54520_, new_n4711_ );
xor  ( new_n54970_, new_n45403_, new_n4292_ );
or   ( new_n54971_, new_n54970_, new_n4709_ );
and  ( new_n54972_, new_n54971_, new_n54969_ );
xor  ( new_n54973_, new_n44183_, new_n7174_ );
or   ( new_n54974_, new_n54973_, new_n7732_ );
nand ( new_n54975_, new_n54595_, new_n7487_ );
and  ( new_n54976_, new_n54975_, new_n54974_ );
nor  ( new_n54977_, new_n54976_, new_n54972_ );
xor  ( new_n54978_, new_n43937_, RIbb2dae0_59 );
and  ( new_n54979_, new_n54978_, new_n9187_ );
and  ( new_n54980_, new_n54525_, new_n9185_ );
nor  ( new_n54981_, new_n54980_, new_n54979_ );
and  ( new_n54982_, new_n54976_, new_n54972_ );
nor  ( new_n54983_, new_n54982_, new_n54981_ );
or   ( new_n54984_, new_n54983_, new_n54977_ );
xnor ( new_n54985_, new_n54697_, new_n54693_ );
xor  ( new_n54986_, new_n54985_, new_n54702_ );
and  ( new_n54987_, new_n54986_, new_n54984_ );
or   ( new_n54988_, new_n54986_, new_n54984_ );
xor  ( new_n54989_, new_n54685_, new_n54684_ );
and  ( new_n54990_, new_n54989_, new_n54988_ );
or   ( new_n54991_, new_n54990_, new_n54987_ );
xnor ( new_n54992_, new_n54687_, new_n54660_ );
xor  ( new_n54993_, new_n54992_, new_n54705_ );
and  ( new_n54994_, new_n54993_, new_n54991_ );
or   ( new_n54995_, new_n54560_, new_n8876_ );
xor  ( new_n54996_, new_n43952_, new_n8254_ );
or   ( new_n54997_, new_n54996_, new_n8874_ );
and  ( new_n54998_, new_n54997_, new_n54995_ );
xor  ( new_n54999_, new_n43894_, new_n10052_ );
or   ( new_n55000_, new_n54999_, new_n21077_ );
or   ( new_n55001_, new_n43799_, new_n10052_ );
or   ( new_n55002_, new_n55001_, RIbb2d888_64 );
and  ( new_n55003_, new_n55002_, new_n55000_ );
nor  ( new_n55004_, new_n55003_, new_n54998_ );
xor  ( new_n55005_, new_n44681_, RIbb2e080_47 );
and  ( new_n55006_, new_n55005_, new_n5917_ );
and  ( new_n55007_, new_n54550_, new_n5915_ );
or   ( new_n55008_, new_n55007_, new_n55006_ );
xor  ( new_n55009_, new_n55003_, new_n54998_ );
and  ( new_n55010_, new_n55009_, new_n55008_ );
nor  ( new_n55011_, new_n55010_, new_n55004_ );
xor  ( new_n55012_, new_n43884_, RIbb2d9f0_61 );
and  ( new_n55013_, new_n55012_, new_n9740_ );
and  ( new_n55014_, new_n54555_, new_n9738_ );
or   ( new_n55015_, new_n55014_, new_n55013_ );
xor  ( new_n55016_, new_n54673_, new_n54672_ );
nand ( new_n55017_, new_n55016_, new_n55015_ );
xor  ( new_n55018_, new_n44506_, RIbb2df90_49 );
and  ( new_n55019_, new_n55018_, new_n6510_ );
and  ( new_n55020_, new_n54725_, new_n6508_ );
nor  ( new_n55021_, new_n55020_, new_n55019_ );
xnor ( new_n55022_, new_n55016_, new_n55015_ );
or   ( new_n55023_, new_n55022_, new_n55021_ );
and  ( new_n55024_, new_n55023_, new_n55017_ );
nor  ( new_n55025_, new_n55024_, new_n55011_ );
xor  ( new_n55026_, new_n55024_, new_n55011_ );
not  ( new_n55027_, new_n55026_ );
or   ( new_n55028_, new_n54566_, new_n8266_ );
xor  ( new_n55029_, new_n43812_, new_n7722_ );
or   ( new_n55030_, new_n55029_, new_n8264_ );
and  ( new_n55031_, new_n55030_, new_n55028_ );
xor  ( new_n55032_, new_n44877_, RIbb2e170_45 );
nand ( new_n55033_, new_n55032_, new_n5373_ );
or   ( new_n55034_, new_n54570_, new_n5606_ );
and  ( new_n55035_, new_n55034_, new_n55033_ );
nor  ( new_n55036_, new_n55035_, new_n55031_ );
and  ( new_n55037_, new_n55035_, new_n55031_ );
xor  ( new_n55038_, new_n45119_, new_n4705_ );
nor  ( new_n55039_, new_n55038_, new_n5207_ );
and  ( new_n55040_, new_n54515_, new_n4958_ );
nor  ( new_n55041_, new_n55040_, new_n55039_ );
nor  ( new_n55042_, new_n55041_, new_n55037_ );
nor  ( new_n55043_, new_n55042_, new_n55036_ );
nor  ( new_n55044_, new_n55043_, new_n55027_ );
nor  ( new_n55045_, new_n55044_, new_n55025_ );
not  ( new_n55046_, new_n55045_ );
xor  ( new_n55047_, new_n54993_, new_n54991_ );
and  ( new_n55048_, new_n55047_, new_n55046_ );
nor  ( new_n55049_, new_n55048_, new_n54994_ );
or   ( new_n55050_, new_n55049_, new_n54968_ );
and  ( new_n55051_, new_n55050_, new_n54967_ );
xnor ( new_n55052_, new_n54602_, new_n54549_ );
xnor ( new_n55053_, new_n54557_, new_n54553_ );
nand ( new_n55054_, new_n55053_, new_n54562_ );
not  ( new_n55055_, new_n54564_ );
or   ( new_n55056_, new_n55055_, new_n54558_ );
and  ( new_n55057_, new_n55056_, new_n55054_ );
xnor ( new_n55058_, new_n54573_, new_n54569_ );
xor  ( new_n55059_, new_n55058_, new_n54580_ );
or   ( new_n55060_, new_n55059_, new_n55057_ );
and  ( new_n55061_, new_n55059_, new_n55057_ );
xor  ( new_n55062_, new_n54522_, new_n54518_ );
not  ( new_n55063_, new_n55062_ );
and  ( new_n55064_, new_n55063_, new_n54528_ );
not  ( new_n55065_, new_n54523_ );
and  ( new_n55066_, new_n54529_, new_n55065_ );
nor  ( new_n55067_, new_n55066_, new_n55064_ );
or   ( new_n55068_, new_n55067_, new_n55061_ );
and  ( new_n55069_, new_n55068_, new_n55060_ );
xnor ( new_n55070_, new_n54530_, new_n54514_ );
xor  ( new_n55071_, new_n55070_, new_n54545_ );
nand ( new_n55072_, new_n55071_, new_n55069_ );
or   ( new_n55073_, new_n55071_, new_n55069_ );
xor  ( new_n55074_, new_n54837_, new_n54836_ );
nand ( new_n55075_, new_n55074_, new_n55073_ );
and  ( new_n55076_, new_n55075_, new_n55072_ );
or   ( new_n55077_, new_n55076_, new_n55052_ );
nand ( new_n55078_, new_n55076_, new_n55052_ );
xnor ( new_n55079_, new_n54582_, new_n54565_ );
xor  ( new_n55080_, new_n55079_, new_n54600_ );
xor  ( new_n55081_, new_n54770_, new_n54768_ );
xor  ( new_n55082_, new_n55081_, new_n54774_ );
nor  ( new_n55083_, new_n55082_, new_n55080_ );
and  ( new_n55084_, new_n55082_, new_n55080_ );
xor  ( new_n55085_, new_n50788_, new_n520_ );
nor  ( new_n55086_, new_n55085_, new_n755_ );
nor  ( new_n55087_, new_n54793_, new_n757_ );
or   ( new_n55088_, new_n55087_, new_n55086_ );
xor  ( new_n55089_, new_n54814_, new_n54813_ );
and  ( new_n55090_, new_n55089_, new_n55088_ );
nor  ( new_n55091_, new_n54797_, new_n899_ );
xor  ( new_n55092_, new_n50115_, new_n745_ );
nor  ( new_n55093_, new_n55092_, new_n897_ );
or   ( new_n55094_, new_n55093_, new_n55091_ );
xor  ( new_n55095_, new_n55089_, new_n55088_ );
and  ( new_n55096_, new_n55095_, new_n55094_ );
or   ( new_n55097_, new_n55096_, new_n55090_ );
xor  ( new_n55098_, new_n54823_, new_n54822_ );
and  ( new_n55099_, new_n55098_, new_n55097_ );
nor  ( new_n55100_, new_n54586_, new_n3463_ );
xor  ( new_n55101_, new_n46137_, RIbb2e620_35 );
and  ( new_n55102_, new_n55101_, new_n3293_ );
nor  ( new_n55103_, new_n55102_, new_n55100_ );
xnor ( new_n55104_, new_n55098_, new_n55097_ );
nor  ( new_n55105_, new_n55104_, new_n55103_ );
or   ( new_n55106_, new_n55105_, new_n55099_ );
xor  ( new_n55107_, new_n54543_, new_n54542_ );
and  ( new_n55108_, new_n55107_, new_n55106_ );
xor  ( new_n55109_, new_n55107_, new_n55106_ );
xnor ( new_n55110_, new_n54592_, new_n54588_ );
xor  ( new_n55111_, new_n55110_, new_n54597_ );
and  ( new_n55112_, new_n55111_, new_n55109_ );
nor  ( new_n55113_, new_n55112_, new_n55108_ );
not  ( new_n55114_, new_n55113_ );
nor  ( new_n55115_, new_n55114_, new_n55084_ );
nor  ( new_n55116_, new_n55115_, new_n55083_ );
nand ( new_n55117_, new_n55116_, new_n55078_ );
and  ( new_n55118_, new_n55117_, new_n55077_ );
nor  ( new_n55119_, new_n55118_, new_n55051_ );
xor  ( new_n55120_, new_n54609_, new_n54608_ );
xor  ( new_n55121_, new_n55118_, new_n55051_ );
and  ( new_n55122_, new_n55121_, new_n55120_ );
or   ( new_n55123_, new_n55122_, new_n55119_ );
xor  ( new_n55124_, new_n54616_, new_n54611_ );
xor  ( new_n55125_, new_n55124_, new_n54712_ );
and  ( new_n55126_, new_n55125_, new_n55123_ );
xor  ( new_n55127_, new_n54751_, new_n54738_ );
xnor ( new_n55128_, new_n54761_, new_n54759_ );
xor  ( new_n55129_, new_n55128_, new_n54776_ );
or   ( new_n55130_, new_n55129_, new_n55127_ );
nand ( new_n55131_, new_n55129_, new_n55127_ );
xor  ( new_n55132_, new_n46789_, new_n2797_ );
or   ( new_n55133_, new_n55132_, new_n3117_ );
or   ( new_n55134_, new_n54885_, new_n3119_ );
and  ( new_n55135_, new_n55134_, new_n55133_ );
xor  ( new_n55136_, new_n48756_, new_n1355_ );
or   ( new_n55137_, new_n55136_, new_n1593_ );
nand ( new_n55138_, new_n54875_, new_n1474_ );
and  ( new_n55139_, new_n55138_, new_n55137_ );
nor  ( new_n55140_, new_n55139_, new_n55135_ );
xor  ( new_n55141_, new_n47640_, new_n1840_ );
nor  ( new_n55142_, new_n55141_, new_n2122_ );
and  ( new_n55143_, new_n54870_, new_n2000_ );
or   ( new_n55144_, new_n55143_, new_n55142_ );
xor  ( new_n55145_, new_n55139_, new_n55135_ );
and  ( new_n55146_, new_n55145_, new_n55144_ );
nor  ( new_n55147_, new_n55146_, new_n55140_ );
not  ( new_n55148_, new_n55147_ );
or   ( new_n55149_, new_n54819_, new_n526_ );
xor  ( new_n55150_, new_n51142_, new_n400_ );
or   ( new_n55151_, new_n55150_, new_n524_ );
and  ( new_n55152_, new_n55151_, new_n55149_ );
nand ( new_n55153_, new_n54892_, new_n1040_ );
xor  ( new_n55154_, new_n49488_, RIbb2eda0_19 );
nand ( new_n55155_, new_n55154_, new_n1042_ );
and  ( new_n55156_, new_n55155_, new_n55153_ );
nor  ( new_n55157_, new_n55156_, new_n55152_ );
and  ( new_n55158_, new_n55101_, new_n3291_ );
xor  ( new_n55159_, new_n46427_, RIbb2e620_35 );
and  ( new_n55160_, new_n55159_, new_n3293_ );
or   ( new_n55161_, new_n55160_, new_n55158_ );
xor  ( new_n55162_, new_n55156_, new_n55152_ );
and  ( new_n55163_, new_n55162_, new_n55161_ );
nor  ( new_n55164_, new_n55163_, new_n55157_ );
not  ( new_n55165_, new_n55164_ );
and  ( new_n55166_, new_n55165_, new_n55148_ );
nor  ( new_n55167_, new_n54810_, new_n320_ );
xor  ( new_n55168_, new_n52908_, RIbb2f340_7 );
nor  ( new_n55169_, new_n55168_, new_n317_ );
or   ( new_n55170_, new_n55169_, new_n55167_ );
xor  ( new_n55171_, new_n54914_, new_n54905_ );
nand ( new_n55172_, new_n55171_, new_n55170_ );
xor  ( new_n55173_, new_n51758_, new_n325_ );
nor  ( new_n55174_, new_n55173_, new_n409_ );
and  ( new_n55175_, new_n54923_, new_n371_ );
or   ( new_n55176_, new_n55175_, new_n55174_ );
xor  ( new_n55177_, new_n55171_, new_n55170_ );
nand ( new_n55178_, new_n55177_, new_n55176_ );
and  ( new_n55179_, new_n55178_, new_n55172_ );
xor  ( new_n55180_, new_n46958_, new_n2421_ );
or   ( new_n55181_, new_n55180_, new_n2807_ );
or   ( new_n55182_, new_n54899_, new_n2809_ );
and  ( new_n55183_, new_n55182_, new_n55181_ );
nor  ( new_n55184_, new_n55183_, new_n55179_ );
xor  ( new_n55185_, new_n47046_, new_n2118_ );
nor  ( new_n55186_, new_n55185_, new_n2425_ );
nor  ( new_n55187_, new_n54929_, new_n2427_ );
or   ( new_n55188_, new_n55187_, new_n55186_ );
xor  ( new_n55189_, new_n55183_, new_n55179_ );
and  ( new_n55190_, new_n55189_, new_n55188_ );
nor  ( new_n55191_, new_n55190_, new_n55184_ );
and  ( new_n55192_, new_n55164_, new_n55147_ );
nor  ( new_n55193_, new_n55192_, new_n55191_ );
nor  ( new_n55194_, new_n55193_, new_n55166_ );
xor  ( new_n55195_, new_n54830_, new_n54825_ );
xor  ( new_n55196_, new_n55195_, new_n54803_ );
nor  ( new_n55197_, new_n55196_, new_n55194_ );
xor  ( new_n55198_, new_n54801_, new_n54800_ );
xor  ( new_n55199_, new_n54878_, new_n54877_ );
and  ( new_n55200_, new_n55199_, new_n55198_ );
xor  ( new_n55201_, new_n46037_, new_n3457_ );
or   ( new_n55202_, new_n55201_, new_n3896_ );
or   ( new_n55203_, new_n54940_, new_n3898_ );
and  ( new_n55204_, new_n55203_, new_n55202_ );
xor  ( new_n55205_, new_n54919_, new_n54915_ );
xor  ( new_n55206_, new_n55205_, new_n54925_ );
nor  ( new_n55207_, new_n55206_, new_n55204_ );
xor  ( new_n55208_, new_n45597_, RIbb2e440_39 );
and  ( new_n55209_, new_n55208_, new_n4034_ );
and  ( new_n55210_, new_n54949_, new_n4032_ );
or   ( new_n55211_, new_n55210_, new_n55209_ );
xor  ( new_n55212_, new_n55206_, new_n55204_ );
and  ( new_n55213_, new_n55212_, new_n55211_ );
or   ( new_n55214_, new_n55213_, new_n55207_ );
xor  ( new_n55215_, new_n55199_, new_n55198_ );
and  ( new_n55216_, new_n55215_, new_n55214_ );
or   ( new_n55217_, new_n55216_, new_n55200_ );
xor  ( new_n55218_, new_n55196_, new_n55194_ );
and  ( new_n55219_, new_n55218_, new_n55217_ );
or   ( new_n55220_, new_n55219_, new_n55197_ );
xor  ( new_n55221_, new_n54745_, new_n54743_ );
xor  ( new_n55222_, new_n55221_, new_n54749_ );
and  ( new_n55223_, new_n55222_, new_n55220_ );
xnor ( new_n55224_, new_n54896_, new_n54880_ );
xor  ( new_n55225_, new_n55224_, new_n54935_ );
xor  ( new_n55226_, new_n49265_, new_n1126_ );
or   ( new_n55227_, new_n55226_, new_n1364_ );
or   ( new_n55228_, new_n54882_, new_n1366_ );
and  ( new_n55229_, new_n55228_, new_n55227_ );
xor  ( new_n55230_, new_n48291_, RIbb2ead0_25 );
nand ( new_n55231_, new_n55230_, new_n1741_ );
or   ( new_n55232_, new_n54865_, new_n1846_ );
and  ( new_n55233_, new_n55232_, new_n55231_ );
nor  ( new_n55234_, new_n55233_, new_n55229_ );
xor  ( new_n55235_, new_n44600_, RIbb2df90_49 );
and  ( new_n55236_, new_n55235_, new_n6510_ );
and  ( new_n55237_, new_n55018_, new_n6508_ );
or   ( new_n55238_, new_n55237_, new_n55236_ );
nand ( new_n55239_, new_n55233_, new_n55229_ );
and  ( new_n55240_, new_n55239_, new_n55238_ );
or   ( new_n55241_, new_n55240_, new_n55234_ );
xnor ( new_n55242_, new_n54888_, new_n54884_ );
nand ( new_n55243_, new_n55242_, new_n54894_ );
not  ( new_n55244_, new_n54895_ );
or   ( new_n55245_, new_n55244_, new_n54889_ );
and  ( new_n55246_, new_n55245_, new_n55243_ );
nand ( new_n55247_, new_n55246_, new_n55241_ );
nor  ( new_n55248_, new_n55246_, new_n55241_ );
xor  ( new_n55249_, new_n54933_, new_n54932_ );
or   ( new_n55250_, new_n55249_, new_n55248_ );
and  ( new_n55251_, new_n55250_, new_n55247_ );
nor  ( new_n55252_, new_n55251_, new_n55225_ );
xor  ( new_n55253_, new_n43985_, new_n8254_ );
or   ( new_n55254_, new_n55253_, new_n8874_ );
or   ( new_n55255_, new_n54996_, new_n8876_ );
and  ( new_n55256_, new_n55255_, new_n55254_ );
nand ( new_n55257_, new_n55012_, new_n9738_ );
xor  ( new_n55258_, new_n43888_, RIbb2d9f0_61 );
nand ( new_n55259_, new_n55258_, new_n9740_ );
and  ( new_n55260_, new_n55259_, new_n55257_ );
or   ( new_n55261_, new_n55260_, new_n55256_ );
xor  ( new_n55262_, new_n44785_, RIbb2e080_47 );
and  ( new_n55263_, new_n55262_, new_n5917_ );
and  ( new_n55264_, new_n55005_, new_n5915_ );
or   ( new_n55265_, new_n55264_, new_n55263_ );
xor  ( new_n55266_, new_n55260_, new_n55256_ );
nand ( new_n55267_, new_n55266_, new_n55265_ );
and  ( new_n55268_, new_n55267_, new_n55261_ );
xor  ( new_n55269_, new_n43914_, RIbb2dcc0_55 );
nand ( new_n55270_, new_n55269_, new_n8042_ );
or   ( new_n55271_, new_n55029_, new_n8266_ );
and  ( new_n55272_, new_n55271_, new_n55270_ );
xor  ( new_n55273_, new_n45204_, new_n4705_ );
or   ( new_n55274_, new_n55273_, new_n5207_ );
or   ( new_n55275_, new_n55038_, new_n5209_ );
and  ( new_n55276_, new_n55275_, new_n55274_ );
nor  ( new_n55277_, new_n55276_, new_n55272_ );
and  ( new_n55278_, new_n55276_, new_n55272_ );
and  ( new_n55279_, new_n55032_, new_n5371_ );
xor  ( new_n55280_, new_n44974_, RIbb2e170_45 );
and  ( new_n55281_, new_n55280_, new_n5373_ );
nor  ( new_n55282_, new_n55281_, new_n55279_ );
nor  ( new_n55283_, new_n55282_, new_n55278_ );
nor  ( new_n55284_, new_n55283_, new_n55277_ );
nor  ( new_n55285_, new_n55284_, new_n55268_ );
xor  ( new_n55286_, new_n44218_, new_n7174_ );
or   ( new_n55287_, new_n55286_, new_n7732_ );
or   ( new_n55288_, new_n54973_, new_n7734_ );
and  ( new_n55289_, new_n55288_, new_n55287_ );
xor  ( new_n55290_, new_n43799_, new_n10052_ );
or   ( new_n55291_, new_n55290_, new_n21077_ );
or   ( new_n55292_, new_n43803_, new_n10052_ );
or   ( new_n55293_, new_n55292_, RIbb2d888_64 );
and  ( new_n55294_, new_n55293_, new_n55291_ );
nor  ( new_n55295_, new_n55294_, new_n55289_ );
xor  ( new_n55296_, new_n45584_, RIbb2e350_41 );
and  ( new_n55297_, new_n55296_, new_n4543_ );
nor  ( new_n55298_, new_n54970_, new_n4711_ );
nor  ( new_n55299_, new_n55298_, new_n55297_ );
not  ( new_n55300_, new_n55299_ );
xor  ( new_n55301_, new_n55294_, new_n55289_ );
and  ( new_n55302_, new_n55301_, new_n55300_ );
nor  ( new_n55303_, new_n55302_, new_n55295_ );
not  ( new_n55304_, new_n55303_ );
xor  ( new_n55305_, new_n55284_, new_n55268_ );
and  ( new_n55306_, new_n55305_, new_n55304_ );
nor  ( new_n55307_, new_n55306_, new_n55285_ );
not  ( new_n55308_, new_n55307_ );
xor  ( new_n55309_, new_n55251_, new_n55225_ );
and  ( new_n55310_, new_n55309_, new_n55308_ );
or   ( new_n55311_, new_n55310_, new_n55252_ );
xor  ( new_n55312_, new_n55222_, new_n55220_ );
and  ( new_n55313_, new_n55312_, new_n55311_ );
nor  ( new_n55314_, new_n55313_, new_n55223_ );
nand ( new_n55315_, new_n55314_, new_n55131_ );
and  ( new_n55316_, new_n55315_, new_n55130_ );
xnor ( new_n55317_, new_n54755_, new_n54753_ );
xor  ( new_n55318_, new_n55317_, new_n54778_ );
and  ( new_n55319_, new_n55318_, new_n55316_ );
xor  ( new_n55320_, new_n55318_, new_n55316_ );
xor  ( new_n55321_, new_n54843_, new_n54841_ );
xor  ( new_n55322_, new_n55321_, new_n54847_ );
and  ( new_n55323_, new_n55322_, new_n55320_ );
nor  ( new_n55324_, new_n55323_, new_n55319_ );
xnor ( new_n55325_, new_n55125_, new_n55123_ );
nor  ( new_n55326_, new_n55325_, new_n55324_ );
or   ( new_n55327_, new_n55326_, new_n55126_ );
or   ( new_n55328_, new_n54632_, new_n54621_ );
or   ( new_n55329_, new_n54711_, new_n54634_ );
and  ( new_n55330_, new_n55329_, new_n55328_ );
nand ( new_n55331_, new_n54854_, new_n54852_ );
nand ( new_n55332_, new_n54857_, new_n54855_ );
and  ( new_n55333_, new_n55332_, new_n55331_ );
xor  ( new_n55334_, new_n55333_, new_n55330_ );
xor  ( new_n55335_, new_n54237_, new_n54235_ );
xor  ( new_n55336_, new_n55335_, new_n55334_ );
xnor ( new_n55337_, new_n55336_, new_n55327_ );
xor  ( new_n55338_, new_n55337_, new_n54863_ );
xnor ( new_n55339_, new_n55325_, new_n55324_ );
xor  ( new_n55340_, new_n54849_, new_n54780_ );
xor  ( new_n55341_, new_n55340_, new_n54858_ );
or   ( new_n55342_, new_n55341_, new_n55339_ );
and  ( new_n55343_, new_n55341_, new_n55339_ );
xor  ( new_n55344_, new_n55121_, new_n55120_ );
xnor ( new_n55345_, new_n54966_, new_n54964_ );
xor  ( new_n55346_, new_n55345_, new_n55049_ );
xor  ( new_n55347_, new_n54784_, new_n54782_ );
xor  ( new_n55348_, new_n55347_, new_n54839_ );
nand ( new_n55349_, new_n55348_, new_n55346_ );
nor  ( new_n55350_, new_n55348_, new_n55346_ );
xnor ( new_n55351_, new_n54962_, new_n54961_ );
xor  ( new_n55352_, new_n54952_, new_n54951_ );
xnor ( new_n55353_, new_n54976_, new_n54972_ );
nand ( new_n55354_, new_n55353_, new_n54981_ );
not  ( new_n55355_, new_n54977_ );
nand ( new_n55356_, new_n54983_, new_n55355_ );
and  ( new_n55357_, new_n55356_, new_n55354_ );
and  ( new_n55358_, new_n55357_, new_n55352_ );
or   ( new_n55359_, new_n55357_, new_n55352_ );
or   ( new_n55360_, new_n54916_, new_n340_ );
xor  ( new_n55361_, new_n52293_, RIbb2f250_9 );
or   ( new_n55362_, new_n55361_, new_n337_ );
and  ( new_n55363_, new_n55362_, new_n55360_ );
nor  ( new_n55364_, new_n55168_, new_n320_ );
xor  ( new_n55365_, new_n53306_, RIbb2f340_7 );
nor  ( new_n55366_, new_n55365_, new_n317_ );
or   ( new_n55367_, new_n55366_, new_n55364_ );
and  ( new_n55368_, new_n53694_, new_n280_ );
nand ( new_n55369_, new_n55368_, new_n55367_ );
xor  ( new_n55370_, new_n52902_, RIbb2f250_9 );
nor  ( new_n55371_, new_n55370_, new_n337_ );
nor  ( new_n55372_, new_n55361_, new_n340_ );
nor  ( new_n55373_, new_n55372_, new_n55371_ );
xnor ( new_n55374_, new_n55368_, new_n55367_ );
or   ( new_n55375_, new_n55374_, new_n55373_ );
and  ( new_n55376_, new_n55375_, new_n55369_ );
or   ( new_n55377_, new_n55376_, new_n55363_ );
nor  ( new_n55378_, new_n55092_, new_n899_ );
xor  ( new_n55379_, new_n50487_, new_n745_ );
nor  ( new_n55380_, new_n55379_, new_n897_ );
or   ( new_n55381_, new_n55380_, new_n55378_ );
xor  ( new_n55382_, new_n55376_, new_n55363_ );
nand ( new_n55383_, new_n55382_, new_n55381_ );
and  ( new_n55384_, new_n55383_, new_n55377_ );
xor  ( new_n55385_, new_n44407_, new_n6635_ );
or   ( new_n55386_, new_n55385_, new_n7184_ );
or   ( new_n55387_, new_n54943_, new_n7186_ );
and  ( new_n55388_, new_n55387_, new_n55386_ );
nor  ( new_n55389_, new_n55388_, new_n55384_ );
and  ( new_n55390_, new_n55388_, new_n55384_ );
xor  ( new_n55391_, new_n43956_, new_n8870_ );
nor  ( new_n55392_, new_n55391_, new_n9422_ );
and  ( new_n55393_, new_n54978_, new_n9185_ );
nor  ( new_n55394_, new_n55393_, new_n55392_ );
nor  ( new_n55395_, new_n55394_, new_n55390_ );
or   ( new_n55396_, new_n55395_, new_n55389_ );
and  ( new_n55397_, new_n55396_, new_n55359_ );
or   ( new_n55398_, new_n55397_, new_n55358_ );
xor  ( new_n55399_, new_n54986_, new_n54984_ );
xor  ( new_n55400_, new_n55399_, new_n54989_ );
nand ( new_n55401_, new_n55400_, new_n55398_ );
or   ( new_n55402_, new_n55400_, new_n55398_ );
xor  ( new_n55403_, new_n55043_, new_n55027_ );
nand ( new_n55404_, new_n55403_, new_n55402_ );
and  ( new_n55405_, new_n55404_, new_n55401_ );
nor  ( new_n55406_, new_n55405_, new_n55351_ );
and  ( new_n55407_, new_n55405_, new_n55351_ );
not  ( new_n55408_, new_n55407_ );
xor  ( new_n55409_, new_n55047_, new_n55046_ );
and  ( new_n55410_, new_n55409_, new_n55408_ );
nor  ( new_n55411_, new_n55410_, new_n55406_ );
or   ( new_n55412_, new_n55411_, new_n55350_ );
nand ( new_n55413_, new_n55412_, new_n55349_ );
nand ( new_n55414_, new_n55413_, new_n55344_ );
xnor ( new_n55415_, new_n55413_, new_n55344_ );
xor  ( new_n55416_, new_n55009_, new_n55008_ );
xnor ( new_n55417_, new_n55035_, new_n55031_ );
nand ( new_n55418_, new_n55417_, new_n55041_ );
not  ( new_n55419_, new_n55042_ );
or   ( new_n55420_, new_n55419_, new_n55036_ );
and  ( new_n55421_, new_n55420_, new_n55418_ );
nor  ( new_n55422_, new_n55421_, new_n55416_ );
nand ( new_n55423_, new_n55421_, new_n55416_ );
xnor ( new_n55424_, new_n55022_, new_n55021_ );
and  ( new_n55425_, new_n55424_, new_n55423_ );
or   ( new_n55426_, new_n55425_, new_n55422_ );
xnor ( new_n55427_, new_n55059_, new_n55057_ );
xor  ( new_n55428_, new_n55427_, new_n55067_ );
nor  ( new_n55429_, new_n55428_, new_n55426_ );
nand ( new_n55430_, new_n55428_, new_n55426_ );
xor  ( new_n55431_, new_n54959_, new_n54958_ );
and  ( new_n55432_, new_n55431_, new_n55430_ );
or   ( new_n55433_, new_n55432_, new_n55429_ );
xor  ( new_n55434_, new_n55071_, new_n55069_ );
xor  ( new_n55435_, new_n55434_, new_n55074_ );
or   ( new_n55436_, new_n55435_, new_n55433_ );
and  ( new_n55437_, new_n55435_, new_n55433_ );
xor  ( new_n55438_, new_n55082_, new_n55080_ );
xor  ( new_n55439_, new_n55438_, new_n55114_ );
or   ( new_n55440_, new_n55439_, new_n55437_ );
and  ( new_n55441_, new_n55440_, new_n55436_ );
xor  ( new_n55442_, new_n55076_, new_n55052_ );
xor  ( new_n55443_, new_n55442_, new_n55116_ );
nand ( new_n55444_, new_n55443_, new_n55441_ );
nor  ( new_n55445_, new_n55443_, new_n55441_ );
xor  ( new_n55446_, new_n55129_, new_n55127_ );
xor  ( new_n55447_, new_n55446_, new_n55314_ );
or   ( new_n55448_, new_n55447_, new_n55445_ );
and  ( new_n55449_, new_n55448_, new_n55444_ );
or   ( new_n55450_, new_n55449_, new_n55415_ );
and  ( new_n55451_, new_n55450_, new_n55414_ );
or   ( new_n55452_, new_n55451_, new_n55343_ );
and  ( new_n55453_, new_n55452_, new_n55342_ );
nor  ( new_n55454_, new_n55453_, new_n55338_ );
xor  ( new_n55455_, new_n55322_, new_n55320_ );
xor  ( new_n55456_, new_n55449_, new_n55415_ );
and  ( new_n55457_, new_n55456_, new_n55455_ );
xnor ( new_n55458_, new_n55104_, new_n55103_ );
xor  ( new_n55459_, new_n46962_, new_n2797_ );
or   ( new_n55460_, new_n55459_, new_n3117_ );
or   ( new_n55461_, new_n55132_, new_n3119_ );
and  ( new_n55462_, new_n55461_, new_n55460_ );
or   ( new_n55463_, new_n55185_, new_n2427_ );
xor  ( new_n55464_, new_n47296_, RIbb2e8f0_29 );
nand ( new_n55465_, new_n55464_, new_n2244_ );
and  ( new_n55466_, new_n55465_, new_n55463_ );
or   ( new_n55467_, new_n55466_, new_n55462_ );
xor  ( new_n55468_, new_n48039_, RIbb2e9e0_27 );
and  ( new_n55469_, new_n55468_, new_n2002_ );
nor  ( new_n55470_, new_n55141_, new_n2124_ );
nor  ( new_n55471_, new_n55470_, new_n55469_ );
not  ( new_n55472_, new_n55471_ );
xor  ( new_n55473_, new_n55466_, new_n55462_ );
nand ( new_n55474_, new_n55473_, new_n55472_ );
and  ( new_n55475_, new_n55474_, new_n55467_ );
or   ( new_n55476_, new_n55150_, new_n526_ );
xor  ( new_n55477_, new_n51446_, RIbb2f070_13 );
nand ( new_n55478_, new_n55477_, new_n456_ );
and  ( new_n55479_, new_n55478_, new_n55476_ );
xor  ( new_n55480_, new_n50894_, new_n520_ );
or   ( new_n55481_, new_n55480_, new_n755_ );
or   ( new_n55482_, new_n55085_, new_n757_ );
and  ( new_n55483_, new_n55482_, new_n55481_ );
or   ( new_n55484_, new_n55483_, new_n55479_ );
xor  ( new_n55485_, new_n49758_, new_n893_ );
nor  ( new_n55486_, new_n55485_, new_n1135_ );
and  ( new_n55487_, new_n55154_, new_n1040_ );
or   ( new_n55488_, new_n55487_, new_n55486_ );
xor  ( new_n55489_, new_n55483_, new_n55479_ );
nand ( new_n55490_, new_n55489_, new_n55488_ );
and  ( new_n55491_, new_n55490_, new_n55484_ );
or   ( new_n55492_, new_n55491_, new_n55475_ );
or   ( new_n55493_, RIbb2f2c8_8, RIbb2f250_9 );
and  ( new_n55494_, new_n53694_, new_n55493_ );
or   ( new_n55495_, new_n55494_, new_n312_ );
or   ( new_n55496_, new_n55365_, new_n320_ );
or   ( new_n55497_, new_n54908_, new_n317_ );
or   ( new_n55498_, new_n55497_, new_n54911_ );
and  ( new_n55499_, new_n55498_, new_n55496_ );
or   ( new_n55500_, new_n55499_, new_n55495_ );
or   ( new_n55501_, new_n55173_, new_n411_ );
xor  ( new_n55502_, new_n52280_, new_n325_ );
or   ( new_n55503_, new_n55502_, new_n409_ );
and  ( new_n55504_, new_n55503_, new_n55501_ );
or   ( new_n55505_, new_n55504_, new_n55500_ );
and  ( new_n55506_, new_n55477_, new_n454_ );
xor  ( new_n55507_, new_n51477_, RIbb2f070_13 );
and  ( new_n55508_, new_n55507_, new_n456_ );
nor  ( new_n55509_, new_n55508_, new_n55506_ );
xnor ( new_n55510_, new_n55504_, new_n55500_ );
or   ( new_n55511_, new_n55510_, new_n55509_ );
and  ( new_n55512_, new_n55511_, new_n55505_ );
or   ( new_n55513_, new_n55180_, new_n2809_ );
xor  ( new_n55514_, new_n47303_, new_n2421_ );
or   ( new_n55515_, new_n55514_, new_n2807_ );
and  ( new_n55516_, new_n55515_, new_n55513_ );
nor  ( new_n55517_, new_n55516_, new_n55512_ );
xor  ( new_n55518_, new_n46619_, new_n3113_ );
nor  ( new_n55519_, new_n55518_, new_n3461_ );
and  ( new_n55520_, new_n55159_, new_n3291_ );
or   ( new_n55521_, new_n55520_, new_n55519_ );
xor  ( new_n55522_, new_n55516_, new_n55512_ );
and  ( new_n55523_, new_n55522_, new_n55521_ );
nor  ( new_n55524_, new_n55523_, new_n55517_ );
and  ( new_n55525_, new_n55491_, new_n55475_ );
or   ( new_n55526_, new_n55525_, new_n55524_ );
and  ( new_n55527_, new_n55526_, new_n55492_ );
nor  ( new_n55528_, new_n55527_, new_n55458_ );
xor  ( new_n55529_, new_n55162_, new_n55161_ );
xor  ( new_n55530_, new_n55095_, new_n55094_ );
and  ( new_n55531_, new_n55530_, new_n55529_ );
or   ( new_n55532_, new_n55226_, new_n1366_ );
xor  ( new_n55533_, new_n49427_, new_n1126_ );
or   ( new_n55534_, new_n55533_, new_n1364_ );
and  ( new_n55535_, new_n55534_, new_n55532_ );
or   ( new_n55536_, new_n55136_, new_n1595_ );
xor  ( new_n55537_, new_n48908_, new_n1355_ );
or   ( new_n55538_, new_n55537_, new_n1593_ );
and  ( new_n55539_, new_n55538_, new_n55536_ );
nor  ( new_n55540_, new_n55539_, new_n55535_ );
xor  ( new_n55541_, new_n48518_, RIbb2ead0_25 );
and  ( new_n55542_, new_n55541_, new_n1741_ );
and  ( new_n55543_, new_n55230_, new_n1739_ );
or   ( new_n55544_, new_n55543_, new_n55542_ );
xor  ( new_n55545_, new_n55539_, new_n55535_ );
and  ( new_n55546_, new_n55545_, new_n55544_ );
nor  ( new_n55547_, new_n55546_, new_n55540_ );
xnor ( new_n55548_, new_n55530_, new_n55529_ );
nor  ( new_n55549_, new_n55548_, new_n55547_ );
or   ( new_n55550_, new_n55549_, new_n55531_ );
xor  ( new_n55551_, new_n55527_, new_n55458_ );
and  ( new_n55552_, new_n55551_, new_n55550_ );
nor  ( new_n55553_, new_n55552_, new_n55528_ );
not  ( new_n55554_, new_n55553_ );
xor  ( new_n55555_, new_n55111_, new_n55109_ );
nand ( new_n55556_, new_n55555_, new_n55554_ );
xor  ( new_n55557_, new_n55555_, new_n55554_ );
xor  ( new_n55558_, new_n55218_, new_n55217_ );
nand ( new_n55559_, new_n55558_, new_n55557_ );
and  ( new_n55560_, new_n55559_, new_n55556_ );
xor  ( new_n55561_, new_n55215_, new_n55214_ );
xnor ( new_n55562_, new_n55246_, new_n55241_ );
xor  ( new_n55563_, new_n55562_, new_n55249_ );
nor  ( new_n55564_, new_n55563_, new_n55561_ );
nand ( new_n55565_, new_n55563_, new_n55561_ );
xor  ( new_n55566_, new_n55301_, new_n55300_ );
xor  ( new_n55567_, new_n55212_, new_n55211_ );
and  ( new_n55568_, new_n55567_, new_n55566_ );
xor  ( new_n55569_, new_n55567_, new_n55566_ );
xor  ( new_n55570_, new_n55266_, new_n55265_ );
and  ( new_n55571_, new_n55570_, new_n55569_ );
nor  ( new_n55572_, new_n55571_, new_n55568_ );
and  ( new_n55573_, new_n55572_, new_n55565_ );
or   ( new_n55574_, new_n55573_, new_n55564_ );
xor  ( new_n55575_, new_n55164_, new_n55148_ );
and  ( new_n55576_, new_n55575_, new_n55191_ );
not  ( new_n55577_, new_n55166_ );
and  ( new_n55578_, new_n55193_, new_n55577_ );
or   ( new_n55579_, new_n55578_, new_n55576_ );
xor  ( new_n55580_, new_n55233_, new_n55229_ );
xor  ( new_n55581_, new_n55580_, new_n55238_ );
xor  ( new_n55582_, new_n55145_, new_n55144_ );
nand ( new_n55583_, new_n55582_, new_n55581_ );
nor  ( new_n55584_, new_n55582_, new_n55581_ );
xor  ( new_n55585_, new_n45738_, new_n4292_ );
or   ( new_n55586_, new_n55585_, new_n4709_ );
nand ( new_n55587_, new_n55296_, new_n4541_ );
and  ( new_n55588_, new_n55587_, new_n55586_ );
or   ( new_n55589_, new_n55286_, new_n7734_ );
xor  ( new_n55590_, new_n44319_, RIbb2ddb0_53 );
nand ( new_n55591_, new_n55590_, new_n7489_ );
and  ( new_n55592_, new_n55591_, new_n55589_ );
nor  ( new_n55593_, new_n55592_, new_n55588_ );
and  ( new_n55594_, new_n55208_, new_n4032_ );
xor  ( new_n55595_, new_n45928_, new_n3892_ );
nor  ( new_n55596_, new_n55595_, new_n4302_ );
or   ( new_n55597_, new_n55596_, new_n55594_ );
xor  ( new_n55598_, new_n55592_, new_n55588_ );
and  ( new_n55599_, new_n55598_, new_n55597_ );
nor  ( new_n55600_, new_n55599_, new_n55593_ );
or   ( new_n55601_, new_n55600_, new_n55584_ );
and  ( new_n55602_, new_n55601_, new_n55583_ );
or   ( new_n55603_, new_n55602_, new_n55579_ );
and  ( new_n55604_, new_n55602_, new_n55579_ );
xor  ( new_n55605_, new_n45403_, new_n4705_ );
or   ( new_n55606_, new_n55605_, new_n5207_ );
or   ( new_n55607_, new_n55273_, new_n5209_ );
and  ( new_n55608_, new_n55607_, new_n55606_ );
xor  ( new_n55609_, new_n43803_, new_n10052_ );
or   ( new_n55610_, new_n55609_, new_n21077_ );
or   ( new_n55611_, new_n43884_, new_n10052_ );
or   ( new_n55612_, new_n55611_, RIbb2d888_64 );
and  ( new_n55613_, new_n55612_, new_n55610_ );
or   ( new_n55614_, new_n55613_, new_n55608_ );
xor  ( new_n55615_, new_n44183_, RIbb2dcc0_55 );
and  ( new_n55616_, new_n55615_, new_n8042_ );
and  ( new_n55617_, new_n55269_, new_n8040_ );
nor  ( new_n55618_, new_n55617_, new_n55616_ );
and  ( new_n55619_, new_n55613_, new_n55608_ );
or   ( new_n55620_, new_n55619_, new_n55618_ );
and  ( new_n55621_, new_n55620_, new_n55614_ );
xor  ( new_n55622_, new_n43812_, new_n8254_ );
or   ( new_n55623_, new_n55622_, new_n8874_ );
or   ( new_n55624_, new_n55253_, new_n8876_ );
and  ( new_n55625_, new_n55624_, new_n55623_ );
xor  ( new_n55626_, new_n45119_, new_n5203_ );
or   ( new_n55627_, new_n55626_, new_n5604_ );
nand ( new_n55628_, new_n55280_, new_n5371_ );
and  ( new_n55629_, new_n55628_, new_n55627_ );
or   ( new_n55630_, new_n55629_, new_n55625_ );
xor  ( new_n55631_, new_n44877_, RIbb2e080_47 );
and  ( new_n55632_, new_n55631_, new_n5917_ );
and  ( new_n55633_, new_n55262_, new_n5915_ );
or   ( new_n55634_, new_n55633_, new_n55632_ );
xor  ( new_n55635_, new_n55629_, new_n55625_ );
nand ( new_n55636_, new_n55635_, new_n55634_ );
and  ( new_n55637_, new_n55636_, new_n55630_ );
nor  ( new_n55638_, new_n55637_, new_n55621_ );
xor  ( new_n55639_, new_n44506_, RIbb2dea0_51 );
nand ( new_n55640_, new_n55639_, new_n6910_ );
or   ( new_n55641_, new_n55385_, new_n7186_ );
and  ( new_n55642_, new_n55641_, new_n55640_ );
or   ( new_n55643_, new_n55201_, new_n3898_ );
xor  ( new_n55644_, new_n46137_, RIbb2e530_37 );
nand ( new_n55645_, new_n55644_, new_n3733_ );
and  ( new_n55646_, new_n55645_, new_n55643_ );
nor  ( new_n55647_, new_n55646_, new_n55642_ );
xor  ( new_n55648_, new_n43952_, new_n8870_ );
nor  ( new_n55649_, new_n55648_, new_n9422_ );
nor  ( new_n55650_, new_n55391_, new_n9424_ );
or   ( new_n55651_, new_n55650_, new_n55649_ );
xor  ( new_n55652_, new_n55646_, new_n55642_ );
and  ( new_n55653_, new_n55652_, new_n55651_ );
or   ( new_n55654_, new_n55653_, new_n55647_ );
xor  ( new_n55655_, new_n55637_, new_n55621_ );
and  ( new_n55656_, new_n55655_, new_n55654_ );
nor  ( new_n55657_, new_n55656_, new_n55638_ );
or   ( new_n55658_, new_n55657_, new_n55604_ );
and  ( new_n55659_, new_n55658_, new_n55603_ );
or   ( new_n55660_, new_n55659_, new_n55574_ );
nand ( new_n55661_, new_n55659_, new_n55574_ );
xor  ( new_n55662_, new_n55309_, new_n55308_ );
nand ( new_n55663_, new_n55662_, new_n55661_ );
and  ( new_n55664_, new_n55663_, new_n55660_ );
nor  ( new_n55665_, new_n55664_, new_n55560_ );
xor  ( new_n55666_, new_n55312_, new_n55311_ );
xor  ( new_n55667_, new_n55664_, new_n55560_ );
and  ( new_n55668_, new_n55667_, new_n55666_ );
or   ( new_n55669_, new_n55668_, new_n55665_ );
xnor ( new_n55670_, new_n55348_, new_n55346_ );
xor  ( new_n55671_, new_n55670_, new_n55411_ );
and  ( new_n55672_, new_n55671_, new_n55669_ );
xor  ( new_n55673_, new_n55305_, new_n55304_ );
xor  ( new_n55674_, new_n55189_, new_n55188_ );
xnor ( new_n55675_, new_n55388_, new_n55384_ );
nand ( new_n55676_, new_n55675_, new_n55394_ );
not  ( new_n55677_, new_n55389_ );
nand ( new_n55678_, new_n55395_, new_n55677_ );
and  ( new_n55679_, new_n55678_, new_n55676_ );
nand ( new_n55680_, new_n55679_, new_n55674_ );
nor  ( new_n55681_, new_n55679_, new_n55674_ );
xor  ( new_n55682_, new_n43937_, RIbb2d9f0_61 );
and  ( new_n55683_, new_n55682_, new_n9740_ );
and  ( new_n55684_, new_n55258_, new_n9738_ );
or   ( new_n55685_, new_n55684_, new_n55683_ );
xor  ( new_n55686_, new_n55177_, new_n55176_ );
and  ( new_n55687_, new_n55686_, new_n55685_ );
xor  ( new_n55688_, new_n44681_, RIbb2df90_49 );
and  ( new_n55689_, new_n55688_, new_n6510_ );
and  ( new_n55690_, new_n55235_, new_n6508_ );
or   ( new_n55691_, new_n55690_, new_n55689_ );
xor  ( new_n55692_, new_n55686_, new_n55685_ );
and  ( new_n55693_, new_n55692_, new_n55691_ );
nor  ( new_n55694_, new_n55693_, new_n55687_ );
or   ( new_n55695_, new_n55694_, new_n55681_ );
nand ( new_n55696_, new_n55695_, new_n55680_ );
and  ( new_n55697_, new_n55696_, new_n55673_ );
xnor ( new_n55698_, new_n55696_, new_n55673_ );
xor  ( new_n55699_, new_n55421_, new_n55416_ );
xor  ( new_n55700_, new_n55699_, new_n55424_ );
nor  ( new_n55701_, new_n55700_, new_n55698_ );
or   ( new_n55702_, new_n55701_, new_n55697_ );
xor  ( new_n55703_, new_n55400_, new_n55398_ );
xor  ( new_n55704_, new_n55703_, new_n55403_ );
nor  ( new_n55705_, new_n55704_, new_n55702_ );
and  ( new_n55706_, new_n55704_, new_n55702_ );
xor  ( new_n55707_, new_n55428_, new_n55426_ );
xor  ( new_n55708_, new_n55707_, new_n55431_ );
nor  ( new_n55709_, new_n55708_, new_n55706_ );
nor  ( new_n55710_, new_n55709_, new_n55705_ );
xor  ( new_n55711_, new_n55405_, new_n55351_ );
xor  ( new_n55712_, new_n55711_, new_n55409_ );
and  ( new_n55713_, new_n55712_, new_n55710_ );
xor  ( new_n55714_, new_n55712_, new_n55710_ );
not  ( new_n55715_, new_n55714_ );
xnor ( new_n55716_, new_n55435_, new_n55433_ );
xor  ( new_n55717_, new_n55716_, new_n55439_ );
nor  ( new_n55718_, new_n55717_, new_n55715_ );
or   ( new_n55719_, new_n55718_, new_n55713_ );
xor  ( new_n55720_, new_n55671_, new_n55669_ );
and  ( new_n55721_, new_n55720_, new_n55719_ );
nor  ( new_n55722_, new_n55721_, new_n55672_ );
xnor ( new_n55723_, new_n55456_, new_n55455_ );
nor  ( new_n55724_, new_n55723_, new_n55722_ );
nor  ( new_n55725_, new_n55724_, new_n55457_ );
xor  ( new_n55726_, new_n55341_, new_n55339_ );
xor  ( new_n55727_, new_n55726_, new_n55451_ );
and  ( new_n55728_, new_n55727_, new_n55725_ );
nor  ( new_n55729_, new_n55727_, new_n55725_ );
xnor ( new_n55730_, new_n55723_, new_n55722_ );
xor  ( new_n55731_, new_n55720_, new_n55719_ );
xnor ( new_n55732_, new_n55443_, new_n55441_ );
xor  ( new_n55733_, new_n55732_, new_n55447_ );
nand ( new_n55734_, new_n55733_, new_n55731_ );
nor  ( new_n55735_, new_n55733_, new_n55731_ );
xnor ( new_n55736_, new_n55558_, new_n55557_ );
xor  ( new_n55737_, new_n50788_, new_n745_ );
or   ( new_n55738_, new_n55737_, new_n897_ );
or   ( new_n55739_, new_n55379_, new_n899_ );
and  ( new_n55740_, new_n55739_, new_n55738_ );
xor  ( new_n55741_, new_n51142_, new_n520_ );
or   ( new_n55742_, new_n55741_, new_n755_ );
or   ( new_n55743_, new_n55480_, new_n757_ );
and  ( new_n55744_, new_n55743_, new_n55742_ );
nor  ( new_n55745_, new_n55744_, new_n55740_ );
nor  ( new_n55746_, new_n55514_, new_n2809_ );
xor  ( new_n55747_, new_n47046_, new_n2421_ );
nor  ( new_n55748_, new_n55747_, new_n2807_ );
nor  ( new_n55749_, new_n55748_, new_n55746_ );
xnor ( new_n55750_, new_n55744_, new_n55740_ );
nor  ( new_n55751_, new_n55750_, new_n55749_ );
or   ( new_n55752_, new_n55751_, new_n55745_ );
xor  ( new_n55753_, new_n55382_, new_n55381_ );
or   ( new_n55754_, new_n55753_, new_n55752_ );
and  ( new_n55755_, new_n55753_, new_n55752_ );
xnor ( new_n55756_, new_n55374_, new_n55373_ );
or   ( new_n55757_, new_n55533_, new_n1366_ );
xor  ( new_n55758_, new_n49488_, new_n1126_ );
or   ( new_n55759_, new_n55758_, new_n1364_ );
and  ( new_n55760_, new_n55759_, new_n55757_ );
and  ( new_n55761_, new_n55760_, new_n55756_ );
nor  ( new_n55762_, new_n55485_, new_n1137_ );
xor  ( new_n55763_, new_n50115_, new_n893_ );
nor  ( new_n55764_, new_n55763_, new_n1135_ );
nor  ( new_n55765_, new_n55764_, new_n55762_ );
nor  ( new_n55766_, new_n55760_, new_n55756_ );
not  ( new_n55767_, new_n55766_ );
and  ( new_n55768_, new_n55767_, new_n55765_ );
nor  ( new_n55769_, new_n55768_, new_n55761_ );
or   ( new_n55770_, new_n55769_, new_n55755_ );
and  ( new_n55771_, new_n55770_, new_n55754_ );
xnor ( new_n55772_, new_n55276_, new_n55272_ );
nand ( new_n55773_, new_n55772_, new_n55282_ );
not  ( new_n55774_, new_n55283_ );
or   ( new_n55775_, new_n55774_, new_n55277_ );
and  ( new_n55776_, new_n55775_, new_n55773_ );
and  ( new_n55777_, new_n55776_, new_n55771_ );
or   ( new_n55778_, new_n55776_, new_n55771_ );
or   ( new_n55779_, new_n55537_, new_n1595_ );
xor  ( new_n55780_, new_n49265_, new_n1355_ );
or   ( new_n55781_, new_n55780_, new_n1593_ );
and  ( new_n55782_, new_n55781_, new_n55779_ );
or   ( new_n55783_, new_n55459_, new_n3119_ );
xor  ( new_n55784_, new_n46958_, new_n2797_ );
or   ( new_n55785_, new_n55784_, new_n3117_ );
and  ( new_n55786_, new_n55785_, new_n55783_ );
nor  ( new_n55787_, new_n55786_, new_n55782_ );
and  ( new_n55788_, new_n55644_, new_n3731_ );
xor  ( new_n55789_, new_n46427_, RIbb2e530_37 );
and  ( new_n55790_, new_n55789_, new_n3733_ );
nor  ( new_n55791_, new_n55790_, new_n55788_ );
and  ( new_n55792_, new_n55786_, new_n55782_ );
nor  ( new_n55793_, new_n55792_, new_n55791_ );
or   ( new_n55794_, new_n55793_, new_n55787_ );
xor  ( new_n55795_, new_n55489_, new_n55488_ );
and  ( new_n55796_, new_n55795_, new_n55794_ );
nor  ( new_n55797_, new_n55795_, new_n55794_ );
nor  ( new_n55798_, new_n55370_, new_n340_ );
xor  ( new_n55799_, new_n52908_, RIbb2f250_9 );
nor  ( new_n55800_, new_n55799_, new_n337_ );
or   ( new_n55801_, new_n55800_, new_n55798_ );
xor  ( new_n55802_, new_n55499_, new_n55495_ );
nand ( new_n55803_, new_n55802_, new_n55801_ );
nor  ( new_n55804_, new_n55502_, new_n411_ );
xor  ( new_n55805_, new_n52293_, RIbb2f160_11 );
nor  ( new_n55806_, new_n55805_, new_n409_ );
or   ( new_n55807_, new_n55806_, new_n55804_ );
xor  ( new_n55808_, new_n55802_, new_n55801_ );
nand ( new_n55809_, new_n55808_, new_n55807_ );
and  ( new_n55810_, new_n55809_, new_n55803_ );
nand ( new_n55811_, new_n55468_, new_n2000_ );
xor  ( new_n55812_, new_n48291_, RIbb2e9e0_27 );
nand ( new_n55813_, new_n55812_, new_n2002_ );
and  ( new_n55814_, new_n55813_, new_n55811_ );
nor  ( new_n55815_, new_n55814_, new_n55810_ );
xor  ( new_n55816_, new_n47640_, new_n2118_ );
nor  ( new_n55817_, new_n55816_, new_n2425_ );
and  ( new_n55818_, new_n55464_, new_n2242_ );
nor  ( new_n55819_, new_n55818_, new_n55817_ );
not  ( new_n55820_, new_n55819_ );
xor  ( new_n55821_, new_n55814_, new_n55810_ );
and  ( new_n55822_, new_n55821_, new_n55820_ );
nor  ( new_n55823_, new_n55822_, new_n55815_ );
nor  ( new_n55824_, new_n55823_, new_n55797_ );
or   ( new_n55825_, new_n55824_, new_n55796_ );
and  ( new_n55826_, new_n55825_, new_n55778_ );
or   ( new_n55827_, new_n55826_, new_n55777_ );
xor  ( new_n55828_, new_n55357_, new_n55352_ );
xor  ( new_n55829_, new_n55828_, new_n55396_ );
nand ( new_n55830_, new_n55829_, new_n55827_ );
nor  ( new_n55831_, new_n55829_, new_n55827_ );
xnor ( new_n55832_, new_n55548_, new_n55547_ );
or   ( new_n55833_, new_n55585_, new_n4711_ );
xor  ( new_n55834_, new_n45597_, RIbb2e350_41 );
nand ( new_n55835_, new_n55834_, new_n4543_ );
and  ( new_n55836_, new_n55835_, new_n55833_ );
or   ( new_n55837_, new_n55595_, new_n4304_ );
xor  ( new_n55838_, new_n46037_, new_n3892_ );
or   ( new_n55839_, new_n55838_, new_n4302_ );
and  ( new_n55840_, new_n55839_, new_n55837_ );
nor  ( new_n55841_, new_n55840_, new_n55836_ );
xor  ( new_n55842_, new_n44407_, RIbb2ddb0_53 );
and  ( new_n55843_, new_n55842_, new_n7489_ );
and  ( new_n55844_, new_n55590_, new_n7487_ );
or   ( new_n55845_, new_n55844_, new_n55843_ );
xor  ( new_n55846_, new_n55840_, new_n55836_ );
and  ( new_n55847_, new_n55846_, new_n55845_ );
or   ( new_n55848_, new_n55847_, new_n55841_ );
xor  ( new_n55849_, new_n55545_, new_n55544_ );
nand ( new_n55850_, new_n55849_, new_n55848_ );
nor  ( new_n55851_, new_n55849_, new_n55848_ );
xnor ( new_n55852_, new_n55510_, new_n55509_ );
xor  ( new_n55853_, new_n43884_, new_n10052_ );
or   ( new_n55854_, new_n55853_, new_n21077_ );
or   ( new_n55855_, new_n43888_, new_n10052_ );
or   ( new_n55856_, new_n55855_, RIbb2d888_64 );
and  ( new_n55857_, new_n55856_, new_n55854_ );
nor  ( new_n55858_, new_n55857_, new_n55852_ );
and  ( new_n55859_, new_n55639_, new_n6908_ );
xor  ( new_n55860_, new_n44600_, RIbb2dea0_51 );
and  ( new_n55861_, new_n55860_, new_n6910_ );
or   ( new_n55862_, new_n55861_, new_n55859_ );
xor  ( new_n55863_, new_n55857_, new_n55852_ );
and  ( new_n55864_, new_n55863_, new_n55862_ );
nor  ( new_n55865_, new_n55864_, new_n55858_ );
or   ( new_n55866_, new_n55865_, new_n55851_ );
and  ( new_n55867_, new_n55866_, new_n55850_ );
nor  ( new_n55868_, new_n55867_, new_n55832_ );
and  ( new_n55869_, new_n55867_, new_n55832_ );
nor  ( new_n55870_, new_n55518_, new_n3463_ );
xor  ( new_n55871_, new_n46789_, new_n3113_ );
nor  ( new_n55872_, new_n55871_, new_n3461_ );
nor  ( new_n55873_, new_n55872_, new_n55870_ );
nand ( new_n55874_, new_n55541_, new_n1739_ );
xor  ( new_n55875_, new_n48756_, RIbb2ead0_25 );
nand ( new_n55876_, new_n55875_, new_n1741_ );
and  ( new_n55877_, new_n55876_, new_n55874_ );
nor  ( new_n55878_, new_n55877_, new_n55873_ );
and  ( new_n55879_, new_n55682_, new_n9738_ );
xor  ( new_n55880_, new_n43956_, new_n9418_ );
nor  ( new_n55881_, new_n55880_, new_n10059_ );
nor  ( new_n55882_, new_n55881_, new_n55879_ );
and  ( new_n55883_, new_n55877_, new_n55873_ );
nor  ( new_n55884_, new_n55883_, new_n55882_ );
or   ( new_n55885_, new_n55884_, new_n55878_ );
xor  ( new_n55886_, new_n55522_, new_n55521_ );
and  ( new_n55887_, new_n55886_, new_n55885_ );
xor  ( new_n55888_, new_n45584_, new_n4705_ );
or   ( new_n55889_, new_n55888_, new_n5207_ );
or   ( new_n55890_, new_n55605_, new_n5209_ );
and  ( new_n55891_, new_n55890_, new_n55889_ );
nand ( new_n55892_, new_n55615_, new_n8040_ );
xor  ( new_n55893_, new_n44218_, new_n7722_ );
or   ( new_n55894_, new_n55893_, new_n8264_ );
and  ( new_n55895_, new_n55894_, new_n55892_ );
nor  ( new_n55896_, new_n55895_, new_n55891_ );
nor  ( new_n55897_, new_n55626_, new_n5606_ );
xor  ( new_n55898_, new_n45204_, RIbb2e170_45 );
and  ( new_n55899_, new_n55898_, new_n5373_ );
or   ( new_n55900_, new_n55899_, new_n55897_ );
xor  ( new_n55901_, new_n55895_, new_n55891_ );
and  ( new_n55902_, new_n55901_, new_n55900_ );
or   ( new_n55903_, new_n55902_, new_n55896_ );
xor  ( new_n55904_, new_n55886_, new_n55885_ );
and  ( new_n55905_, new_n55904_, new_n55903_ );
nor  ( new_n55906_, new_n55905_, new_n55887_ );
nor  ( new_n55907_, new_n55906_, new_n55869_ );
nor  ( new_n55908_, new_n55907_, new_n55868_ );
or   ( new_n55909_, new_n55908_, new_n55831_ );
and  ( new_n55910_, new_n55909_, new_n55830_ );
nor  ( new_n55911_, new_n55910_, new_n55736_ );
xor  ( new_n55912_, new_n55551_, new_n55550_ );
xnor ( new_n55913_, new_n55602_, new_n55579_ );
xor  ( new_n55914_, new_n55913_, new_n55657_ );
and  ( new_n55915_, new_n55914_, new_n55912_ );
xnor ( new_n55916_, new_n55491_, new_n55475_ );
xor  ( new_n55917_, new_n55916_, new_n55524_ );
xnor ( new_n55918_, new_n55679_, new_n55674_ );
xor  ( new_n55919_, new_n55918_, new_n55694_ );
and  ( new_n55920_, new_n55919_, new_n55917_ );
xor  ( new_n55921_, new_n55473_, new_n55472_ );
not  ( new_n55922_, new_n55921_ );
xor  ( new_n55923_, new_n43914_, new_n8254_ );
or   ( new_n55924_, new_n55923_, new_n8874_ );
or   ( new_n55925_, new_n55622_, new_n8876_ );
and  ( new_n55926_, new_n55925_, new_n55924_ );
xor  ( new_n55927_, new_n44974_, RIbb2e080_47 );
nand ( new_n55928_, new_n55927_, new_n5917_ );
nand ( new_n55929_, new_n55631_, new_n5915_ );
and  ( new_n55930_, new_n55929_, new_n55928_ );
or   ( new_n55931_, new_n55930_, new_n55926_ );
xor  ( new_n55932_, new_n44785_, RIbb2df90_49 );
and  ( new_n55933_, new_n55932_, new_n6510_ );
and  ( new_n55934_, new_n55688_, new_n6508_ );
nor  ( new_n55935_, new_n55934_, new_n55933_ );
and  ( new_n55936_, new_n55930_, new_n55926_ );
or   ( new_n55937_, new_n55936_, new_n55935_ );
and  ( new_n55938_, new_n55937_, new_n55931_ );
nor  ( new_n55939_, new_n55938_, new_n55922_ );
xor  ( new_n55940_, new_n55938_, new_n55922_ );
xor  ( new_n55941_, new_n55635_, new_n55634_ );
and  ( new_n55942_, new_n55941_, new_n55940_ );
or   ( new_n55943_, new_n55942_, new_n55939_ );
xor  ( new_n55944_, new_n55919_, new_n55917_ );
and  ( new_n55945_, new_n55944_, new_n55943_ );
or   ( new_n55946_, new_n55945_, new_n55920_ );
xor  ( new_n55947_, new_n55914_, new_n55912_ );
and  ( new_n55948_, new_n55947_, new_n55946_ );
nor  ( new_n55949_, new_n55948_, new_n55915_ );
xnor ( new_n55950_, new_n55910_, new_n55736_ );
nor  ( new_n55951_, new_n55950_, new_n55949_ );
or   ( new_n55952_, new_n55951_, new_n55911_ );
xor  ( new_n55953_, new_n55667_, new_n55666_ );
and  ( new_n55954_, new_n55953_, new_n55952_ );
nor  ( new_n55955_, new_n55953_, new_n55952_ );
xor  ( new_n55956_, new_n55717_, new_n55715_ );
not  ( new_n55957_, new_n55956_ );
nor  ( new_n55958_, new_n55957_, new_n55955_ );
nor  ( new_n55959_, new_n55958_, new_n55954_ );
or   ( new_n55960_, new_n55959_, new_n55735_ );
and  ( new_n55961_, new_n55960_, new_n55734_ );
and  ( new_n55962_, new_n55961_, new_n55730_ );
xnor ( new_n55963_, new_n55950_, new_n55949_ );
xnor ( new_n55964_, new_n55570_, new_n55569_ );
xnor ( new_n55965_, new_n55613_, new_n55608_ );
xor  ( new_n55966_, new_n55965_, new_n55618_ );
xor  ( new_n55967_, new_n55598_, new_n55597_ );
nand ( new_n55968_, new_n55967_, new_n55966_ );
nor  ( new_n55969_, new_n55967_, new_n55966_ );
xor  ( new_n55970_, new_n55753_, new_n55752_ );
xnor ( new_n55971_, new_n55970_, new_n55769_ );
or   ( new_n55972_, new_n55971_, new_n55969_ );
and  ( new_n55973_, new_n55972_, new_n55968_ );
nor  ( new_n55974_, new_n55973_, new_n55964_ );
and  ( new_n55975_, new_n55973_, new_n55964_ );
xor  ( new_n55976_, new_n55795_, new_n55794_ );
xor  ( new_n55977_, new_n55976_, new_n55823_ );
xor  ( new_n55978_, new_n47303_, new_n2797_ );
or   ( new_n55979_, new_n55978_, new_n3117_ );
or   ( new_n55980_, new_n55784_, new_n3119_ );
and  ( new_n55981_, new_n55980_, new_n55979_ );
xor  ( new_n55982_, new_n46962_, new_n3113_ );
or   ( new_n55983_, new_n55982_, new_n3461_ );
or   ( new_n55984_, new_n55871_, new_n3463_ );
and  ( new_n55985_, new_n55984_, new_n55983_ );
nor  ( new_n55986_, new_n55985_, new_n55981_ );
xor  ( new_n55987_, new_n48908_, new_n1583_ );
nor  ( new_n55988_, new_n55987_, new_n1844_ );
and  ( new_n55989_, new_n55875_, new_n1739_ );
nor  ( new_n55990_, new_n55989_, new_n55988_ );
xnor ( new_n55991_, new_n55985_, new_n55981_ );
nor  ( new_n55992_, new_n55991_, new_n55990_ );
nor  ( new_n55993_, new_n55992_, new_n55986_ );
not  ( new_n55994_, new_n55993_ );
or   ( new_n55995_, new_n55780_, new_n1595_ );
xor  ( new_n55996_, new_n49427_, RIbb2ebc0_23 );
nand ( new_n55997_, new_n55996_, new_n1476_ );
and  ( new_n55998_, new_n55997_, new_n55995_ );
nand ( new_n55999_, new_n55789_, new_n3731_ );
xor  ( new_n56000_, new_n46619_, new_n3457_ );
or   ( new_n56001_, new_n56000_, new_n3896_ );
and  ( new_n56002_, new_n56001_, new_n55999_ );
nor  ( new_n56003_, new_n56002_, new_n55998_ );
and  ( new_n56004_, new_n55812_, new_n2000_ );
xor  ( new_n56005_, new_n48518_, RIbb2e9e0_27 );
and  ( new_n56006_, new_n56005_, new_n2002_ );
or   ( new_n56007_, new_n56006_, new_n56004_ );
xor  ( new_n56008_, new_n56002_, new_n55998_ );
and  ( new_n56009_, new_n56008_, new_n56007_ );
nor  ( new_n56010_, new_n56009_, new_n56003_ );
not  ( new_n56011_, new_n56010_ );
and  ( new_n56012_, new_n56011_, new_n55994_ );
and  ( new_n56013_, new_n56010_, new_n55993_ );
or   ( new_n56014_, new_n55816_, new_n2427_ );
xor  ( new_n56015_, new_n48039_, new_n2118_ );
or   ( new_n56016_, new_n56015_, new_n2425_ );
and  ( new_n56017_, new_n56016_, new_n56014_ );
xor  ( new_n56018_, new_n47296_, new_n2421_ );
or   ( new_n56019_, new_n56018_, new_n2807_ );
or   ( new_n56020_, new_n55747_, new_n2809_ );
and  ( new_n56021_, new_n56020_, new_n56019_ );
nor  ( new_n56022_, new_n56021_, new_n56017_ );
xor  ( new_n56023_, new_n53306_, RIbb2f250_9 );
nor  ( new_n56024_, new_n56023_, new_n340_ );
nand ( new_n56025_, new_n53694_, RIbb2f250_9 );
nor  ( new_n56026_, new_n53694_, RIbb2f250_9 );
nor  ( new_n56027_, new_n56026_, new_n337_ );
and  ( new_n56028_, new_n56027_, new_n56025_ );
or   ( new_n56029_, new_n56028_, new_n56024_ );
or   ( new_n56030_, new_n53695_, new_n13844_ );
and  ( new_n56031_, new_n56030_, new_n331_ );
nand ( new_n56032_, new_n56031_, new_n56029_ );
xor  ( new_n56033_, new_n51758_, new_n400_ );
or   ( new_n56034_, new_n56033_, new_n526_ );
xor  ( new_n56035_, new_n52280_, new_n400_ );
or   ( new_n56036_, new_n56035_, new_n524_ );
and  ( new_n56037_, new_n56036_, new_n56034_ );
nor  ( new_n56038_, new_n56037_, new_n56032_ );
xor  ( new_n56039_, new_n51446_, RIbb2ef80_15 );
and  ( new_n56040_, new_n56039_, new_n660_ );
xor  ( new_n56041_, new_n51477_, RIbb2ef80_15 );
and  ( new_n56042_, new_n56041_, new_n662_ );
nor  ( new_n56043_, new_n56042_, new_n56040_ );
xnor ( new_n56044_, new_n56037_, new_n56032_ );
nor  ( new_n56045_, new_n56044_, new_n56043_ );
nor  ( new_n56046_, new_n56045_, new_n56038_ );
and  ( new_n56047_, new_n56021_, new_n56017_ );
nor  ( new_n56048_, new_n56047_, new_n56046_ );
nor  ( new_n56049_, new_n56048_, new_n56022_ );
nor  ( new_n56050_, new_n56049_, new_n56013_ );
nor  ( new_n56051_, new_n56050_, new_n56012_ );
nor  ( new_n56052_, new_n56051_, new_n55977_ );
xor  ( new_n56053_, new_n55821_, new_n55820_ );
xnor ( new_n56054_, new_n55786_, new_n55782_ );
nand ( new_n56055_, new_n56054_, new_n55791_ );
not  ( new_n56056_, new_n55787_ );
nand ( new_n56057_, new_n55793_, new_n56056_ );
and  ( new_n56058_, new_n56057_, new_n56055_ );
and  ( new_n56059_, new_n56058_, new_n56053_ );
xnor ( new_n56060_, new_n56058_, new_n56053_ );
xor  ( new_n56061_, new_n45403_, new_n5203_ );
or   ( new_n56062_, new_n56061_, new_n5604_ );
nand ( new_n56063_, new_n55898_, new_n5371_ );
and  ( new_n56064_, new_n56063_, new_n56062_ );
xor  ( new_n56065_, new_n44183_, RIbb2dbd0_57 );
nand ( new_n56066_, new_n56065_, new_n8651_ );
or   ( new_n56067_, new_n55923_, new_n8876_ );
and  ( new_n56068_, new_n56067_, new_n56066_ );
nor  ( new_n56069_, new_n56068_, new_n56064_ );
and  ( new_n56070_, new_n56068_, new_n56064_ );
xor  ( new_n56071_, new_n45119_, new_n5594_ );
nor  ( new_n56072_, new_n56071_, new_n6173_ );
and  ( new_n56073_, new_n55927_, new_n5915_ );
nor  ( new_n56074_, new_n56073_, new_n56072_ );
nor  ( new_n56075_, new_n56074_, new_n56070_ );
nor  ( new_n56076_, new_n56075_, new_n56069_ );
nor  ( new_n56077_, new_n56076_, new_n56060_ );
nor  ( new_n56078_, new_n56077_, new_n56059_ );
and  ( new_n56079_, new_n56051_, new_n55977_ );
nor  ( new_n56080_, new_n56079_, new_n56078_ );
nor  ( new_n56081_, new_n56080_, new_n56052_ );
nor  ( new_n56082_, new_n56081_, new_n55975_ );
or   ( new_n56083_, new_n56082_, new_n55974_ );
xnor ( new_n56084_, new_n55829_, new_n55827_ );
xor  ( new_n56085_, new_n56084_, new_n55908_ );
nand ( new_n56086_, new_n56085_, new_n56083_ );
nor  ( new_n56087_, new_n56085_, new_n56083_ );
xnor ( new_n56088_, new_n55750_, new_n55749_ );
xor  ( new_n56089_, new_n55760_, new_n55756_ );
xor  ( new_n56090_, new_n56089_, new_n55765_ );
nor  ( new_n56091_, new_n56090_, new_n56088_ );
nor  ( new_n56092_, new_n55880_, new_n10061_ );
xor  ( new_n56093_, new_n43952_, new_n9418_ );
nor  ( new_n56094_, new_n56093_, new_n10059_ );
or   ( new_n56095_, new_n56094_, new_n56092_ );
xor  ( new_n56096_, new_n55808_, new_n55807_ );
and  ( new_n56097_, new_n56096_, new_n56095_ );
and  ( new_n56098_, new_n55932_, new_n6508_ );
xor  ( new_n56099_, new_n44877_, RIbb2df90_49 );
and  ( new_n56100_, new_n56099_, new_n6510_ );
or   ( new_n56101_, new_n56100_, new_n56098_ );
xor  ( new_n56102_, new_n56096_, new_n56095_ );
and  ( new_n56103_, new_n56102_, new_n56101_ );
nor  ( new_n56104_, new_n56103_, new_n56097_ );
and  ( new_n56105_, new_n56090_, new_n56088_ );
nor  ( new_n56106_, new_n56105_, new_n56104_ );
or   ( new_n56107_, new_n56106_, new_n56091_ );
xor  ( new_n56108_, new_n44319_, RIbb2dcc0_55 );
nand ( new_n56109_, new_n56108_, new_n8042_ );
or   ( new_n56110_, new_n55893_, new_n8266_ );
and  ( new_n56111_, new_n56110_, new_n56109_ );
or   ( new_n56112_, new_n55888_, new_n5209_ );
xor  ( new_n56113_, new_n45738_, new_n4705_ );
or   ( new_n56114_, new_n56113_, new_n5207_ );
and  ( new_n56115_, new_n56114_, new_n56112_ );
nor  ( new_n56116_, new_n56115_, new_n56111_ );
and  ( new_n56117_, new_n56115_, new_n56111_ );
xor  ( new_n56118_, new_n45928_, new_n4292_ );
nor  ( new_n56119_, new_n56118_, new_n4709_ );
and  ( new_n56120_, new_n55834_, new_n4541_ );
nor  ( new_n56121_, new_n56120_, new_n56119_ );
nor  ( new_n56122_, new_n56121_, new_n56117_ );
nor  ( new_n56123_, new_n56122_, new_n56116_ );
or   ( new_n56124_, new_n55838_, new_n4304_ );
xor  ( new_n56125_, new_n46137_, RIbb2e440_39 );
nand ( new_n56126_, new_n56125_, new_n4034_ );
and  ( new_n56127_, new_n56126_, new_n56124_ );
xor  ( new_n56128_, new_n44681_, RIbb2dea0_51 );
nand ( new_n56129_, new_n56128_, new_n6910_ );
nand ( new_n56130_, new_n55860_, new_n6908_ );
and  ( new_n56131_, new_n56130_, new_n56129_ );
or   ( new_n56132_, new_n56131_, new_n56127_ );
and  ( new_n56133_, new_n55842_, new_n7487_ );
xor  ( new_n56134_, new_n44506_, RIbb2ddb0_53 );
and  ( new_n56135_, new_n56134_, new_n7489_ );
nor  ( new_n56136_, new_n56135_, new_n56133_ );
and  ( new_n56137_, new_n56131_, new_n56127_ );
or   ( new_n56138_, new_n56137_, new_n56136_ );
and  ( new_n56139_, new_n56138_, new_n56132_ );
nand ( new_n56140_, new_n56139_, new_n56123_ );
nor  ( new_n56141_, new_n56139_, new_n56123_ );
xor  ( new_n56142_, new_n55877_, new_n55873_ );
not  ( new_n56143_, new_n56142_ );
and  ( new_n56144_, new_n56143_, new_n55882_ );
not  ( new_n56145_, new_n55878_ );
and  ( new_n56146_, new_n55884_, new_n56145_ );
nor  ( new_n56147_, new_n56146_, new_n56144_ );
or   ( new_n56148_, new_n56147_, new_n56141_ );
and  ( new_n56149_, new_n56148_, new_n56140_ );
and  ( new_n56150_, new_n56149_, new_n56107_ );
xor  ( new_n56151_, new_n55941_, new_n55940_ );
xor  ( new_n56152_, new_n56149_, new_n56107_ );
and  ( new_n56153_, new_n56152_, new_n56151_ );
or   ( new_n56154_, new_n56153_, new_n56150_ );
xor  ( new_n56155_, new_n55776_, new_n55771_ );
xor  ( new_n56156_, new_n56155_, new_n55825_ );
nand ( new_n56157_, new_n56156_, new_n56154_ );
nor  ( new_n56158_, new_n56156_, new_n56154_ );
xor  ( new_n56159_, new_n55867_, new_n55832_ );
xor  ( new_n56160_, new_n56159_, new_n55906_ );
or   ( new_n56161_, new_n56160_, new_n56158_ );
and  ( new_n56162_, new_n56161_, new_n56157_ );
or   ( new_n56163_, new_n56162_, new_n56087_ );
and  ( new_n56164_, new_n56163_, new_n56086_ );
or   ( new_n56165_, new_n56164_, new_n55963_ );
xor  ( new_n56166_, new_n56164_, new_n55963_ );
xor  ( new_n56167_, new_n55904_, new_n55903_ );
xnor ( new_n56168_, new_n55849_, new_n55848_ );
xor  ( new_n56169_, new_n56168_, new_n55865_ );
and  ( new_n56170_, new_n56169_, new_n56167_ );
xor  ( new_n56171_, new_n49758_, new_n1126_ );
nor  ( new_n56172_, new_n56171_, new_n1366_ );
xor  ( new_n56173_, new_n50115_, new_n1126_ );
nor  ( new_n56174_, new_n56173_, new_n1364_ );
or   ( new_n56175_, new_n56174_, new_n56172_ );
xor  ( new_n56176_, new_n52902_, RIbb2f160_11 );
nor  ( new_n56177_, new_n56176_, new_n409_ );
nor  ( new_n56178_, new_n55805_, new_n411_ );
or   ( new_n56179_, new_n56178_, new_n56177_ );
nor  ( new_n56180_, new_n55799_, new_n340_ );
nor  ( new_n56181_, new_n56023_, new_n337_ );
or   ( new_n56182_, new_n56181_, new_n56180_ );
and  ( new_n56183_, new_n53694_, new_n314_ );
xor  ( new_n56184_, new_n56183_, new_n56182_ );
xor  ( new_n56185_, new_n56184_, new_n56179_ );
nand ( new_n56186_, new_n56185_, new_n56175_ );
xor  ( new_n56187_, new_n50487_, new_n893_ );
nor  ( new_n56188_, new_n56187_, new_n1137_ );
xor  ( new_n56189_, new_n50788_, new_n893_ );
nor  ( new_n56190_, new_n56189_, new_n1135_ );
or   ( new_n56191_, new_n56190_, new_n56188_ );
xor  ( new_n56192_, new_n56185_, new_n56175_ );
nand ( new_n56193_, new_n56192_, new_n56191_ );
and  ( new_n56194_, new_n56193_, new_n56186_ );
xor  ( new_n56195_, new_n43888_, new_n10052_ );
or   ( new_n56196_, new_n56195_, new_n21077_ );
or   ( new_n56197_, new_n43937_, new_n10052_ );
or   ( new_n56198_, new_n56197_, RIbb2d888_64 );
and  ( new_n56199_, new_n56198_, new_n56196_ );
nor  ( new_n56200_, new_n56199_, new_n56194_ );
xor  ( new_n56201_, new_n43985_, RIbb2dae0_59 );
and  ( new_n56202_, new_n56201_, new_n9185_ );
xor  ( new_n56203_, new_n43812_, RIbb2dae0_59 );
and  ( new_n56204_, new_n56203_, new_n9187_ );
or   ( new_n56205_, new_n56204_, new_n56202_ );
xor  ( new_n56206_, new_n56199_, new_n56194_ );
and  ( new_n56207_, new_n56206_, new_n56205_ );
nor  ( new_n56208_, new_n56207_, new_n56200_ );
not  ( new_n56209_, new_n56208_ );
xor  ( new_n56210_, new_n55863_, new_n55862_ );
and  ( new_n56211_, new_n56210_, new_n56209_ );
xor  ( new_n56212_, new_n56210_, new_n56209_ );
xnor ( new_n56213_, new_n55930_, new_n55926_ );
xor  ( new_n56214_, new_n56213_, new_n55935_ );
and  ( new_n56215_, new_n56214_, new_n56212_ );
nor  ( new_n56216_, new_n56215_, new_n56211_ );
not  ( new_n56217_, new_n56216_ );
xor  ( new_n56218_, new_n56169_, new_n56167_ );
and  ( new_n56219_, new_n56218_, new_n56217_ );
or   ( new_n56220_, new_n56219_, new_n56170_ );
xor  ( new_n56221_, new_n55944_, new_n55943_ );
and  ( new_n56222_, new_n56221_, new_n56220_ );
xor  ( new_n56223_, new_n55901_, new_n55900_ );
xor  ( new_n56224_, new_n55846_, new_n55845_ );
and  ( new_n56225_, new_n56224_, new_n56223_ );
nor  ( new_n56226_, new_n56187_, new_n1135_ );
nor  ( new_n56227_, new_n55763_, new_n1137_ );
nor  ( new_n56228_, new_n56227_, new_n56226_ );
nand ( new_n56229_, new_n55507_, new_n454_ );
or   ( new_n56230_, new_n56033_, new_n524_ );
and  ( new_n56231_, new_n56230_, new_n56229_ );
nand ( new_n56232_, new_n56183_, new_n56182_ );
nand ( new_n56233_, new_n56184_, new_n56179_ );
and  ( new_n56234_, new_n56233_, new_n56232_ );
xnor ( new_n56235_, new_n56234_, new_n56231_ );
xnor ( new_n56236_, new_n56235_, new_n56228_ );
xor  ( new_n56237_, new_n50894_, new_n745_ );
nor  ( new_n56238_, new_n56237_, new_n899_ );
xor  ( new_n56239_, new_n51142_, new_n745_ );
nor  ( new_n56240_, new_n56239_, new_n897_ );
nor  ( new_n56241_, new_n56240_, new_n56238_ );
or   ( new_n56242_, new_n56018_, new_n2809_ );
xor  ( new_n56243_, new_n47640_, new_n2421_ );
or   ( new_n56244_, new_n56243_, new_n2807_ );
and  ( new_n56245_, new_n56244_, new_n56242_ );
nor  ( new_n56246_, new_n56245_, new_n56241_ );
and  ( new_n56247_, new_n56245_, new_n56241_ );
and  ( new_n56248_, new_n55996_, new_n1474_ );
xor  ( new_n56249_, new_n49488_, RIbb2ebc0_23 );
and  ( new_n56250_, new_n56249_, new_n1476_ );
nor  ( new_n56251_, new_n56250_, new_n56248_ );
nor  ( new_n56252_, new_n56251_, new_n56247_ );
nor  ( new_n56253_, new_n56252_, new_n56246_ );
nor  ( new_n56254_, new_n56253_, new_n56236_ );
or   ( new_n56255_, new_n56015_, new_n2427_ );
xor  ( new_n56256_, new_n48291_, new_n2118_ );
or   ( new_n56257_, new_n56256_, new_n2425_ );
and  ( new_n56258_, new_n56257_, new_n56255_ );
or   ( new_n56259_, new_n55987_, new_n1846_ );
xor  ( new_n56260_, new_n49265_, new_n1583_ );
or   ( new_n56261_, new_n56260_, new_n1844_ );
and  ( new_n56262_, new_n56261_, new_n56259_ );
nor  ( new_n56263_, new_n56262_, new_n56258_ );
and  ( new_n56264_, new_n56005_, new_n2000_ );
xor  ( new_n56265_, new_n48756_, RIbb2e9e0_27 );
and  ( new_n56266_, new_n56265_, new_n2002_ );
nor  ( new_n56267_, new_n56266_, new_n56264_ );
xnor ( new_n56268_, new_n56262_, new_n56258_ );
nor  ( new_n56269_, new_n56268_, new_n56267_ );
nor  ( new_n56270_, new_n56269_, new_n56263_ );
not  ( new_n56271_, new_n56270_ );
xor  ( new_n56272_, new_n56253_, new_n56236_ );
and  ( new_n56273_, new_n56272_, new_n56271_ );
or   ( new_n56274_, new_n56273_, new_n56254_ );
xor  ( new_n56275_, new_n56224_, new_n56223_ );
and  ( new_n56276_, new_n56275_, new_n56274_ );
nor  ( new_n56277_, new_n56276_, new_n56225_ );
not  ( new_n56278_, new_n56277_ );
or   ( new_n56279_, new_n56234_, new_n56231_ );
or   ( new_n56280_, new_n56235_, new_n56228_ );
and  ( new_n56281_, new_n56280_, new_n56279_ );
or   ( new_n56282_, new_n55758_, new_n1366_ );
or   ( new_n56283_, new_n56171_, new_n1364_ );
and  ( new_n56284_, new_n56283_, new_n56282_ );
or   ( new_n56285_, new_n55737_, new_n899_ );
or   ( new_n56286_, new_n56237_, new_n897_ );
and  ( new_n56287_, new_n56286_, new_n56285_ );
or   ( new_n56288_, new_n56287_, new_n56284_ );
nor  ( new_n56289_, new_n55741_, new_n757_ );
and  ( new_n56290_, new_n56039_, new_n662_ );
nor  ( new_n56291_, new_n56290_, new_n56289_ );
and  ( new_n56292_, new_n56287_, new_n56284_ );
or   ( new_n56293_, new_n56292_, new_n56291_ );
and  ( new_n56294_, new_n56293_, new_n56288_ );
nor  ( new_n56295_, new_n56294_, new_n56281_ );
and  ( new_n56296_, new_n56201_, new_n9187_ );
nor  ( new_n56297_, new_n55648_, new_n9424_ );
or   ( new_n56298_, new_n56297_, new_n56296_ );
xor  ( new_n56299_, new_n56294_, new_n56281_ );
and  ( new_n56300_, new_n56299_, new_n56298_ );
or   ( new_n56301_, new_n56300_, new_n56295_ );
xor  ( new_n56302_, new_n55692_, new_n55691_ );
xor  ( new_n56303_, new_n56302_, new_n56301_ );
xor  ( new_n56304_, new_n55652_, new_n55651_ );
xor  ( new_n56305_, new_n56304_, new_n56303_ );
and  ( new_n56306_, new_n56305_, new_n56278_ );
xor  ( new_n56307_, new_n56305_, new_n56278_ );
xnor ( new_n56308_, new_n55967_, new_n55966_ );
xor  ( new_n56309_, new_n56308_, new_n55971_ );
and  ( new_n56310_, new_n56309_, new_n56307_ );
nor  ( new_n56311_, new_n56310_, new_n56306_ );
not  ( new_n56312_, new_n56311_ );
xor  ( new_n56313_, new_n56221_, new_n56220_ );
and  ( new_n56314_, new_n56313_, new_n56312_ );
or   ( new_n56315_, new_n56314_, new_n56222_ );
xor  ( new_n56316_, new_n55947_, new_n55946_ );
or   ( new_n56317_, new_n56316_, new_n56315_ );
and  ( new_n56318_, new_n56302_, new_n56301_ );
and  ( new_n56319_, new_n56304_, new_n56303_ );
nor  ( new_n56320_, new_n56319_, new_n56318_ );
not  ( new_n56321_, new_n56320_ );
xnor ( new_n56322_, new_n55582_, new_n55581_ );
xor  ( new_n56323_, new_n56322_, new_n55600_ );
and  ( new_n56324_, new_n56323_, new_n56321_ );
xor  ( new_n56325_, new_n56323_, new_n56321_ );
xor  ( new_n56326_, new_n55655_, new_n55654_ );
and  ( new_n56327_, new_n56326_, new_n56325_ );
or   ( new_n56328_, new_n56327_, new_n56324_ );
xor  ( new_n56329_, new_n55700_, new_n55698_ );
xnor ( new_n56330_, new_n55563_, new_n55561_ );
xor  ( new_n56331_, new_n56330_, new_n55572_ );
xor  ( new_n56332_, new_n56331_, new_n56329_ );
xor  ( new_n56333_, new_n56332_, new_n56328_ );
and  ( new_n56334_, new_n56316_, new_n56315_ );
or   ( new_n56335_, new_n56334_, new_n56333_ );
and  ( new_n56336_, new_n56335_, new_n56317_ );
nand ( new_n56337_, new_n56336_, new_n56166_ );
and  ( new_n56338_, new_n56337_, new_n56165_ );
and  ( new_n56339_, new_n56331_, new_n56329_ );
and  ( new_n56340_, new_n56332_, new_n56328_ );
or   ( new_n56341_, new_n56340_, new_n56339_ );
xor  ( new_n56342_, new_n55659_, new_n55574_ );
xor  ( new_n56343_, new_n56342_, new_n55662_ );
nand ( new_n56344_, new_n56343_, new_n56341_ );
nor  ( new_n56345_, new_n56343_, new_n56341_ );
xor  ( new_n56346_, new_n55704_, new_n55702_ );
xnor ( new_n56347_, new_n56346_, new_n55708_ );
or   ( new_n56348_, new_n56347_, new_n56345_ );
and  ( new_n56349_, new_n56348_, new_n56344_ );
nor  ( new_n56350_, new_n56349_, new_n56338_ );
and  ( new_n56351_, new_n56349_, new_n56338_ );
xor  ( new_n56352_, new_n55953_, new_n55952_ );
xor  ( new_n56353_, new_n56352_, new_n55956_ );
not  ( new_n56354_, new_n56353_ );
nor  ( new_n56355_, new_n56354_, new_n56351_ );
nor  ( new_n56356_, new_n56355_, new_n56350_ );
xor  ( new_n56357_, new_n55733_, new_n55731_ );
xnor ( new_n56358_, new_n56357_, new_n55959_ );
not  ( new_n56359_, new_n56358_ );
and  ( new_n56360_, new_n56359_, new_n56356_ );
not  ( new_n56361_, new_n56360_ );
xor  ( new_n56362_, new_n56349_, new_n56338_ );
xor  ( new_n56363_, new_n56362_, new_n56354_ );
xor  ( new_n56364_, new_n56336_, new_n56166_ );
xnor ( new_n56365_, new_n56343_, new_n56341_ );
xor  ( new_n56366_, new_n56365_, new_n56347_ );
nand ( new_n56367_, new_n56366_, new_n56364_ );
nor  ( new_n56368_, new_n56366_, new_n56364_ );
xor  ( new_n56369_, new_n56085_, new_n56083_ );
xor  ( new_n56370_, new_n56369_, new_n56162_ );
xnor ( new_n56371_, new_n56326_, new_n56325_ );
xor  ( new_n56372_, new_n55973_, new_n55964_ );
xor  ( new_n56373_, new_n56372_, new_n56081_ );
or   ( new_n56374_, new_n56373_, new_n56371_ );
and  ( new_n56375_, new_n56373_, new_n56371_ );
xor  ( new_n56376_, new_n56287_, new_n56284_ );
xnor ( new_n56377_, new_n56376_, new_n56291_ );
xor  ( new_n56378_, new_n56008_, new_n56007_ );
and  ( new_n56379_, new_n56378_, new_n56377_ );
xnor ( new_n56380_, new_n56378_, new_n56377_ );
or   ( new_n56381_, new_n55978_, new_n3119_ );
xor  ( new_n56382_, new_n47046_, new_n2797_ );
or   ( new_n56383_, new_n56382_, new_n3117_ );
and  ( new_n56384_, new_n56383_, new_n56381_ );
or   ( new_n56385_, new_n56000_, new_n3898_ );
xor  ( new_n56386_, new_n46789_, new_n3457_ );
or   ( new_n56387_, new_n56386_, new_n3896_ );
and  ( new_n56388_, new_n56387_, new_n56385_ );
nor  ( new_n56389_, new_n56388_, new_n56384_ );
and  ( new_n56390_, new_n56125_, new_n4032_ );
xor  ( new_n56391_, new_n46427_, RIbb2e440_39 );
and  ( new_n56392_, new_n56391_, new_n4034_ );
nor  ( new_n56393_, new_n56392_, new_n56390_ );
and  ( new_n56394_, new_n56388_, new_n56384_ );
nor  ( new_n56395_, new_n56394_, new_n56393_ );
nor  ( new_n56396_, new_n56395_, new_n56389_ );
nor  ( new_n56397_, new_n56396_, new_n56380_ );
nor  ( new_n56398_, new_n56397_, new_n56379_ );
xnor ( new_n56399_, new_n56299_, new_n56298_ );
or   ( new_n56400_, new_n56399_, new_n56398_ );
xnor ( new_n56401_, new_n56399_, new_n56398_ );
xnor ( new_n56402_, new_n56044_, new_n56043_ );
xor  ( new_n56403_, new_n43937_, new_n10052_ );
or   ( new_n56404_, new_n56403_, new_n21077_ );
or   ( new_n56405_, new_n43956_, new_n10052_ );
or   ( new_n56406_, new_n56405_, RIbb2d888_64 );
and  ( new_n56407_, new_n56406_, new_n56404_ );
or   ( new_n56408_, new_n56407_, new_n56402_ );
and  ( new_n56409_, new_n56128_, new_n6908_ );
xor  ( new_n56410_, new_n44785_, RIbb2dea0_51 );
and  ( new_n56411_, new_n56410_, new_n6910_ );
or   ( new_n56412_, new_n56411_, new_n56409_ );
xor  ( new_n56413_, new_n56407_, new_n56402_ );
nand ( new_n56414_, new_n56413_, new_n56412_ );
and  ( new_n56415_, new_n56414_, new_n56408_ );
xor  ( new_n56416_, new_n43914_, RIbb2dae0_59 );
nand ( new_n56417_, new_n56416_, new_n9187_ );
nand ( new_n56418_, new_n56203_, new_n9185_ );
and  ( new_n56419_, new_n56418_, new_n56417_ );
xor  ( new_n56420_, new_n46037_, new_n4292_ );
or   ( new_n56421_, new_n56420_, new_n4709_ );
or   ( new_n56422_, new_n56118_, new_n4711_ );
and  ( new_n56423_, new_n56422_, new_n56421_ );
or   ( new_n56424_, new_n56423_, new_n56419_ );
xor  ( new_n56425_, new_n44600_, RIbb2ddb0_53 );
and  ( new_n56426_, new_n56425_, new_n7489_ );
and  ( new_n56427_, new_n56134_, new_n7487_ );
nor  ( new_n56428_, new_n56427_, new_n56426_ );
xnor ( new_n56429_, new_n56423_, new_n56419_ );
or   ( new_n56430_, new_n56429_, new_n56428_ );
and  ( new_n56431_, new_n56430_, new_n56424_ );
or   ( new_n56432_, new_n56431_, new_n56415_ );
or   ( new_n56433_, new_n56071_, new_n6175_ );
xor  ( new_n56434_, new_n45204_, new_n5594_ );
or   ( new_n56435_, new_n56434_, new_n6173_ );
and  ( new_n56436_, new_n56435_, new_n56433_ );
nand ( new_n56437_, new_n56099_, new_n6508_ );
xor  ( new_n56438_, new_n44974_, RIbb2df90_49 );
nand ( new_n56439_, new_n56438_, new_n6510_ );
and  ( new_n56440_, new_n56439_, new_n56437_ );
nor  ( new_n56441_, new_n56440_, new_n56436_ );
and  ( new_n56442_, new_n56065_, new_n8649_ );
xor  ( new_n56443_, new_n44218_, RIbb2dbd0_57 );
and  ( new_n56444_, new_n56443_, new_n8651_ );
nor  ( new_n56445_, new_n56444_, new_n56442_ );
xnor ( new_n56446_, new_n56440_, new_n56436_ );
nor  ( new_n56447_, new_n56446_, new_n56445_ );
nor  ( new_n56448_, new_n56447_, new_n56441_ );
and  ( new_n56449_, new_n56431_, new_n56415_ );
or   ( new_n56450_, new_n56449_, new_n56448_ );
and  ( new_n56451_, new_n56450_, new_n56432_ );
or   ( new_n56452_, new_n56451_, new_n56401_ );
and  ( new_n56453_, new_n56452_, new_n56400_ );
xor  ( new_n56454_, new_n56102_, new_n56101_ );
xnor ( new_n56455_, new_n56131_, new_n56127_ );
xor  ( new_n56456_, new_n56455_, new_n56136_ );
and  ( new_n56457_, new_n56456_, new_n56454_ );
xor  ( new_n56458_, new_n56456_, new_n56454_ );
xnor ( new_n56459_, new_n56115_, new_n56111_ );
nand ( new_n56460_, new_n56459_, new_n56121_ );
not  ( new_n56461_, new_n56122_ );
or   ( new_n56462_, new_n56461_, new_n56116_ );
and  ( new_n56463_, new_n56462_, new_n56460_ );
and  ( new_n56464_, new_n56463_, new_n56458_ );
or   ( new_n56465_, new_n56464_, new_n56457_ );
xor  ( new_n56466_, new_n56076_, new_n56060_ );
nand ( new_n56467_, new_n56466_, new_n56465_ );
nor  ( new_n56468_, new_n56466_, new_n56465_ );
nor  ( new_n56469_, new_n56176_, new_n411_ );
xor  ( new_n56470_, new_n52908_, RIbb2f160_11 );
nor  ( new_n56471_, new_n56470_, new_n409_ );
or   ( new_n56472_, new_n56471_, new_n56469_ );
xor  ( new_n56473_, new_n56031_, new_n56029_ );
nand ( new_n56474_, new_n56473_, new_n56472_ );
nor  ( new_n56475_, new_n56035_, new_n526_ );
xor  ( new_n56476_, new_n52293_, RIbb2f070_13 );
nor  ( new_n56477_, new_n56476_, new_n524_ );
or   ( new_n56478_, new_n56477_, new_n56475_ );
xor  ( new_n56479_, new_n56473_, new_n56472_ );
nand ( new_n56480_, new_n56479_, new_n56478_ );
and  ( new_n56481_, new_n56480_, new_n56474_ );
or   ( new_n56482_, new_n55982_, new_n3463_ );
xor  ( new_n56483_, new_n46958_, RIbb2e620_35 );
nand ( new_n56484_, new_n56483_, new_n3293_ );
and  ( new_n56485_, new_n56484_, new_n56482_ );
nor  ( new_n56486_, new_n56485_, new_n56481_ );
nor  ( new_n56487_, new_n56093_, new_n10061_ );
xor  ( new_n56488_, new_n43985_, RIbb2d9f0_61 );
and  ( new_n56489_, new_n56488_, new_n9740_ );
nor  ( new_n56490_, new_n56489_, new_n56487_ );
not  ( new_n56491_, new_n56490_ );
xor  ( new_n56492_, new_n56485_, new_n56481_ );
and  ( new_n56493_, new_n56492_, new_n56491_ );
nor  ( new_n56494_, new_n56493_, new_n56486_ );
not  ( new_n56495_, new_n56494_ );
xor  ( new_n56496_, new_n56206_, new_n56205_ );
and  ( new_n56497_, new_n56496_, new_n56495_ );
xor  ( new_n56498_, new_n56496_, new_n56495_ );
xnor ( new_n56499_, new_n56068_, new_n56064_ );
nand ( new_n56500_, new_n56499_, new_n56074_ );
not  ( new_n56501_, new_n56075_ );
or   ( new_n56502_, new_n56501_, new_n56069_ );
and  ( new_n56503_, new_n56502_, new_n56500_ );
and  ( new_n56504_, new_n56503_, new_n56498_ );
nor  ( new_n56505_, new_n56504_, new_n56497_ );
or   ( new_n56506_, new_n56505_, new_n56468_ );
and  ( new_n56507_, new_n56506_, new_n56467_ );
nor  ( new_n56508_, new_n56507_, new_n56453_ );
and  ( new_n56509_, new_n56507_, new_n56453_ );
xor  ( new_n56510_, new_n56010_, new_n55994_ );
and  ( new_n56511_, new_n56510_, new_n56049_ );
not  ( new_n56512_, new_n56012_ );
and  ( new_n56513_, new_n56050_, new_n56512_ );
or   ( new_n56514_, new_n56513_, new_n56511_ );
xnor ( new_n56515_, new_n55991_, new_n55990_ );
xor  ( new_n56516_, new_n45597_, new_n4705_ );
or   ( new_n56517_, new_n56516_, new_n5207_ );
or   ( new_n56518_, new_n56113_, new_n5209_ );
and  ( new_n56519_, new_n56518_, new_n56517_ );
or   ( new_n56520_, new_n56061_, new_n5606_ );
xor  ( new_n56521_, new_n45584_, new_n5203_ );
or   ( new_n56522_, new_n56521_, new_n5604_ );
and  ( new_n56523_, new_n56522_, new_n56520_ );
or   ( new_n56524_, new_n56523_, new_n56519_ );
xor  ( new_n56525_, new_n44407_, RIbb2dcc0_55 );
and  ( new_n56526_, new_n56525_, new_n8042_ );
and  ( new_n56527_, new_n56108_, new_n8040_ );
nor  ( new_n56528_, new_n56527_, new_n56526_ );
and  ( new_n56529_, new_n56523_, new_n56519_ );
or   ( new_n56530_, new_n56529_, new_n56528_ );
and  ( new_n56531_, new_n56530_, new_n56524_ );
or   ( new_n56532_, new_n56531_, new_n56515_ );
nand ( new_n56533_, new_n56531_, new_n56515_ );
xor  ( new_n56534_, new_n56021_, new_n56017_ );
xnor ( new_n56535_, new_n56534_, new_n56046_ );
nand ( new_n56536_, new_n56535_, new_n56533_ );
and  ( new_n56537_, new_n56536_, new_n56532_ );
and  ( new_n56538_, new_n56537_, new_n56514_ );
nor  ( new_n56539_, new_n56537_, new_n56514_ );
not  ( new_n56540_, new_n56539_ );
xor  ( new_n56541_, new_n56090_, new_n56088_ );
xor  ( new_n56542_, new_n56541_, new_n56104_ );
and  ( new_n56543_, new_n56542_, new_n56540_ );
nor  ( new_n56544_, new_n56543_, new_n56538_ );
not  ( new_n56545_, new_n56544_ );
nor  ( new_n56546_, new_n56545_, new_n56509_ );
nor  ( new_n56547_, new_n56546_, new_n56508_ );
or   ( new_n56548_, new_n56547_, new_n56375_ );
and  ( new_n56549_, new_n56548_, new_n56374_ );
nor  ( new_n56550_, new_n56549_, new_n56370_ );
and  ( new_n56551_, new_n56549_, new_n56370_ );
xnor ( new_n56552_, new_n56152_, new_n56151_ );
xor  ( new_n56553_, new_n56051_, new_n55977_ );
xor  ( new_n56554_, new_n56553_, new_n56078_ );
nor  ( new_n56555_, new_n56554_, new_n56552_ );
nand ( new_n56556_, new_n56554_, new_n56552_ );
xor  ( new_n56557_, new_n56218_, new_n56217_ );
and  ( new_n56558_, new_n56557_, new_n56556_ );
or   ( new_n56559_, new_n56558_, new_n56555_ );
xnor ( new_n56560_, new_n56156_, new_n56154_ );
xor  ( new_n56561_, new_n56560_, new_n56160_ );
and  ( new_n56562_, new_n56561_, new_n56559_ );
nor  ( new_n56563_, new_n56561_, new_n56559_ );
not  ( new_n56564_, new_n56563_ );
xor  ( new_n56565_, new_n56313_, new_n56312_ );
and  ( new_n56566_, new_n56565_, new_n56564_ );
nor  ( new_n56567_, new_n56566_, new_n56562_ );
nor  ( new_n56568_, new_n56567_, new_n56551_ );
nor  ( new_n56569_, new_n56568_, new_n56550_ );
or   ( new_n56570_, new_n56569_, new_n56368_ );
and  ( new_n56571_, new_n56570_, new_n56367_ );
nor  ( new_n56572_, new_n56571_, new_n56363_ );
and  ( new_n56573_, new_n56571_, new_n56363_ );
xor  ( new_n56574_, new_n56316_, new_n56315_ );
xor  ( new_n56575_, new_n56574_, new_n56333_ );
xnor ( new_n56576_, new_n56549_, new_n56370_ );
xor  ( new_n56577_, new_n56576_, new_n56567_ );
nor  ( new_n56578_, new_n56577_, new_n56575_ );
xnor ( new_n56579_, new_n56214_, new_n56212_ );
xnor ( new_n56580_, new_n56139_, new_n56123_ );
xor  ( new_n56581_, new_n56580_, new_n56147_ );
or   ( new_n56582_, new_n56581_, new_n56579_ );
xor  ( new_n56583_, new_n56275_, new_n56274_ );
xor  ( new_n56584_, new_n56581_, new_n56579_ );
nand ( new_n56585_, new_n56584_, new_n56583_ );
and  ( new_n56586_, new_n56585_, new_n56582_ );
xor  ( new_n56587_, new_n56272_, new_n56271_ );
xor  ( new_n56588_, new_n56396_, new_n56380_ );
nand ( new_n56589_, new_n56588_, new_n56587_ );
xnor ( new_n56590_, new_n56588_, new_n56587_ );
xor  ( new_n56591_, new_n44877_, new_n6635_ );
or   ( new_n56592_, new_n56591_, new_n7184_ );
nand ( new_n56593_, new_n56410_, new_n6908_ );
and  ( new_n56594_, new_n56593_, new_n56592_ );
xor  ( new_n56595_, new_n44681_, RIbb2ddb0_53 );
nand ( new_n56596_, new_n56595_, new_n7489_ );
nand ( new_n56597_, new_n56425_, new_n7487_ );
and  ( new_n56598_, new_n56597_, new_n56596_ );
nor  ( new_n56599_, new_n56598_, new_n56594_ );
and  ( new_n56600_, new_n56598_, new_n56594_ );
xor  ( new_n56601_, new_n44183_, RIbb2dae0_59 );
and  ( new_n56602_, new_n56601_, new_n9187_ );
and  ( new_n56603_, new_n56416_, new_n9185_ );
nor  ( new_n56604_, new_n56603_, new_n56602_ );
nor  ( new_n56605_, new_n56604_, new_n56600_ );
or   ( new_n56606_, new_n56605_, new_n56599_ );
xnor ( new_n56607_, new_n56388_, new_n56384_ );
nand ( new_n56608_, new_n56607_, new_n56393_ );
not  ( new_n56609_, new_n56395_ );
or   ( new_n56610_, new_n56609_, new_n56389_ );
and  ( new_n56611_, new_n56610_, new_n56608_ );
nand ( new_n56612_, new_n56611_, new_n56606_ );
or   ( new_n56613_, new_n56611_, new_n56606_ );
xor  ( new_n56614_, new_n56492_, new_n56491_ );
nand ( new_n56615_, new_n56614_, new_n56613_ );
and  ( new_n56616_, new_n56615_, new_n56612_ );
or   ( new_n56617_, new_n56616_, new_n56590_ );
and  ( new_n56618_, new_n56617_, new_n56589_ );
xor  ( new_n56619_, new_n49758_, new_n1355_ );
or   ( new_n56620_, new_n56619_, new_n1593_ );
nand ( new_n56621_, new_n56249_, new_n1474_ );
and  ( new_n56622_, new_n56621_, new_n56620_ );
or   ( new_n56623_, new_n56189_, new_n1137_ );
xor  ( new_n56624_, new_n50894_, new_n893_ );
or   ( new_n56625_, new_n56624_, new_n1135_ );
and  ( new_n56626_, new_n56625_, new_n56623_ );
or   ( new_n56627_, new_n56626_, new_n56622_ );
nor  ( new_n56628_, new_n56239_, new_n899_ );
xor  ( new_n56629_, new_n51446_, RIbb2ee90_17 );
and  ( new_n56630_, new_n56629_, new_n822_ );
nor  ( new_n56631_, new_n56630_, new_n56628_ );
xnor ( new_n56632_, new_n56626_, new_n56622_ );
or   ( new_n56633_, new_n56632_, new_n56631_ );
and  ( new_n56634_, new_n56633_, new_n56627_ );
nor  ( new_n56635_, new_n56470_, new_n411_ );
xor  ( new_n56636_, new_n53306_, RIbb2f160_11 );
nor  ( new_n56637_, new_n56636_, new_n409_ );
or   ( new_n56638_, new_n56637_, new_n56635_ );
and  ( new_n56639_, new_n53694_, new_n334_ );
nand ( new_n56640_, new_n56639_, new_n56638_ );
xor  ( new_n56641_, new_n52902_, RIbb2f070_13 );
nor  ( new_n56642_, new_n56641_, new_n524_ );
nor  ( new_n56643_, new_n56476_, new_n526_ );
or   ( new_n56644_, new_n56643_, new_n56642_ );
xor  ( new_n56645_, new_n56639_, new_n56638_ );
nand ( new_n56646_, new_n56645_, new_n56644_ );
and  ( new_n56647_, new_n56646_, new_n56640_ );
xor  ( new_n56648_, new_n51758_, new_n520_ );
or   ( new_n56649_, new_n56648_, new_n755_ );
nand ( new_n56650_, new_n56041_, new_n660_ );
and  ( new_n56651_, new_n56650_, new_n56649_ );
or   ( new_n56652_, new_n56651_, new_n56647_ );
nor  ( new_n56653_, new_n56173_, new_n1366_ );
xor  ( new_n56654_, new_n50487_, new_n1126_ );
nor  ( new_n56655_, new_n56654_, new_n1364_ );
or   ( new_n56656_, new_n56655_, new_n56653_ );
xor  ( new_n56657_, new_n56651_, new_n56647_ );
nand ( new_n56658_, new_n56657_, new_n56656_ );
and  ( new_n56659_, new_n56658_, new_n56652_ );
or   ( new_n56660_, new_n56659_, new_n56634_ );
xor  ( new_n56661_, new_n48518_, new_n2118_ );
or   ( new_n56662_, new_n56661_, new_n2425_ );
or   ( new_n56663_, new_n56256_, new_n2427_ );
and  ( new_n56664_, new_n56663_, new_n56662_ );
or   ( new_n56665_, new_n56243_, new_n2809_ );
xor  ( new_n56666_, new_n48039_, new_n2421_ );
or   ( new_n56667_, new_n56666_, new_n2807_ );
and  ( new_n56668_, new_n56667_, new_n56665_ );
nor  ( new_n56669_, new_n56668_, new_n56664_ );
xor  ( new_n56670_, new_n48908_, new_n1840_ );
nor  ( new_n56671_, new_n56670_, new_n2122_ );
and  ( new_n56672_, new_n56265_, new_n2000_ );
or   ( new_n56673_, new_n56672_, new_n56671_ );
xor  ( new_n56674_, new_n56668_, new_n56664_ );
and  ( new_n56675_, new_n56674_, new_n56673_ );
nor  ( new_n56676_, new_n56675_, new_n56669_ );
not  ( new_n56677_, new_n56676_ );
xor  ( new_n56678_, new_n56659_, new_n56634_ );
nand ( new_n56679_, new_n56678_, new_n56677_ );
and  ( new_n56680_, new_n56679_, new_n56660_ );
xnor ( new_n56681_, new_n56245_, new_n56241_ );
and  ( new_n56682_, new_n56681_, new_n56251_ );
not  ( new_n56683_, new_n56246_ );
and  ( new_n56684_, new_n56252_, new_n56683_ );
or   ( new_n56685_, new_n56684_, new_n56682_ );
or   ( new_n56686_, new_n56382_, new_n3119_ );
xor  ( new_n56687_, new_n47296_, new_n2797_ );
or   ( new_n56688_, new_n56687_, new_n3117_ );
and  ( new_n56689_, new_n56688_, new_n56686_ );
nand ( new_n56690_, new_n56391_, new_n4032_ );
xor  ( new_n56691_, new_n46619_, new_n3892_ );
or   ( new_n56692_, new_n56691_, new_n4302_ );
and  ( new_n56693_, new_n56692_, new_n56690_ );
or   ( new_n56694_, new_n56693_, new_n56689_ );
nor  ( new_n56695_, new_n56260_, new_n1846_ );
xor  ( new_n56696_, new_n49427_, RIbb2ead0_25 );
and  ( new_n56697_, new_n56696_, new_n1741_ );
nor  ( new_n56698_, new_n56697_, new_n56695_ );
and  ( new_n56699_, new_n56693_, new_n56689_ );
or   ( new_n56700_, new_n56699_, new_n56698_ );
and  ( new_n56701_, new_n56700_, new_n56694_ );
or   ( new_n56702_, new_n56701_, new_n56685_ );
and  ( new_n56703_, new_n56701_, new_n56685_ );
nor  ( new_n56704_, new_n56386_, new_n3898_ );
xor  ( new_n56705_, new_n46962_, new_n3457_ );
nor  ( new_n56706_, new_n56705_, new_n3896_ );
or   ( new_n56707_, new_n56706_, new_n56704_ );
xor  ( new_n56708_, new_n56479_, new_n56478_ );
and  ( new_n56709_, new_n56708_, new_n56707_ );
xor  ( new_n56710_, new_n47303_, new_n3113_ );
nor  ( new_n56711_, new_n56710_, new_n3461_ );
and  ( new_n56712_, new_n56483_, new_n3291_ );
or   ( new_n56713_, new_n56712_, new_n56711_ );
xor  ( new_n56714_, new_n56708_, new_n56707_ );
and  ( new_n56715_, new_n56714_, new_n56713_ );
nor  ( new_n56716_, new_n56715_, new_n56709_ );
or   ( new_n56717_, new_n56716_, new_n56703_ );
and  ( new_n56718_, new_n56717_, new_n56702_ );
or   ( new_n56719_, new_n56718_, new_n56680_ );
and  ( new_n56720_, new_n56718_, new_n56680_ );
or   ( new_n56721_, new_n56521_, new_n5606_ );
xor  ( new_n56722_, new_n45738_, new_n5203_ );
or   ( new_n56723_, new_n56722_, new_n5604_ );
and  ( new_n56724_, new_n56723_, new_n56721_ );
xor  ( new_n56725_, new_n45403_, new_n5594_ );
or   ( new_n56726_, new_n56725_, new_n6173_ );
or   ( new_n56727_, new_n56434_, new_n6175_ );
and  ( new_n56728_, new_n56727_, new_n56726_ );
nor  ( new_n56729_, new_n56728_, new_n56724_ );
nand ( new_n56730_, new_n56728_, new_n56724_ );
xor  ( new_n56731_, new_n44319_, RIbb2dbd0_57 );
and  ( new_n56732_, new_n56731_, new_n8651_ );
and  ( new_n56733_, new_n56443_, new_n8649_ );
or   ( new_n56734_, new_n56733_, new_n56732_ );
and  ( new_n56735_, new_n56734_, new_n56730_ );
or   ( new_n56736_, new_n56735_, new_n56729_ );
xor  ( new_n56737_, new_n56192_, new_n56191_ );
and  ( new_n56738_, new_n56737_, new_n56736_ );
nor  ( new_n56739_, new_n53695_, new_n43906_ );
or   ( new_n56740_, new_n56739_, new_n328_ );
or   ( new_n56741_, new_n56636_, new_n411_ );
and  ( new_n56742_, new_n43905_, RIbb2f160_11 );
and  ( new_n56743_, new_n53694_, RIbb2f070_13 );
nor  ( new_n56744_, new_n56743_, new_n56742_ );
and  ( new_n56745_, RIbb2f0e8_12, new_n325_ );
nor  ( new_n56746_, new_n53694_, RIbb2f070_13 );
nor  ( new_n56747_, new_n56746_, new_n56745_ );
or   ( new_n56748_, new_n56747_, new_n56744_ );
and  ( new_n56749_, new_n56748_, new_n56741_ );
or   ( new_n56750_, new_n56749_, new_n56740_ );
or   ( new_n56751_, new_n56648_, new_n757_ );
xor  ( new_n56752_, new_n52280_, new_n520_ );
or   ( new_n56753_, new_n56752_, new_n755_ );
and  ( new_n56754_, new_n56753_, new_n56751_ );
or   ( new_n56755_, new_n56754_, new_n56750_ );
and  ( new_n56756_, new_n56629_, new_n820_ );
xor  ( new_n56757_, new_n51477_, RIbb2ee90_17 );
and  ( new_n56758_, new_n56757_, new_n822_ );
or   ( new_n56759_, new_n56758_, new_n56756_ );
xor  ( new_n56760_, new_n56754_, new_n56750_ );
nand ( new_n56761_, new_n56760_, new_n56759_ );
and  ( new_n56762_, new_n56761_, new_n56755_ );
xor  ( new_n56763_, new_n43812_, RIbb2d9f0_61 );
nand ( new_n56764_, new_n56763_, new_n9740_ );
nand ( new_n56765_, new_n56488_, new_n9738_ );
and  ( new_n56766_, new_n56765_, new_n56764_ );
nor  ( new_n56767_, new_n56766_, new_n56762_ );
and  ( new_n56768_, new_n56438_, new_n6508_ );
xor  ( new_n56769_, new_n45119_, new_n6163_ );
nor  ( new_n56770_, new_n56769_, new_n6645_ );
nor  ( new_n56771_, new_n56770_, new_n56768_ );
not  ( new_n56772_, new_n56771_ );
xor  ( new_n56773_, new_n56766_, new_n56762_ );
and  ( new_n56774_, new_n56773_, new_n56772_ );
or   ( new_n56775_, new_n56774_, new_n56767_ );
xor  ( new_n56776_, new_n56737_, new_n56736_ );
and  ( new_n56777_, new_n56776_, new_n56775_ );
nor  ( new_n56778_, new_n56777_, new_n56738_ );
or   ( new_n56779_, new_n56778_, new_n56720_ );
and  ( new_n56780_, new_n56779_, new_n56719_ );
or   ( new_n56781_, new_n56780_, new_n56618_ );
and  ( new_n56782_, new_n56780_, new_n56618_ );
xor  ( new_n56783_, new_n56537_, new_n56514_ );
xor  ( new_n56784_, new_n56783_, new_n56542_ );
or   ( new_n56785_, new_n56784_, new_n56782_ );
and  ( new_n56786_, new_n56785_, new_n56781_ );
nor  ( new_n56787_, new_n56786_, new_n56586_ );
xor  ( new_n56788_, new_n56309_, new_n56307_ );
xor  ( new_n56789_, new_n56786_, new_n56586_ );
and  ( new_n56790_, new_n56789_, new_n56788_ );
nor  ( new_n56791_, new_n56790_, new_n56787_ );
not  ( new_n56792_, new_n56791_ );
xnor ( new_n56793_, new_n56373_, new_n56371_ );
xor  ( new_n56794_, new_n56793_, new_n56547_ );
nor  ( new_n56795_, new_n56794_, new_n56792_ );
xor  ( new_n56796_, new_n56794_, new_n56792_ );
xnor ( new_n56797_, new_n56554_, new_n56552_ );
xor  ( new_n56798_, new_n56797_, new_n56557_ );
xor  ( new_n56799_, new_n56507_, new_n56453_ );
xor  ( new_n56800_, new_n56799_, new_n56545_ );
or   ( new_n56801_, new_n56800_, new_n56798_ );
nand ( new_n56802_, new_n56800_, new_n56798_ );
xor  ( new_n56803_, new_n56451_, new_n56401_ );
xnor ( new_n56804_, new_n56466_, new_n56465_ );
xor  ( new_n56805_, new_n56804_, new_n56505_ );
nor  ( new_n56806_, new_n56805_, new_n56803_ );
and  ( new_n56807_, new_n56805_, new_n56803_ );
not  ( new_n56808_, new_n56807_ );
xnor ( new_n56809_, new_n56268_, new_n56267_ );
or   ( new_n56810_, new_n56420_, new_n4711_ );
xor  ( new_n56811_, new_n46137_, RIbb2e350_41 );
nand ( new_n56812_, new_n56811_, new_n4543_ );
and  ( new_n56813_, new_n56812_, new_n56810_ );
or   ( new_n56814_, new_n56516_, new_n5209_ );
xor  ( new_n56815_, new_n45928_, new_n4705_ );
or   ( new_n56816_, new_n56815_, new_n5207_ );
and  ( new_n56817_, new_n56816_, new_n56814_ );
or   ( new_n56818_, new_n56817_, new_n56813_ );
and  ( new_n56819_, new_n56817_, new_n56813_ );
and  ( new_n56820_, new_n56525_, new_n8040_ );
xor  ( new_n56821_, new_n44506_, RIbb2dcc0_55 );
and  ( new_n56822_, new_n56821_, new_n8042_ );
nor  ( new_n56823_, new_n56822_, new_n56820_ );
or   ( new_n56824_, new_n56823_, new_n56819_ );
and  ( new_n56825_, new_n56824_, new_n56818_ );
nor  ( new_n56826_, new_n56825_, new_n56809_ );
nand ( new_n56827_, new_n56825_, new_n56809_ );
xor  ( new_n56828_, new_n56413_, new_n56412_ );
and  ( new_n56829_, new_n56828_, new_n56827_ );
or   ( new_n56830_, new_n56829_, new_n56826_ );
xnor ( new_n56831_, new_n56446_, new_n56445_ );
xor  ( new_n56832_, new_n50115_, new_n1355_ );
nor  ( new_n56833_, new_n56832_, new_n1593_ );
nor  ( new_n56834_, new_n56619_, new_n1595_ );
or   ( new_n56835_, new_n56834_, new_n56833_ );
xor  ( new_n56836_, new_n56645_, new_n56644_ );
and  ( new_n56837_, new_n56836_, new_n56835_ );
xor  ( new_n56838_, new_n50788_, new_n1126_ );
nor  ( new_n56839_, new_n56838_, new_n1364_ );
nor  ( new_n56840_, new_n56654_, new_n1366_ );
or   ( new_n56841_, new_n56840_, new_n56839_ );
xor  ( new_n56842_, new_n56836_, new_n56835_ );
and  ( new_n56843_, new_n56842_, new_n56841_ );
nor  ( new_n56844_, new_n56843_, new_n56837_ );
xnor ( new_n56845_, new_n56657_, new_n56656_ );
or   ( new_n56846_, new_n56845_, new_n56844_ );
xnor ( new_n56847_, new_n56845_, new_n56844_ );
xor  ( new_n56848_, new_n43956_, new_n10052_ );
or   ( new_n56849_, new_n56848_, new_n21077_ );
or   ( new_n56850_, new_n43952_, new_n10052_ );
or   ( new_n56851_, new_n56850_, RIbb2d888_64 );
and  ( new_n56852_, new_n56851_, new_n56849_ );
or   ( new_n56853_, new_n56852_, new_n56847_ );
and  ( new_n56854_, new_n56853_, new_n56846_ );
nand ( new_n56855_, new_n56854_, new_n56831_ );
nor  ( new_n56856_, new_n56854_, new_n56831_ );
xor  ( new_n56857_, new_n56523_, new_n56519_ );
xnor ( new_n56858_, new_n56857_, new_n56528_ );
or   ( new_n56859_, new_n56858_, new_n56856_ );
and  ( new_n56860_, new_n56859_, new_n56855_ );
and  ( new_n56861_, new_n56860_, new_n56830_ );
xor  ( new_n56862_, new_n56860_, new_n56830_ );
xnor ( new_n56863_, new_n56431_, new_n56415_ );
xor  ( new_n56864_, new_n56863_, new_n56448_ );
and  ( new_n56865_, new_n56864_, new_n56862_ );
nor  ( new_n56866_, new_n56865_, new_n56861_ );
and  ( new_n56867_, new_n56866_, new_n56808_ );
nor  ( new_n56868_, new_n56867_, new_n56806_ );
nand ( new_n56869_, new_n56868_, new_n56802_ );
and  ( new_n56870_, new_n56869_, new_n56801_ );
and  ( new_n56871_, new_n56870_, new_n56796_ );
nor  ( new_n56872_, new_n56871_, new_n56795_ );
not  ( new_n56873_, new_n56872_ );
xor  ( new_n56874_, new_n56577_, new_n56575_ );
and  ( new_n56875_, new_n56874_, new_n56873_ );
nor  ( new_n56876_, new_n56875_, new_n56578_ );
xor  ( new_n56877_, new_n56366_, new_n56364_ );
xnor ( new_n56878_, new_n56877_, new_n56569_ );
and  ( new_n56879_, new_n56878_, new_n56876_ );
nor  ( new_n56880_, new_n56878_, new_n56876_ );
xor  ( new_n56881_, new_n56874_, new_n56873_ );
xnor ( new_n56882_, new_n56870_, new_n56796_ );
xor  ( new_n56883_, new_n56561_, new_n56559_ );
xor  ( new_n56884_, new_n56883_, new_n56565_ );
nand ( new_n56885_, new_n56884_, new_n56882_ );
nor  ( new_n56886_, new_n56884_, new_n56882_ );
xnor ( new_n56887_, new_n56789_, new_n56788_ );
xor  ( new_n56888_, new_n56780_, new_n56618_ );
xor  ( new_n56889_, new_n56888_, new_n56784_ );
xor  ( new_n56890_, new_n56805_, new_n56803_ );
xor  ( new_n56891_, new_n56890_, new_n56866_ );
or   ( new_n56892_, new_n56891_, new_n56889_ );
and  ( new_n56893_, new_n56891_, new_n56889_ );
xor  ( new_n56894_, new_n56616_, new_n56590_ );
xor  ( new_n56895_, new_n56864_, new_n56862_ );
nor  ( new_n56896_, new_n56895_, new_n56894_ );
nand ( new_n56897_, new_n56895_, new_n56894_ );
xnor ( new_n56898_, new_n56693_, new_n56689_ );
xor  ( new_n56899_, new_n56898_, new_n56698_ );
xor  ( new_n56900_, new_n56728_, new_n56724_ );
xor  ( new_n56901_, new_n56900_, new_n56734_ );
or   ( new_n56902_, new_n56901_, new_n56899_ );
and  ( new_n56903_, new_n56901_, new_n56899_ );
xor  ( new_n56904_, new_n56674_, new_n56673_ );
or   ( new_n56905_, new_n56904_, new_n56903_ );
and  ( new_n56906_, new_n56905_, new_n56902_ );
xor  ( new_n56907_, new_n56825_, new_n56809_ );
xor  ( new_n56908_, new_n56907_, new_n56828_ );
and  ( new_n56909_, new_n56908_, new_n56906_ );
nor  ( new_n56910_, new_n56908_, new_n56906_ );
xor  ( new_n56911_, new_n56598_, new_n56594_ );
xor  ( new_n56912_, new_n56911_, new_n56604_ );
xor  ( new_n56913_, new_n44218_, new_n8870_ );
or   ( new_n56914_, new_n56913_, new_n9422_ );
nand ( new_n56915_, new_n56601_, new_n9185_ );
and  ( new_n56916_, new_n56915_, new_n56914_ );
xor  ( new_n56917_, new_n44974_, RIbb2dea0_51 );
nand ( new_n56918_, new_n56917_, new_n6910_ );
or   ( new_n56919_, new_n56591_, new_n7186_ );
and  ( new_n56920_, new_n56919_, new_n56918_ );
or   ( new_n56921_, new_n56920_, new_n56916_ );
xor  ( new_n56922_, new_n51142_, new_n893_ );
or   ( new_n56923_, new_n56922_, new_n1137_ );
xor  ( new_n56924_, new_n51446_, RIbb2eda0_19 );
nand ( new_n56925_, new_n56924_, new_n1042_ );
and  ( new_n56926_, new_n56925_, new_n56923_ );
xor  ( new_n56927_, new_n49758_, new_n1583_ );
or   ( new_n56928_, new_n56927_, new_n1844_ );
xor  ( new_n56929_, new_n49488_, RIbb2ead0_25 );
nand ( new_n56930_, new_n56929_, new_n1739_ );
and  ( new_n56931_, new_n56930_, new_n56928_ );
nor  ( new_n56932_, new_n56931_, new_n56926_ );
xor  ( new_n56933_, new_n50894_, new_n1126_ );
nor  ( new_n56934_, new_n56933_, new_n1364_ );
nor  ( new_n56935_, new_n56838_, new_n1366_ );
or   ( new_n56936_, new_n56935_, new_n56934_ );
xor  ( new_n56937_, new_n56931_, new_n56926_ );
and  ( new_n56938_, new_n56937_, new_n56936_ );
nor  ( new_n56939_, new_n56938_, new_n56932_ );
and  ( new_n56940_, new_n56920_, new_n56916_ );
or   ( new_n56941_, new_n56940_, new_n56939_ );
and  ( new_n56942_, new_n56941_, new_n56921_ );
nor  ( new_n56943_, new_n56942_, new_n56912_ );
and  ( new_n56944_, new_n56942_, new_n56912_ );
not  ( new_n56945_, new_n56944_ );
xor  ( new_n56946_, new_n56773_, new_n56772_ );
and  ( new_n56947_, new_n56946_, new_n56945_ );
nor  ( new_n56948_, new_n56947_, new_n56943_ );
nor  ( new_n56949_, new_n56948_, new_n56910_ );
nor  ( new_n56950_, new_n56949_, new_n56909_ );
and  ( new_n56951_, new_n56950_, new_n56897_ );
or   ( new_n56952_, new_n56951_, new_n56896_ );
or   ( new_n56953_, new_n56952_, new_n56893_ );
and  ( new_n56954_, new_n56953_, new_n56892_ );
nor  ( new_n56955_, new_n56954_, new_n56887_ );
and  ( new_n56956_, new_n56954_, new_n56887_ );
xnor ( new_n56957_, new_n56429_, new_n56428_ );
xnor ( new_n56958_, new_n56632_, new_n56631_ );
or   ( new_n56959_, new_n56922_, new_n1135_ );
or   ( new_n56960_, new_n56624_, new_n1137_ );
and  ( new_n56961_, new_n56960_, new_n56959_ );
xor  ( new_n56962_, new_n48291_, new_n2421_ );
or   ( new_n56963_, new_n56962_, new_n2807_ );
or   ( new_n56964_, new_n56666_, new_n2809_ );
and  ( new_n56965_, new_n56964_, new_n56963_ );
or   ( new_n56966_, new_n56965_, new_n56961_ );
and  ( new_n56967_, new_n56696_, new_n1739_ );
and  ( new_n56968_, new_n56929_, new_n1741_ );
nor  ( new_n56969_, new_n56968_, new_n56967_ );
and  ( new_n56970_, new_n56965_, new_n56961_ );
or   ( new_n56971_, new_n56970_, new_n56969_ );
and  ( new_n56972_, new_n56971_, new_n56966_ );
or   ( new_n56973_, new_n56972_, new_n56958_ );
and  ( new_n56974_, new_n56972_, new_n56958_ );
xor  ( new_n56975_, new_n47640_, new_n2797_ );
or   ( new_n56976_, new_n56975_, new_n3117_ );
or   ( new_n56977_, new_n56687_, new_n3119_ );
and  ( new_n56978_, new_n56977_, new_n56976_ );
xor  ( new_n56979_, new_n48756_, new_n2118_ );
or   ( new_n56980_, new_n56979_, new_n2425_ );
or   ( new_n56981_, new_n56661_, new_n2427_ );
and  ( new_n56982_, new_n56981_, new_n56980_ );
or   ( new_n56983_, new_n56982_, new_n56978_ );
nor  ( new_n56984_, new_n56670_, new_n2124_ );
xor  ( new_n56985_, new_n49265_, new_n1840_ );
nor  ( new_n56986_, new_n56985_, new_n2122_ );
nor  ( new_n56987_, new_n56986_, new_n56984_ );
and  ( new_n56988_, new_n56982_, new_n56978_ );
or   ( new_n56989_, new_n56988_, new_n56987_ );
and  ( new_n56990_, new_n56989_, new_n56983_ );
or   ( new_n56991_, new_n56990_, new_n56974_ );
and  ( new_n56992_, new_n56991_, new_n56973_ );
and  ( new_n56993_, new_n56992_, new_n56957_ );
xor  ( new_n56994_, new_n56678_, new_n56677_ );
nor  ( new_n56995_, new_n56992_, new_n56957_ );
nor  ( new_n56996_, new_n56995_, new_n56994_ );
nor  ( new_n56997_, new_n56996_, new_n56993_ );
xor  ( new_n56998_, new_n56531_, new_n56515_ );
xor  ( new_n56999_, new_n56998_, new_n56535_ );
and  ( new_n57000_, new_n56999_, new_n56997_ );
xor  ( new_n57001_, new_n56999_, new_n56997_ );
xor  ( new_n57002_, new_n56463_, new_n56458_ );
and  ( new_n57003_, new_n57002_, new_n57001_ );
or   ( new_n57004_, new_n57003_, new_n57000_ );
xor  ( new_n57005_, new_n56584_, new_n56583_ );
and  ( new_n57006_, new_n57005_, new_n57004_ );
nor  ( new_n57007_, new_n57005_, new_n57004_ );
xor  ( new_n57008_, new_n56503_, new_n56498_ );
xnor ( new_n57009_, new_n56718_, new_n56680_ );
xor  ( new_n57010_, new_n57009_, new_n56778_ );
and  ( new_n57011_, new_n57010_, new_n57008_ );
xnor ( new_n57012_, new_n57010_, new_n57008_ );
xor  ( new_n57013_, new_n46789_, new_n3892_ );
or   ( new_n57014_, new_n57013_, new_n4302_ );
or   ( new_n57015_, new_n56691_, new_n4304_ );
and  ( new_n57016_, new_n57015_, new_n57014_ );
xor  ( new_n57017_, new_n46958_, RIbb2e530_37 );
nand ( new_n57018_, new_n57017_, new_n3733_ );
or   ( new_n57019_, new_n56705_, new_n3898_ );
and  ( new_n57020_, new_n57019_, new_n57018_ );
or   ( new_n57021_, new_n57020_, new_n57016_ );
and  ( new_n57022_, new_n56811_, new_n4541_ );
xor  ( new_n57023_, new_n46427_, RIbb2e350_41 );
and  ( new_n57024_, new_n57023_, new_n4543_ );
or   ( new_n57025_, new_n57024_, new_n57022_ );
xor  ( new_n57026_, new_n57020_, new_n57016_ );
nand ( new_n57027_, new_n57026_, new_n57025_ );
and  ( new_n57028_, new_n57027_, new_n57021_ );
nor  ( new_n57029_, new_n56641_, new_n526_ );
xor  ( new_n57030_, new_n52908_, RIbb2f070_13 );
nor  ( new_n57031_, new_n57030_, new_n524_ );
or   ( new_n57032_, new_n57031_, new_n57029_ );
xor  ( new_n57033_, new_n56749_, new_n56740_ );
nand ( new_n57034_, new_n57033_, new_n57032_ );
xor  ( new_n57035_, new_n51758_, new_n745_ );
nor  ( new_n57036_, new_n57035_, new_n897_ );
and  ( new_n57037_, new_n56757_, new_n820_ );
or   ( new_n57038_, new_n57037_, new_n57036_ );
xor  ( new_n57039_, new_n57033_, new_n57032_ );
nand ( new_n57040_, new_n57039_, new_n57038_ );
and  ( new_n57041_, new_n57040_, new_n57034_ );
xor  ( new_n57042_, new_n47046_, new_n3113_ );
or   ( new_n57043_, new_n57042_, new_n3461_ );
or   ( new_n57044_, new_n56710_, new_n3463_ );
and  ( new_n57045_, new_n57044_, new_n57043_ );
or   ( new_n57046_, new_n57045_, new_n57041_ );
and  ( new_n57047_, new_n56763_, new_n9738_ );
xor  ( new_n57048_, new_n43914_, RIbb2d9f0_61 );
and  ( new_n57049_, new_n57048_, new_n9740_ );
or   ( new_n57050_, new_n57049_, new_n57047_ );
xor  ( new_n57051_, new_n57045_, new_n57041_ );
nand ( new_n57052_, new_n57051_, new_n57050_ );
and  ( new_n57053_, new_n57052_, new_n57046_ );
nor  ( new_n57054_, new_n57053_, new_n57028_ );
or   ( new_n57055_, new_n56725_, new_n6175_ );
xor  ( new_n57056_, new_n45584_, new_n5594_ );
or   ( new_n57057_, new_n57056_, new_n6173_ );
and  ( new_n57058_, new_n57057_, new_n57055_ );
xor  ( new_n57059_, new_n45204_, RIbb2df90_49 );
nand ( new_n57060_, new_n57059_, new_n6510_ );
or   ( new_n57061_, new_n56769_, new_n6647_ );
and  ( new_n57062_, new_n57061_, new_n57060_ );
nor  ( new_n57063_, new_n57062_, new_n57058_ );
and  ( new_n57064_, new_n56731_, new_n8649_ );
xor  ( new_n57065_, new_n44407_, RIbb2dbd0_57 );
and  ( new_n57066_, new_n57065_, new_n8651_ );
or   ( new_n57067_, new_n57066_, new_n57064_ );
xor  ( new_n57068_, new_n57062_, new_n57058_ );
and  ( new_n57069_, new_n57068_, new_n57067_ );
nor  ( new_n57070_, new_n57069_, new_n57063_ );
not  ( new_n57071_, new_n57070_ );
xor  ( new_n57072_, new_n57053_, new_n57028_ );
and  ( new_n57073_, new_n57072_, new_n57071_ );
or   ( new_n57074_, new_n57073_, new_n57054_ );
xnor ( new_n57075_, new_n56701_, new_n56685_ );
xor  ( new_n57076_, new_n57075_, new_n56716_ );
nand ( new_n57077_, new_n57076_, new_n57074_ );
nor  ( new_n57078_, new_n57076_, new_n57074_ );
xor  ( new_n57079_, new_n45597_, RIbb2e170_45 );
nand ( new_n57080_, new_n57079_, new_n5373_ );
or   ( new_n57081_, new_n56722_, new_n5606_ );
and  ( new_n57082_, new_n57081_, new_n57080_ );
nand ( new_n57083_, new_n56821_, new_n8040_ );
xor  ( new_n57084_, new_n44600_, new_n7722_ );
or   ( new_n57085_, new_n57084_, new_n8264_ );
and  ( new_n57086_, new_n57085_, new_n57083_ );
nor  ( new_n57087_, new_n57086_, new_n57082_ );
xor  ( new_n57088_, new_n46037_, new_n4705_ );
nor  ( new_n57089_, new_n57088_, new_n5207_ );
nor  ( new_n57090_, new_n56815_, new_n5209_ );
or   ( new_n57091_, new_n57090_, new_n57089_ );
xor  ( new_n57092_, new_n57086_, new_n57082_ );
and  ( new_n57093_, new_n57092_, new_n57091_ );
or   ( new_n57094_, new_n57093_, new_n57087_ );
xor  ( new_n57095_, new_n56714_, new_n56713_ );
and  ( new_n57096_, new_n57095_, new_n57094_ );
nor  ( new_n57097_, new_n57095_, new_n57094_ );
xor  ( new_n57098_, new_n43952_, RIbb2d900_63 );
and  ( new_n57099_, new_n57098_, RIbb2d888_64 );
and  ( new_n57100_, new_n21077_, RIbb2d900_63 );
and  ( new_n57101_, new_n57100_, new_n44139_ );
or   ( new_n57102_, new_n57101_, new_n57099_ );
xor  ( new_n57103_, new_n56760_, new_n56759_ );
and  ( new_n57104_, new_n57103_, new_n57102_ );
and  ( new_n57105_, new_n56595_, new_n7487_ );
xor  ( new_n57106_, new_n44785_, RIbb2ddb0_53 );
and  ( new_n57107_, new_n57106_, new_n7489_ );
or   ( new_n57108_, new_n57107_, new_n57105_ );
xor  ( new_n57109_, new_n57103_, new_n57102_ );
and  ( new_n57110_, new_n57109_, new_n57108_ );
nor  ( new_n57111_, new_n57110_, new_n57104_ );
nor  ( new_n57112_, new_n57111_, new_n57097_ );
nor  ( new_n57113_, new_n57112_, new_n57096_ );
or   ( new_n57114_, new_n57113_, new_n57078_ );
and  ( new_n57115_, new_n57114_, new_n57077_ );
nor  ( new_n57116_, new_n57115_, new_n57012_ );
nor  ( new_n57117_, new_n57116_, new_n57011_ );
nor  ( new_n57118_, new_n57117_, new_n57007_ );
nor  ( new_n57119_, new_n57118_, new_n57006_ );
nor  ( new_n57120_, new_n57119_, new_n56956_ );
nor  ( new_n57121_, new_n57120_, new_n56955_ );
or   ( new_n57122_, new_n57121_, new_n56886_ );
and  ( new_n57123_, new_n57122_, new_n56885_ );
nor  ( new_n57124_, new_n57123_, new_n56881_ );
and  ( new_n57125_, new_n57123_, new_n56881_ );
xor  ( new_n57126_, new_n56884_, new_n56882_ );
xnor ( new_n57127_, new_n57126_, new_n57121_ );
not  ( new_n57128_, new_n57127_ );
xor  ( new_n57129_, new_n57002_, new_n57001_ );
not  ( new_n57130_, new_n57129_ );
xor  ( new_n57131_, new_n56776_, new_n56775_ );
xor  ( new_n57132_, new_n56611_, new_n56606_ );
xor  ( new_n57133_, new_n57132_, new_n56614_ );
nand ( new_n57134_, new_n57133_, new_n57131_ );
nor  ( new_n57135_, new_n57133_, new_n57131_ );
nor  ( new_n57136_, new_n57042_, new_n3463_ );
xor  ( new_n57137_, new_n47296_, RIbb2e620_35 );
and  ( new_n57138_, new_n57137_, new_n3293_ );
or   ( new_n57139_, new_n57138_, new_n57136_ );
xor  ( new_n57140_, new_n57039_, new_n57038_ );
and  ( new_n57141_, new_n57140_, new_n57139_ );
xor  ( new_n57142_, new_n47303_, new_n3457_ );
nor  ( new_n57143_, new_n57142_, new_n3896_ );
and  ( new_n57144_, new_n57017_, new_n3731_ );
or   ( new_n57145_, new_n57144_, new_n57143_ );
xor  ( new_n57146_, new_n57140_, new_n57139_ );
and  ( new_n57147_, new_n57146_, new_n57145_ );
nor  ( new_n57148_, new_n57147_, new_n57141_ );
not  ( new_n57149_, new_n57148_ );
xor  ( new_n57150_, new_n56842_, new_n56841_ );
and  ( new_n57151_, new_n57150_, new_n57149_ );
xor  ( new_n57152_, new_n57150_, new_n57149_ );
xnor ( new_n57153_, new_n56965_, new_n56961_ );
xor  ( new_n57154_, new_n57153_, new_n56969_ );
and  ( new_n57155_, new_n57154_, new_n57152_ );
nor  ( new_n57156_, new_n57155_, new_n57151_ );
not  ( new_n57157_, new_n57156_ );
xor  ( new_n57158_, new_n56852_, new_n56847_ );
nand ( new_n57159_, new_n57158_, new_n57157_ );
xor  ( new_n57160_, new_n57158_, new_n57157_ );
xnor ( new_n57161_, new_n56817_, new_n56813_ );
xor  ( new_n57162_, new_n57161_, new_n56823_ );
nand ( new_n57163_, new_n57162_, new_n57160_ );
and  ( new_n57164_, new_n57163_, new_n57159_ );
or   ( new_n57165_, new_n57164_, new_n57135_ );
and  ( new_n57166_, new_n57165_, new_n57134_ );
nor  ( new_n57167_, new_n57166_, new_n57130_ );
xor  ( new_n57168_, new_n57166_, new_n57130_ );
xnor ( new_n57169_, new_n56992_, new_n56957_ );
xor  ( new_n57170_, new_n57169_, new_n56994_ );
xnor ( new_n57171_, new_n56854_, new_n56831_ );
xor  ( new_n57172_, new_n57171_, new_n56858_ );
or   ( new_n57173_, new_n57172_, new_n57170_ );
and  ( new_n57174_, new_n57172_, new_n57170_ );
xor  ( new_n57175_, new_n56972_, new_n56958_ );
xor  ( new_n57176_, new_n57175_, new_n56990_ );
or   ( new_n57177_, new_n56752_, new_n757_ );
xor  ( new_n57178_, new_n52293_, RIbb2ef80_15 );
or   ( new_n57179_, new_n57178_, new_n755_ );
and  ( new_n57180_, new_n57179_, new_n57177_ );
nor  ( new_n57181_, new_n57030_, new_n526_ );
xor  ( new_n57182_, new_n53306_, RIbb2f070_13 );
nor  ( new_n57183_, new_n57182_, new_n524_ );
or   ( new_n57184_, new_n57183_, new_n57181_ );
and  ( new_n57185_, new_n53694_, new_n371_ );
nand ( new_n57186_, new_n57185_, new_n57184_ );
nor  ( new_n57187_, new_n57178_, new_n757_ );
xor  ( new_n57188_, new_n52902_, RIbb2ef80_15 );
nor  ( new_n57189_, new_n57188_, new_n755_ );
or   ( new_n57190_, new_n57189_, new_n57187_ );
xor  ( new_n57191_, new_n57185_, new_n57184_ );
nand ( new_n57192_, new_n57191_, new_n57190_ );
and  ( new_n57193_, new_n57192_, new_n57186_ );
or   ( new_n57194_, new_n57193_, new_n57180_ );
xor  ( new_n57195_, new_n50487_, new_n1355_ );
nor  ( new_n57196_, new_n57195_, new_n1593_ );
nor  ( new_n57197_, new_n56832_, new_n1595_ );
or   ( new_n57198_, new_n57197_, new_n57196_ );
xor  ( new_n57199_, new_n57193_, new_n57180_ );
nand ( new_n57200_, new_n57199_, new_n57198_ );
and  ( new_n57201_, new_n57200_, new_n57194_ );
xor  ( new_n57202_, new_n48518_, new_n2421_ );
or   ( new_n57203_, new_n57202_, new_n2807_ );
or   ( new_n57204_, new_n56962_, new_n2809_ );
and  ( new_n57205_, new_n57204_, new_n57203_ );
xor  ( new_n57206_, new_n48908_, new_n2118_ );
or   ( new_n57207_, new_n57206_, new_n2425_ );
or   ( new_n57208_, new_n56979_, new_n2427_ );
and  ( new_n57209_, new_n57208_, new_n57207_ );
or   ( new_n57210_, new_n57209_, new_n57205_ );
nor  ( new_n57211_, new_n56985_, new_n2124_ );
xor  ( new_n57212_, new_n49427_, RIbb2e9e0_27 );
and  ( new_n57213_, new_n57212_, new_n2002_ );
nor  ( new_n57214_, new_n57213_, new_n57211_ );
and  ( new_n57215_, new_n57209_, new_n57205_ );
or   ( new_n57216_, new_n57215_, new_n57214_ );
and  ( new_n57217_, new_n57216_, new_n57210_ );
or   ( new_n57218_, new_n57217_, new_n57201_ );
and  ( new_n57219_, new_n57217_, new_n57201_ );
or   ( new_n57220_, new_n56975_, new_n3119_ );
xor  ( new_n57221_, new_n48039_, RIbb2e710_33 );
nand ( new_n57222_, new_n57221_, new_n2930_ );
and  ( new_n57223_, new_n57222_, new_n57220_ );
xor  ( new_n57224_, new_n46962_, new_n3892_ );
or   ( new_n57225_, new_n57224_, new_n4302_ );
or   ( new_n57226_, new_n57013_, new_n4304_ );
and  ( new_n57227_, new_n57226_, new_n57225_ );
nor  ( new_n57228_, new_n57227_, new_n57223_ );
xor  ( new_n57229_, new_n46619_, new_n4292_ );
nor  ( new_n57230_, new_n57229_, new_n4709_ );
and  ( new_n57231_, new_n57023_, new_n4541_ );
nor  ( new_n57232_, new_n57231_, new_n57230_ );
and  ( new_n57233_, new_n57227_, new_n57223_ );
nor  ( new_n57234_, new_n57233_, new_n57232_ );
nor  ( new_n57235_, new_n57234_, new_n57228_ );
or   ( new_n57236_, new_n57235_, new_n57219_ );
and  ( new_n57237_, new_n57236_, new_n57218_ );
nor  ( new_n57238_, new_n57237_, new_n57176_ );
and  ( new_n57239_, new_n57237_, new_n57176_ );
and  ( new_n57240_, new_n53694_, new_n43969_ );
or   ( new_n57241_, new_n57240_, new_n403_ );
or   ( new_n57242_, new_n57182_, new_n526_ );
or   ( new_n57243_, new_n56743_, new_n524_ );
or   ( new_n57244_, new_n57243_, new_n56746_ );
and  ( new_n57245_, new_n57244_, new_n57242_ );
or   ( new_n57246_, new_n57245_, new_n57241_ );
xor  ( new_n57247_, new_n52280_, new_n745_ );
or   ( new_n57248_, new_n57247_, new_n897_ );
or   ( new_n57249_, new_n57035_, new_n899_ );
and  ( new_n57250_, new_n57249_, new_n57248_ );
or   ( new_n57251_, new_n57250_, new_n57246_ );
and  ( new_n57252_, new_n56924_, new_n1040_ );
xor  ( new_n57253_, new_n51477_, RIbb2eda0_19 );
and  ( new_n57254_, new_n57253_, new_n1042_ );
or   ( new_n57255_, new_n57254_, new_n57252_ );
xor  ( new_n57256_, new_n57250_, new_n57246_ );
nand ( new_n57257_, new_n57256_, new_n57255_ );
and  ( new_n57258_, new_n57257_, new_n57251_ );
xor  ( new_n57259_, new_n44183_, new_n9418_ );
or   ( new_n57260_, new_n57259_, new_n10059_ );
nand ( new_n57261_, new_n57048_, new_n9738_ );
and  ( new_n57262_, new_n57261_, new_n57260_ );
or   ( new_n57263_, new_n57262_, new_n57258_ );
xor  ( new_n57264_, new_n45403_, new_n6163_ );
nor  ( new_n57265_, new_n57264_, new_n6645_ );
and  ( new_n57266_, new_n57059_, new_n6508_ );
or   ( new_n57267_, new_n57266_, new_n57265_ );
xor  ( new_n57268_, new_n57262_, new_n57258_ );
nand ( new_n57269_, new_n57268_, new_n57267_ );
and  ( new_n57270_, new_n57269_, new_n57263_ );
nand ( new_n57271_, new_n57065_, new_n8649_ );
xor  ( new_n57272_, new_n44506_, new_n8254_ );
or   ( new_n57273_, new_n57272_, new_n8874_ );
and  ( new_n57274_, new_n57273_, new_n57271_ );
xor  ( new_n57275_, new_n45738_, RIbb2e080_47 );
nand ( new_n57276_, new_n57275_, new_n5917_ );
or   ( new_n57277_, new_n57056_, new_n6175_ );
and  ( new_n57278_, new_n57277_, new_n57276_ );
or   ( new_n57279_, new_n57278_, new_n57274_ );
xor  ( new_n57280_, new_n45928_, new_n5203_ );
nor  ( new_n57281_, new_n57280_, new_n5604_ );
and  ( new_n57282_, new_n57079_, new_n5371_ );
or   ( new_n57283_, new_n57282_, new_n57281_ );
xor  ( new_n57284_, new_n57278_, new_n57274_ );
nand ( new_n57285_, new_n57284_, new_n57283_ );
and  ( new_n57286_, new_n57285_, new_n57279_ );
nor  ( new_n57287_, new_n57286_, new_n57270_ );
and  ( new_n57288_, new_n57286_, new_n57270_ );
or   ( new_n57289_, new_n57088_, new_n5209_ );
xor  ( new_n57290_, new_n46137_, RIbb2e260_43 );
nand ( new_n57291_, new_n57290_, new_n4960_ );
and  ( new_n57292_, new_n57291_, new_n57289_ );
xor  ( new_n57293_, new_n44681_, new_n7722_ );
or   ( new_n57294_, new_n57293_, new_n8264_ );
or   ( new_n57295_, new_n57084_, new_n8266_ );
and  ( new_n57296_, new_n57295_, new_n57294_ );
nor  ( new_n57297_, new_n57296_, new_n57292_ );
xor  ( new_n57298_, new_n44877_, RIbb2ddb0_53 );
and  ( new_n57299_, new_n57298_, new_n7489_ );
and  ( new_n57300_, new_n57106_, new_n7487_ );
nor  ( new_n57301_, new_n57300_, new_n57299_ );
and  ( new_n57302_, new_n57296_, new_n57292_ );
nor  ( new_n57303_, new_n57302_, new_n57301_ );
nor  ( new_n57304_, new_n57303_, new_n57297_ );
nor  ( new_n57305_, new_n57304_, new_n57288_ );
nor  ( new_n57306_, new_n57305_, new_n57287_ );
nor  ( new_n57307_, new_n57306_, new_n57239_ );
nor  ( new_n57308_, new_n57307_, new_n57238_ );
or   ( new_n57309_, new_n57308_, new_n57174_ );
nand ( new_n57310_, new_n57309_, new_n57173_ );
and  ( new_n57311_, new_n57310_, new_n57168_ );
or   ( new_n57312_, new_n57311_, new_n57167_ );
xnor ( new_n57313_, new_n57005_, new_n57004_ );
xor  ( new_n57314_, new_n57313_, new_n57117_ );
or   ( new_n57315_, new_n57314_, new_n57312_ );
and  ( new_n57316_, new_n57314_, new_n57312_ );
xor  ( new_n57317_, new_n57115_, new_n57012_ );
xnor ( new_n57318_, new_n56895_, new_n56894_ );
xor  ( new_n57319_, new_n57318_, new_n56950_ );
nor  ( new_n57320_, new_n57319_, new_n57317_ );
and  ( new_n57321_, new_n57319_, new_n57317_ );
not  ( new_n57322_, new_n57321_ );
xor  ( new_n57323_, new_n44319_, RIbb2dae0_59 );
nand ( new_n57324_, new_n57323_, new_n9187_ );
or   ( new_n57325_, new_n56913_, new_n9424_ );
and  ( new_n57326_, new_n57325_, new_n57324_ );
and  ( new_n57327_, new_n43985_, RIbb2d888_64 );
and  ( new_n57328_, new_n43812_, new_n21077_ );
or   ( new_n57329_, new_n57328_, new_n10052_ );
or   ( new_n57330_, new_n57329_, new_n57327_ );
nand ( new_n57331_, new_n57327_, new_n10052_ );
and  ( new_n57332_, new_n57331_, new_n57330_ );
nor  ( new_n57333_, new_n57332_, new_n57326_ );
and  ( new_n57334_, new_n56917_, new_n6908_ );
xor  ( new_n57335_, new_n45119_, new_n6635_ );
nor  ( new_n57336_, new_n57335_, new_n7184_ );
nor  ( new_n57337_, new_n57336_, new_n57334_ );
xnor ( new_n57338_, new_n57332_, new_n57326_ );
nor  ( new_n57339_, new_n57338_, new_n57337_ );
or   ( new_n57340_, new_n57339_, new_n57333_ );
xor  ( new_n57341_, new_n57026_, new_n57025_ );
and  ( new_n57342_, new_n57341_, new_n57340_ );
or   ( new_n57343_, new_n57341_, new_n57340_ );
xor  ( new_n57344_, new_n57051_, new_n57050_ );
and  ( new_n57345_, new_n57344_, new_n57343_ );
or   ( new_n57346_, new_n57345_, new_n57342_ );
xor  ( new_n57347_, new_n56901_, new_n56899_ );
xor  ( new_n57348_, new_n57347_, new_n56904_ );
or   ( new_n57349_, new_n57348_, new_n57346_ );
and  ( new_n57350_, new_n57348_, new_n57346_ );
xor  ( new_n57351_, new_n57095_, new_n57094_ );
xnor ( new_n57352_, new_n57351_, new_n57111_ );
or   ( new_n57353_, new_n57352_, new_n57350_ );
and  ( new_n57354_, new_n57353_, new_n57349_ );
xnor ( new_n57355_, new_n57076_, new_n57074_ );
xor  ( new_n57356_, new_n57355_, new_n57113_ );
and  ( new_n57357_, new_n57356_, new_n57354_ );
xor  ( new_n57358_, new_n57356_, new_n57354_ );
xnor ( new_n57359_, new_n56908_, new_n56906_ );
xor  ( new_n57360_, new_n57359_, new_n56948_ );
and  ( new_n57361_, new_n57360_, new_n57358_ );
nor  ( new_n57362_, new_n57361_, new_n57357_ );
and  ( new_n57363_, new_n57362_, new_n57322_ );
nor  ( new_n57364_, new_n57363_, new_n57320_ );
or   ( new_n57365_, new_n57364_, new_n57316_ );
and  ( new_n57366_, new_n57365_, new_n57315_ );
xnor ( new_n57367_, new_n56954_, new_n56887_ );
xor  ( new_n57368_, new_n57367_, new_n57119_ );
nand ( new_n57369_, new_n57368_, new_n57366_ );
nor  ( new_n57370_, new_n57368_, new_n57366_ );
xor  ( new_n57371_, new_n56800_, new_n56798_ );
xor  ( new_n57372_, new_n57371_, new_n56868_ );
not  ( new_n57373_, new_n57372_ );
or   ( new_n57374_, new_n57373_, new_n57370_ );
and  ( new_n57375_, new_n57374_, new_n57369_ );
and  ( new_n57376_, new_n57375_, new_n57128_ );
nor  ( new_n57377_, new_n57375_, new_n57128_ );
xor  ( new_n57378_, new_n57368_, new_n57366_ );
xor  ( new_n57379_, new_n57378_, new_n57373_ );
xor  ( new_n57380_, new_n56891_, new_n56889_ );
xor  ( new_n57381_, new_n57380_, new_n56952_ );
xnor ( new_n57382_, new_n57310_, new_n57168_ );
xor  ( new_n57383_, new_n57072_, new_n57071_ );
not  ( new_n57384_, new_n57383_ );
xor  ( new_n57385_, new_n57092_, new_n57091_ );
xor  ( new_n57386_, new_n57109_, new_n57108_ );
nand ( new_n57387_, new_n57386_, new_n57385_ );
nor  ( new_n57388_, new_n57386_, new_n57385_ );
nor  ( new_n57389_, new_n56927_, new_n1846_ );
xor  ( new_n57390_, new_n50115_, new_n1583_ );
nor  ( new_n57391_, new_n57390_, new_n1844_ );
or   ( new_n57392_, new_n57391_, new_n57389_ );
xor  ( new_n57393_, new_n57191_, new_n57190_ );
and  ( new_n57394_, new_n57393_, new_n57392_ );
and  ( new_n57395_, new_n57212_, new_n2000_ );
xor  ( new_n57396_, new_n49488_, RIbb2e9e0_27 );
and  ( new_n57397_, new_n57396_, new_n2002_ );
nor  ( new_n57398_, new_n57397_, new_n57395_ );
not  ( new_n57399_, new_n57398_ );
xor  ( new_n57400_, new_n57393_, new_n57392_ );
and  ( new_n57401_, new_n57400_, new_n57399_ );
nor  ( new_n57402_, new_n57401_, new_n57394_ );
not  ( new_n57403_, new_n57402_ );
xor  ( new_n57404_, new_n57199_, new_n57198_ );
and  ( new_n57405_, new_n57404_, new_n57403_ );
xor  ( new_n57406_, new_n57404_, new_n57403_ );
not  ( new_n57407_, new_n57406_ );
xor  ( new_n57408_, new_n50788_, new_n1355_ );
or   ( new_n57409_, new_n57408_, new_n1593_ );
or   ( new_n57410_, new_n57195_, new_n1595_ );
and  ( new_n57411_, new_n57410_, new_n57409_ );
xor  ( new_n57412_, new_n51142_, new_n1126_ );
or   ( new_n57413_, new_n57412_, new_n1364_ );
or   ( new_n57414_, new_n56933_, new_n1366_ );
and  ( new_n57415_, new_n57414_, new_n57413_ );
or   ( new_n57416_, new_n57415_, new_n57411_ );
and  ( new_n57417_, new_n57415_, new_n57411_ );
xor  ( new_n57418_, new_n48291_, RIbb2e710_33 );
and  ( new_n57419_, new_n57418_, new_n2930_ );
and  ( new_n57420_, new_n57221_, new_n2928_ );
nor  ( new_n57421_, new_n57420_, new_n57419_ );
or   ( new_n57422_, new_n57421_, new_n57417_ );
and  ( new_n57423_, new_n57422_, new_n57416_ );
nor  ( new_n57424_, new_n57423_, new_n57407_ );
nor  ( new_n57425_, new_n57424_, new_n57405_ );
or   ( new_n57426_, new_n57425_, new_n57388_ );
and  ( new_n57427_, new_n57426_, new_n57387_ );
or   ( new_n57428_, new_n57427_, new_n57384_ );
xor  ( new_n57429_, new_n57427_, new_n57384_ );
not  ( new_n57430_, new_n57429_ );
xor  ( new_n57431_, new_n57068_, new_n57067_ );
xnor ( new_n57432_, new_n56982_, new_n56978_ );
xor  ( new_n57433_, new_n57432_, new_n56987_ );
nand ( new_n57434_, new_n57433_, new_n57431_ );
or   ( new_n57435_, new_n57433_, new_n57431_ );
xor  ( new_n57436_, new_n56920_, new_n56916_ );
xnor ( new_n57437_, new_n57436_, new_n56939_ );
nand ( new_n57438_, new_n57437_, new_n57435_ );
and  ( new_n57439_, new_n57438_, new_n57434_ );
or   ( new_n57440_, new_n57439_, new_n57430_ );
and  ( new_n57441_, new_n57440_, new_n57428_ );
xor  ( new_n57442_, new_n57133_, new_n57131_ );
xor  ( new_n57443_, new_n57442_, new_n57164_ );
or   ( new_n57444_, new_n57443_, new_n57441_ );
and  ( new_n57445_, new_n57443_, new_n57441_ );
xor  ( new_n57446_, new_n48756_, new_n2421_ );
or   ( new_n57447_, new_n57446_, new_n2807_ );
or   ( new_n57448_, new_n57202_, new_n2809_ );
and  ( new_n57449_, new_n57448_, new_n57447_ );
xor  ( new_n57450_, new_n49265_, new_n2118_ );
or   ( new_n57451_, new_n57450_, new_n2425_ );
or   ( new_n57452_, new_n57206_, new_n2427_ );
and  ( new_n57453_, new_n57452_, new_n57451_ );
nor  ( new_n57454_, new_n57453_, new_n57449_ );
and  ( new_n57455_, new_n57290_, new_n4958_ );
xor  ( new_n57456_, new_n46427_, RIbb2e260_43 );
and  ( new_n57457_, new_n57456_, new_n4960_ );
or   ( new_n57458_, new_n57457_, new_n57455_ );
xor  ( new_n57459_, new_n57453_, new_n57449_ );
and  ( new_n57460_, new_n57459_, new_n57458_ );
or   ( new_n57461_, new_n57460_, new_n57454_ );
xor  ( new_n57462_, new_n56937_, new_n56936_ );
and  ( new_n57463_, new_n57462_, new_n57461_ );
xor  ( new_n57464_, new_n46958_, RIbb2e440_39 );
nand ( new_n57465_, new_n57464_, new_n4034_ );
or   ( new_n57466_, new_n57224_, new_n4304_ );
and  ( new_n57467_, new_n57466_, new_n57465_ );
or   ( new_n57468_, new_n57229_, new_n4711_ );
xor  ( new_n57469_, new_n46789_, new_n4292_ );
or   ( new_n57470_, new_n57469_, new_n4709_ );
and  ( new_n57471_, new_n57470_, new_n57468_ );
nor  ( new_n57472_, new_n57471_, new_n57467_ );
xor  ( new_n57473_, new_n47046_, new_n3457_ );
nor  ( new_n57474_, new_n57473_, new_n3896_ );
nor  ( new_n57475_, new_n57142_, new_n3898_ );
nor  ( new_n57476_, new_n57475_, new_n57474_ );
not  ( new_n57477_, new_n57476_ );
xor  ( new_n57478_, new_n57471_, new_n57467_ );
and  ( new_n57479_, new_n57478_, new_n57477_ );
or   ( new_n57480_, new_n57479_, new_n57472_ );
xor  ( new_n57481_, new_n57462_, new_n57461_ );
and  ( new_n57482_, new_n57481_, new_n57480_ );
nor  ( new_n57483_, new_n57482_, new_n57463_ );
xnor ( new_n57484_, new_n57217_, new_n57201_ );
xnor ( new_n57485_, new_n57484_, new_n57235_ );
nor  ( new_n57486_, new_n57485_, new_n57483_ );
xnor ( new_n57487_, new_n57485_, new_n57483_ );
xor  ( new_n57488_, new_n57146_, new_n57145_ );
xnor ( new_n57489_, new_n57209_, new_n57205_ );
xor  ( new_n57490_, new_n57489_, new_n57214_ );
nand ( new_n57491_, new_n57490_, new_n57488_ );
or   ( new_n57492_, new_n57490_, new_n57488_ );
xor  ( new_n57493_, new_n57227_, new_n57223_ );
xnor ( new_n57494_, new_n57493_, new_n57232_ );
nand ( new_n57495_, new_n57494_, new_n57492_ );
and  ( new_n57496_, new_n57495_, new_n57491_ );
nor  ( new_n57497_, new_n57496_, new_n57487_ );
or   ( new_n57498_, new_n57497_, new_n57486_ );
xor  ( new_n57499_, new_n56942_, new_n56912_ );
xor  ( new_n57500_, new_n57499_, new_n56946_ );
nor  ( new_n57501_, new_n57500_, new_n57498_ );
nand ( new_n57502_, new_n57500_, new_n57498_ );
xnor ( new_n57503_, new_n57162_, new_n57160_ );
and  ( new_n57504_, new_n57503_, new_n57502_ );
or   ( new_n57505_, new_n57504_, new_n57501_ );
or   ( new_n57506_, new_n57505_, new_n57445_ );
and  ( new_n57507_, new_n57506_, new_n57444_ );
or   ( new_n57508_, new_n57507_, new_n57382_ );
and  ( new_n57509_, new_n57507_, new_n57382_ );
xor  ( new_n57510_, new_n57172_, new_n57170_ );
xnor ( new_n57511_, new_n57510_, new_n57308_ );
not  ( new_n57512_, new_n57511_ );
xnor ( new_n57513_, new_n57154_, new_n57152_ );
xor  ( new_n57514_, new_n44785_, RIbb2dcc0_55 );
nand ( new_n57515_, new_n57514_, new_n8042_ );
or   ( new_n57516_, new_n57293_, new_n8266_ );
and  ( new_n57517_, new_n57516_, new_n57515_ );
or   ( new_n57518_, new_n57259_, new_n10061_ );
xor  ( new_n57519_, new_n44218_, new_n9418_ );
or   ( new_n57520_, new_n57519_, new_n10059_ );
and  ( new_n57521_, new_n57520_, new_n57518_ );
or   ( new_n57522_, new_n57521_, new_n57517_ );
xor  ( new_n57523_, new_n46037_, new_n5203_ );
nor  ( new_n57524_, new_n57523_, new_n5604_ );
nor  ( new_n57525_, new_n57280_, new_n5606_ );
nor  ( new_n57526_, new_n57525_, new_n57524_ );
and  ( new_n57527_, new_n57521_, new_n57517_ );
or   ( new_n57528_, new_n57527_, new_n57526_ );
and  ( new_n57529_, new_n57528_, new_n57522_ );
xor  ( new_n57530_, new_n44600_, new_n8254_ );
or   ( new_n57531_, new_n57530_, new_n8874_ );
or   ( new_n57532_, new_n57272_, new_n8876_ );
and  ( new_n57533_, new_n57532_, new_n57531_ );
xor  ( new_n57534_, new_n45584_, RIbb2df90_49 );
nand ( new_n57535_, new_n57534_, new_n6510_ );
or   ( new_n57536_, new_n57264_, new_n6647_ );
and  ( new_n57537_, new_n57536_, new_n57535_ );
or   ( new_n57538_, new_n57537_, new_n57533_ );
xor  ( new_n57539_, new_n45597_, RIbb2e080_47 );
and  ( new_n57540_, new_n57539_, new_n5917_ );
and  ( new_n57541_, new_n57275_, new_n5915_ );
nor  ( new_n57542_, new_n57541_, new_n57540_ );
and  ( new_n57543_, new_n57537_, new_n57533_ );
or   ( new_n57544_, new_n57543_, new_n57542_ );
and  ( new_n57545_, new_n57544_, new_n57538_ );
or   ( new_n57546_, new_n57545_, new_n57529_ );
xor  ( new_n57547_, new_n44974_, RIbb2ddb0_53 );
and  ( new_n57548_, new_n57547_, new_n7489_ );
and  ( new_n57549_, new_n57298_, new_n7487_ );
or   ( new_n57550_, new_n57549_, new_n57548_ );
xor  ( new_n57551_, new_n57256_, new_n57255_ );
and  ( new_n57552_, new_n57551_, new_n57550_ );
xor  ( new_n57553_, new_n44407_, RIbb2dae0_59 );
and  ( new_n57554_, new_n57553_, new_n9187_ );
and  ( new_n57555_, new_n57323_, new_n9185_ );
nor  ( new_n57556_, new_n57555_, new_n57554_ );
not  ( new_n57557_, new_n57556_ );
xor  ( new_n57558_, new_n57551_, new_n57550_ );
and  ( new_n57559_, new_n57558_, new_n57557_ );
nor  ( new_n57560_, new_n57559_, new_n57552_ );
and  ( new_n57561_, new_n57545_, new_n57529_ );
or   ( new_n57562_, new_n57561_, new_n57560_ );
and  ( new_n57563_, new_n57562_, new_n57546_ );
nor  ( new_n57564_, new_n57563_, new_n57513_ );
xnor ( new_n57565_, new_n57338_, new_n57337_ );
or   ( new_n57566_, new_n57335_, new_n7186_ );
xor  ( new_n57567_, new_n45204_, new_n6635_ );
or   ( new_n57568_, new_n57567_, new_n7184_ );
and  ( new_n57569_, new_n57568_, new_n57566_ );
xor  ( new_n57570_, new_n50894_, new_n1355_ );
or   ( new_n57571_, new_n57570_, new_n1593_ );
or   ( new_n57572_, new_n57408_, new_n1595_ );
and  ( new_n57573_, new_n57572_, new_n57571_ );
or   ( new_n57574_, new_n57390_, new_n1846_ );
xor  ( new_n57575_, new_n50487_, new_n1583_ );
or   ( new_n57576_, new_n57575_, new_n1844_ );
and  ( new_n57577_, new_n57576_, new_n57574_ );
or   ( new_n57578_, new_n57577_, new_n57573_ );
or   ( new_n57579_, new_n57412_, new_n1366_ );
xor  ( new_n57580_, new_n51446_, new_n1126_ );
or   ( new_n57581_, new_n57580_, new_n1364_ );
and  ( new_n57582_, new_n57581_, new_n57579_ );
and  ( new_n57583_, new_n57577_, new_n57573_ );
or   ( new_n57584_, new_n57583_, new_n57582_ );
and  ( new_n57585_, new_n57584_, new_n57578_ );
or   ( new_n57586_, new_n57585_, new_n57569_ );
or   ( new_n57587_, new_n57247_, new_n899_ );
xor  ( new_n57588_, new_n52293_, RIbb2ee90_17 );
or   ( new_n57589_, new_n57588_, new_n897_ );
and  ( new_n57590_, new_n57589_, new_n57587_ );
xor  ( new_n57591_, new_n52908_, RIbb2ef80_15 );
nor  ( new_n57592_, new_n57591_, new_n757_ );
xor  ( new_n57593_, new_n53306_, RIbb2ef80_15 );
nor  ( new_n57594_, new_n57593_, new_n755_ );
or   ( new_n57595_, new_n57594_, new_n57592_ );
and  ( new_n57596_, new_n53694_, new_n454_ );
nand ( new_n57597_, new_n57596_, new_n57595_ );
xor  ( new_n57598_, new_n52902_, RIbb2ee90_17 );
nor  ( new_n57599_, new_n57598_, new_n897_ );
nor  ( new_n57600_, new_n57588_, new_n899_ );
or   ( new_n57601_, new_n57600_, new_n57599_ );
xor  ( new_n57602_, new_n57596_, new_n57595_ );
nand ( new_n57603_, new_n57602_, new_n57601_ );
and  ( new_n57604_, new_n57603_, new_n57597_ );
nor  ( new_n57605_, new_n57604_, new_n57590_ );
xor  ( new_n57606_, new_n49758_, new_n1840_ );
nor  ( new_n57607_, new_n57606_, new_n2122_ );
and  ( new_n57608_, new_n57396_, new_n2000_ );
or   ( new_n57609_, new_n57608_, new_n57607_ );
xor  ( new_n57610_, new_n57604_, new_n57590_ );
and  ( new_n57611_, new_n57610_, new_n57609_ );
nor  ( new_n57612_, new_n57611_, new_n57605_ );
and  ( new_n57613_, new_n57585_, new_n57569_ );
or   ( new_n57614_, new_n57613_, new_n57612_ );
and  ( new_n57615_, new_n57614_, new_n57586_ );
nor  ( new_n57616_, new_n57615_, new_n57565_ );
xor  ( new_n57617_, new_n57615_, new_n57565_ );
xnor ( new_n57618_, new_n57296_, new_n57292_ );
xor  ( new_n57619_, new_n57618_, new_n57301_ );
and  ( new_n57620_, new_n57619_, new_n57617_ );
or   ( new_n57621_, new_n57620_, new_n57616_ );
xor  ( new_n57622_, new_n57563_, new_n57513_ );
and  ( new_n57623_, new_n57622_, new_n57621_ );
or   ( new_n57624_, new_n57623_, new_n57564_ );
xnor ( new_n57625_, new_n57237_, new_n57176_ );
xor  ( new_n57626_, new_n57625_, new_n57306_ );
nand ( new_n57627_, new_n57626_, new_n57624_ );
nor  ( new_n57628_, new_n57626_, new_n57624_ );
nor  ( new_n57629_, new_n57188_, new_n757_ );
nor  ( new_n57630_, new_n57591_, new_n755_ );
or   ( new_n57631_, new_n57630_, new_n57629_ );
xor  ( new_n57632_, new_n57245_, new_n57241_ );
and  ( new_n57633_, new_n57632_, new_n57631_ );
and  ( new_n57634_, new_n57253_, new_n1040_ );
xor  ( new_n57635_, new_n51758_, new_n893_ );
nor  ( new_n57636_, new_n57635_, new_n1135_ );
or   ( new_n57637_, new_n57636_, new_n57634_ );
xor  ( new_n57638_, new_n57632_, new_n57631_ );
and  ( new_n57639_, new_n57638_, new_n57637_ );
nor  ( new_n57640_, new_n57639_, new_n57633_ );
xor  ( new_n57641_, new_n47640_, new_n3113_ );
or   ( new_n57642_, new_n57641_, new_n3461_ );
nand ( new_n57643_, new_n57137_, new_n3291_ );
and  ( new_n57644_, new_n57643_, new_n57642_ );
nor  ( new_n57645_, new_n57644_, new_n57640_ );
xor  ( new_n57646_, new_n57644_, new_n57640_ );
and  ( new_n57647_, new_n43812_, RIbb2d888_64 );
or   ( new_n57648_, new_n57647_, RIbb2d900_63 );
nand ( new_n57649_, new_n57647_, RIbb2d900_63 );
or   ( new_n57650_, new_n44191_, RIbb2d888_64 );
and  ( new_n57651_, new_n57650_, new_n57649_ );
and  ( new_n57652_, new_n57651_, new_n57648_ );
and  ( new_n57653_, new_n57652_, new_n57646_ );
or   ( new_n57654_, new_n57653_, new_n57645_ );
xor  ( new_n57655_, new_n57284_, new_n57283_ );
and  ( new_n57656_, new_n57655_, new_n57654_ );
xor  ( new_n57657_, new_n57655_, new_n57654_ );
xor  ( new_n57658_, new_n57268_, new_n57267_ );
and  ( new_n57659_, new_n57658_, new_n57657_ );
nor  ( new_n57660_, new_n57659_, new_n57656_ );
not  ( new_n57661_, new_n57660_ );
xnor ( new_n57662_, new_n57286_, new_n57270_ );
xor  ( new_n57663_, new_n57662_, new_n57304_ );
and  ( new_n57664_, new_n57663_, new_n57661_ );
xor  ( new_n57665_, new_n57663_, new_n57661_ );
xor  ( new_n57666_, new_n57341_, new_n57340_ );
xor  ( new_n57667_, new_n57666_, new_n57344_ );
and  ( new_n57668_, new_n57667_, new_n57665_ );
nor  ( new_n57669_, new_n57668_, new_n57664_ );
or   ( new_n57670_, new_n57669_, new_n57628_ );
and  ( new_n57671_, new_n57670_, new_n57627_ );
or   ( new_n57672_, new_n57671_, new_n57512_ );
xor  ( new_n57673_, new_n57671_, new_n57512_ );
xor  ( new_n57674_, new_n57360_, new_n57358_ );
nand ( new_n57675_, new_n57674_, new_n57673_ );
and  ( new_n57676_, new_n57675_, new_n57672_ );
or   ( new_n57677_, new_n57676_, new_n57509_ );
and  ( new_n57678_, new_n57677_, new_n57508_ );
or   ( new_n57679_, new_n57678_, new_n57381_ );
and  ( new_n57680_, new_n57678_, new_n57381_ );
xor  ( new_n57681_, new_n57314_, new_n57312_ );
xnor ( new_n57682_, new_n57681_, new_n57364_ );
or   ( new_n57683_, new_n57682_, new_n57680_ );
and  ( new_n57684_, new_n57683_, new_n57679_ );
nor  ( new_n57685_, new_n57684_, new_n57379_ );
and  ( new_n57686_, new_n57684_, new_n57379_ );
xor  ( new_n57687_, new_n57507_, new_n57382_ );
xor  ( new_n57688_, new_n57687_, new_n57676_ );
xor  ( new_n57689_, new_n57319_, new_n57317_ );
xor  ( new_n57690_, new_n57689_, new_n57362_ );
nor  ( new_n57691_, new_n57690_, new_n57688_ );
and  ( new_n57692_, new_n57690_, new_n57688_ );
xor  ( new_n57693_, new_n57439_, new_n57430_ );
xor  ( new_n57694_, new_n57423_, new_n57407_ );
not  ( new_n57695_, new_n57694_ );
or   ( new_n57696_, new_n57450_, new_n2427_ );
xor  ( new_n57697_, new_n49427_, RIbb2e8f0_29 );
nand ( new_n57698_, new_n57697_, new_n2244_ );
and  ( new_n57699_, new_n57698_, new_n57696_ );
xor  ( new_n57700_, new_n48908_, new_n2421_ );
or   ( new_n57701_, new_n57700_, new_n2807_ );
or   ( new_n57702_, new_n57446_, new_n2809_ );
and  ( new_n57703_, new_n57702_, new_n57701_ );
or   ( new_n57704_, new_n57703_, new_n57699_ );
and  ( new_n57705_, new_n57418_, new_n2928_ );
xor  ( new_n57706_, new_n48518_, RIbb2e710_33 );
and  ( new_n57707_, new_n57706_, new_n2930_ );
nor  ( new_n57708_, new_n57707_, new_n57705_ );
and  ( new_n57709_, new_n57703_, new_n57699_ );
or   ( new_n57710_, new_n57709_, new_n57708_ );
and  ( new_n57711_, new_n57710_, new_n57704_ );
xor  ( new_n57712_, new_n46619_, new_n4705_ );
or   ( new_n57713_, new_n57712_, new_n5207_ );
nand ( new_n57714_, new_n57456_, new_n4958_ );
and  ( new_n57715_, new_n57714_, new_n57713_ );
xor  ( new_n57716_, new_n46962_, new_n4292_ );
or   ( new_n57717_, new_n57716_, new_n4709_ );
or   ( new_n57718_, new_n57469_, new_n4711_ );
and  ( new_n57719_, new_n57718_, new_n57717_ );
or   ( new_n57720_, new_n57719_, new_n57715_ );
and  ( new_n57721_, new_n57464_, new_n4032_ );
xor  ( new_n57722_, new_n47303_, new_n3892_ );
nor  ( new_n57723_, new_n57722_, new_n4302_ );
nor  ( new_n57724_, new_n57723_, new_n57721_ );
and  ( new_n57725_, new_n57719_, new_n57715_ );
or   ( new_n57726_, new_n57725_, new_n57724_ );
and  ( new_n57727_, new_n57726_, new_n57720_ );
or   ( new_n57728_, new_n57727_, new_n57711_ );
nor  ( new_n57729_, new_n57473_, new_n3898_ );
xor  ( new_n57730_, new_n47296_, RIbb2e530_37 );
and  ( new_n57731_, new_n57730_, new_n3733_ );
or   ( new_n57732_, new_n57731_, new_n57729_ );
xor  ( new_n57733_, new_n57638_, new_n57637_ );
nor  ( new_n57734_, new_n57733_, new_n57732_ );
nand ( new_n57735_, new_n57733_, new_n57732_ );
nor  ( new_n57736_, new_n57593_, new_n757_ );
and  ( new_n57737_, new_n44211_, RIbb2ef80_15 );
and  ( new_n57738_, new_n53694_, RIbb2ee90_17 );
or   ( new_n57739_, new_n57738_, new_n57737_ );
and  ( new_n57740_, RIbb2ef08_16, new_n520_ );
nor  ( new_n57741_, new_n53694_, RIbb2ee90_17 );
or   ( new_n57742_, new_n57741_, new_n57740_ );
and  ( new_n57743_, new_n57742_, new_n57739_ );
or   ( new_n57744_, new_n57743_, new_n57736_ );
or   ( new_n57745_, new_n53695_, new_n44212_ );
and  ( new_n57746_, new_n57745_, new_n522_ );
nand ( new_n57747_, new_n57746_, new_n57744_ );
or   ( new_n57748_, new_n57635_, new_n1137_ );
xor  ( new_n57749_, new_n52280_, new_n893_ );
or   ( new_n57750_, new_n57749_, new_n1135_ );
and  ( new_n57751_, new_n57750_, new_n57748_ );
and  ( new_n57752_, new_n57751_, new_n57747_ );
or   ( new_n57753_, new_n57751_, new_n57747_ );
xor  ( new_n57754_, new_n51477_, RIbb2ecb0_21 );
nand ( new_n57755_, new_n57754_, new_n1253_ );
or   ( new_n57756_, new_n57580_, new_n1366_ );
and  ( new_n57757_, new_n57756_, new_n57755_ );
and  ( new_n57758_, new_n57757_, new_n57753_ );
or   ( new_n57759_, new_n57758_, new_n57752_ );
and  ( new_n57760_, new_n57759_, new_n57735_ );
or   ( new_n57761_, new_n57760_, new_n57734_ );
and  ( new_n57762_, new_n57727_, new_n57711_ );
or   ( new_n57763_, new_n57762_, new_n57761_ );
and  ( new_n57764_, new_n57763_, new_n57728_ );
nor  ( new_n57765_, new_n57764_, new_n57695_ );
xor  ( new_n57766_, new_n57764_, new_n57695_ );
xor  ( new_n57767_, new_n57481_, new_n57480_ );
and  ( new_n57768_, new_n57767_, new_n57766_ );
or   ( new_n57769_, new_n57768_, new_n57765_ );
xor  ( new_n57770_, new_n57433_, new_n57431_ );
xor  ( new_n57771_, new_n57770_, new_n57437_ );
nand ( new_n57772_, new_n57771_, new_n57769_ );
nor  ( new_n57773_, new_n57771_, new_n57769_ );
xor  ( new_n57774_, new_n57386_, new_n57385_ );
xor  ( new_n57775_, new_n57774_, new_n57425_ );
or   ( new_n57776_, new_n57775_, new_n57773_ );
nand ( new_n57777_, new_n57776_, new_n57772_ );
nand ( new_n57778_, new_n57777_, new_n57693_ );
xnor ( new_n57779_, new_n57777_, new_n57693_ );
xnor ( new_n57780_, new_n57348_, new_n57346_ );
xor  ( new_n57781_, new_n57780_, new_n57352_ );
or   ( new_n57782_, new_n57781_, new_n57779_ );
and  ( new_n57783_, new_n57782_, new_n57778_ );
xor  ( new_n57784_, new_n57443_, new_n57441_ );
xor  ( new_n57785_, new_n57784_, new_n57505_ );
nor  ( new_n57786_, new_n57785_, new_n57783_ );
xor  ( new_n57787_, new_n57674_, new_n57673_ );
not  ( new_n57788_, new_n57787_ );
and  ( new_n57789_, new_n57785_, new_n57783_ );
nor  ( new_n57790_, new_n57789_, new_n57788_ );
nor  ( new_n57791_, new_n57790_, new_n57786_ );
nor  ( new_n57792_, new_n57791_, new_n57692_ );
nor  ( new_n57793_, new_n57792_, new_n57691_ );
not  ( new_n57794_, new_n57793_ );
xnor ( new_n57795_, new_n57678_, new_n57381_ );
xor  ( new_n57796_, new_n57795_, new_n57682_ );
nor  ( new_n57797_, new_n57796_, new_n57794_ );
and  ( new_n57798_, new_n57796_, new_n57794_ );
xor  ( new_n57799_, new_n57667_, new_n57665_ );
xor  ( new_n57800_, new_n57622_, new_n57621_ );
and  ( new_n57801_, new_n57800_, new_n57799_ );
xnor ( new_n57802_, new_n57800_, new_n57799_ );
xor  ( new_n57803_, new_n57658_, new_n57657_ );
xor  ( new_n57804_, new_n57619_, new_n57617_ );
nand ( new_n57805_, new_n57804_, new_n57803_ );
nor  ( new_n57806_, new_n57804_, new_n57803_ );
xor  ( new_n57807_, new_n57577_, new_n57573_ );
xor  ( new_n57808_, new_n57807_, new_n57582_ );
xor  ( new_n57809_, new_n50115_, new_n1840_ );
or   ( new_n57810_, new_n57809_, new_n2122_ );
or   ( new_n57811_, new_n57606_, new_n2124_ );
and  ( new_n57812_, new_n57811_, new_n57810_ );
xor  ( new_n57813_, new_n50788_, new_n1583_ );
or   ( new_n57814_, new_n57813_, new_n1844_ );
or   ( new_n57815_, new_n57575_, new_n1846_ );
and  ( new_n57816_, new_n57815_, new_n57814_ );
nor  ( new_n57817_, new_n57816_, new_n57812_ );
xor  ( new_n57818_, new_n46137_, RIbb2e170_45 );
and  ( new_n57819_, new_n57818_, new_n5371_ );
xor  ( new_n57820_, new_n46427_, RIbb2e170_45 );
and  ( new_n57821_, new_n57820_, new_n5373_ );
nor  ( new_n57822_, new_n57821_, new_n57819_ );
and  ( new_n57823_, new_n57816_, new_n57812_ );
nor  ( new_n57824_, new_n57823_, new_n57822_ );
nor  ( new_n57825_, new_n57824_, new_n57817_ );
or   ( new_n57826_, new_n57825_, new_n57808_ );
nor  ( new_n57827_, new_n57598_, new_n899_ );
xor  ( new_n57828_, new_n52908_, RIbb2ee90_17 );
nor  ( new_n57829_, new_n57828_, new_n897_ );
or   ( new_n57830_, new_n57829_, new_n57827_ );
xor  ( new_n57831_, new_n57746_, new_n57744_ );
nand ( new_n57832_, new_n57831_, new_n57830_ );
nor  ( new_n57833_, new_n57749_, new_n1137_ );
xor  ( new_n57834_, new_n52293_, RIbb2eda0_19 );
nor  ( new_n57835_, new_n57834_, new_n1135_ );
or   ( new_n57836_, new_n57835_, new_n57833_ );
xor  ( new_n57837_, new_n57831_, new_n57830_ );
nand ( new_n57838_, new_n57837_, new_n57836_ );
and  ( new_n57839_, new_n57838_, new_n57832_ );
xor  ( new_n57840_, new_n48291_, new_n3113_ );
or   ( new_n57841_, new_n57840_, new_n3461_ );
xor  ( new_n57842_, new_n48039_, new_n3113_ );
or   ( new_n57843_, new_n57842_, new_n3463_ );
and  ( new_n57844_, new_n57843_, new_n57841_ );
nor  ( new_n57845_, new_n57844_, new_n57839_ );
xor  ( new_n57846_, new_n45738_, RIbb2df90_49 );
and  ( new_n57847_, new_n57846_, new_n6508_ );
xor  ( new_n57848_, new_n45597_, RIbb2df90_49 );
and  ( new_n57849_, new_n57848_, new_n6510_ );
or   ( new_n57850_, new_n57849_, new_n57847_ );
xor  ( new_n57851_, new_n57844_, new_n57839_ );
and  ( new_n57852_, new_n57851_, new_n57850_ );
nor  ( new_n57853_, new_n57852_, new_n57845_ );
xnor ( new_n57854_, new_n57825_, new_n57808_ );
or   ( new_n57855_, new_n57854_, new_n57853_ );
and  ( new_n57856_, new_n57855_, new_n57826_ );
xor  ( new_n57857_, new_n57727_, new_n57711_ );
xor  ( new_n57858_, new_n57857_, new_n57761_ );
nor  ( new_n57859_, new_n57858_, new_n57856_ );
and  ( new_n57860_, new_n57858_, new_n57856_ );
xor  ( new_n57861_, new_n57400_, new_n57399_ );
or   ( new_n57862_, new_n57641_, new_n3463_ );
or   ( new_n57863_, new_n57842_, new_n3461_ );
and  ( new_n57864_, new_n57863_, new_n57862_ );
and  ( new_n57865_, new_n43914_, RIbb2d888_64 );
and  ( new_n57866_, new_n44183_, new_n21077_ );
or   ( new_n57867_, new_n57866_, new_n10052_ );
or   ( new_n57868_, new_n57867_, new_n57865_ );
nand ( new_n57869_, new_n57865_, new_n10052_ );
and  ( new_n57870_, new_n57869_, new_n57868_ );
nor  ( new_n57871_, new_n57870_, new_n57864_ );
and  ( new_n57872_, new_n57846_, new_n6510_ );
and  ( new_n57873_, new_n57534_, new_n6508_ );
or   ( new_n57874_, new_n57873_, new_n57872_ );
xor  ( new_n57875_, new_n57870_, new_n57864_ );
and  ( new_n57876_, new_n57875_, new_n57874_ );
or   ( new_n57877_, new_n57876_, new_n57871_ );
xnor ( new_n57878_, new_n57415_, new_n57411_ );
xor  ( new_n57879_, new_n57878_, new_n57421_ );
xor  ( new_n57880_, new_n57879_, new_n57877_ );
xor  ( new_n57881_, new_n57880_, new_n57861_ );
not  ( new_n57882_, new_n57881_ );
nor  ( new_n57883_, new_n57882_, new_n57860_ );
nor  ( new_n57884_, new_n57883_, new_n57859_ );
or   ( new_n57885_, new_n57884_, new_n57806_ );
and  ( new_n57886_, new_n57885_, new_n57805_ );
nor  ( new_n57887_, new_n57886_, new_n57802_ );
or   ( new_n57888_, new_n57887_, new_n57801_ );
xor  ( new_n57889_, new_n57781_, new_n57779_ );
nor  ( new_n57890_, new_n57889_, new_n57888_ );
and  ( new_n57891_, new_n57889_, new_n57888_ );
xor  ( new_n57892_, new_n57478_, new_n57477_ );
xor  ( new_n57893_, new_n57459_, new_n57458_ );
xnor ( new_n57894_, new_n57893_, new_n57892_ );
nand ( new_n57895_, new_n57553_, new_n9185_ );
xor  ( new_n57896_, new_n44506_, new_n8870_ );
or   ( new_n57897_, new_n57896_, new_n9422_ );
and  ( new_n57898_, new_n57897_, new_n57895_ );
or   ( new_n57899_, new_n57567_, new_n7186_ );
xor  ( new_n57900_, new_n45403_, new_n6635_ );
or   ( new_n57901_, new_n57900_, new_n7184_ );
and  ( new_n57902_, new_n57901_, new_n57899_ );
nand ( new_n57903_, new_n57902_, new_n57898_ );
nor  ( new_n57904_, new_n57902_, new_n57898_ );
xor  ( new_n57905_, new_n57610_, new_n57609_ );
or   ( new_n57906_, new_n57905_, new_n57904_ );
and  ( new_n57907_, new_n57906_, new_n57903_ );
xor  ( new_n57908_, new_n57907_, new_n57894_ );
xnor ( new_n57909_, new_n57719_, new_n57715_ );
xor  ( new_n57910_, new_n57909_, new_n57724_ );
xnor ( new_n57911_, new_n57703_, new_n57699_ );
xor  ( new_n57912_, new_n57911_, new_n57708_ );
nand ( new_n57913_, new_n57912_, new_n57910_ );
nor  ( new_n57914_, new_n57912_, new_n57910_ );
xor  ( new_n57915_, new_n45928_, new_n5594_ );
or   ( new_n57916_, new_n57915_, new_n6175_ );
xor  ( new_n57917_, new_n46037_, new_n5594_ );
or   ( new_n57918_, new_n57917_, new_n6173_ );
and  ( new_n57919_, new_n57918_, new_n57916_ );
xor  ( new_n57920_, new_n44785_, new_n8254_ );
or   ( new_n57921_, new_n57920_, new_n8874_ );
xor  ( new_n57922_, new_n44681_, new_n8254_ );
or   ( new_n57923_, new_n57922_, new_n8876_ );
and  ( new_n57924_, new_n57923_, new_n57921_ );
nor  ( new_n57925_, new_n57924_, new_n57919_ );
xor  ( new_n57926_, new_n45204_, RIbb2ddb0_53 );
and  ( new_n57927_, new_n57926_, new_n7489_ );
xor  ( new_n57928_, new_n45119_, new_n7174_ );
nor  ( new_n57929_, new_n57928_, new_n7734_ );
nor  ( new_n57930_, new_n57929_, new_n57927_ );
and  ( new_n57931_, new_n57924_, new_n57919_ );
nor  ( new_n57932_, new_n57931_, new_n57930_ );
nor  ( new_n57933_, new_n57932_, new_n57925_ );
or   ( new_n57934_, new_n57933_, new_n57914_ );
and  ( new_n57935_, new_n57934_, new_n57913_ );
or   ( new_n57936_, new_n57935_, new_n57908_ );
and  ( new_n57937_, new_n57935_, new_n57908_ );
xor  ( new_n57938_, new_n57875_, new_n57874_ );
and  ( new_n57939_, new_n57514_, new_n8040_ );
xor  ( new_n57940_, new_n44877_, RIbb2dcc0_55 );
and  ( new_n57941_, new_n57940_, new_n8042_ );
or   ( new_n57942_, new_n57941_, new_n57939_ );
xor  ( new_n57943_, new_n44319_, new_n9418_ );
or   ( new_n57944_, new_n57943_, new_n10059_ );
or   ( new_n57945_, new_n57519_, new_n10061_ );
and  ( new_n57946_, new_n57945_, new_n57944_ );
nand ( new_n57947_, new_n57547_, new_n7487_ );
or   ( new_n57948_, new_n57928_, new_n7732_ );
and  ( new_n57949_, new_n57948_, new_n57947_ );
xor  ( new_n57950_, new_n57949_, new_n57946_ );
xor  ( new_n57951_, new_n57950_, new_n57942_ );
and  ( new_n57952_, new_n57951_, new_n57938_ );
nor  ( new_n57953_, new_n57951_, new_n57938_ );
not  ( new_n57954_, new_n57953_ );
nor  ( new_n57955_, new_n57523_, new_n5606_ );
and  ( new_n57956_, new_n57818_, new_n5373_ );
nor  ( new_n57957_, new_n57956_, new_n57955_ );
or   ( new_n57958_, new_n57922_, new_n8874_ );
or   ( new_n57959_, new_n57530_, new_n8876_ );
and  ( new_n57960_, new_n57959_, new_n57958_ );
or   ( new_n57961_, new_n57915_, new_n6173_ );
nand ( new_n57962_, new_n57539_, new_n5915_ );
and  ( new_n57963_, new_n57962_, new_n57961_ );
xor  ( new_n57964_, new_n57963_, new_n57960_ );
xnor ( new_n57965_, new_n57964_, new_n57957_ );
and  ( new_n57966_, new_n57965_, new_n57954_ );
nor  ( new_n57967_, new_n57966_, new_n57952_ );
or   ( new_n57968_, new_n57967_, new_n57937_ );
and  ( new_n57969_, new_n57968_, new_n57936_ );
xnor ( new_n57970_, new_n57521_, new_n57517_ );
xor  ( new_n57971_, new_n57970_, new_n57526_ );
xnor ( new_n57972_, new_n57537_, new_n57533_ );
xor  ( new_n57973_, new_n57972_, new_n57542_ );
nor  ( new_n57974_, new_n57973_, new_n57971_ );
and  ( new_n57975_, new_n57973_, new_n57971_ );
xor  ( new_n57976_, new_n57558_, new_n57557_ );
nor  ( new_n57977_, new_n57976_, new_n57975_ );
nor  ( new_n57978_, new_n57977_, new_n57974_ );
or   ( new_n57979_, new_n57893_, new_n57892_ );
and  ( new_n57980_, new_n57893_, new_n57892_ );
or   ( new_n57981_, new_n57907_, new_n57980_ );
and  ( new_n57982_, new_n57981_, new_n57979_ );
xor  ( new_n57983_, new_n57490_, new_n57488_ );
xor  ( new_n57984_, new_n57983_, new_n57494_ );
xnor ( new_n57985_, new_n57984_, new_n57982_ );
xor  ( new_n57986_, new_n57985_, new_n57978_ );
nand ( new_n57987_, new_n57986_, new_n57969_ );
nor  ( new_n57988_, new_n57986_, new_n57969_ );
and  ( new_n57989_, new_n57697_, new_n2242_ );
xor  ( new_n57990_, new_n49488_, RIbb2e8f0_29 );
and  ( new_n57991_, new_n57990_, new_n2244_ );
or   ( new_n57992_, new_n57991_, new_n57989_ );
xor  ( new_n57993_, new_n51142_, new_n1355_ );
nor  ( new_n57994_, new_n57993_, new_n1593_ );
nor  ( new_n57995_, new_n57570_, new_n1595_ );
or   ( new_n57996_, new_n57995_, new_n57994_ );
xor  ( new_n57997_, new_n57602_, new_n57601_ );
xor  ( new_n57998_, new_n57997_, new_n57996_ );
xor  ( new_n57999_, new_n57998_, new_n57992_ );
xnor ( new_n58000_, new_n57816_, new_n57812_ );
nand ( new_n58001_, new_n58000_, new_n57822_ );
not  ( new_n58002_, new_n57824_ );
or   ( new_n58003_, new_n58002_, new_n57817_ );
and  ( new_n58004_, new_n58003_, new_n58001_ );
and  ( new_n58005_, new_n58004_, new_n57999_ );
and  ( new_n58006_, new_n53694_, new_n44376_ );
or   ( new_n58007_, new_n58006_, new_n748_ );
xor  ( new_n58008_, new_n53306_, RIbb2ee90_17 );
or   ( new_n58009_, new_n58008_, new_n899_ );
or   ( new_n58010_, new_n57738_, new_n897_ );
or   ( new_n58011_, new_n58010_, new_n57741_ );
and  ( new_n58012_, new_n58011_, new_n58009_ );
or   ( new_n58013_, new_n58012_, new_n58007_ );
xor  ( new_n58014_, new_n51758_, new_n1126_ );
or   ( new_n58015_, new_n58014_, new_n1366_ );
xor  ( new_n58016_, new_n52280_, new_n1126_ );
or   ( new_n58017_, new_n58016_, new_n1364_ );
and  ( new_n58018_, new_n58017_, new_n58015_ );
or   ( new_n58019_, new_n58018_, new_n58013_ );
xor  ( new_n58020_, new_n51446_, RIbb2ebc0_23 );
and  ( new_n58021_, new_n58020_, new_n1474_ );
xor  ( new_n58022_, new_n51477_, RIbb2ebc0_23 );
and  ( new_n58023_, new_n58022_, new_n1476_ );
or   ( new_n58024_, new_n58023_, new_n58021_ );
xor  ( new_n58025_, new_n58018_, new_n58013_ );
nand ( new_n58026_, new_n58025_, new_n58024_ );
and  ( new_n58027_, new_n58026_, new_n58019_ );
xor  ( new_n58028_, new_n47296_, RIbb2e440_39 );
nand ( new_n58029_, new_n58028_, new_n4034_ );
xor  ( new_n58030_, new_n47046_, new_n3892_ );
or   ( new_n58031_, new_n58030_, new_n4304_ );
and  ( new_n58032_, new_n58031_, new_n58029_ );
nor  ( new_n58033_, new_n58032_, new_n58027_ );
xor  ( new_n58034_, new_n48039_, RIbb2e530_37 );
and  ( new_n58035_, new_n58034_, new_n3733_ );
xor  ( new_n58036_, new_n47640_, new_n3457_ );
nor  ( new_n58037_, new_n58036_, new_n3898_ );
nor  ( new_n58038_, new_n58037_, new_n58035_ );
not  ( new_n58039_, new_n58038_ );
xor  ( new_n58040_, new_n58032_, new_n58027_ );
and  ( new_n58041_, new_n58040_, new_n58039_ );
or   ( new_n58042_, new_n58041_, new_n58033_ );
xor  ( new_n58043_, new_n58004_, new_n57999_ );
and  ( new_n58044_, new_n58043_, new_n58042_ );
or   ( new_n58045_, new_n58044_, new_n58005_ );
xor  ( new_n58046_, new_n57902_, new_n57898_ );
xor  ( new_n58047_, new_n58046_, new_n57905_ );
or   ( new_n58048_, new_n58047_, new_n58045_ );
nand ( new_n58049_, new_n58047_, new_n58045_ );
or   ( new_n58050_, new_n57993_, new_n1595_ );
nand ( new_n58051_, new_n58020_, new_n1476_ );
and  ( new_n58052_, new_n58051_, new_n58050_ );
or   ( new_n58053_, new_n57809_, new_n2124_ );
xor  ( new_n58054_, new_n50487_, new_n1840_ );
or   ( new_n58055_, new_n58054_, new_n2122_ );
and  ( new_n58056_, new_n58055_, new_n58053_ );
nor  ( new_n58057_, new_n58056_, new_n58052_ );
xor  ( new_n58058_, new_n50894_, new_n1583_ );
nor  ( new_n58059_, new_n58058_, new_n1844_ );
nor  ( new_n58060_, new_n57813_, new_n1846_ );
nor  ( new_n58061_, new_n58060_, new_n58059_ );
and  ( new_n58062_, new_n58056_, new_n58052_ );
nor  ( new_n58063_, new_n58062_, new_n58061_ );
nor  ( new_n58064_, new_n58063_, new_n58057_ );
nor  ( new_n58065_, new_n57828_, new_n899_ );
nor  ( new_n58066_, new_n58008_, new_n897_ );
or   ( new_n58067_, new_n58066_, new_n58065_ );
and  ( new_n58068_, new_n53694_, new_n660_ );
nand ( new_n58069_, new_n58068_, new_n58067_ );
xor  ( new_n58070_, new_n52902_, RIbb2eda0_19 );
nor  ( new_n58071_, new_n58070_, new_n1135_ );
nor  ( new_n58072_, new_n57834_, new_n1137_ );
or   ( new_n58073_, new_n58072_, new_n58071_ );
xor  ( new_n58074_, new_n58068_, new_n58067_ );
nand ( new_n58075_, new_n58074_, new_n58073_ );
and  ( new_n58076_, new_n58075_, new_n58069_ );
nand ( new_n58077_, new_n57990_, new_n2242_ );
xor  ( new_n58078_, new_n49758_, new_n2118_ );
or   ( new_n58079_, new_n58078_, new_n2425_ );
and  ( new_n58080_, new_n58079_, new_n58077_ );
or   ( new_n58081_, new_n58080_, new_n58076_ );
nor  ( new_n58082_, new_n58014_, new_n1364_ );
and  ( new_n58083_, new_n57754_, new_n1251_ );
nor  ( new_n58084_, new_n58083_, new_n58082_ );
and  ( new_n58085_, new_n58080_, new_n58076_ );
or   ( new_n58086_, new_n58085_, new_n58084_ );
and  ( new_n58087_, new_n58086_, new_n58081_ );
nor  ( new_n58088_, new_n58087_, new_n58064_ );
and  ( new_n58089_, new_n58087_, new_n58064_ );
xor  ( new_n58090_, new_n47303_, new_n4292_ );
nor  ( new_n58091_, new_n58090_, new_n4709_ );
xor  ( new_n58092_, new_n46958_, RIbb2e350_41 );
and  ( new_n58093_, new_n58092_, new_n4541_ );
or   ( new_n58094_, new_n58093_, new_n58091_ );
xor  ( new_n58095_, new_n57837_, new_n57836_ );
and  ( new_n58096_, new_n58095_, new_n58094_ );
xor  ( new_n58097_, new_n48908_, new_n2797_ );
nor  ( new_n58098_, new_n58097_, new_n3117_ );
xor  ( new_n58099_, new_n48756_, RIbb2e710_33 );
and  ( new_n58100_, new_n58099_, new_n2928_ );
or   ( new_n58101_, new_n58100_, new_n58098_ );
xor  ( new_n58102_, new_n58095_, new_n58094_ );
and  ( new_n58103_, new_n58102_, new_n58101_ );
nor  ( new_n58104_, new_n58103_, new_n58096_ );
nor  ( new_n58105_, new_n58104_, new_n58089_ );
nor  ( new_n58106_, new_n58105_, new_n58088_ );
nand ( new_n58107_, new_n58106_, new_n58049_ );
and  ( new_n58108_, new_n58107_, new_n58048_ );
xor  ( new_n58109_, new_n57973_, new_n57971_ );
xor  ( new_n58110_, new_n58109_, new_n57976_ );
nor  ( new_n58111_, new_n58110_, new_n58108_ );
nor  ( new_n58112_, new_n57949_, new_n57946_ );
and  ( new_n58113_, new_n57950_, new_n57942_ );
nor  ( new_n58114_, new_n58113_, new_n58112_ );
not  ( new_n58115_, new_n58114_ );
xnor ( new_n58116_, new_n57652_, new_n57646_ );
or   ( new_n58117_, new_n57963_, new_n57960_ );
and  ( new_n58118_, new_n57963_, new_n57960_ );
or   ( new_n58119_, new_n58118_, new_n57957_ );
and  ( new_n58120_, new_n58119_, new_n58117_ );
xor  ( new_n58121_, new_n58120_, new_n58116_ );
xor  ( new_n58122_, new_n58121_, new_n58115_ );
and  ( new_n58123_, new_n58110_, new_n58108_ );
nor  ( new_n58124_, new_n58123_, new_n58122_ );
nor  ( new_n58125_, new_n58124_, new_n58111_ );
or   ( new_n58126_, new_n58125_, new_n57988_ );
and  ( new_n58127_, new_n58126_, new_n57987_ );
xnor ( new_n58128_, new_n57771_, new_n57769_ );
xor  ( new_n58129_, new_n58128_, new_n57775_ );
nor  ( new_n58130_, new_n58129_, new_n58127_ );
and  ( new_n58131_, new_n58129_, new_n58127_ );
xnor ( new_n58132_, new_n57767_, new_n57766_ );
and  ( new_n58133_, new_n57997_, new_n57996_ );
and  ( new_n58134_, new_n57998_, new_n57992_ );
nor  ( new_n58135_, new_n58134_, new_n58133_ );
nand ( new_n58136_, new_n57730_, new_n3731_ );
or   ( new_n58137_, new_n58036_, new_n3896_ );
and  ( new_n58138_, new_n58137_, new_n58136_ );
nand ( new_n58139_, new_n58092_, new_n4543_ );
or   ( new_n58140_, new_n57716_, new_n4711_ );
and  ( new_n58141_, new_n58140_, new_n58139_ );
or   ( new_n58142_, new_n58141_, new_n58138_ );
nor  ( new_n58143_, new_n57722_, new_n4304_ );
nor  ( new_n58144_, new_n58030_, new_n4302_ );
nor  ( new_n58145_, new_n58144_, new_n58143_ );
and  ( new_n58146_, new_n58141_, new_n58138_ );
or   ( new_n58147_, new_n58146_, new_n58145_ );
and  ( new_n58148_, new_n58147_, new_n58142_ );
nor  ( new_n58149_, new_n58148_, new_n58135_ );
xnor ( new_n58150_, new_n58148_, new_n58135_ );
xor  ( new_n58151_, new_n46789_, new_n4705_ );
or   ( new_n58152_, new_n58151_, new_n5207_ );
or   ( new_n58153_, new_n57712_, new_n5209_ );
and  ( new_n58154_, new_n58153_, new_n58152_ );
xor  ( new_n58155_, new_n49265_, new_n2421_ );
or   ( new_n58156_, new_n58155_, new_n2807_ );
or   ( new_n58157_, new_n57700_, new_n2809_ );
and  ( new_n58158_, new_n58157_, new_n58156_ );
or   ( new_n58159_, new_n58158_, new_n58154_ );
and  ( new_n58160_, new_n57706_, new_n2928_ );
and  ( new_n58161_, new_n58099_, new_n2930_ );
nor  ( new_n58162_, new_n58161_, new_n58160_ );
and  ( new_n58163_, new_n58158_, new_n58154_ );
or   ( new_n58164_, new_n58163_, new_n58162_ );
and  ( new_n58165_, new_n58164_, new_n58159_ );
nor  ( new_n58166_, new_n58165_, new_n58150_ );
or   ( new_n58167_, new_n58166_, new_n58149_ );
xnor ( new_n58168_, new_n57585_, new_n57569_ );
xor  ( new_n58169_, new_n58168_, new_n57612_ );
nand ( new_n58170_, new_n58169_, new_n58167_ );
nor  ( new_n58171_, new_n58169_, new_n58167_ );
or   ( new_n58172_, new_n57943_, new_n10061_ );
xor  ( new_n58173_, new_n44407_, new_n9418_ );
or   ( new_n58174_, new_n58173_, new_n10059_ );
and  ( new_n58175_, new_n58174_, new_n58172_ );
and  ( new_n58176_, new_n44183_, RIbb2d888_64 );
and  ( new_n58177_, new_n44218_, new_n21077_ );
or   ( new_n58178_, new_n58177_, new_n10052_ );
or   ( new_n58179_, new_n58178_, new_n58176_ );
nand ( new_n58180_, new_n58176_, new_n10052_ );
and  ( new_n58181_, new_n58180_, new_n58179_ );
or   ( new_n58182_, new_n58181_, new_n58175_ );
xor  ( new_n58183_, new_n44974_, RIbb2dcc0_55 );
and  ( new_n58184_, new_n58183_, new_n8042_ );
and  ( new_n58185_, new_n57940_, new_n8040_ );
or   ( new_n58186_, new_n58185_, new_n58184_ );
xor  ( new_n58187_, new_n58181_, new_n58175_ );
nand ( new_n58188_, new_n58187_, new_n58186_ );
and  ( new_n58189_, new_n58188_, new_n58182_ );
xor  ( new_n58190_, new_n57733_, new_n57732_ );
xor  ( new_n58191_, new_n58190_, new_n57759_ );
nor  ( new_n58192_, new_n58191_, new_n58189_ );
or   ( new_n58193_, new_n57896_, new_n9424_ );
xor  ( new_n58194_, new_n44600_, new_n8870_ );
or   ( new_n58195_, new_n58194_, new_n9422_ );
and  ( new_n58196_, new_n58195_, new_n58193_ );
xor  ( new_n58197_, new_n57751_, new_n57747_ );
xor  ( new_n58198_, new_n58197_, new_n57757_ );
nor  ( new_n58199_, new_n58198_, new_n58196_ );
xor  ( new_n58200_, new_n45584_, RIbb2dea0_51 );
and  ( new_n58201_, new_n58200_, new_n6910_ );
nor  ( new_n58202_, new_n57900_, new_n7186_ );
or   ( new_n58203_, new_n58202_, new_n58201_ );
xor  ( new_n58204_, new_n58198_, new_n58196_ );
and  ( new_n58205_, new_n58204_, new_n58203_ );
nor  ( new_n58206_, new_n58205_, new_n58199_ );
not  ( new_n58207_, new_n58206_ );
xor  ( new_n58208_, new_n58191_, new_n58189_ );
and  ( new_n58209_, new_n58208_, new_n58207_ );
nor  ( new_n58210_, new_n58209_, new_n58192_ );
or   ( new_n58211_, new_n58210_, new_n58171_ );
and  ( new_n58212_, new_n58211_, new_n58170_ );
nor  ( new_n58213_, new_n58212_, new_n58132_ );
xor  ( new_n58214_, new_n58212_, new_n58132_ );
or   ( new_n58215_, new_n58120_, new_n58116_ );
nand ( new_n58216_, new_n58121_, new_n58115_ );
and  ( new_n58217_, new_n58216_, new_n58215_ );
nand ( new_n58218_, new_n57879_, new_n57877_ );
or   ( new_n58219_, new_n57879_, new_n57877_ );
nand ( new_n58220_, new_n58219_, new_n57861_ );
and  ( new_n58221_, new_n58220_, new_n58218_ );
xor  ( new_n58222_, new_n58221_, new_n58217_ );
xnor ( new_n58223_, new_n57545_, new_n57529_ );
xor  ( new_n58224_, new_n58223_, new_n57560_ );
xor  ( new_n58225_, new_n58224_, new_n58222_ );
and  ( new_n58226_, new_n58225_, new_n58214_ );
nor  ( new_n58227_, new_n58226_, new_n58213_ );
not  ( new_n58228_, new_n58227_ );
nor  ( new_n58229_, new_n58228_, new_n58131_ );
nor  ( new_n58230_, new_n58229_, new_n58130_ );
nor  ( new_n58231_, new_n58230_, new_n57891_ );
nor  ( new_n58232_, new_n58231_, new_n57890_ );
not  ( new_n58233_, new_n58232_ );
xor  ( new_n58234_, new_n57496_, new_n57487_ );
or   ( new_n58235_, new_n57984_, new_n57982_ );
and  ( new_n58236_, new_n57984_, new_n57982_ );
or   ( new_n58237_, new_n58236_, new_n57978_ );
and  ( new_n58238_, new_n58237_, new_n58235_ );
nand ( new_n58239_, new_n58238_, new_n58234_ );
nor  ( new_n58240_, new_n58221_, new_n58217_ );
and  ( new_n58241_, new_n58224_, new_n58222_ );
or   ( new_n58242_, new_n58241_, new_n58240_ );
xor  ( new_n58243_, new_n58238_, new_n58234_ );
nand ( new_n58244_, new_n58243_, new_n58242_ );
and  ( new_n58245_, new_n58244_, new_n58239_ );
xor  ( new_n58246_, new_n57500_, new_n57498_ );
xor  ( new_n58247_, new_n58246_, new_n57503_ );
or   ( new_n58248_, new_n58247_, new_n58245_ );
and  ( new_n58249_, new_n58247_, new_n58245_ );
xor  ( new_n58250_, new_n57626_, new_n57624_ );
xnor ( new_n58251_, new_n58250_, new_n57669_ );
not  ( new_n58252_, new_n58251_ );
or   ( new_n58253_, new_n58252_, new_n58249_ );
and  ( new_n58254_, new_n58253_, new_n58248_ );
and  ( new_n58255_, new_n58254_, new_n58233_ );
xor  ( new_n58256_, new_n58254_, new_n58233_ );
xor  ( new_n58257_, new_n57785_, new_n57783_ );
xor  ( new_n58258_, new_n58257_, new_n57788_ );
and  ( new_n58259_, new_n58258_, new_n58256_ );
nor  ( new_n58260_, new_n58259_, new_n58255_ );
xnor ( new_n58261_, new_n57690_, new_n57688_ );
xor  ( new_n58262_, new_n58261_, new_n57791_ );
nor  ( new_n58263_, new_n58262_, new_n58260_ );
and  ( new_n58264_, new_n58262_, new_n58260_ );
xor  ( new_n58265_, new_n58258_, new_n58256_ );
xor  ( new_n58266_, new_n58243_, new_n58242_ );
xor  ( new_n58267_, new_n57886_, new_n57802_ );
and  ( new_n58268_, new_n58267_, new_n58266_ );
xnor ( new_n58269_, new_n57804_, new_n57803_ );
xor  ( new_n58270_, new_n58269_, new_n57884_ );
xnor ( new_n58271_, new_n57854_, new_n57853_ );
xnor ( new_n58272_, new_n58141_, new_n58138_ );
xor  ( new_n58273_, new_n58272_, new_n58145_ );
xnor ( new_n58274_, new_n58158_, new_n58154_ );
xor  ( new_n58275_, new_n58274_, new_n58162_ );
nand ( new_n58276_, new_n58275_, new_n58273_ );
nor  ( new_n58277_, new_n58275_, new_n58273_ );
or   ( new_n58278_, new_n57917_, new_n6175_ );
xor  ( new_n58279_, new_n46137_, RIbb2e080_47 );
nand ( new_n58280_, new_n58279_, new_n5917_ );
and  ( new_n58281_, new_n58280_, new_n58278_ );
and  ( new_n58282_, new_n44218_, RIbb2d888_64 );
and  ( new_n58283_, new_n44319_, new_n21077_ );
or   ( new_n58284_, new_n58283_, new_n10052_ );
or   ( new_n58285_, new_n58284_, new_n58282_ );
nand ( new_n58286_, new_n58282_, new_n10052_ );
and  ( new_n58287_, new_n58286_, new_n58285_ );
nor  ( new_n58288_, new_n58287_, new_n58281_ );
and  ( new_n58289_, new_n58287_, new_n58281_ );
xor  ( new_n58290_, new_n45119_, new_n7722_ );
nor  ( new_n58291_, new_n58290_, new_n8264_ );
and  ( new_n58292_, new_n58183_, new_n8040_ );
nor  ( new_n58293_, new_n58292_, new_n58291_ );
nor  ( new_n58294_, new_n58293_, new_n58289_ );
nor  ( new_n58295_, new_n58294_, new_n58288_ );
or   ( new_n58296_, new_n58295_, new_n58277_ );
and  ( new_n58297_, new_n58296_, new_n58276_ );
nor  ( new_n58298_, new_n58297_, new_n58271_ );
or   ( new_n58299_, new_n58155_, new_n2809_ );
xor  ( new_n58300_, new_n49427_, new_n2421_ );
or   ( new_n58301_, new_n58300_, new_n2807_ );
and  ( new_n58302_, new_n58301_, new_n58299_ );
nand ( new_n58303_, new_n57820_, new_n5371_ );
xor  ( new_n58304_, new_n46619_, new_n5203_ );
or   ( new_n58305_, new_n58304_, new_n5604_ );
and  ( new_n58306_, new_n58305_, new_n58303_ );
nor  ( new_n58307_, new_n58306_, new_n58302_ );
nor  ( new_n58308_, new_n58151_, new_n5209_ );
xor  ( new_n58309_, new_n46962_, new_n4705_ );
nor  ( new_n58310_, new_n58309_, new_n5207_ );
or   ( new_n58311_, new_n58310_, new_n58308_ );
xor  ( new_n58312_, new_n58306_, new_n58302_ );
and  ( new_n58313_, new_n58312_, new_n58311_ );
or   ( new_n58314_, new_n58313_, new_n58307_ );
xor  ( new_n58315_, new_n57851_, new_n57850_ );
and  ( new_n58316_, new_n58315_, new_n58314_ );
xor  ( new_n58317_, new_n44681_, new_n8870_ );
or   ( new_n58318_, new_n58317_, new_n9422_ );
or   ( new_n58319_, new_n58194_, new_n9424_ );
and  ( new_n58320_, new_n58319_, new_n58318_ );
xor  ( new_n58321_, new_n44506_, new_n9418_ );
or   ( new_n58322_, new_n58321_, new_n10059_ );
or   ( new_n58323_, new_n58173_, new_n10061_ );
and  ( new_n58324_, new_n58323_, new_n58322_ );
nor  ( new_n58325_, new_n58324_, new_n58320_ );
xor  ( new_n58326_, new_n45403_, new_n7174_ );
nor  ( new_n58327_, new_n58326_, new_n7732_ );
and  ( new_n58328_, new_n57926_, new_n7487_ );
or   ( new_n58329_, new_n58328_, new_n58327_ );
xor  ( new_n58330_, new_n58324_, new_n58320_ );
and  ( new_n58331_, new_n58330_, new_n58329_ );
or   ( new_n58332_, new_n58331_, new_n58325_ );
xor  ( new_n58333_, new_n58315_, new_n58314_ );
and  ( new_n58334_, new_n58333_, new_n58332_ );
nor  ( new_n58335_, new_n58334_, new_n58316_ );
xnor ( new_n58336_, new_n58297_, new_n58271_ );
nor  ( new_n58337_, new_n58336_, new_n58335_ );
or   ( new_n58338_, new_n58337_, new_n58298_ );
xnor ( new_n58339_, new_n58169_, new_n58167_ );
xor  ( new_n58340_, new_n58339_, new_n58210_ );
or   ( new_n58341_, new_n58340_, new_n58338_ );
nand ( new_n58342_, new_n58340_, new_n58338_ );
xor  ( new_n58343_, new_n57858_, new_n57856_ );
xor  ( new_n58344_, new_n58343_, new_n57882_ );
nand ( new_n58345_, new_n58344_, new_n58342_ );
and  ( new_n58346_, new_n58345_, new_n58341_ );
and  ( new_n58347_, new_n58346_, new_n58270_ );
xor  ( new_n58348_, new_n58225_, new_n58214_ );
xor  ( new_n58349_, new_n58346_, new_n58270_ );
and  ( new_n58350_, new_n58349_, new_n58348_ );
nor  ( new_n58351_, new_n58350_, new_n58347_ );
not  ( new_n58352_, new_n58351_ );
xor  ( new_n58353_, new_n58267_, new_n58266_ );
and  ( new_n58354_, new_n58353_, new_n58352_ );
or   ( new_n58355_, new_n58354_, new_n58268_ );
xor  ( new_n58356_, new_n57889_, new_n57888_ );
xor  ( new_n58357_, new_n58356_, new_n58230_ );
nand ( new_n58358_, new_n58357_, new_n58355_ );
nor  ( new_n58359_, new_n58357_, new_n58355_ );
xor  ( new_n58360_, new_n58247_, new_n58245_ );
xor  ( new_n58361_, new_n58360_, new_n58252_ );
or   ( new_n58362_, new_n58361_, new_n58359_ );
and  ( new_n58363_, new_n58362_, new_n58358_ );
and  ( new_n58364_, new_n58363_, new_n58265_ );
xor  ( new_n58365_, new_n58353_, new_n58352_ );
xor  ( new_n58366_, new_n58129_, new_n58127_ );
xor  ( new_n58367_, new_n58366_, new_n58228_ );
and  ( new_n58368_, new_n58367_, new_n58365_ );
xor  ( new_n58369_, new_n58367_, new_n58365_ );
not  ( new_n58370_, new_n58369_ );
xor  ( new_n58371_, new_n58165_, new_n58150_ );
xnor ( new_n58372_, new_n57912_, new_n57910_ );
xor  ( new_n58373_, new_n58372_, new_n57933_ );
nor  ( new_n58374_, new_n58373_, new_n58371_ );
and  ( new_n58375_, new_n58373_, new_n58371_ );
xor  ( new_n58376_, new_n58208_, new_n58207_ );
nor  ( new_n58377_, new_n58376_, new_n58375_ );
nor  ( new_n58378_, new_n58377_, new_n58374_ );
xor  ( new_n58379_, new_n58204_, new_n58203_ );
xnor ( new_n58380_, new_n57924_, new_n57919_ );
xor  ( new_n58381_, new_n58380_, new_n57930_ );
and  ( new_n58382_, new_n58381_, new_n58379_ );
or   ( new_n58383_, new_n58304_, new_n5606_ );
xor  ( new_n58384_, new_n46789_, new_n5203_ );
or   ( new_n58385_, new_n58384_, new_n5604_ );
and  ( new_n58386_, new_n58385_, new_n58383_ );
xor  ( new_n58387_, new_n46958_, RIbb2e260_43 );
nand ( new_n58388_, new_n58387_, new_n4960_ );
or   ( new_n58389_, new_n58309_, new_n5209_ );
and  ( new_n58390_, new_n58389_, new_n58388_ );
nor  ( new_n58391_, new_n58390_, new_n58386_ );
and  ( new_n58392_, new_n58279_, new_n5915_ );
xor  ( new_n58393_, new_n46427_, RIbb2e080_47 );
and  ( new_n58394_, new_n58393_, new_n5917_ );
or   ( new_n58395_, new_n58394_, new_n58392_ );
xor  ( new_n58396_, new_n58390_, new_n58386_ );
and  ( new_n58397_, new_n58396_, new_n58395_ );
nor  ( new_n58398_, new_n58397_, new_n58391_ );
not  ( new_n58399_, new_n58398_ );
xnor ( new_n58400_, new_n58056_, new_n58052_ );
nand ( new_n58401_, new_n58400_, new_n58061_ );
not  ( new_n58402_, new_n58063_ );
or   ( new_n58403_, new_n58402_, new_n58057_ );
and  ( new_n58404_, new_n58403_, new_n58401_ );
and  ( new_n58405_, new_n58404_, new_n58399_ );
xor  ( new_n58406_, new_n58404_, new_n58399_ );
nor  ( new_n58407_, new_n58070_, new_n1137_ );
xor  ( new_n58408_, new_n52908_, RIbb2eda0_19 );
nor  ( new_n58409_, new_n58408_, new_n1135_ );
or   ( new_n58410_, new_n58409_, new_n58407_ );
xor  ( new_n58411_, new_n58012_, new_n58007_ );
nand ( new_n58412_, new_n58411_, new_n58410_ );
and  ( new_n58413_, new_n58022_, new_n1474_ );
xor  ( new_n58414_, new_n51758_, new_n1355_ );
nor  ( new_n58415_, new_n58414_, new_n1593_ );
or   ( new_n58416_, new_n58415_, new_n58413_ );
xor  ( new_n58417_, new_n58411_, new_n58410_ );
nand ( new_n58418_, new_n58417_, new_n58416_ );
and  ( new_n58419_, new_n58418_, new_n58412_ );
or   ( new_n58420_, new_n58090_, new_n4711_ );
xor  ( new_n58421_, new_n47046_, new_n4292_ );
or   ( new_n58422_, new_n58421_, new_n4709_ );
and  ( new_n58423_, new_n58422_, new_n58420_ );
or   ( new_n58424_, new_n58423_, new_n58419_ );
xor  ( new_n58425_, new_n47640_, new_n3892_ );
nor  ( new_n58426_, new_n58425_, new_n4302_ );
and  ( new_n58427_, new_n58028_, new_n4032_ );
nor  ( new_n58428_, new_n58427_, new_n58426_ );
and  ( new_n58429_, new_n58423_, new_n58419_ );
or   ( new_n58430_, new_n58429_, new_n58428_ );
nand ( new_n58431_, new_n58430_, new_n58424_ );
and  ( new_n58432_, new_n58431_, new_n58406_ );
nor  ( new_n58433_, new_n58432_, new_n58405_ );
not  ( new_n58434_, new_n58433_ );
xor  ( new_n58435_, new_n58381_, new_n58379_ );
and  ( new_n58436_, new_n58435_, new_n58434_ );
or   ( new_n58437_, new_n58436_, new_n58382_ );
xor  ( new_n58438_, new_n57951_, new_n57938_ );
xor  ( new_n58439_, new_n58438_, new_n57965_ );
or   ( new_n58440_, new_n58439_, new_n58437_ );
nand ( new_n58441_, new_n58439_, new_n58437_ );
or   ( new_n58442_, new_n57840_, new_n3463_ );
xor  ( new_n58443_, new_n48518_, new_n3113_ );
or   ( new_n58444_, new_n58443_, new_n3461_ );
and  ( new_n58445_, new_n58444_, new_n58442_ );
xor  ( new_n58446_, new_n44877_, RIbb2dbd0_57 );
nand ( new_n58447_, new_n58446_, new_n8651_ );
or   ( new_n58448_, new_n57920_, new_n8876_ );
and  ( new_n58449_, new_n58448_, new_n58447_ );
nor  ( new_n58450_, new_n58449_, new_n58445_ );
xor  ( new_n58451_, new_n45928_, new_n6163_ );
nor  ( new_n58452_, new_n58451_, new_n6645_ );
and  ( new_n58453_, new_n57848_, new_n6508_ );
or   ( new_n58454_, new_n58453_, new_n58452_ );
xor  ( new_n58455_, new_n58449_, new_n58445_ );
and  ( new_n58456_, new_n58455_, new_n58454_ );
or   ( new_n58457_, new_n58456_, new_n58450_ );
xor  ( new_n58458_, new_n58187_, new_n58186_ );
and  ( new_n58459_, new_n58458_, new_n58457_ );
nor  ( new_n58460_, new_n58458_, new_n58457_ );
xor  ( new_n58461_, new_n50788_, new_n1840_ );
nor  ( new_n58462_, new_n58461_, new_n2122_ );
nor  ( new_n58463_, new_n58054_, new_n2124_ );
or   ( new_n58464_, new_n58463_, new_n58462_ );
xor  ( new_n58465_, new_n58074_, new_n58073_ );
and  ( new_n58466_, new_n58465_, new_n58464_ );
nor  ( new_n58467_, new_n58058_, new_n1846_ );
xor  ( new_n58468_, new_n51142_, new_n1583_ );
nor  ( new_n58469_, new_n58468_, new_n1844_ );
or   ( new_n58470_, new_n58469_, new_n58467_ );
xor  ( new_n58471_, new_n58465_, new_n58464_ );
and  ( new_n58472_, new_n58471_, new_n58470_ );
or   ( new_n58473_, new_n58472_, new_n58466_ );
xnor ( new_n58474_, new_n58080_, new_n58076_ );
xor  ( new_n58475_, new_n58474_, new_n58084_ );
and  ( new_n58476_, new_n58475_, new_n58473_ );
xor  ( new_n58477_, new_n45738_, RIbb2dea0_51 );
and  ( new_n58478_, new_n58477_, new_n6910_ );
and  ( new_n58479_, new_n58200_, new_n6908_ );
nor  ( new_n58480_, new_n58479_, new_n58478_ );
not  ( new_n58481_, new_n58480_ );
xor  ( new_n58482_, new_n58475_, new_n58473_ );
and  ( new_n58483_, new_n58482_, new_n58481_ );
nor  ( new_n58484_, new_n58483_, new_n58476_ );
nor  ( new_n58485_, new_n58484_, new_n58460_ );
nor  ( new_n58486_, new_n58485_, new_n58459_ );
nand ( new_n58487_, new_n58486_, new_n58441_ );
and  ( new_n58488_, new_n58487_, new_n58440_ );
nand ( new_n58489_, new_n58488_, new_n58378_ );
xor  ( new_n58490_, new_n58488_, new_n58378_ );
xnor ( new_n58491_, new_n57935_, new_n57908_ );
xor  ( new_n58492_, new_n58491_, new_n57967_ );
nand ( new_n58493_, new_n58492_, new_n58490_ );
and  ( new_n58494_, new_n58493_, new_n58489_ );
xnor ( new_n58495_, new_n57986_, new_n57969_ );
xor  ( new_n58496_, new_n58495_, new_n58125_ );
or   ( new_n58497_, new_n58496_, new_n58494_ );
and  ( new_n58498_, new_n58496_, new_n58494_ );
xor  ( new_n58499_, new_n58043_, new_n58042_ );
xnor ( new_n58500_, new_n58087_, new_n58064_ );
xor  ( new_n58501_, new_n58500_, new_n58104_ );
and  ( new_n58502_, new_n58501_, new_n58499_ );
xor  ( new_n58503_, new_n58040_, new_n58039_ );
xor  ( new_n58504_, new_n58102_, new_n58101_ );
and  ( new_n58505_, new_n58504_, new_n58503_ );
xor  ( new_n58506_, new_n58504_, new_n58503_ );
xor  ( new_n58507_, new_n44600_, RIbb2d9f0_61 );
nand ( new_n58508_, new_n58507_, new_n9740_ );
or   ( new_n58509_, new_n58321_, new_n10061_ );
and  ( new_n58510_, new_n58509_, new_n58508_ );
or   ( new_n58511_, new_n58290_, new_n8266_ );
xor  ( new_n58512_, new_n45204_, new_n7722_ );
or   ( new_n58513_, new_n58512_, new_n8264_ );
and  ( new_n58514_, new_n58513_, new_n58511_ );
or   ( new_n58515_, new_n58514_, new_n58510_ );
and  ( new_n58516_, new_n58446_, new_n8649_ );
xor  ( new_n58517_, new_n44974_, RIbb2dbd0_57 );
and  ( new_n58518_, new_n58517_, new_n8651_ );
nor  ( new_n58519_, new_n58518_, new_n58516_ );
and  ( new_n58520_, new_n58514_, new_n58510_ );
or   ( new_n58521_, new_n58520_, new_n58519_ );
nand ( new_n58522_, new_n58521_, new_n58515_ );
and  ( new_n58523_, new_n58522_, new_n58506_ );
or   ( new_n58524_, new_n58523_, new_n58505_ );
xor  ( new_n58525_, new_n58501_, new_n58499_ );
and  ( new_n58526_, new_n58525_, new_n58524_ );
nor  ( new_n58527_, new_n58526_, new_n58502_ );
xor  ( new_n58528_, new_n58047_, new_n58045_ );
xor  ( new_n58529_, new_n58528_, new_n58106_ );
and  ( new_n58530_, new_n58529_, new_n58527_ );
xor  ( new_n58531_, new_n58529_, new_n58527_ );
xor  ( new_n58532_, new_n50115_, new_n2118_ );
or   ( new_n58533_, new_n58532_, new_n2425_ );
or   ( new_n58534_, new_n58078_, new_n2427_ );
and  ( new_n58535_, new_n58534_, new_n58533_ );
or   ( new_n58536_, new_n58300_, new_n2809_ );
xor  ( new_n58537_, new_n49488_, RIbb2e800_31 );
nand ( new_n58538_, new_n58537_, new_n2615_ );
and  ( new_n58539_, new_n58538_, new_n58536_ );
nor  ( new_n58540_, new_n58539_, new_n58535_ );
nor  ( new_n58541_, new_n58097_, new_n3119_ );
xor  ( new_n58542_, new_n49265_, new_n2797_ );
nor  ( new_n58543_, new_n58542_, new_n3117_ );
or   ( new_n58544_, new_n58543_, new_n58541_ );
xor  ( new_n58545_, new_n58539_, new_n58535_ );
and  ( new_n58546_, new_n58545_, new_n58544_ );
nor  ( new_n58547_, new_n58546_, new_n58540_ );
xor  ( new_n58548_, new_n48756_, new_n3113_ );
or   ( new_n58549_, new_n58548_, new_n3461_ );
or   ( new_n58550_, new_n58443_, new_n3463_ );
and  ( new_n58551_, new_n58550_, new_n58549_ );
nand ( new_n58552_, new_n58034_, new_n3731_ );
xor  ( new_n58553_, new_n48291_, new_n3457_ );
or   ( new_n58554_, new_n58553_, new_n3896_ );
and  ( new_n58555_, new_n58554_, new_n58552_ );
nor  ( new_n58556_, new_n58555_, new_n58551_ );
and  ( new_n58557_, new_n58555_, new_n58551_ );
nor  ( new_n58558_, new_n58451_, new_n6647_ );
xor  ( new_n58559_, new_n46037_, new_n6163_ );
nor  ( new_n58560_, new_n58559_, new_n6645_ );
nor  ( new_n58561_, new_n58560_, new_n58558_ );
nor  ( new_n58562_, new_n58561_, new_n58557_ );
nor  ( new_n58563_, new_n58562_, new_n58556_ );
nor  ( new_n58564_, new_n58563_, new_n58547_ );
xor  ( new_n58565_, new_n58025_, new_n58024_ );
and  ( new_n58566_, new_n44319_, RIbb2d888_64 );
or   ( new_n58567_, new_n58566_, RIbb2d900_63 );
nand ( new_n58568_, new_n58566_, RIbb2d900_63 );
or   ( new_n58569_, new_n44587_, RIbb2d888_64 );
and  ( new_n58570_, new_n58569_, new_n58568_ );
and  ( new_n58571_, new_n58570_, new_n58567_ );
and  ( new_n58572_, new_n58571_, new_n58565_ );
nor  ( new_n58573_, new_n58326_, new_n7734_ );
xor  ( new_n58574_, new_n45584_, RIbb2ddb0_53 );
and  ( new_n58575_, new_n58574_, new_n7489_ );
or   ( new_n58576_, new_n58575_, new_n58573_ );
xor  ( new_n58577_, new_n58571_, new_n58565_ );
and  ( new_n58578_, new_n58577_, new_n58576_ );
nor  ( new_n58579_, new_n58578_, new_n58572_ );
not  ( new_n58580_, new_n58579_ );
and  ( new_n58581_, new_n58563_, new_n58547_ );
not  ( new_n58582_, new_n58581_ );
and  ( new_n58583_, new_n58582_, new_n58580_ );
nor  ( new_n58584_, new_n58583_, new_n58564_ );
xor  ( new_n58585_, new_n58330_, new_n58329_ );
xor  ( new_n58586_, new_n58312_, new_n58311_ );
nand ( new_n58587_, new_n58586_, new_n58585_ );
nor  ( new_n58588_, new_n58586_, new_n58585_ );
or   ( new_n58589_, new_n58016_, new_n1366_ );
xor  ( new_n58590_, new_n52293_, RIbb2ecb0_21 );
or   ( new_n58591_, new_n58590_, new_n1364_ );
and  ( new_n58592_, new_n58591_, new_n58589_ );
nor  ( new_n58593_, new_n58408_, new_n1137_ );
xor  ( new_n58594_, new_n53306_, RIbb2eda0_19 );
nor  ( new_n58595_, new_n58594_, new_n1135_ );
or   ( new_n58596_, new_n58595_, new_n58593_ );
and  ( new_n58597_, new_n53694_, new_n820_ );
nand ( new_n58598_, new_n58597_, new_n58596_ );
nor  ( new_n58599_, new_n58590_, new_n1366_ );
xor  ( new_n58600_, new_n52902_, RIbb2ecb0_21 );
nor  ( new_n58601_, new_n58600_, new_n1364_ );
or   ( new_n58602_, new_n58601_, new_n58599_ );
xor  ( new_n58603_, new_n58597_, new_n58596_ );
nand ( new_n58604_, new_n58603_, new_n58602_ );
and  ( new_n58605_, new_n58604_, new_n58598_ );
or   ( new_n58606_, new_n58605_, new_n58592_ );
nor  ( new_n58607_, new_n58461_, new_n2124_ );
xor  ( new_n58608_, new_n50894_, new_n1840_ );
nor  ( new_n58609_, new_n58608_, new_n2122_ );
or   ( new_n58610_, new_n58609_, new_n58607_ );
xor  ( new_n58611_, new_n58605_, new_n58592_ );
nand ( new_n58612_, new_n58611_, new_n58610_ );
and  ( new_n58613_, new_n58612_, new_n58606_ );
xor  ( new_n58614_, new_n44785_, RIbb2dae0_59 );
nand ( new_n58615_, new_n58614_, new_n9187_ );
or   ( new_n58616_, new_n58317_, new_n9424_ );
and  ( new_n58617_, new_n58616_, new_n58615_ );
or   ( new_n58618_, new_n58617_, new_n58613_ );
and  ( new_n58619_, new_n58477_, new_n6908_ );
xor  ( new_n58620_, new_n45597_, RIbb2dea0_51 );
and  ( new_n58621_, new_n58620_, new_n6910_ );
or   ( new_n58622_, new_n58621_, new_n58619_ );
xor  ( new_n58623_, new_n58617_, new_n58613_ );
nand ( new_n58624_, new_n58623_, new_n58622_ );
and  ( new_n58625_, new_n58624_, new_n58618_ );
or   ( new_n58626_, new_n58625_, new_n58588_ );
and  ( new_n58627_, new_n58626_, new_n58587_ );
or   ( new_n58628_, new_n58627_, new_n58584_ );
and  ( new_n58629_, new_n58627_, new_n58584_ );
xor  ( new_n58630_, new_n58275_, new_n58273_ );
xnor ( new_n58631_, new_n58630_, new_n58295_ );
not  ( new_n58632_, new_n58631_ );
or   ( new_n58633_, new_n58632_, new_n58629_ );
and  ( new_n58634_, new_n58633_, new_n58628_ );
and  ( new_n58635_, new_n58634_, new_n58531_ );
or   ( new_n58636_, new_n58635_, new_n58530_ );
xnor ( new_n58637_, new_n58110_, new_n58108_ );
xor  ( new_n58638_, new_n58637_, new_n58122_ );
and  ( new_n58639_, new_n58638_, new_n58636_ );
or   ( new_n58640_, new_n58638_, new_n58636_ );
xor  ( new_n58641_, new_n58340_, new_n58338_ );
xor  ( new_n58642_, new_n58641_, new_n58344_ );
and  ( new_n58643_, new_n58642_, new_n58640_ );
or   ( new_n58644_, new_n58643_, new_n58639_ );
or   ( new_n58645_, new_n58644_, new_n58498_ );
and  ( new_n58646_, new_n58645_, new_n58497_ );
nor  ( new_n58647_, new_n58646_, new_n58370_ );
nor  ( new_n58648_, new_n58647_, new_n58368_ );
not  ( new_n58649_, new_n58648_ );
xor  ( new_n58650_, new_n58357_, new_n58355_ );
xnor ( new_n58651_, new_n58650_, new_n58361_ );
and  ( new_n58652_, new_n58651_, new_n58649_ );
xor  ( new_n58653_, new_n58623_, new_n58622_ );
xor  ( new_n58654_, new_n58577_, new_n58576_ );
xor  ( new_n58655_, new_n58654_, new_n58653_ );
xnor ( new_n58656_, new_n58514_, new_n58510_ );
xor  ( new_n58657_, new_n58656_, new_n58519_ );
xor  ( new_n58658_, new_n58657_, new_n58655_ );
xor  ( new_n58659_, new_n50788_, new_n2118_ );
nor  ( new_n58660_, new_n58659_, new_n2425_ );
xor  ( new_n58661_, new_n50487_, new_n2118_ );
nor  ( new_n58662_, new_n58661_, new_n2427_ );
or   ( new_n58663_, new_n58662_, new_n58660_ );
xor  ( new_n58664_, new_n58603_, new_n58602_ );
and  ( new_n58665_, new_n58664_, new_n58663_ );
xor  ( new_n58666_, new_n51142_, new_n1840_ );
nor  ( new_n58667_, new_n58666_, new_n2122_ );
nor  ( new_n58668_, new_n58608_, new_n2124_ );
or   ( new_n58669_, new_n58668_, new_n58667_ );
xor  ( new_n58670_, new_n58664_, new_n58663_ );
and  ( new_n58671_, new_n58670_, new_n58669_ );
or   ( new_n58672_, new_n58671_, new_n58665_ );
xor  ( new_n58673_, new_n58611_, new_n58610_ );
xor  ( new_n58674_, new_n58673_, new_n58672_ );
and  ( new_n58675_, new_n58537_, new_n2613_ );
xor  ( new_n58676_, new_n49758_, new_n2421_ );
nor  ( new_n58677_, new_n58676_, new_n2807_ );
or   ( new_n58678_, new_n58677_, new_n58675_ );
or   ( new_n58679_, new_n58532_, new_n2427_ );
or   ( new_n58680_, new_n58661_, new_n2425_ );
and  ( new_n58681_, new_n58680_, new_n58679_ );
or   ( new_n58682_, new_n58468_, new_n1846_ );
xor  ( new_n58683_, new_n51446_, new_n1583_ );
or   ( new_n58684_, new_n58683_, new_n1844_ );
and  ( new_n58685_, new_n58684_, new_n58682_ );
xor  ( new_n58686_, new_n58685_, new_n58681_ );
xor  ( new_n58687_, new_n58686_, new_n58678_ );
xor  ( new_n58688_, new_n58687_, new_n58674_ );
and  ( new_n58689_, new_n44506_, new_n21077_ );
not  ( new_n58690_, new_n58689_ );
and  ( new_n58691_, new_n44407_, RIbb2d888_64 );
nor  ( new_n58692_, new_n58691_, new_n10052_ );
and  ( new_n58693_, new_n58692_, new_n58690_ );
and  ( new_n58694_, new_n58691_, new_n10052_ );
nor  ( new_n58695_, new_n58694_, new_n58693_ );
or   ( new_n58696_, new_n58512_, new_n8266_ );
xor  ( new_n58697_, new_n45403_, new_n7722_ );
or   ( new_n58698_, new_n58697_, new_n8264_ );
and  ( new_n58699_, new_n58698_, new_n58696_ );
nand ( new_n58700_, new_n58517_, new_n8649_ );
xor  ( new_n58701_, new_n45119_, new_n8254_ );
or   ( new_n58702_, new_n58701_, new_n8874_ );
and  ( new_n58703_, new_n58702_, new_n58700_ );
xnor ( new_n58704_, new_n58703_, new_n58699_ );
xor  ( new_n58705_, new_n58704_, new_n58695_ );
or   ( new_n58706_, new_n58705_, new_n58688_ );
xor  ( new_n58707_, new_n46619_, new_n5594_ );
nor  ( new_n58708_, new_n58707_, new_n6175_ );
xor  ( new_n58709_, new_n46789_, new_n5594_ );
nor  ( new_n58710_, new_n58709_, new_n6173_ );
or   ( new_n58711_, new_n58710_, new_n58708_ );
or   ( new_n58712_, new_n58676_, new_n2809_ );
xor  ( new_n58713_, new_n50115_, new_n2421_ );
or   ( new_n58714_, new_n58713_, new_n2807_ );
and  ( new_n58715_, new_n58714_, new_n58712_ );
xor  ( new_n58716_, new_n49427_, RIbb2e710_33 );
nand ( new_n58717_, new_n58716_, new_n2928_ );
xor  ( new_n58718_, new_n49488_, new_n2797_ );
or   ( new_n58719_, new_n58718_, new_n3117_ );
and  ( new_n58720_, new_n58719_, new_n58717_ );
xor  ( new_n58721_, new_n58720_, new_n58715_ );
xor  ( new_n58722_, new_n58721_, new_n58711_ );
xor  ( new_n58723_, new_n58670_, new_n58669_ );
and  ( new_n58724_, new_n58723_, new_n58722_ );
and  ( new_n58725_, new_n53694_, new_n44802_ );
or   ( new_n58726_, new_n58725_, new_n1129_ );
xor  ( new_n58727_, new_n53306_, RIbb2ecb0_21 );
or   ( new_n58728_, new_n58727_, new_n1366_ );
nor  ( new_n58729_, new_n53694_, RIbb2ecb0_21 );
and  ( new_n58730_, new_n53694_, RIbb2ecb0_21 );
or   ( new_n58731_, new_n58730_, new_n1364_ );
or   ( new_n58732_, new_n58731_, new_n58729_ );
and  ( new_n58733_, new_n58732_, new_n58728_ );
or   ( new_n58734_, new_n58733_, new_n58726_ );
xor  ( new_n58735_, new_n52280_, new_n1583_ );
or   ( new_n58736_, new_n58735_, new_n1844_ );
xor  ( new_n58737_, new_n51758_, new_n1583_ );
or   ( new_n58738_, new_n58737_, new_n1846_ );
and  ( new_n58739_, new_n58738_, new_n58736_ );
or   ( new_n58740_, new_n58739_, new_n58734_ );
xor  ( new_n58741_, new_n51446_, RIbb2e9e0_27 );
and  ( new_n58742_, new_n58741_, new_n2000_ );
xor  ( new_n58743_, new_n51477_, RIbb2e9e0_27 );
and  ( new_n58744_, new_n58743_, new_n2002_ );
or   ( new_n58745_, new_n58744_, new_n58742_ );
xor  ( new_n58746_, new_n58739_, new_n58734_ );
nand ( new_n58747_, new_n58746_, new_n58745_ );
and  ( new_n58748_, new_n58747_, new_n58740_ );
xor  ( new_n58749_, new_n48291_, new_n3892_ );
or   ( new_n58750_, new_n58749_, new_n4304_ );
xor  ( new_n58751_, new_n48518_, new_n3892_ );
or   ( new_n58752_, new_n58751_, new_n4302_ );
and  ( new_n58753_, new_n58752_, new_n58750_ );
nor  ( new_n58754_, new_n58753_, new_n58748_ );
xor  ( new_n58755_, new_n48756_, RIbb2e530_37 );
and  ( new_n58756_, new_n58755_, new_n3731_ );
xor  ( new_n58757_, new_n48908_, new_n3457_ );
nor  ( new_n58758_, new_n58757_, new_n3896_ );
nor  ( new_n58759_, new_n58758_, new_n58756_ );
not  ( new_n58760_, new_n58759_ );
xor  ( new_n58761_, new_n58753_, new_n58748_ );
and  ( new_n58762_, new_n58761_, new_n58760_ );
or   ( new_n58763_, new_n58762_, new_n58754_ );
xor  ( new_n58764_, new_n58723_, new_n58722_ );
and  ( new_n58765_, new_n58764_, new_n58763_ );
or   ( new_n58766_, new_n58765_, new_n58724_ );
and  ( new_n58767_, new_n58705_, new_n58688_ );
or   ( new_n58768_, new_n58767_, new_n58766_ );
and  ( new_n58769_, new_n58768_, new_n58706_ );
nand ( new_n58770_, new_n58769_, new_n58658_ );
or   ( new_n58771_, new_n58720_, new_n58715_ );
nand ( new_n58772_, new_n58721_, new_n58711_ );
and  ( new_n58773_, new_n58772_, new_n58771_ );
nor  ( new_n58774_, new_n58600_, new_n1366_ );
xor  ( new_n58775_, new_n52908_, RIbb2ecb0_21 );
nor  ( new_n58776_, new_n58775_, new_n1364_ );
or   ( new_n58777_, new_n58776_, new_n58774_ );
and  ( new_n58778_, new_n53694_, new_n44565_ );
or   ( new_n58779_, new_n58778_, new_n896_ );
or   ( new_n58780_, new_n58594_, new_n1137_ );
and  ( new_n58781_, new_n44563_, RIbb2eda0_19 );
nor  ( new_n58782_, new_n58730_, new_n58781_ );
and  ( new_n58783_, RIbb2ed28_20, new_n893_ );
nor  ( new_n58784_, new_n58729_, new_n58783_ );
or   ( new_n58785_, new_n58784_, new_n58782_ );
and  ( new_n58786_, new_n58785_, new_n58780_ );
xor  ( new_n58787_, new_n58786_, new_n58779_ );
nand ( new_n58788_, new_n58787_, new_n58777_ );
xor  ( new_n58789_, new_n51477_, RIbb2ead0_25 );
and  ( new_n58790_, new_n58789_, new_n1739_ );
nor  ( new_n58791_, new_n58737_, new_n1844_ );
or   ( new_n58792_, new_n58791_, new_n58790_ );
xor  ( new_n58793_, new_n58787_, new_n58777_ );
nand ( new_n58794_, new_n58793_, new_n58792_ );
and  ( new_n58795_, new_n58794_, new_n58788_ );
or   ( new_n58796_, new_n58749_, new_n4302_ );
xor  ( new_n58797_, new_n48039_, new_n3892_ );
or   ( new_n58798_, new_n58797_, new_n4304_ );
and  ( new_n58799_, new_n58798_, new_n58796_ );
or   ( new_n58800_, new_n58799_, new_n58795_ );
xor  ( new_n58801_, new_n47296_, RIbb2e350_41 );
and  ( new_n58802_, new_n58801_, new_n4541_ );
xor  ( new_n58803_, new_n47640_, new_n4292_ );
nor  ( new_n58804_, new_n58803_, new_n4709_ );
nor  ( new_n58805_, new_n58804_, new_n58802_ );
not  ( new_n58806_, new_n58805_ );
xor  ( new_n58807_, new_n58799_, new_n58795_ );
nand ( new_n58808_, new_n58807_, new_n58806_ );
and  ( new_n58809_, new_n58808_, new_n58800_ );
xor  ( new_n58810_, new_n47046_, new_n4705_ );
or   ( new_n58811_, new_n58810_, new_n5207_ );
xor  ( new_n58812_, new_n47303_, new_n4705_ );
or   ( new_n58813_, new_n58812_, new_n5209_ );
and  ( new_n58814_, new_n58813_, new_n58811_ );
xor  ( new_n58815_, new_n46427_, new_n6163_ );
or   ( new_n58816_, new_n58815_, new_n6645_ );
xor  ( new_n58817_, new_n46137_, new_n6163_ );
or   ( new_n58818_, new_n58817_, new_n6647_ );
and  ( new_n58819_, new_n58818_, new_n58816_ );
or   ( new_n58820_, new_n58819_, new_n58814_ );
xor  ( new_n58821_, new_n46962_, new_n5203_ );
nor  ( new_n58822_, new_n58821_, new_n5606_ );
xor  ( new_n58823_, new_n46958_, RIbb2e170_45 );
and  ( new_n58824_, new_n58823_, new_n5373_ );
or   ( new_n58825_, new_n58824_, new_n58822_ );
xor  ( new_n58826_, new_n58819_, new_n58814_ );
nand ( new_n58827_, new_n58826_, new_n58825_ );
and  ( new_n58828_, new_n58827_, new_n58820_ );
xor  ( new_n58829_, new_n58828_, new_n58809_ );
xor  ( new_n58830_, new_n58829_, new_n58773_ );
xor  ( new_n58831_, new_n48039_, RIbb2e350_41 );
and  ( new_n58832_, new_n58831_, new_n4543_ );
nor  ( new_n58833_, new_n58803_, new_n4711_ );
or   ( new_n58834_, new_n58833_, new_n58832_ );
xor  ( new_n58835_, new_n58793_, new_n58792_ );
nand ( new_n58836_, new_n58835_, new_n58834_ );
nor  ( new_n58837_, new_n58810_, new_n5209_ );
xor  ( new_n58838_, new_n47296_, RIbb2e260_43 );
and  ( new_n58839_, new_n58838_, new_n4960_ );
nor  ( new_n58840_, new_n58839_, new_n58837_ );
not  ( new_n58841_, new_n58840_ );
xor  ( new_n58842_, new_n58835_, new_n58834_ );
nand ( new_n58843_, new_n58842_, new_n58841_ );
and  ( new_n58844_, new_n58843_, new_n58836_ );
xor  ( new_n58845_, new_n46962_, new_n5594_ );
or   ( new_n58846_, new_n58845_, new_n6173_ );
or   ( new_n58847_, new_n58709_, new_n6175_ );
and  ( new_n58848_, new_n58847_, new_n58846_ );
xor  ( new_n58849_, new_n46619_, new_n6163_ );
or   ( new_n58850_, new_n58849_, new_n6645_ );
or   ( new_n58851_, new_n58815_, new_n6647_ );
and  ( new_n58852_, new_n58851_, new_n58850_ );
or   ( new_n58853_, new_n58852_, new_n58848_ );
and  ( new_n58854_, new_n58823_, new_n5371_ );
xor  ( new_n58855_, new_n47303_, new_n5203_ );
nor  ( new_n58856_, new_n58855_, new_n5604_ );
nor  ( new_n58857_, new_n58856_, new_n58854_ );
and  ( new_n58858_, new_n58852_, new_n58848_ );
or   ( new_n58859_, new_n58858_, new_n58857_ );
and  ( new_n58860_, new_n58859_, new_n58853_ );
or   ( new_n58861_, new_n58860_, new_n58844_ );
and  ( new_n58862_, new_n58860_, new_n58844_ );
xor  ( new_n58863_, new_n45204_, RIbb2dbd0_57 );
and  ( new_n58864_, new_n58863_, new_n8649_ );
xor  ( new_n58865_, new_n45403_, new_n8254_ );
nor  ( new_n58866_, new_n58865_, new_n8874_ );
nor  ( new_n58867_, new_n58866_, new_n58864_ );
xor  ( new_n58868_, new_n49265_, new_n3113_ );
nor  ( new_n58869_, new_n58868_, new_n3463_ );
xor  ( new_n58870_, new_n49427_, RIbb2e620_35 );
and  ( new_n58871_, new_n58870_, new_n3293_ );
nor  ( new_n58872_, new_n58871_, new_n58869_ );
nor  ( new_n58873_, new_n58872_, new_n58867_ );
and  ( new_n58874_, new_n58872_, new_n58867_ );
and  ( new_n58875_, new_n44600_, RIbb2d888_64 );
not  ( new_n58876_, new_n58875_ );
and  ( new_n58877_, new_n44681_, new_n21077_ );
nor  ( new_n58878_, new_n58877_, new_n10052_ );
and  ( new_n58879_, new_n58878_, new_n58876_ );
and  ( new_n58880_, new_n58875_, new_n10052_ );
nor  ( new_n58881_, new_n58880_, new_n58879_ );
nor  ( new_n58882_, new_n58881_, new_n58874_ );
nor  ( new_n58883_, new_n58882_, new_n58873_ );
or   ( new_n58884_, new_n58883_, new_n58862_ );
and  ( new_n58885_, new_n58884_, new_n58861_ );
nor  ( new_n58886_, new_n58885_, new_n58830_ );
xor  ( new_n58887_, new_n58807_, new_n58806_ );
xor  ( new_n58888_, new_n58826_, new_n58825_ );
and  ( new_n58889_, new_n58888_, new_n58887_ );
xnor ( new_n58890_, new_n58888_, new_n58887_ );
xor  ( new_n58891_, new_n44785_, RIbb2d9f0_61 );
nand ( new_n58892_, new_n58891_, new_n9738_ );
xor  ( new_n58893_, new_n44877_, RIbb2d9f0_61 );
nand ( new_n58894_, new_n58893_, new_n9740_ );
and  ( new_n58895_, new_n58894_, new_n58892_ );
xor  ( new_n58896_, new_n45738_, RIbb2dcc0_55 );
nand ( new_n58897_, new_n58896_, new_n8042_ );
xor  ( new_n58898_, new_n45584_, new_n7722_ );
or   ( new_n58899_, new_n58898_, new_n8266_ );
and  ( new_n58900_, new_n58899_, new_n58897_ );
nor  ( new_n58901_, new_n58900_, new_n58895_ );
and  ( new_n58902_, new_n58900_, new_n58895_ );
xor  ( new_n58903_, new_n45597_, RIbb2ddb0_53 );
and  ( new_n58904_, new_n58903_, new_n7487_ );
xor  ( new_n58905_, new_n45928_, new_n7174_ );
nor  ( new_n58906_, new_n58905_, new_n7732_ );
nor  ( new_n58907_, new_n58906_, new_n58904_ );
nor  ( new_n58908_, new_n58907_, new_n58902_ );
nor  ( new_n58909_, new_n58908_, new_n58901_ );
nor  ( new_n58910_, new_n58909_, new_n58890_ );
or   ( new_n58911_, new_n58910_, new_n58889_ );
xor  ( new_n58912_, new_n58885_, new_n58830_ );
and  ( new_n58913_, new_n58912_, new_n58911_ );
or   ( new_n58914_, new_n58913_, new_n58886_ );
xor  ( new_n58915_, new_n58769_, new_n58658_ );
nand ( new_n58916_, new_n58915_, new_n58914_ );
and  ( new_n58917_, new_n58916_, new_n58770_ );
nand ( new_n58918_, new_n58654_, new_n58653_ );
nand ( new_n58919_, new_n58657_, new_n58655_ );
and  ( new_n58920_, new_n58919_, new_n58918_ );
xnor ( new_n58921_, new_n58522_, new_n58506_ );
xor  ( new_n58922_, new_n58482_, new_n58481_ );
xor  ( new_n58923_, new_n58455_, new_n58454_ );
xnor ( new_n58924_, new_n58287_, new_n58281_ );
xor  ( new_n58925_, new_n58924_, new_n58293_ );
xnor ( new_n58926_, new_n58925_, new_n58923_ );
xor  ( new_n58927_, new_n58926_, new_n58922_ );
xor  ( new_n58928_, new_n58927_, new_n58921_ );
xor  ( new_n58929_, new_n58928_, new_n58920_ );
or   ( new_n58930_, new_n58929_, new_n58917_ );
and  ( new_n58931_, new_n58673_, new_n58672_ );
and  ( new_n58932_, new_n58687_, new_n58674_ );
nor  ( new_n58933_, new_n58932_, new_n58931_ );
or   ( new_n58934_, new_n58828_, new_n58809_ );
and  ( new_n58935_, new_n58828_, new_n58809_ );
or   ( new_n58936_, new_n58935_, new_n58773_ );
and  ( new_n58937_, new_n58936_, new_n58934_ );
xor  ( new_n58938_, new_n58937_, new_n58933_ );
not  ( new_n58939_, new_n58938_ );
or   ( new_n58940_, new_n58414_, new_n1595_ );
xor  ( new_n58941_, new_n52280_, new_n1355_ );
or   ( new_n58942_, new_n58941_, new_n1593_ );
and  ( new_n58943_, new_n58942_, new_n58940_ );
or   ( new_n58944_, new_n58683_, new_n1846_ );
nand ( new_n58945_, new_n58789_, new_n1741_ );
and  ( new_n58946_, new_n58945_, new_n58944_ );
nand ( new_n58947_, new_n58946_, new_n58943_ );
nor  ( new_n58948_, new_n58786_, new_n58779_ );
nor  ( new_n58949_, new_n58946_, new_n58943_ );
or   ( new_n58950_, new_n58949_, new_n58948_ );
and  ( new_n58951_, new_n58950_, new_n58947_ );
or   ( new_n58952_, new_n58425_, new_n4304_ );
or   ( new_n58953_, new_n58797_, new_n4302_ );
and  ( new_n58954_, new_n58953_, new_n58952_ );
or   ( new_n58955_, new_n58553_, new_n3898_ );
xor  ( new_n58956_, new_n48518_, RIbb2e530_37 );
nand ( new_n58957_, new_n58956_, new_n3733_ );
and  ( new_n58958_, new_n58957_, new_n58955_ );
xor  ( new_n58959_, new_n58958_, new_n58954_ );
xor  ( new_n58960_, new_n58959_, new_n58951_ );
nor  ( new_n58961_, new_n58542_, new_n3119_ );
and  ( new_n58962_, new_n58716_, new_n2930_ );
nor  ( new_n58963_, new_n58962_, new_n58961_ );
or   ( new_n58964_, new_n58821_, new_n5604_ );
or   ( new_n58965_, new_n58384_, new_n5606_ );
and  ( new_n58966_, new_n58965_, new_n58964_ );
or   ( new_n58967_, new_n58707_, new_n6173_ );
nand ( new_n58968_, new_n58393_, new_n5915_ );
and  ( new_n58969_, new_n58968_, new_n58967_ );
xnor ( new_n58970_, new_n58969_, new_n58966_ );
xor  ( new_n58971_, new_n58970_, new_n58963_ );
nand ( new_n58972_, new_n58971_, new_n58960_ );
nor  ( new_n58973_, new_n58971_, new_n58960_ );
and  ( new_n58974_, new_n58801_, new_n4543_ );
nor  ( new_n58975_, new_n58421_, new_n4711_ );
nor  ( new_n58976_, new_n58975_, new_n58974_ );
and  ( new_n58977_, new_n58387_, new_n4958_ );
nor  ( new_n58978_, new_n58812_, new_n5207_ );
or   ( new_n58979_, new_n58978_, new_n58977_ );
xor  ( new_n58980_, new_n58417_, new_n58416_ );
xnor ( new_n58981_, new_n58980_, new_n58979_ );
xnor ( new_n58982_, new_n58981_, new_n58976_ );
or   ( new_n58983_, new_n58982_, new_n58973_ );
and  ( new_n58984_, new_n58983_, new_n58972_ );
xor  ( new_n58985_, new_n58984_, new_n58939_ );
or   ( new_n58986_, new_n58868_, new_n3461_ );
xor  ( new_n58987_, new_n48908_, new_n3113_ );
or   ( new_n58988_, new_n58987_, new_n3463_ );
and  ( new_n58989_, new_n58988_, new_n58986_ );
nand ( new_n58990_, new_n58863_, new_n8651_ );
or   ( new_n58991_, new_n58701_, new_n8876_ );
and  ( new_n58992_, new_n58991_, new_n58990_ );
or   ( new_n58993_, new_n58992_, new_n58989_ );
and  ( new_n58994_, new_n58956_, new_n3731_ );
and  ( new_n58995_, new_n58755_, new_n3733_ );
nor  ( new_n58996_, new_n58995_, new_n58994_ );
xnor ( new_n58997_, new_n58992_, new_n58989_ );
or   ( new_n58998_, new_n58997_, new_n58996_ );
and  ( new_n58999_, new_n58998_, new_n58993_ );
xor  ( new_n59000_, new_n44974_, RIbb2dae0_59 );
nand ( new_n59001_, new_n59000_, new_n9187_ );
xor  ( new_n59002_, new_n44877_, RIbb2dae0_59 );
nand ( new_n59003_, new_n59002_, new_n9185_ );
and  ( new_n59004_, new_n59003_, new_n59001_ );
xnor ( new_n59005_, new_n58946_, new_n58943_ );
xor  ( new_n59006_, new_n59005_, new_n58948_ );
or   ( new_n59007_, new_n59006_, new_n59004_ );
and  ( new_n59008_, new_n59006_, new_n59004_ );
and  ( new_n59009_, new_n58903_, new_n7489_ );
xor  ( new_n59010_, new_n45738_, RIbb2ddb0_53 );
and  ( new_n59011_, new_n59010_, new_n7487_ );
nor  ( new_n59012_, new_n59011_, new_n59009_ );
or   ( new_n59013_, new_n59012_, new_n59008_ );
and  ( new_n59014_, new_n59013_, new_n59007_ );
nor  ( new_n59015_, new_n59014_, new_n58999_ );
or   ( new_n59016_, new_n58697_, new_n8266_ );
or   ( new_n59017_, new_n58898_, new_n8264_ );
and  ( new_n59018_, new_n59017_, new_n59016_ );
and  ( new_n59019_, new_n44506_, RIbb2d888_64 );
and  ( new_n59020_, new_n44600_, new_n21077_ );
or   ( new_n59021_, new_n59020_, new_n10052_ );
or   ( new_n59022_, new_n59021_, new_n59019_ );
nand ( new_n59023_, new_n59019_, new_n10052_ );
and  ( new_n59024_, new_n59023_, new_n59022_ );
nor  ( new_n59025_, new_n59024_, new_n59018_ );
and  ( new_n59026_, new_n58891_, new_n9740_ );
xor  ( new_n59027_, new_n44681_, RIbb2d9f0_61 );
and  ( new_n59028_, new_n59027_, new_n9738_ );
nor  ( new_n59029_, new_n59028_, new_n59026_ );
not  ( new_n59030_, new_n59029_ );
xor  ( new_n59031_, new_n59024_, new_n59018_ );
and  ( new_n59032_, new_n59031_, new_n59030_ );
or   ( new_n59033_, new_n59032_, new_n59025_ );
xor  ( new_n59034_, new_n59014_, new_n58999_ );
and  ( new_n59035_, new_n59034_, new_n59033_ );
or   ( new_n59036_, new_n59035_, new_n59015_ );
and  ( new_n59037_, new_n58980_, new_n58979_ );
nor  ( new_n59038_, new_n58981_, new_n58976_ );
nor  ( new_n59039_, new_n59038_, new_n59037_ );
xnor ( new_n59040_, new_n58471_, new_n58470_ );
xnor ( new_n59041_, new_n59040_, new_n59039_ );
or   ( new_n59042_, new_n58969_, new_n58966_ );
and  ( new_n59043_, new_n58969_, new_n58966_ );
or   ( new_n59044_, new_n59043_, new_n58963_ );
and  ( new_n59045_, new_n59044_, new_n59042_ );
xor  ( new_n59046_, new_n59045_, new_n59041_ );
nor  ( new_n59047_, new_n58685_, new_n58681_ );
and  ( new_n59048_, new_n58686_, new_n58678_ );
or   ( new_n59049_, new_n59048_, new_n59047_ );
xor  ( new_n59050_, new_n58545_, new_n58544_ );
xor  ( new_n59051_, new_n59050_, new_n59049_ );
nand ( new_n59052_, new_n58958_, new_n58954_ );
nor  ( new_n59053_, new_n58958_, new_n58954_ );
or   ( new_n59054_, new_n59053_, new_n58951_ );
and  ( new_n59055_, new_n59054_, new_n59052_ );
xor  ( new_n59056_, new_n59055_, new_n59051_ );
xor  ( new_n59057_, new_n59056_, new_n59046_ );
xor  ( new_n59058_, new_n59057_, new_n59036_ );
and  ( new_n59059_, new_n59058_, new_n58985_ );
xor  ( new_n59060_, new_n59058_, new_n58985_ );
xor  ( new_n59061_, new_n59034_, new_n59033_ );
xnor ( new_n59062_, new_n58997_, new_n58996_ );
and  ( new_n59063_, new_n59000_, new_n9185_ );
xor  ( new_n59064_, new_n45119_, new_n8870_ );
nor  ( new_n59065_, new_n59064_, new_n9422_ );
or   ( new_n59066_, new_n59065_, new_n59063_ );
nor  ( new_n59067_, new_n58659_, new_n2427_ );
xor  ( new_n59068_, new_n50894_, new_n2118_ );
nor  ( new_n59069_, new_n59068_, new_n2425_ );
or   ( new_n59070_, new_n59069_, new_n59067_ );
or   ( new_n59071_, new_n58941_, new_n1595_ );
xor  ( new_n59072_, new_n52293_, RIbb2ebc0_23 );
or   ( new_n59073_, new_n59072_, new_n1593_ );
and  ( new_n59074_, new_n59073_, new_n59071_ );
nor  ( new_n59075_, new_n58775_, new_n1366_ );
nor  ( new_n59076_, new_n58727_, new_n1364_ );
or   ( new_n59077_, new_n59076_, new_n59075_ );
and  ( new_n59078_, new_n53694_, new_n1040_ );
nand ( new_n59079_, new_n59078_, new_n59077_ );
xor  ( new_n59080_, new_n52902_, RIbb2ebc0_23 );
nor  ( new_n59081_, new_n59080_, new_n1593_ );
nor  ( new_n59082_, new_n59072_, new_n1595_ );
or   ( new_n59083_, new_n59082_, new_n59081_ );
xor  ( new_n59084_, new_n59078_, new_n59077_ );
nand ( new_n59085_, new_n59084_, new_n59083_ );
and  ( new_n59086_, new_n59085_, new_n59079_ );
xor  ( new_n59087_, new_n59086_, new_n59074_ );
xor  ( new_n59088_, new_n59087_, new_n59070_ );
nand ( new_n59089_, new_n59088_, new_n59066_ );
xor  ( new_n59090_, new_n46037_, new_n6635_ );
nor  ( new_n59091_, new_n59090_, new_n7186_ );
xor  ( new_n59092_, new_n46137_, RIbb2dea0_51 );
and  ( new_n59093_, new_n59092_, new_n6910_ );
nor  ( new_n59094_, new_n59093_, new_n59091_ );
not  ( new_n59095_, new_n59094_ );
xor  ( new_n59096_, new_n59088_, new_n59066_ );
nand ( new_n59097_, new_n59096_, new_n59095_ );
and  ( new_n59098_, new_n59097_, new_n59089_ );
nand ( new_n59099_, new_n59098_, new_n59062_ );
xor  ( new_n59100_, new_n59031_, new_n59030_ );
nor  ( new_n59101_, new_n59098_, new_n59062_ );
or   ( new_n59102_, new_n59101_, new_n59100_ );
and  ( new_n59103_, new_n59102_, new_n59099_ );
nand ( new_n59104_, new_n59103_, new_n59061_ );
nor  ( new_n59105_, new_n59103_, new_n59061_ );
xor  ( new_n59106_, new_n58971_, new_n58960_ );
xor  ( new_n59107_, new_n59106_, new_n58982_ );
or   ( new_n59108_, new_n59107_, new_n59105_ );
nand ( new_n59109_, new_n59108_, new_n59104_ );
and  ( new_n59110_, new_n59109_, new_n59060_ );
or   ( new_n59111_, new_n59110_, new_n59059_ );
xor  ( new_n59112_, new_n58929_, new_n58917_ );
nand ( new_n59113_, new_n59112_, new_n59111_ );
and  ( new_n59114_, new_n59113_, new_n58930_ );
nor  ( new_n59115_, new_n58937_, new_n58933_ );
nor  ( new_n59116_, new_n58984_, new_n58939_ );
nor  ( new_n59117_, new_n59116_, new_n59115_ );
xor  ( new_n59118_, new_n58586_, new_n58585_ );
xor  ( new_n59119_, new_n59118_, new_n58625_ );
xor  ( new_n59120_, new_n59119_, new_n59117_ );
and  ( new_n59121_, new_n59050_, new_n59049_ );
and  ( new_n59122_, new_n59055_, new_n59051_ );
nor  ( new_n59123_, new_n59122_, new_n59121_ );
nor  ( new_n59124_, new_n59040_, new_n59039_ );
nor  ( new_n59125_, new_n59045_, new_n59041_ );
nor  ( new_n59126_, new_n59125_, new_n59124_ );
nand ( new_n59127_, new_n58620_, new_n6908_ );
xor  ( new_n59128_, new_n45928_, new_n6635_ );
or   ( new_n59129_, new_n59128_, new_n7184_ );
and  ( new_n59130_, new_n59129_, new_n59127_ );
nand ( new_n59131_, new_n58574_, new_n7487_ );
nand ( new_n59132_, new_n59010_, new_n7489_ );
and  ( new_n59133_, new_n59132_, new_n59131_ );
nor  ( new_n59134_, new_n59133_, new_n59130_ );
and  ( new_n59135_, new_n58614_, new_n9185_ );
and  ( new_n59136_, new_n59002_, new_n9187_ );
nor  ( new_n59137_, new_n59136_, new_n59135_ );
and  ( new_n59138_, new_n59133_, new_n59130_ );
nor  ( new_n59139_, new_n59138_, new_n59137_ );
nor  ( new_n59140_, new_n59139_, new_n59134_ );
or   ( new_n59141_, new_n58703_, new_n58699_ );
and  ( new_n59142_, new_n58703_, new_n58699_ );
or   ( new_n59143_, new_n59142_, new_n58695_ );
and  ( new_n59144_, new_n59143_, new_n59141_ );
nor  ( new_n59145_, new_n59144_, new_n59140_ );
or   ( new_n59146_, new_n58548_, new_n3463_ );
or   ( new_n59147_, new_n58987_, new_n3461_ );
and  ( new_n59148_, new_n59147_, new_n59146_ );
or   ( new_n59149_, new_n58559_, new_n6647_ );
or   ( new_n59150_, new_n58817_, new_n6645_ );
and  ( new_n59151_, new_n59150_, new_n59149_ );
nor  ( new_n59152_, new_n59151_, new_n59148_ );
and  ( new_n59153_, new_n58507_, new_n9738_ );
and  ( new_n59154_, new_n59027_, new_n9740_ );
nor  ( new_n59155_, new_n59154_, new_n59153_ );
not  ( new_n59156_, new_n59155_ );
xor  ( new_n59157_, new_n59151_, new_n59148_ );
and  ( new_n59158_, new_n59157_, new_n59156_ );
or   ( new_n59159_, new_n59158_, new_n59152_ );
xor  ( new_n59160_, new_n59144_, new_n59140_ );
and  ( new_n59161_, new_n59160_, new_n59159_ );
nor  ( new_n59162_, new_n59161_, new_n59145_ );
xnor ( new_n59163_, new_n59162_, new_n59126_ );
nand ( new_n59164_, new_n59163_, new_n59123_ );
nor  ( new_n59165_, new_n59162_, new_n59126_ );
and  ( new_n59166_, new_n59162_, new_n59126_ );
nor  ( new_n59167_, new_n59166_, new_n59123_ );
not  ( new_n59168_, new_n59167_ );
or   ( new_n59169_, new_n59168_, new_n59165_ );
and  ( new_n59170_, new_n59169_, new_n59164_ );
xnor ( new_n59171_, new_n59170_, new_n59120_ );
xor  ( new_n59172_, new_n58563_, new_n58547_ );
nor  ( new_n59173_, new_n59172_, new_n58580_ );
not  ( new_n59174_, new_n58564_ );
and  ( new_n59175_, new_n58583_, new_n59174_ );
nor  ( new_n59176_, new_n59175_, new_n59173_ );
xnor ( new_n59177_, new_n58431_, new_n58406_ );
xor  ( new_n59178_, new_n58396_, new_n58395_ );
xnor ( new_n59179_, new_n58555_, new_n58551_ );
xor  ( new_n59180_, new_n59179_, new_n58561_ );
nand ( new_n59181_, new_n59180_, new_n59178_ );
or   ( new_n59182_, new_n59180_, new_n59178_ );
xor  ( new_n59183_, new_n58423_, new_n58419_ );
xnor ( new_n59184_, new_n59183_, new_n58428_ );
nand ( new_n59185_, new_n59184_, new_n59182_ );
and  ( new_n59186_, new_n59185_, new_n59181_ );
xor  ( new_n59187_, new_n59186_, new_n59177_ );
xor  ( new_n59188_, new_n59187_, new_n59176_ );
and  ( new_n59189_, new_n59056_, new_n59046_ );
and  ( new_n59190_, new_n59057_, new_n59036_ );
or   ( new_n59191_, new_n59190_, new_n59189_ );
xor  ( new_n59192_, new_n59160_, new_n59159_ );
xor  ( new_n59193_, new_n59180_, new_n59178_ );
xor  ( new_n59194_, new_n59193_, new_n59184_ );
or   ( new_n59195_, new_n59194_, new_n59192_ );
nand ( new_n59196_, new_n59194_, new_n59192_ );
xor  ( new_n59197_, new_n59157_, new_n59156_ );
not  ( new_n59198_, new_n59197_ );
or   ( new_n59199_, new_n59128_, new_n7186_ );
or   ( new_n59200_, new_n59090_, new_n7184_ );
and  ( new_n59201_, new_n59200_, new_n59199_ );
or   ( new_n59202_, new_n59086_, new_n59074_ );
nand ( new_n59203_, new_n59087_, new_n59070_ );
and  ( new_n59204_, new_n59203_, new_n59202_ );
or   ( new_n59205_, new_n59204_, new_n59201_ );
and  ( new_n59206_, new_n59204_, new_n59201_ );
xor  ( new_n59207_, new_n49758_, new_n2797_ );
or   ( new_n59208_, new_n59207_, new_n3117_ );
or   ( new_n59209_, new_n58718_, new_n3119_ );
and  ( new_n59210_, new_n59209_, new_n59208_ );
xor  ( new_n59211_, new_n50487_, new_n2421_ );
or   ( new_n59212_, new_n59211_, new_n2807_ );
or   ( new_n59213_, new_n58713_, new_n2809_ );
and  ( new_n59214_, new_n59213_, new_n59212_ );
nor  ( new_n59215_, new_n59214_, new_n59210_ );
nor  ( new_n59216_, new_n58666_, new_n2124_ );
and  ( new_n59217_, new_n58741_, new_n2002_ );
nor  ( new_n59218_, new_n59217_, new_n59216_ );
and  ( new_n59219_, new_n59214_, new_n59210_ );
nor  ( new_n59220_, new_n59219_, new_n59218_ );
nor  ( new_n59221_, new_n59220_, new_n59215_ );
or   ( new_n59222_, new_n59221_, new_n59206_ );
and  ( new_n59223_, new_n59222_, new_n59205_ );
nor  ( new_n59224_, new_n59223_, new_n59198_ );
xor  ( new_n59225_, new_n59223_, new_n59198_ );
xnor ( new_n59226_, new_n59133_, new_n59130_ );
nand ( new_n59227_, new_n59226_, new_n59137_ );
not  ( new_n59228_, new_n59139_ );
or   ( new_n59229_, new_n59228_, new_n59134_ );
and  ( new_n59230_, new_n59229_, new_n59227_ );
and  ( new_n59231_, new_n59230_, new_n59225_ );
nor  ( new_n59232_, new_n59231_, new_n59224_ );
nand ( new_n59233_, new_n59232_, new_n59196_ );
and  ( new_n59234_, new_n59233_, new_n59195_ );
xnor ( new_n59235_, new_n59234_, new_n59191_ );
xor  ( new_n59236_, new_n59235_, new_n59188_ );
or   ( new_n59237_, new_n59236_, new_n59171_ );
xnor ( new_n59238_, new_n59230_, new_n59225_ );
xnor ( new_n59239_, new_n59006_, new_n59004_ );
xor  ( new_n59240_, new_n59239_, new_n59012_ );
xnor ( new_n59241_, new_n59204_, new_n59201_ );
xor  ( new_n59242_, new_n59241_, new_n59221_ );
nand ( new_n59243_, new_n59242_, new_n59240_ );
nor  ( new_n59244_, new_n59211_, new_n2809_ );
xor  ( new_n59245_, new_n50788_, new_n2421_ );
nor  ( new_n59246_, new_n59245_, new_n2807_ );
or   ( new_n59247_, new_n59246_, new_n59244_ );
xor  ( new_n59248_, new_n59084_, new_n59083_ );
and  ( new_n59249_, new_n59248_, new_n59247_ );
nor  ( new_n59250_, new_n59207_, new_n3119_ );
xor  ( new_n59251_, new_n50115_, new_n2797_ );
nor  ( new_n59252_, new_n59251_, new_n3117_ );
nor  ( new_n59253_, new_n59252_, new_n59250_ );
not  ( new_n59254_, new_n59253_ );
xor  ( new_n59255_, new_n59248_, new_n59247_ );
and  ( new_n59256_, new_n59255_, new_n59254_ );
nor  ( new_n59257_, new_n59256_, new_n59249_ );
not  ( new_n59258_, new_n59257_ );
xnor ( new_n59259_, new_n59214_, new_n59210_ );
xor  ( new_n59260_, new_n59259_, new_n59218_ );
and  ( new_n59261_, new_n59260_, new_n59258_ );
xor  ( new_n59262_, new_n59260_, new_n59258_ );
nand ( new_n59263_, new_n58838_, new_n4958_ );
xor  ( new_n59264_, new_n47640_, new_n4705_ );
or   ( new_n59265_, new_n59264_, new_n5207_ );
and  ( new_n59266_, new_n59265_, new_n59263_ );
or   ( new_n59267_, new_n58845_, new_n6175_ );
xor  ( new_n59268_, new_n46958_, new_n5594_ );
or   ( new_n59269_, new_n59268_, new_n6173_ );
and  ( new_n59270_, new_n59269_, new_n59267_ );
nor  ( new_n59271_, new_n59270_, new_n59266_ );
and  ( new_n59272_, new_n59270_, new_n59266_ );
nor  ( new_n59273_, new_n58855_, new_n5606_ );
xor  ( new_n59274_, new_n47046_, new_n5203_ );
nor  ( new_n59275_, new_n59274_, new_n5604_ );
nor  ( new_n59276_, new_n59275_, new_n59273_ );
nor  ( new_n59277_, new_n59276_, new_n59272_ );
or   ( new_n59278_, new_n59277_, new_n59271_ );
and  ( new_n59279_, new_n59278_, new_n59262_ );
nor  ( new_n59280_, new_n59279_, new_n59261_ );
nor  ( new_n59281_, new_n59242_, new_n59240_ );
or   ( new_n59282_, new_n59281_, new_n59280_ );
and  ( new_n59283_, new_n59282_, new_n59243_ );
nor  ( new_n59284_, new_n59283_, new_n59238_ );
xor  ( new_n59285_, new_n59283_, new_n59238_ );
nand ( new_n59286_, new_n58870_, new_n3291_ );
xor  ( new_n59287_, new_n49488_, RIbb2e620_35 );
nand ( new_n59288_, new_n59287_, new_n3293_ );
and  ( new_n59289_, new_n59288_, new_n59286_ );
or   ( new_n59290_, new_n59068_, new_n2427_ );
xor  ( new_n59291_, new_n51142_, new_n2118_ );
or   ( new_n59292_, new_n59291_, new_n2425_ );
and  ( new_n59293_, new_n59292_, new_n59290_ );
nor  ( new_n59294_, new_n59293_, new_n59289_ );
nor  ( new_n59295_, new_n58849_, new_n6647_ );
xor  ( new_n59296_, new_n46789_, new_n6163_ );
nor  ( new_n59297_, new_n59296_, new_n6645_ );
nor  ( new_n59298_, new_n59297_, new_n59295_ );
and  ( new_n59299_, new_n59293_, new_n59289_ );
nor  ( new_n59300_, new_n59299_, new_n59298_ );
nor  ( new_n59301_, new_n59300_, new_n59294_ );
nor  ( new_n59302_, new_n59080_, new_n1595_ );
xor  ( new_n59303_, new_n52908_, RIbb2ebc0_23 );
nor  ( new_n59304_, new_n59303_, new_n1593_ );
or   ( new_n59305_, new_n59304_, new_n59302_ );
xor  ( new_n59306_, new_n58733_, new_n58726_ );
nand ( new_n59307_, new_n59306_, new_n59305_ );
xor  ( new_n59308_, new_n51758_, new_n1840_ );
nor  ( new_n59309_, new_n59308_, new_n2122_ );
and  ( new_n59310_, new_n58743_, new_n2000_ );
or   ( new_n59311_, new_n59310_, new_n59309_ );
xor  ( new_n59312_, new_n59306_, new_n59305_ );
nand ( new_n59313_, new_n59312_, new_n59311_ );
and  ( new_n59314_, new_n59313_, new_n59307_ );
xor  ( new_n59315_, new_n48756_, RIbb2e440_39 );
nand ( new_n59316_, new_n59315_, new_n4034_ );
or   ( new_n59317_, new_n58751_, new_n4304_ );
and  ( new_n59318_, new_n59317_, new_n59316_ );
or   ( new_n59319_, new_n59318_, new_n59314_ );
and  ( new_n59320_, new_n59092_, new_n6908_ );
xor  ( new_n59321_, new_n46427_, RIbb2dea0_51 );
and  ( new_n59322_, new_n59321_, new_n6910_ );
or   ( new_n59323_, new_n59322_, new_n59320_ );
xor  ( new_n59324_, new_n59318_, new_n59314_ );
nand ( new_n59325_, new_n59324_, new_n59323_ );
and  ( new_n59326_, new_n59325_, new_n59319_ );
nor  ( new_n59327_, new_n59326_, new_n59301_ );
and  ( new_n59328_, new_n58893_, new_n9738_ );
xor  ( new_n59329_, new_n44974_, RIbb2d9f0_61 );
and  ( new_n59330_, new_n59329_, new_n9740_ );
or   ( new_n59331_, new_n59330_, new_n59328_ );
xor  ( new_n59332_, new_n58746_, new_n58745_ );
and  ( new_n59333_, new_n59332_, new_n59331_ );
and  ( new_n59334_, new_n58896_, new_n8040_ );
xor  ( new_n59335_, new_n45597_, RIbb2dcc0_55 );
and  ( new_n59336_, new_n59335_, new_n8042_ );
or   ( new_n59337_, new_n59336_, new_n59334_ );
xor  ( new_n59338_, new_n59332_, new_n59331_ );
and  ( new_n59339_, new_n59338_, new_n59337_ );
nor  ( new_n59340_, new_n59339_, new_n59333_ );
xnor ( new_n59341_, new_n59326_, new_n59301_ );
nor  ( new_n59342_, new_n59341_, new_n59340_ );
or   ( new_n59343_, new_n59342_, new_n59327_ );
xnor ( new_n59344_, new_n58860_, new_n58844_ );
xor  ( new_n59345_, new_n59344_, new_n58883_ );
or   ( new_n59346_, new_n59345_, new_n59343_ );
nand ( new_n59347_, new_n59345_, new_n59343_ );
xor  ( new_n59348_, new_n45204_, RIbb2dae0_59 );
and  ( new_n59349_, new_n59348_, new_n9187_ );
nor  ( new_n59350_, new_n59064_, new_n9424_ );
or   ( new_n59351_, new_n59350_, new_n59349_ );
and  ( new_n59352_, new_n44681_, RIbb2d888_64 );
or   ( new_n59353_, new_n59352_, RIbb2d900_63 );
nand ( new_n59354_, new_n59352_, RIbb2d900_63 );
or   ( new_n59355_, new_n44944_, RIbb2d888_64 );
and  ( new_n59356_, new_n59355_, new_n59354_ );
and  ( new_n59357_, new_n59356_, new_n59353_ );
nand ( new_n59358_, new_n59357_, new_n59351_ );
nor  ( new_n59359_, new_n59357_, new_n59351_ );
nor  ( new_n59360_, new_n58905_, new_n7734_ );
xor  ( new_n59361_, new_n46037_, new_n7174_ );
nor  ( new_n59362_, new_n59361_, new_n7732_ );
nor  ( new_n59363_, new_n59362_, new_n59360_ );
or   ( new_n59364_, new_n59363_, new_n59359_ );
and  ( new_n59365_, new_n59364_, new_n59358_ );
xor  ( new_n59366_, new_n45584_, new_n8254_ );
or   ( new_n59367_, new_n59366_, new_n8874_ );
or   ( new_n59368_, new_n58865_, new_n8876_ );
and  ( new_n59369_, new_n59368_, new_n59367_ );
nand ( new_n59370_, new_n58831_, new_n4541_ );
xor  ( new_n59371_, new_n48291_, new_n4292_ );
or   ( new_n59372_, new_n59371_, new_n4709_ );
and  ( new_n59373_, new_n59372_, new_n59370_ );
or   ( new_n59374_, new_n59373_, new_n59369_ );
xor  ( new_n59375_, new_n49265_, new_n3457_ );
nor  ( new_n59376_, new_n59375_, new_n3896_ );
nor  ( new_n59377_, new_n58757_, new_n3898_ );
nor  ( new_n59378_, new_n59377_, new_n59376_ );
and  ( new_n59379_, new_n59373_, new_n59369_ );
or   ( new_n59380_, new_n59379_, new_n59378_ );
and  ( new_n59381_, new_n59380_, new_n59374_ );
nor  ( new_n59382_, new_n59381_, new_n59365_ );
and  ( new_n59383_, new_n59381_, new_n59365_ );
xor  ( new_n59384_, new_n58842_, new_n58841_ );
not  ( new_n59385_, new_n59384_ );
nor  ( new_n59386_, new_n59385_, new_n59383_ );
nor  ( new_n59387_, new_n59386_, new_n59382_ );
nand ( new_n59388_, new_n59387_, new_n59347_ );
and  ( new_n59389_, new_n59388_, new_n59346_ );
and  ( new_n59390_, new_n59389_, new_n59285_ );
nor  ( new_n59391_, new_n59390_, new_n59284_ );
xor  ( new_n59392_, new_n59194_, new_n59192_ );
xor  ( new_n59393_, new_n59392_, new_n59232_ );
nor  ( new_n59394_, new_n59393_, new_n59391_ );
xor  ( new_n59395_, new_n59393_, new_n59391_ );
xor  ( new_n59396_, new_n58915_, new_n58914_ );
and  ( new_n59397_, new_n59396_, new_n59395_ );
or   ( new_n59398_, new_n59397_, new_n59394_ );
xor  ( new_n59399_, new_n59236_, new_n59171_ );
nand ( new_n59400_, new_n59399_, new_n59398_ );
and  ( new_n59401_, new_n59400_, new_n59237_ );
nor  ( new_n59402_, new_n59401_, new_n59114_ );
xor  ( new_n59403_, new_n59401_, new_n59114_ );
nor  ( new_n59404_, new_n59119_, new_n59117_ );
and  ( new_n59405_, new_n59170_, new_n59120_ );
nor  ( new_n59406_, new_n59405_, new_n59404_ );
xor  ( new_n59407_, new_n58435_, new_n58434_ );
xor  ( new_n59408_, new_n58333_, new_n58332_ );
or   ( new_n59409_, new_n58925_, new_n58923_ );
and  ( new_n59410_, new_n58925_, new_n58923_ );
or   ( new_n59411_, new_n59410_, new_n58922_ );
and  ( new_n59412_, new_n59411_, new_n59409_ );
xnor ( new_n59413_, new_n59412_, new_n59408_ );
xor  ( new_n59414_, new_n59413_, new_n59407_ );
xor  ( new_n59415_, new_n59414_, new_n59406_ );
or   ( new_n59416_, new_n59234_, new_n59191_ );
and  ( new_n59417_, new_n59234_, new_n59191_ );
or   ( new_n59418_, new_n59417_, new_n59188_ );
and  ( new_n59419_, new_n59418_, new_n59416_ );
xor  ( new_n59420_, new_n59419_, new_n59415_ );
xor  ( new_n59421_, new_n58627_, new_n58584_ );
xor  ( new_n59422_, new_n59421_, new_n58632_ );
or   ( new_n59423_, new_n59186_, new_n59177_ );
nand ( new_n59424_, new_n59186_, new_n59177_ );
nand ( new_n59425_, new_n59424_, new_n59176_ );
and  ( new_n59426_, new_n59425_, new_n59423_ );
xnor ( new_n59427_, new_n59426_, new_n59422_ );
or   ( new_n59428_, new_n58927_, new_n58921_ );
and  ( new_n59429_, new_n58927_, new_n58921_ );
or   ( new_n59430_, new_n59429_, new_n58920_ );
and  ( new_n59431_, new_n59430_, new_n59428_ );
xor  ( new_n59432_, new_n59431_, new_n59427_ );
or   ( new_n59433_, new_n59167_, new_n59165_ );
xor  ( new_n59434_, new_n58525_, new_n58524_ );
xnor ( new_n59435_, new_n58458_, new_n58457_ );
xor  ( new_n59436_, new_n59435_, new_n58484_ );
xor  ( new_n59437_, new_n59436_, new_n59434_ );
xor  ( new_n59438_, new_n59437_, new_n59433_ );
xor  ( new_n59439_, new_n59438_, new_n59432_ );
xor  ( new_n59440_, new_n59439_, new_n59420_ );
and  ( new_n59441_, new_n59440_, new_n59403_ );
nor  ( new_n59442_, new_n59441_, new_n59402_ );
not  ( new_n59443_, new_n59442_ );
nor  ( new_n59444_, new_n59414_, new_n59406_ );
and  ( new_n59445_, new_n59419_, new_n59415_ );
nor  ( new_n59446_, new_n59445_, new_n59444_ );
not  ( new_n59447_, new_n59446_ );
nor  ( new_n59448_, new_n59426_, new_n59422_ );
nor  ( new_n59449_, new_n59431_, new_n59427_ );
or   ( new_n59450_, new_n59449_, new_n59448_ );
nor  ( new_n59451_, new_n59412_, new_n59408_ );
and  ( new_n59452_, new_n59412_, new_n59408_ );
nor  ( new_n59453_, new_n59452_, new_n59407_ );
nor  ( new_n59454_, new_n59453_, new_n59451_ );
xnor ( new_n59455_, new_n58336_, new_n58335_ );
xnor ( new_n59456_, new_n58373_, new_n58371_ );
xor  ( new_n59457_, new_n59456_, new_n58376_ );
xor  ( new_n59458_, new_n59457_, new_n59455_ );
xor  ( new_n59459_, new_n59458_, new_n59454_ );
xor  ( new_n59460_, new_n59459_, new_n59450_ );
xor  ( new_n59461_, new_n59460_, new_n59447_ );
xor  ( new_n59462_, new_n58439_, new_n58437_ );
xor  ( new_n59463_, new_n59462_, new_n58486_ );
xnor ( new_n59464_, new_n58634_, new_n58531_ );
or   ( new_n59465_, new_n59436_, new_n59434_ );
and  ( new_n59466_, new_n59436_, new_n59434_ );
or   ( new_n59467_, new_n59466_, new_n59433_ );
and  ( new_n59468_, new_n59467_, new_n59465_ );
xor  ( new_n59469_, new_n59468_, new_n59464_ );
xnor ( new_n59470_, new_n59469_, new_n59463_ );
xnor ( new_n59471_, new_n59470_, new_n59461_ );
nand ( new_n59472_, new_n59438_, new_n59432_ );
or   ( new_n59473_, new_n59438_, new_n59432_ );
nand ( new_n59474_, new_n59473_, new_n59420_ );
and  ( new_n59475_, new_n59474_, new_n59472_ );
xor  ( new_n59476_, new_n59475_, new_n59471_ );
and  ( new_n59477_, new_n59476_, new_n59443_ );
nor  ( new_n59478_, new_n59476_, new_n59443_ );
xnor ( new_n59479_, new_n59109_, new_n59060_ );
xor  ( new_n59480_, new_n58912_, new_n58911_ );
xor  ( new_n59481_, new_n58705_, new_n58688_ );
xor  ( new_n59482_, new_n59481_, new_n58766_ );
nand ( new_n59483_, new_n59482_, new_n59480_ );
nor  ( new_n59484_, new_n59482_, new_n59480_ );
xor  ( new_n59485_, new_n58909_, new_n58890_ );
xor  ( new_n59486_, new_n58764_, new_n58763_ );
nand ( new_n59487_, new_n59486_, new_n59485_ );
nor  ( new_n59488_, new_n59486_, new_n59485_ );
xor  ( new_n59489_, new_n58761_, new_n58760_ );
xnor ( new_n59490_, new_n58852_, new_n58848_ );
xor  ( new_n59491_, new_n59490_, new_n58857_ );
nand ( new_n59492_, new_n59491_, new_n59489_ );
xor  ( new_n59493_, new_n59491_, new_n59489_ );
xnor ( new_n59494_, new_n58872_, new_n58867_ );
xor  ( new_n59495_, new_n59494_, new_n58881_ );
nand ( new_n59496_, new_n59495_, new_n59493_ );
and  ( new_n59497_, new_n59496_, new_n59492_ );
or   ( new_n59498_, new_n59497_, new_n59488_ );
and  ( new_n59499_, new_n59498_, new_n59487_ );
or   ( new_n59500_, new_n59499_, new_n59484_ );
and  ( new_n59501_, new_n59500_, new_n59483_ );
nor  ( new_n59502_, new_n59501_, new_n59479_ );
xor  ( new_n59503_, new_n59096_, new_n59095_ );
xnor ( new_n59504_, new_n58900_, new_n58895_ );
nand ( new_n59505_, new_n59504_, new_n58907_ );
not  ( new_n59506_, new_n58908_ );
or   ( new_n59507_, new_n59506_, new_n58901_ );
and  ( new_n59508_, new_n59507_, new_n59505_ );
nand ( new_n59509_, new_n59508_, new_n59503_ );
xor  ( new_n59510_, new_n59508_, new_n59503_ );
not  ( new_n59511_, new_n59510_ );
or   ( new_n59512_, new_n58735_, new_n1846_ );
xor  ( new_n59513_, new_n52293_, RIbb2ead0_25 );
or   ( new_n59514_, new_n59513_, new_n1844_ );
and  ( new_n59515_, new_n59514_, new_n59512_ );
nor  ( new_n59516_, new_n59303_, new_n1595_ );
xor  ( new_n59517_, new_n53306_, RIbb2ebc0_23 );
nor  ( new_n59518_, new_n59517_, new_n1593_ );
or   ( new_n59519_, new_n59518_, new_n59516_ );
and  ( new_n59520_, new_n53694_, new_n1251_ );
nand ( new_n59521_, new_n59520_, new_n59519_ );
nor  ( new_n59522_, new_n59513_, new_n1846_ );
xor  ( new_n59523_, new_n52902_, RIbb2ead0_25 );
nor  ( new_n59524_, new_n59523_, new_n1844_ );
or   ( new_n59525_, new_n59524_, new_n59522_ );
xor  ( new_n59526_, new_n59520_, new_n59519_ );
nand ( new_n59527_, new_n59526_, new_n59525_ );
and  ( new_n59528_, new_n59527_, new_n59521_ );
nor  ( new_n59529_, new_n59528_, new_n59515_ );
nor  ( new_n59530_, new_n59251_, new_n3119_ );
xor  ( new_n59531_, new_n50487_, new_n2797_ );
nor  ( new_n59532_, new_n59531_, new_n3117_ );
or   ( new_n59533_, new_n59532_, new_n59530_ );
xor  ( new_n59534_, new_n59528_, new_n59515_ );
and  ( new_n59535_, new_n59534_, new_n59533_ );
nor  ( new_n59536_, new_n59535_, new_n59529_ );
not  ( new_n59537_, new_n59536_ );
and  ( new_n59538_, new_n59321_, new_n6908_ );
xor  ( new_n59539_, new_n46619_, new_n6635_ );
nor  ( new_n59540_, new_n59539_, new_n7184_ );
or   ( new_n59541_, new_n59540_, new_n59538_ );
xor  ( new_n59542_, new_n59312_, new_n59311_ );
and  ( new_n59543_, new_n59542_, new_n59541_ );
nor  ( new_n59544_, new_n59264_, new_n5209_ );
xor  ( new_n59545_, new_n48039_, RIbb2e260_43 );
and  ( new_n59546_, new_n59545_, new_n4960_ );
or   ( new_n59547_, new_n59546_, new_n59544_ );
xor  ( new_n59548_, new_n59542_, new_n59541_ );
and  ( new_n59549_, new_n59548_, new_n59547_ );
nor  ( new_n59550_, new_n59549_, new_n59543_ );
not  ( new_n59551_, new_n59550_ );
and  ( new_n59552_, new_n59551_, new_n59537_ );
and  ( new_n59553_, new_n59550_, new_n59536_ );
or   ( new_n59554_, new_n59245_, new_n2809_ );
xor  ( new_n59555_, new_n50894_, new_n2421_ );
or   ( new_n59556_, new_n59555_, new_n2807_ );
and  ( new_n59557_, new_n59556_, new_n59554_ );
or   ( new_n59558_, new_n59291_, new_n2427_ );
xor  ( new_n59559_, new_n51446_, RIbb2e8f0_29 );
nand ( new_n59560_, new_n59559_, new_n2244_ );
and  ( new_n59561_, new_n59560_, new_n59558_ );
nor  ( new_n59562_, new_n59561_, new_n59557_ );
and  ( new_n59563_, new_n59287_, new_n3291_ );
xor  ( new_n59564_, new_n49758_, new_n3113_ );
nor  ( new_n59565_, new_n59564_, new_n3461_ );
or   ( new_n59566_, new_n59565_, new_n59563_ );
xor  ( new_n59567_, new_n59561_, new_n59557_ );
and  ( new_n59568_, new_n59567_, new_n59566_ );
nor  ( new_n59569_, new_n59568_, new_n59562_ );
nor  ( new_n59570_, new_n59569_, new_n59553_ );
nor  ( new_n59571_, new_n59570_, new_n59552_ );
or   ( new_n59572_, new_n59571_, new_n59511_ );
and  ( new_n59573_, new_n59572_, new_n59509_ );
xnor ( new_n59574_, new_n59098_, new_n59062_ );
xor  ( new_n59575_, new_n59574_, new_n59100_ );
nor  ( new_n59576_, new_n59575_, new_n59573_ );
and  ( new_n59577_, new_n59575_, new_n59573_ );
xor  ( new_n59578_, new_n59242_, new_n59240_ );
xor  ( new_n59579_, new_n59578_, new_n59280_ );
nor  ( new_n59580_, new_n59579_, new_n59577_ );
nor  ( new_n59581_, new_n59580_, new_n59576_ );
xor  ( new_n59582_, new_n59103_, new_n59061_ );
xor  ( new_n59583_, new_n59582_, new_n59107_ );
nor  ( new_n59584_, new_n59583_, new_n59581_ );
xor  ( new_n59585_, new_n59583_, new_n59581_ );
xor  ( new_n59586_, new_n59389_, new_n59285_ );
and  ( new_n59587_, new_n59586_, new_n59585_ );
nor  ( new_n59588_, new_n59587_, new_n59584_ );
not  ( new_n59589_, new_n59588_ );
xor  ( new_n59590_, new_n59501_, new_n59479_ );
and  ( new_n59591_, new_n59590_, new_n59589_ );
or   ( new_n59592_, new_n59591_, new_n59502_ );
xor  ( new_n59593_, new_n59112_, new_n59111_ );
and  ( new_n59594_, new_n59593_, new_n59592_ );
xor  ( new_n59595_, new_n59593_, new_n59592_ );
xor  ( new_n59596_, new_n59399_, new_n59398_ );
and  ( new_n59597_, new_n59596_, new_n59595_ );
nor  ( new_n59598_, new_n59597_, new_n59594_ );
not  ( new_n59599_, new_n59598_ );
xor  ( new_n59600_, new_n59440_, new_n59403_ );
and  ( new_n59601_, new_n59600_, new_n59599_ );
nor  ( new_n59602_, new_n59600_, new_n59599_ );
xnor ( new_n59603_, new_n59396_, new_n59395_ );
xor  ( new_n59604_, new_n59482_, new_n59480_ );
xor  ( new_n59605_, new_n59604_, new_n59499_ );
xnor ( new_n59606_, new_n59341_, new_n59340_ );
xor  ( new_n59607_, new_n47303_, new_n5594_ );
or   ( new_n59608_, new_n59607_, new_n6173_ );
or   ( new_n59609_, new_n59268_, new_n6175_ );
and  ( new_n59610_, new_n59609_, new_n59608_ );
or   ( new_n59611_, new_n59274_, new_n5606_ );
xor  ( new_n59612_, new_n47296_, RIbb2e170_45 );
nand ( new_n59613_, new_n59612_, new_n5373_ );
and  ( new_n59614_, new_n59613_, new_n59611_ );
nor  ( new_n59615_, new_n59614_, new_n59610_ );
nor  ( new_n59616_, new_n59296_, new_n6647_ );
xor  ( new_n59617_, new_n46962_, new_n6163_ );
nor  ( new_n59618_, new_n59617_, new_n6645_ );
or   ( new_n59619_, new_n59618_, new_n59616_ );
xor  ( new_n59620_, new_n59614_, new_n59610_ );
and  ( new_n59621_, new_n59620_, new_n59619_ );
or   ( new_n59622_, new_n59621_, new_n59615_ );
xnor ( new_n59623_, new_n59293_, new_n59289_ );
nand ( new_n59624_, new_n59623_, new_n59298_ );
not  ( new_n59625_, new_n59300_ );
or   ( new_n59626_, new_n59625_, new_n59294_ );
and  ( new_n59627_, new_n59626_, new_n59624_ );
nand ( new_n59628_, new_n59627_, new_n59622_ );
or   ( new_n59629_, new_n59627_, new_n59622_ );
xor  ( new_n59630_, new_n59255_, new_n59254_ );
nand ( new_n59631_, new_n59630_, new_n59629_ );
and  ( new_n59632_, new_n59631_, new_n59628_ );
nor  ( new_n59633_, new_n59632_, new_n59606_ );
and  ( new_n59634_, new_n53694_, new_n44833_ );
or   ( new_n59635_, new_n59634_, new_n1358_ );
or   ( new_n59636_, new_n59517_, new_n1595_ );
and  ( new_n59637_, new_n44831_, RIbb2ebc0_23 );
and  ( new_n59638_, new_n53694_, RIbb2ead0_25 );
nor  ( new_n59639_, new_n59638_, new_n59637_ );
and  ( new_n59640_, RIbb2eb48_24, new_n1355_ );
nor  ( new_n59641_, new_n53694_, RIbb2ead0_25 );
nor  ( new_n59642_, new_n59641_, new_n59640_ );
or   ( new_n59643_, new_n59642_, new_n59639_ );
and  ( new_n59644_, new_n59643_, new_n59636_ );
or   ( new_n59645_, new_n59644_, new_n59635_ );
or   ( new_n59646_, new_n59308_, new_n2124_ );
xor  ( new_n59647_, new_n52280_, new_n1840_ );
or   ( new_n59648_, new_n59647_, new_n2122_ );
and  ( new_n59649_, new_n59648_, new_n59646_ );
or   ( new_n59650_, new_n59649_, new_n59645_ );
and  ( new_n59651_, new_n59559_, new_n2242_ );
xor  ( new_n59652_, new_n51477_, RIbb2e8f0_29 );
and  ( new_n59653_, new_n59652_, new_n2244_ );
or   ( new_n59654_, new_n59653_, new_n59651_ );
xor  ( new_n59655_, new_n59649_, new_n59645_ );
nand ( new_n59656_, new_n59655_, new_n59654_ );
and  ( new_n59657_, new_n59656_, new_n59650_ );
or   ( new_n59658_, new_n59371_, new_n4711_ );
xor  ( new_n59659_, new_n48518_, new_n4292_ );
or   ( new_n59660_, new_n59659_, new_n4709_ );
and  ( new_n59661_, new_n59660_, new_n59658_ );
nor  ( new_n59662_, new_n59661_, new_n59657_ );
xor  ( new_n59663_, new_n48908_, new_n3892_ );
nor  ( new_n59664_, new_n59663_, new_n4302_ );
and  ( new_n59665_, new_n59315_, new_n4032_ );
nor  ( new_n59666_, new_n59665_, new_n59664_ );
xnor ( new_n59667_, new_n59661_, new_n59657_ );
nor  ( new_n59668_, new_n59667_, new_n59666_ );
or   ( new_n59669_, new_n59668_, new_n59662_ );
xor  ( new_n59670_, new_n59324_, new_n59323_ );
and  ( new_n59671_, new_n59670_, new_n59669_ );
nor  ( new_n59672_, new_n59361_, new_n7734_ );
xor  ( new_n59673_, new_n46137_, RIbb2ddb0_53 );
and  ( new_n59674_, new_n59673_, new_n7489_ );
nor  ( new_n59675_, new_n59674_, new_n59672_ );
xor  ( new_n59676_, new_n45928_, new_n7722_ );
or   ( new_n59677_, new_n59676_, new_n8264_ );
nand ( new_n59678_, new_n59335_, new_n8040_ );
and  ( new_n59679_, new_n59678_, new_n59677_ );
nor  ( new_n59680_, new_n59679_, new_n59675_ );
xnor ( new_n59681_, new_n59679_, new_n59675_ );
and  ( new_n59682_, new_n44785_, RIbb2d888_64 );
and  ( new_n59683_, new_n44877_, new_n21077_ );
or   ( new_n59684_, new_n59683_, new_n10052_ );
or   ( new_n59685_, new_n59684_, new_n59682_ );
nand ( new_n59686_, new_n59682_, new_n10052_ );
and  ( new_n59687_, new_n59686_, new_n59685_ );
nor  ( new_n59688_, new_n59687_, new_n59681_ );
nor  ( new_n59689_, new_n59688_, new_n59680_ );
not  ( new_n59690_, new_n59689_ );
xor  ( new_n59691_, new_n59670_, new_n59669_ );
and  ( new_n59692_, new_n59691_, new_n59690_ );
nor  ( new_n59693_, new_n59692_, new_n59671_ );
not  ( new_n59694_, new_n59693_ );
xor  ( new_n59695_, new_n59632_, new_n59606_ );
and  ( new_n59696_, new_n59695_, new_n59694_ );
nor  ( new_n59697_, new_n59696_, new_n59633_ );
not  ( new_n59698_, new_n59697_ );
xor  ( new_n59699_, new_n59345_, new_n59343_ );
xor  ( new_n59700_, new_n59699_, new_n59387_ );
not  ( new_n59701_, new_n59700_ );
and  ( new_n59702_, new_n59701_, new_n59698_ );
and  ( new_n59703_, new_n59700_, new_n59697_ );
xnor ( new_n59704_, new_n59278_, new_n59262_ );
xnor ( new_n59705_, new_n59270_, new_n59266_ );
nand ( new_n59706_, new_n59705_, new_n59276_ );
not  ( new_n59707_, new_n59277_ );
or   ( new_n59708_, new_n59707_, new_n59271_ );
and  ( new_n59709_, new_n59708_, new_n59706_ );
xnor ( new_n59710_, new_n59373_, new_n59369_ );
xor  ( new_n59711_, new_n59710_, new_n59378_ );
nand ( new_n59712_, new_n59711_, new_n59709_ );
nor  ( new_n59713_, new_n59711_, new_n59709_ );
or   ( new_n59714_, new_n59375_, new_n3898_ );
xor  ( new_n59715_, new_n49427_, RIbb2e530_37 );
nand ( new_n59716_, new_n59715_, new_n3733_ );
and  ( new_n59717_, new_n59716_, new_n59714_ );
or   ( new_n59718_, new_n59366_, new_n8876_ );
xor  ( new_n59719_, new_n45738_, RIbb2dbd0_57 );
nand ( new_n59720_, new_n59719_, new_n8651_ );
and  ( new_n59721_, new_n59720_, new_n59718_ );
or   ( new_n59722_, new_n59721_, new_n59717_ );
xor  ( new_n59723_, new_n45119_, new_n9418_ );
nor  ( new_n59724_, new_n59723_, new_n10059_ );
and  ( new_n59725_, new_n59329_, new_n9738_ );
or   ( new_n59726_, new_n59725_, new_n59724_ );
xor  ( new_n59727_, new_n59721_, new_n59717_ );
nand ( new_n59728_, new_n59727_, new_n59726_ );
and  ( new_n59729_, new_n59728_, new_n59722_ );
or   ( new_n59730_, new_n59729_, new_n59713_ );
and  ( new_n59731_, new_n59730_, new_n59712_ );
nor  ( new_n59732_, new_n59731_, new_n59704_ );
xor  ( new_n59733_, new_n59731_, new_n59704_ );
xor  ( new_n59734_, new_n59338_, new_n59337_ );
xnor ( new_n59735_, new_n59357_, new_n59351_ );
xor  ( new_n59736_, new_n59735_, new_n59363_ );
or   ( new_n59737_, new_n59736_, new_n59734_ );
nand ( new_n59738_, new_n59736_, new_n59734_ );
xor  ( new_n59739_, new_n45403_, new_n8870_ );
nor  ( new_n59740_, new_n59739_, new_n9422_ );
and  ( new_n59741_, new_n59348_, new_n9185_ );
or   ( new_n59742_, new_n59741_, new_n59740_ );
xor  ( new_n59743_, new_n59534_, new_n59533_ );
and  ( new_n59744_, new_n59743_, new_n59742_ );
xor  ( new_n59745_, new_n50788_, new_n2797_ );
nor  ( new_n59746_, new_n59745_, new_n3117_ );
nor  ( new_n59747_, new_n59531_, new_n3119_ );
or   ( new_n59748_, new_n59747_, new_n59746_ );
xor  ( new_n59749_, new_n59526_, new_n59525_ );
and  ( new_n59750_, new_n59749_, new_n59748_ );
and  ( new_n59751_, new_n59715_, new_n3731_ );
xor  ( new_n59752_, new_n49488_, RIbb2e530_37 );
and  ( new_n59753_, new_n59752_, new_n3733_ );
or   ( new_n59754_, new_n59753_, new_n59751_ );
xor  ( new_n59755_, new_n59749_, new_n59748_ );
and  ( new_n59756_, new_n59755_, new_n59754_ );
nor  ( new_n59757_, new_n59756_, new_n59750_ );
xnor ( new_n59758_, new_n59743_, new_n59742_ );
nor  ( new_n59759_, new_n59758_, new_n59757_ );
nor  ( new_n59760_, new_n59759_, new_n59744_ );
nand ( new_n59761_, new_n59760_, new_n59738_ );
and  ( new_n59762_, new_n59761_, new_n59737_ );
and  ( new_n59763_, new_n59762_, new_n59733_ );
nor  ( new_n59764_, new_n59763_, new_n59732_ );
nor  ( new_n59765_, new_n59764_, new_n59703_ );
nor  ( new_n59766_, new_n59765_, new_n59702_ );
or   ( new_n59767_, new_n59766_, new_n59605_ );
and  ( new_n59768_, new_n59766_, new_n59605_ );
xnor ( new_n59769_, new_n59495_, new_n59493_ );
xor  ( new_n59770_, new_n59381_, new_n59365_ );
xor  ( new_n59771_, new_n59770_, new_n59385_ );
or   ( new_n59772_, new_n59771_, new_n59769_ );
xor  ( new_n59773_, new_n59571_, new_n59511_ );
xor  ( new_n59774_, new_n59771_, new_n59769_ );
nand ( new_n59775_, new_n59774_, new_n59773_ );
and  ( new_n59776_, new_n59775_, new_n59772_ );
xor  ( new_n59777_, new_n59486_, new_n59485_ );
xor  ( new_n59778_, new_n59777_, new_n59497_ );
nor  ( new_n59779_, new_n59778_, new_n59776_ );
and  ( new_n59780_, new_n59778_, new_n59776_ );
xor  ( new_n59781_, new_n59575_, new_n59573_ );
xnor ( new_n59782_, new_n59781_, new_n59579_ );
not  ( new_n59783_, new_n59782_ );
nor  ( new_n59784_, new_n59783_, new_n59780_ );
nor  ( new_n59785_, new_n59784_, new_n59779_ );
or   ( new_n59786_, new_n59785_, new_n59768_ );
and  ( new_n59787_, new_n59786_, new_n59767_ );
nor  ( new_n59788_, new_n59787_, new_n59603_ );
xor  ( new_n59789_, new_n59590_, new_n59589_ );
xor  ( new_n59790_, new_n59787_, new_n59603_ );
and  ( new_n59791_, new_n59790_, new_n59789_ );
nor  ( new_n59792_, new_n59791_, new_n59788_ );
not  ( new_n59793_, new_n59792_ );
xor  ( new_n59794_, new_n59596_, new_n59595_ );
and  ( new_n59795_, new_n59794_, new_n59793_ );
nor  ( new_n59796_, new_n59794_, new_n59793_ );
xor  ( new_n59797_, new_n59790_, new_n59789_ );
not  ( new_n59798_, new_n59797_ );
xnor ( new_n59799_, new_n59586_, new_n59585_ );
xor  ( new_n59800_, new_n59695_, new_n59694_ );
xor  ( new_n59801_, new_n51142_, new_n2421_ );
or   ( new_n59802_, new_n59801_, new_n2807_ );
or   ( new_n59803_, new_n59555_, new_n2809_ );
and  ( new_n59804_, new_n59803_, new_n59802_ );
or   ( new_n59805_, new_n59564_, new_n3463_ );
xor  ( new_n59806_, new_n50115_, new_n3113_ );
or   ( new_n59807_, new_n59806_, new_n3461_ );
and  ( new_n59808_, new_n59807_, new_n59805_ );
nor  ( new_n59809_, new_n59808_, new_n59804_ );
nor  ( new_n59810_, new_n59617_, new_n6647_ );
xor  ( new_n59811_, new_n46958_, RIbb2df90_49 );
and  ( new_n59812_, new_n59811_, new_n6510_ );
nor  ( new_n59813_, new_n59812_, new_n59810_ );
and  ( new_n59814_, new_n59808_, new_n59804_ );
nor  ( new_n59815_, new_n59814_, new_n59813_ );
or   ( new_n59816_, new_n59815_, new_n59809_ );
xor  ( new_n59817_, new_n59567_, new_n59566_ );
and  ( new_n59818_, new_n59817_, new_n59816_ );
nor  ( new_n59819_, new_n59523_, new_n1846_ );
xor  ( new_n59820_, new_n52908_, RIbb2ead0_25 );
nor  ( new_n59821_, new_n59820_, new_n1844_ );
or   ( new_n59822_, new_n59821_, new_n59819_ );
xor  ( new_n59823_, new_n59644_, new_n59635_ );
nand ( new_n59824_, new_n59823_, new_n59822_ );
nor  ( new_n59825_, new_n59647_, new_n2124_ );
xor  ( new_n59826_, new_n52293_, RIbb2e9e0_27 );
nor  ( new_n59827_, new_n59826_, new_n2122_ );
or   ( new_n59828_, new_n59827_, new_n59825_ );
xor  ( new_n59829_, new_n59823_, new_n59822_ );
nand ( new_n59830_, new_n59829_, new_n59828_ );
and  ( new_n59831_, new_n59830_, new_n59824_ );
xor  ( new_n59832_, new_n48756_, RIbb2e350_41 );
nand ( new_n59833_, new_n59832_, new_n4543_ );
or   ( new_n59834_, new_n59659_, new_n4711_ );
and  ( new_n59835_, new_n59834_, new_n59833_ );
nor  ( new_n59836_, new_n59835_, new_n59831_ );
nor  ( new_n59837_, new_n59663_, new_n4304_ );
xor  ( new_n59838_, new_n49265_, new_n3892_ );
nor  ( new_n59839_, new_n59838_, new_n4302_ );
or   ( new_n59840_, new_n59839_, new_n59837_ );
xor  ( new_n59841_, new_n59835_, new_n59831_ );
and  ( new_n59842_, new_n59841_, new_n59840_ );
nor  ( new_n59843_, new_n59842_, new_n59836_ );
xnor ( new_n59844_, new_n59817_, new_n59816_ );
nor  ( new_n59845_, new_n59844_, new_n59843_ );
or   ( new_n59846_, new_n59845_, new_n59818_ );
xor  ( new_n59847_, new_n59550_, new_n59537_ );
nand ( new_n59848_, new_n59847_, new_n59569_ );
or   ( new_n59849_, new_n59569_, new_n59553_ );
or   ( new_n59850_, new_n59849_, new_n59552_ );
and  ( new_n59851_, new_n59850_, new_n59848_ );
or   ( new_n59852_, new_n59851_, new_n59846_ );
and  ( new_n59853_, new_n59851_, new_n59846_ );
xor  ( new_n59854_, new_n59627_, new_n59622_ );
xor  ( new_n59855_, new_n59854_, new_n59630_ );
or   ( new_n59856_, new_n59855_, new_n59853_ );
and  ( new_n59857_, new_n59856_, new_n59852_ );
and  ( new_n59858_, new_n59857_, new_n59800_ );
xor  ( new_n59859_, new_n59857_, new_n59800_ );
xor  ( new_n59860_, new_n59762_, new_n59733_ );
and  ( new_n59861_, new_n59860_, new_n59859_ );
or   ( new_n59862_, new_n59861_, new_n59858_ );
xor  ( new_n59863_, new_n59700_, new_n59698_ );
nand ( new_n59864_, new_n59863_, new_n59764_ );
or   ( new_n59865_, new_n59764_, new_n59703_ );
or   ( new_n59866_, new_n59865_, new_n59702_ );
and  ( new_n59867_, new_n59866_, new_n59864_ );
nand ( new_n59868_, new_n59867_, new_n59862_ );
nor  ( new_n59869_, new_n59867_, new_n59862_ );
xor  ( new_n59870_, new_n48291_, RIbb2e260_43 );
nand ( new_n59871_, new_n59870_, new_n4960_ );
nand ( new_n59872_, new_n59545_, new_n4958_ );
and  ( new_n59873_, new_n59872_, new_n59871_ );
xor  ( new_n59874_, new_n47046_, new_n5594_ );
or   ( new_n59875_, new_n59874_, new_n6173_ );
or   ( new_n59876_, new_n59607_, new_n6175_ );
and  ( new_n59877_, new_n59876_, new_n59875_ );
nor  ( new_n59878_, new_n59877_, new_n59873_ );
xor  ( new_n59879_, new_n47640_, new_n5203_ );
nor  ( new_n59880_, new_n59879_, new_n5604_ );
and  ( new_n59881_, new_n59612_, new_n5371_ );
nor  ( new_n59882_, new_n59881_, new_n59880_ );
and  ( new_n59883_, new_n59877_, new_n59873_ );
nor  ( new_n59884_, new_n59883_, new_n59882_ );
nor  ( new_n59885_, new_n59884_, new_n59878_ );
not  ( new_n59886_, new_n59885_ );
xor  ( new_n59887_, new_n59548_, new_n59547_ );
nand ( new_n59888_, new_n59887_, new_n59886_ );
xor  ( new_n59889_, new_n59887_, new_n59886_ );
xor  ( new_n59890_, new_n59620_, new_n59619_ );
nand ( new_n59891_, new_n59890_, new_n59889_ );
and  ( new_n59892_, new_n59891_, new_n59888_ );
xnor ( new_n59893_, new_n59667_, new_n59666_ );
or   ( new_n59894_, new_n59539_, new_n7186_ );
xor  ( new_n59895_, new_n46789_, new_n6635_ );
or   ( new_n59896_, new_n59895_, new_n7184_ );
and  ( new_n59897_, new_n59896_, new_n59894_ );
nand ( new_n59898_, new_n59673_, new_n7487_ );
xor  ( new_n59899_, new_n46427_, RIbb2ddb0_53 );
nand ( new_n59900_, new_n59899_, new_n7489_ );
and  ( new_n59901_, new_n59900_, new_n59898_ );
nor  ( new_n59902_, new_n59901_, new_n59897_ );
xor  ( new_n59903_, new_n45597_, RIbb2dbd0_57 );
and  ( new_n59904_, new_n59903_, new_n8651_ );
and  ( new_n59905_, new_n59719_, new_n8649_ );
nor  ( new_n59906_, new_n59905_, new_n59904_ );
and  ( new_n59907_, new_n59901_, new_n59897_ );
nor  ( new_n59908_, new_n59907_, new_n59906_ );
nor  ( new_n59909_, new_n59908_, new_n59902_ );
or   ( new_n59910_, new_n59909_, new_n59893_ );
xor  ( new_n59911_, new_n46037_, new_n7722_ );
nor  ( new_n59912_, new_n59911_, new_n8264_ );
nor  ( new_n59913_, new_n59676_, new_n8266_ );
or   ( new_n59914_, new_n59913_, new_n59912_ );
xor  ( new_n59915_, new_n59655_, new_n59654_ );
and  ( new_n59916_, new_n59915_, new_n59914_ );
xor  ( new_n59917_, new_n45204_, RIbb2d9f0_61 );
and  ( new_n59918_, new_n59917_, new_n9740_ );
nor  ( new_n59919_, new_n59723_, new_n10061_ );
or   ( new_n59920_, new_n59919_, new_n59918_ );
xor  ( new_n59921_, new_n59915_, new_n59914_ );
and  ( new_n59922_, new_n59921_, new_n59920_ );
nor  ( new_n59923_, new_n59922_, new_n59916_ );
not  ( new_n59924_, new_n59923_ );
xor  ( new_n59925_, new_n59909_, new_n59893_ );
nand ( new_n59926_, new_n59925_, new_n59924_ );
and  ( new_n59927_, new_n59926_, new_n59910_ );
or   ( new_n59928_, new_n59927_, new_n59892_ );
xor  ( new_n59929_, new_n59727_, new_n59726_ );
xor  ( new_n59930_, new_n59687_, new_n59681_ );
and  ( new_n59931_, new_n59930_, new_n59929_ );
nor  ( new_n59932_, new_n59820_, new_n1846_ );
xor  ( new_n59933_, new_n53306_, RIbb2ead0_25 );
nor  ( new_n59934_, new_n59933_, new_n1844_ );
or   ( new_n59935_, new_n59934_, new_n59932_ );
and  ( new_n59936_, new_n53694_, new_n1474_ );
nand ( new_n59937_, new_n59936_, new_n59935_ );
xor  ( new_n59938_, new_n52902_, RIbb2e9e0_27 );
nor  ( new_n59939_, new_n59938_, new_n2122_ );
nor  ( new_n59940_, new_n59826_, new_n2124_ );
or   ( new_n59941_, new_n59940_, new_n59939_ );
xor  ( new_n59942_, new_n59936_, new_n59935_ );
nand ( new_n59943_, new_n59942_, new_n59941_ );
and  ( new_n59944_, new_n59943_, new_n59937_ );
xor  ( new_n59945_, new_n51758_, new_n2118_ );
or   ( new_n59946_, new_n59945_, new_n2425_ );
nand ( new_n59947_, new_n59652_, new_n2242_ );
and  ( new_n59948_, new_n59947_, new_n59946_ );
or   ( new_n59949_, new_n59948_, new_n59944_ );
xor  ( new_n59950_, new_n49758_, new_n3457_ );
nor  ( new_n59951_, new_n59950_, new_n3896_ );
and  ( new_n59952_, new_n59752_, new_n3731_ );
or   ( new_n59953_, new_n59952_, new_n59951_ );
xor  ( new_n59954_, new_n59948_, new_n59944_ );
nand ( new_n59955_, new_n59954_, new_n59953_ );
and  ( new_n59956_, new_n59955_, new_n59949_ );
and  ( new_n59957_, new_n44877_, RIbb2d888_64 );
and  ( new_n59958_, new_n44974_, new_n21077_ );
or   ( new_n59959_, new_n59958_, new_n10052_ );
or   ( new_n59960_, new_n59959_, new_n59957_ );
nand ( new_n59961_, new_n59957_, new_n10052_ );
and  ( new_n59962_, new_n59961_, new_n59960_ );
nor  ( new_n59963_, new_n59962_, new_n59956_ );
xor  ( new_n59964_, new_n45584_, RIbb2dae0_59 );
and  ( new_n59965_, new_n59964_, new_n9187_ );
nor  ( new_n59966_, new_n59739_, new_n9424_ );
or   ( new_n59967_, new_n59966_, new_n59965_ );
xor  ( new_n59968_, new_n59962_, new_n59956_ );
and  ( new_n59969_, new_n59968_, new_n59967_ );
or   ( new_n59970_, new_n59969_, new_n59963_ );
xor  ( new_n59971_, new_n59930_, new_n59929_ );
and  ( new_n59972_, new_n59971_, new_n59970_ );
or   ( new_n59973_, new_n59972_, new_n59931_ );
xor  ( new_n59974_, new_n59927_, new_n59892_ );
nand ( new_n59975_, new_n59974_, new_n59973_ );
and  ( new_n59976_, new_n59975_, new_n59928_ );
xor  ( new_n59977_, new_n59691_, new_n59690_ );
not  ( new_n59978_, new_n59977_ );
xor  ( new_n59979_, new_n59711_, new_n59709_ );
xor  ( new_n59980_, new_n59979_, new_n59729_ );
or   ( new_n59981_, new_n59980_, new_n59978_ );
xor  ( new_n59982_, new_n59980_, new_n59978_ );
not  ( new_n59983_, new_n59982_ );
xnor ( new_n59984_, new_n59758_, new_n59757_ );
or   ( new_n59985_, new_n59801_, new_n2809_ );
xor  ( new_n59986_, new_n51446_, RIbb2e800_31 );
nand ( new_n59987_, new_n59986_, new_n2615_ );
and  ( new_n59988_, new_n59987_, new_n59985_ );
xor  ( new_n59989_, new_n50894_, new_n2797_ );
or   ( new_n59990_, new_n59989_, new_n3117_ );
or   ( new_n59991_, new_n59745_, new_n3119_ );
and  ( new_n59992_, new_n59991_, new_n59990_ );
nor  ( new_n59993_, new_n59992_, new_n59988_ );
xor  ( new_n59994_, new_n50487_, new_n3113_ );
nor  ( new_n59995_, new_n59994_, new_n3461_ );
nor  ( new_n59996_, new_n59806_, new_n3463_ );
or   ( new_n59997_, new_n59996_, new_n59995_ );
xor  ( new_n59998_, new_n59992_, new_n59988_ );
and  ( new_n59999_, new_n59998_, new_n59997_ );
or   ( new_n60000_, new_n59999_, new_n59993_ );
xnor ( new_n60001_, new_n59808_, new_n59804_ );
nand ( new_n60002_, new_n60001_, new_n59813_ );
not  ( new_n60003_, new_n59809_ );
nand ( new_n60004_, new_n59815_, new_n60003_ );
and  ( new_n60005_, new_n60004_, new_n60002_ );
nand ( new_n60006_, new_n60005_, new_n60000_ );
nor  ( new_n60007_, new_n60005_, new_n60000_ );
xor  ( new_n60008_, new_n47296_, RIbb2e080_47 );
and  ( new_n60009_, new_n60008_, new_n5917_ );
nor  ( new_n60010_, new_n59874_, new_n6175_ );
or   ( new_n60011_, new_n60010_, new_n60009_ );
xor  ( new_n60012_, new_n59829_, new_n59828_ );
and  ( new_n60013_, new_n60012_, new_n60011_ );
xor  ( new_n60014_, new_n47303_, new_n6163_ );
nor  ( new_n60015_, new_n60014_, new_n6645_ );
and  ( new_n60016_, new_n59811_, new_n6508_ );
nor  ( new_n60017_, new_n60016_, new_n60015_ );
xnor ( new_n60018_, new_n60012_, new_n60011_ );
nor  ( new_n60019_, new_n60018_, new_n60017_ );
nor  ( new_n60020_, new_n60019_, new_n60013_ );
or   ( new_n60021_, new_n60020_, new_n60007_ );
and  ( new_n60022_, new_n60021_, new_n60006_ );
or   ( new_n60023_, new_n60022_, new_n59984_ );
and  ( new_n60024_, new_n60022_, new_n59984_ );
xor  ( new_n60025_, new_n48518_, RIbb2e260_43 );
and  ( new_n60026_, new_n60025_, new_n4960_ );
and  ( new_n60027_, new_n59870_, new_n4958_ );
nor  ( new_n60028_, new_n60027_, new_n60026_ );
xor  ( new_n60029_, new_n48039_, new_n5203_ );
or   ( new_n60030_, new_n60029_, new_n5604_ );
or   ( new_n60031_, new_n59879_, new_n5606_ );
and  ( new_n60032_, new_n60031_, new_n60030_ );
nor  ( new_n60033_, new_n60032_, new_n60028_ );
xor  ( new_n60034_, new_n48908_, new_n4292_ );
nor  ( new_n60035_, new_n60034_, new_n4709_ );
and  ( new_n60036_, new_n59832_, new_n4541_ );
nor  ( new_n60037_, new_n60036_, new_n60035_ );
and  ( new_n60038_, new_n60032_, new_n60028_ );
nor  ( new_n60039_, new_n60038_, new_n60037_ );
or   ( new_n60040_, new_n60039_, new_n60033_ );
xor  ( new_n60041_, new_n59755_, new_n59754_ );
and  ( new_n60042_, new_n60041_, new_n60040_ );
nor  ( new_n60043_, new_n60041_, new_n60040_ );
and  ( new_n60044_, new_n53694_, new_n45123_ );
or   ( new_n60045_, new_n60044_, new_n1586_ );
or   ( new_n60046_, new_n59933_, new_n1846_ );
or   ( new_n60047_, new_n59638_, new_n1844_ );
or   ( new_n60048_, new_n60047_, new_n59641_ );
and  ( new_n60049_, new_n60048_, new_n60046_ );
or   ( new_n60050_, new_n60049_, new_n60045_ );
or   ( new_n60051_, new_n59945_, new_n2427_ );
xor  ( new_n60052_, new_n52280_, new_n2118_ );
or   ( new_n60053_, new_n60052_, new_n2425_ );
and  ( new_n60054_, new_n60053_, new_n60051_ );
or   ( new_n60055_, new_n60054_, new_n60050_ );
and  ( new_n60056_, new_n59986_, new_n2613_ );
xor  ( new_n60057_, new_n51477_, RIbb2e800_31 );
and  ( new_n60058_, new_n60057_, new_n2615_ );
nor  ( new_n60059_, new_n60058_, new_n60056_ );
xnor ( new_n60060_, new_n60054_, new_n60050_ );
or   ( new_n60061_, new_n60060_, new_n60059_ );
and  ( new_n60062_, new_n60061_, new_n60055_ );
or   ( new_n60063_, new_n59838_, new_n4304_ );
xor  ( new_n60064_, new_n49427_, RIbb2e440_39 );
nand ( new_n60065_, new_n60064_, new_n4034_ );
and  ( new_n60066_, new_n60065_, new_n60063_ );
nor  ( new_n60067_, new_n60066_, new_n60062_ );
xor  ( new_n60068_, new_n46619_, new_n7174_ );
nor  ( new_n60069_, new_n60068_, new_n7732_ );
and  ( new_n60070_, new_n59899_, new_n7487_ );
nor  ( new_n60071_, new_n60070_, new_n60069_ );
not  ( new_n60072_, new_n60071_ );
xor  ( new_n60073_, new_n60066_, new_n60062_ );
and  ( new_n60074_, new_n60073_, new_n60072_ );
nor  ( new_n60075_, new_n60074_, new_n60067_ );
nor  ( new_n60076_, new_n60075_, new_n60043_ );
nor  ( new_n60077_, new_n60076_, new_n60042_ );
or   ( new_n60078_, new_n60077_, new_n60024_ );
and  ( new_n60079_, new_n60078_, new_n60023_ );
or   ( new_n60080_, new_n60079_, new_n59983_ );
and  ( new_n60081_, new_n60080_, new_n59981_ );
nor  ( new_n60082_, new_n60081_, new_n59976_ );
and  ( new_n60083_, new_n60081_, new_n59976_ );
xor  ( new_n60084_, new_n59774_, new_n59773_ );
not  ( new_n60085_, new_n60084_ );
nor  ( new_n60086_, new_n60085_, new_n60083_ );
nor  ( new_n60087_, new_n60086_, new_n60082_ );
or   ( new_n60088_, new_n60087_, new_n59869_ );
and  ( new_n60089_, new_n60088_, new_n59868_ );
or   ( new_n60090_, new_n60089_, new_n59799_ );
and  ( new_n60091_, new_n60089_, new_n59799_ );
xor  ( new_n60092_, new_n59766_, new_n59605_ );
xnor ( new_n60093_, new_n60092_, new_n59785_ );
not  ( new_n60094_, new_n60093_ );
or   ( new_n60095_, new_n60094_, new_n60091_ );
and  ( new_n60096_, new_n60095_, new_n60090_ );
nor  ( new_n60097_, new_n60096_, new_n59798_ );
and  ( new_n60098_, new_n60096_, new_n59798_ );
xor  ( new_n60099_, new_n60073_, new_n60072_ );
xnor ( new_n60100_, new_n60018_, new_n60017_ );
xor  ( new_n60101_, new_n46137_, RIbb2dcc0_55 );
nand ( new_n60102_, new_n60101_, new_n8040_ );
xor  ( new_n60103_, new_n46427_, RIbb2dcc0_55 );
nand ( new_n60104_, new_n60103_, new_n8042_ );
and  ( new_n60105_, new_n60104_, new_n60102_ );
xor  ( new_n60106_, new_n46958_, new_n6635_ );
or   ( new_n60107_, new_n60106_, new_n7184_ );
xor  ( new_n60108_, new_n46962_, new_n6635_ );
or   ( new_n60109_, new_n60108_, new_n7186_ );
and  ( new_n60110_, new_n60109_, new_n60107_ );
or   ( new_n60111_, new_n60110_, new_n60105_ );
xor  ( new_n60112_, new_n46037_, new_n8254_ );
nor  ( new_n60113_, new_n60112_, new_n8874_ );
xor  ( new_n60114_, new_n45928_, new_n8254_ );
nor  ( new_n60115_, new_n60114_, new_n8876_ );
or   ( new_n60116_, new_n60115_, new_n60113_ );
xor  ( new_n60117_, new_n60110_, new_n60105_ );
nand ( new_n60118_, new_n60117_, new_n60116_ );
and  ( new_n60119_, new_n60118_, new_n60111_ );
xor  ( new_n60120_, new_n60119_, new_n60100_ );
xor  ( new_n60121_, new_n60120_, new_n60099_ );
xor  ( new_n60122_, new_n49265_, new_n4292_ );
or   ( new_n60123_, new_n60122_, new_n4711_ );
xor  ( new_n60124_, new_n49427_, RIbb2e350_41 );
nand ( new_n60125_, new_n60124_, new_n4543_ );
and  ( new_n60126_, new_n60125_, new_n60123_ );
or   ( new_n60127_, new_n60106_, new_n7186_ );
xor  ( new_n60128_, new_n47303_, new_n6635_ );
or   ( new_n60129_, new_n60128_, new_n7184_ );
and  ( new_n60130_, new_n60129_, new_n60127_ );
or   ( new_n60131_, new_n60130_, new_n60126_ );
xor  ( new_n60132_, new_n46789_, new_n7174_ );
nor  ( new_n60133_, new_n60132_, new_n7734_ );
xor  ( new_n60134_, new_n46962_, new_n7174_ );
nor  ( new_n60135_, new_n60134_, new_n7732_ );
nor  ( new_n60136_, new_n60135_, new_n60133_ );
xnor ( new_n60137_, new_n60130_, new_n60126_ );
or   ( new_n60138_, new_n60137_, new_n60136_ );
and  ( new_n60139_, new_n60138_, new_n60131_ );
xor  ( new_n60140_, new_n48039_, RIbb2e080_47 );
and  ( new_n60141_, new_n60140_, new_n5917_ );
xor  ( new_n60142_, new_n47640_, new_n5594_ );
nor  ( new_n60143_, new_n60142_, new_n6175_ );
or   ( new_n60144_, new_n60143_, new_n60141_ );
nor  ( new_n60145_, new_n60052_, new_n2427_ );
xor  ( new_n60146_, new_n52293_, RIbb2e8f0_29 );
nor  ( new_n60147_, new_n60146_, new_n2425_ );
or   ( new_n60148_, new_n60147_, new_n60145_ );
nor  ( new_n60149_, new_n59938_, new_n2124_ );
xor  ( new_n60150_, new_n52908_, RIbb2e9e0_27 );
nor  ( new_n60151_, new_n60150_, new_n2122_ );
or   ( new_n60152_, new_n60151_, new_n60149_ );
xor  ( new_n60153_, new_n60049_, new_n60045_ );
xor  ( new_n60154_, new_n60153_, new_n60152_ );
xor  ( new_n60155_, new_n60154_, new_n60148_ );
nand ( new_n60156_, new_n60155_, new_n60144_ );
xor  ( new_n60157_, new_n47046_, new_n6163_ );
nor  ( new_n60158_, new_n60157_, new_n6647_ );
xor  ( new_n60159_, new_n47296_, RIbb2df90_49 );
and  ( new_n60160_, new_n60159_, new_n6510_ );
or   ( new_n60161_, new_n60160_, new_n60158_ );
xor  ( new_n60162_, new_n60155_, new_n60144_ );
nand ( new_n60163_, new_n60162_, new_n60161_ );
and  ( new_n60164_, new_n60163_, new_n60156_ );
or   ( new_n60165_, new_n60164_, new_n60139_ );
xor  ( new_n60166_, new_n60117_, new_n60116_ );
xor  ( new_n60167_, new_n60164_, new_n60139_ );
nand ( new_n60168_, new_n60167_, new_n60166_ );
and  ( new_n60169_, new_n60168_, new_n60165_ );
xnor ( new_n60170_, new_n60060_, new_n60059_ );
xor  ( new_n60171_, new_n45119_, new_n10052_ );
or   ( new_n60172_, new_n60171_, new_n21077_ );
not  ( new_n60173_, new_n57100_ );
or   ( new_n60174_, new_n60173_, new_n45204_ );
and  ( new_n60175_, new_n60174_, new_n60172_ );
or   ( new_n60176_, new_n60175_, new_n60170_ );
xor  ( new_n60177_, new_n45584_, RIbb2d9f0_61 );
and  ( new_n60178_, new_n60177_, new_n9740_ );
xor  ( new_n60179_, new_n45403_, new_n9418_ );
nor  ( new_n60180_, new_n60179_, new_n10061_ );
or   ( new_n60181_, new_n60180_, new_n60178_ );
xor  ( new_n60182_, new_n60175_, new_n60170_ );
nand ( new_n60183_, new_n60182_, new_n60181_ );
and  ( new_n60184_, new_n60183_, new_n60176_ );
xnor ( new_n60185_, new_n60032_, new_n60028_ );
and  ( new_n60186_, new_n60185_, new_n60037_ );
or   ( new_n60187_, new_n60038_, new_n60037_ );
nor  ( new_n60188_, new_n60187_, new_n60033_ );
or   ( new_n60189_, new_n60188_, new_n60186_ );
xor  ( new_n60190_, new_n45597_, RIbb2dae0_59 );
nand ( new_n60191_, new_n60190_, new_n9187_ );
xor  ( new_n60192_, new_n45738_, RIbb2dae0_59 );
nand ( new_n60193_, new_n60192_, new_n9185_ );
and  ( new_n60194_, new_n60193_, new_n60191_ );
xor  ( new_n60195_, new_n51142_, new_n2797_ );
or   ( new_n60196_, new_n60195_, new_n3119_ );
xor  ( new_n60197_, new_n51446_, RIbb2e710_33 );
nand ( new_n60198_, new_n60197_, new_n2930_ );
and  ( new_n60199_, new_n60198_, new_n60196_ );
xor  ( new_n60200_, new_n50115_, new_n3457_ );
or   ( new_n60201_, new_n60200_, new_n3898_ );
xor  ( new_n60202_, new_n50487_, new_n3457_ );
or   ( new_n60203_, new_n60202_, new_n3896_ );
and  ( new_n60204_, new_n60203_, new_n60201_ );
or   ( new_n60205_, new_n60204_, new_n60199_ );
xor  ( new_n60206_, new_n50894_, new_n3113_ );
nor  ( new_n60207_, new_n60206_, new_n3461_ );
xor  ( new_n60208_, new_n50788_, new_n3113_ );
nor  ( new_n60209_, new_n60208_, new_n3463_ );
or   ( new_n60210_, new_n60209_, new_n60207_ );
xor  ( new_n60211_, new_n60204_, new_n60199_ );
nand ( new_n60212_, new_n60211_, new_n60210_ );
and  ( new_n60213_, new_n60212_, new_n60205_ );
or   ( new_n60214_, new_n60213_, new_n60194_ );
xor  ( new_n60215_, new_n51758_, new_n2421_ );
or   ( new_n60216_, new_n60215_, new_n2807_ );
nand ( new_n60217_, new_n60057_, new_n2613_ );
and  ( new_n60218_, new_n60217_, new_n60216_ );
nor  ( new_n60219_, new_n60150_, new_n2124_ );
xor  ( new_n60220_, new_n53306_, RIbb2e9e0_27 );
nor  ( new_n60221_, new_n60220_, new_n2122_ );
or   ( new_n60222_, new_n60221_, new_n60219_ );
and  ( new_n60223_, new_n53694_, new_n1739_ );
nand ( new_n60224_, new_n60223_, new_n60222_ );
xor  ( new_n60225_, new_n52902_, RIbb2e8f0_29 );
nor  ( new_n60226_, new_n60225_, new_n2425_ );
nor  ( new_n60227_, new_n60146_, new_n2427_ );
or   ( new_n60228_, new_n60227_, new_n60226_ );
xor  ( new_n60229_, new_n60223_, new_n60222_ );
nand ( new_n60230_, new_n60229_, new_n60228_ );
and  ( new_n60231_, new_n60230_, new_n60224_ );
nor  ( new_n60232_, new_n60231_, new_n60218_ );
xor  ( new_n60233_, new_n49488_, RIbb2e440_39 );
and  ( new_n60234_, new_n60233_, new_n4032_ );
xor  ( new_n60235_, new_n49758_, new_n3892_ );
nor  ( new_n60236_, new_n60235_, new_n4302_ );
or   ( new_n60237_, new_n60236_, new_n60234_ );
xor  ( new_n60238_, new_n60231_, new_n60218_ );
and  ( new_n60239_, new_n60238_, new_n60237_ );
nor  ( new_n60240_, new_n60239_, new_n60232_ );
and  ( new_n60241_, new_n60213_, new_n60194_ );
or   ( new_n60242_, new_n60241_, new_n60240_ );
and  ( new_n60243_, new_n60242_, new_n60214_ );
xor  ( new_n60244_, new_n60243_, new_n60189_ );
xor  ( new_n60245_, new_n60244_, new_n60184_ );
xor  ( new_n60246_, new_n60245_, new_n60169_ );
xor  ( new_n60247_, new_n60246_, new_n60121_ );
not  ( new_n60248_, new_n60247_ );
and  ( new_n60249_, new_n53694_, new_n45443_ );
or   ( new_n60250_, new_n60249_, new_n1843_ );
or   ( new_n60251_, new_n60220_, new_n2124_ );
and  ( new_n60252_, new_n45441_, RIbb2e9e0_27 );
and  ( new_n60253_, new_n53694_, RIbb2e8f0_29 );
nor  ( new_n60254_, new_n60253_, new_n60252_ );
and  ( new_n60255_, RIbb2e968_28, new_n1840_ );
nor  ( new_n60256_, new_n53694_, RIbb2e8f0_29 );
nor  ( new_n60257_, new_n60256_, new_n60255_ );
or   ( new_n60258_, new_n60257_, new_n60254_ );
and  ( new_n60259_, new_n60258_, new_n60251_ );
or   ( new_n60260_, new_n60259_, new_n60250_ );
or   ( new_n60261_, new_n60215_, new_n2809_ );
xor  ( new_n60262_, new_n52280_, new_n2421_ );
or   ( new_n60263_, new_n60262_, new_n2807_ );
and  ( new_n60264_, new_n60263_, new_n60261_ );
or   ( new_n60265_, new_n60264_, new_n60260_ );
and  ( new_n60266_, new_n60197_, new_n2928_ );
xor  ( new_n60267_, new_n51477_, RIbb2e710_33 );
and  ( new_n60268_, new_n60267_, new_n2930_ );
nor  ( new_n60269_, new_n60268_, new_n60266_ );
xnor ( new_n60270_, new_n60264_, new_n60260_ );
or   ( new_n60271_, new_n60270_, new_n60269_ );
and  ( new_n60272_, new_n60271_, new_n60265_ );
xor  ( new_n60273_, new_n48756_, RIbb2e260_43 );
nand ( new_n60274_, new_n60273_, new_n4958_ );
xor  ( new_n60275_, new_n48908_, new_n4705_ );
or   ( new_n60276_, new_n60275_, new_n5207_ );
and  ( new_n60277_, new_n60276_, new_n60274_ );
nor  ( new_n60278_, new_n60277_, new_n60272_ );
xor  ( new_n60279_, new_n48518_, RIbb2e170_45 );
and  ( new_n60280_, new_n60279_, new_n5373_ );
xor  ( new_n60281_, new_n48291_, RIbb2e170_45 );
and  ( new_n60282_, new_n60281_, new_n5371_ );
or   ( new_n60283_, new_n60282_, new_n60280_ );
xor  ( new_n60284_, new_n60277_, new_n60272_ );
and  ( new_n60285_, new_n60284_, new_n60283_ );
nor  ( new_n60286_, new_n60285_, new_n60278_ );
not  ( new_n60287_, new_n60286_ );
nor  ( new_n60288_, new_n60157_, new_n6645_ );
nor  ( new_n60289_, new_n60014_, new_n6647_ );
or   ( new_n60290_, new_n60289_, new_n60288_ );
or   ( new_n60291_, new_n60208_, new_n3461_ );
or   ( new_n60292_, new_n59994_, new_n3463_ );
and  ( new_n60293_, new_n60292_, new_n60291_ );
or   ( new_n60294_, new_n60200_, new_n3896_ );
or   ( new_n60295_, new_n59950_, new_n3898_ );
and  ( new_n60296_, new_n60295_, new_n60294_ );
xor  ( new_n60297_, new_n60296_, new_n60293_ );
xor  ( new_n60298_, new_n60297_, new_n60290_ );
and  ( new_n60299_, new_n60064_, new_n4032_ );
and  ( new_n60300_, new_n60233_, new_n4034_ );
or   ( new_n60301_, new_n60300_, new_n60299_ );
nor  ( new_n60302_, new_n59989_, new_n3119_ );
nor  ( new_n60303_, new_n60195_, new_n3117_ );
or   ( new_n60304_, new_n60303_, new_n60302_ );
xor  ( new_n60305_, new_n59942_, new_n59941_ );
xor  ( new_n60306_, new_n60305_, new_n60304_ );
xor  ( new_n60307_, new_n60306_, new_n60301_ );
xor  ( new_n60308_, new_n60307_, new_n60298_ );
xor  ( new_n60309_, new_n60308_, new_n60287_ );
xor  ( new_n60310_, new_n60167_, new_n60166_ );
nand ( new_n60311_, new_n60310_, new_n60309_ );
xor  ( new_n60312_, new_n60310_, new_n60309_ );
xor  ( new_n60313_, new_n60284_, new_n60283_ );
and  ( new_n60314_, new_n60103_, new_n8040_ );
xor  ( new_n60315_, new_n46619_, new_n7722_ );
nor  ( new_n60316_, new_n60315_, new_n8264_ );
nor  ( new_n60317_, new_n60316_, new_n60314_ );
or   ( new_n60318_, new_n60112_, new_n8876_ );
xor  ( new_n60319_, new_n46137_, new_n8254_ );
or   ( new_n60320_, new_n60319_, new_n8874_ );
and  ( new_n60321_, new_n60320_, new_n60318_ );
and  ( new_n60322_, new_n45722_, new_n10052_ );
and  ( new_n60323_, new_n45204_, RIbb2d900_63 );
or   ( new_n60324_, new_n60323_, new_n21077_ );
or   ( new_n60325_, new_n60324_, new_n60322_ );
or   ( new_n60326_, new_n45403_, new_n10052_ );
or   ( new_n60327_, new_n60326_, RIbb2d888_64 );
and  ( new_n60328_, new_n60327_, new_n60325_ );
xnor ( new_n60329_, new_n60328_, new_n60321_ );
xor  ( new_n60330_, new_n60329_, new_n60317_ );
or   ( new_n60331_, new_n60330_, new_n60313_ );
and  ( new_n60332_, new_n60330_, new_n60313_ );
and  ( new_n60333_, new_n60190_, new_n9185_ );
xor  ( new_n60334_, new_n45928_, new_n8870_ );
nor  ( new_n60335_, new_n60334_, new_n9422_ );
nor  ( new_n60336_, new_n60335_, new_n60333_ );
not  ( new_n60337_, new_n60336_ );
xor  ( new_n60338_, new_n45738_, RIbb2d9f0_61 );
and  ( new_n60339_, new_n60338_, new_n9740_ );
and  ( new_n60340_, new_n60177_, new_n9738_ );
or   ( new_n60341_, new_n60340_, new_n60339_ );
xor  ( new_n60342_, new_n60238_, new_n60237_ );
xor  ( new_n60343_, new_n60342_, new_n60341_ );
xor  ( new_n60344_, new_n60343_, new_n60337_ );
or   ( new_n60345_, new_n60344_, new_n60332_ );
and  ( new_n60346_, new_n60345_, new_n60331_ );
nand ( new_n60347_, new_n60346_, new_n60312_ );
and  ( new_n60348_, new_n60347_, new_n60311_ );
nor  ( new_n60349_, new_n60132_, new_n7732_ );
nor  ( new_n60350_, new_n60068_, new_n7734_ );
nor  ( new_n60351_, new_n60350_, new_n60349_ );
not  ( new_n60352_, new_n60351_ );
nand ( new_n60353_, new_n60153_, new_n60152_ );
nand ( new_n60354_, new_n60154_, new_n60148_ );
and  ( new_n60355_, new_n60354_, new_n60353_ );
or   ( new_n60356_, new_n60122_, new_n4709_ );
or   ( new_n60357_, new_n60034_, new_n4711_ );
and  ( new_n60358_, new_n60357_, new_n60356_ );
xor  ( new_n60359_, new_n60358_, new_n60355_ );
xor  ( new_n60360_, new_n60359_, new_n60352_ );
and  ( new_n60361_, new_n60273_, new_n4960_ );
and  ( new_n60362_, new_n60025_, new_n4958_ );
or   ( new_n60363_, new_n60362_, new_n60361_ );
nand ( new_n60364_, new_n60281_, new_n5373_ );
or   ( new_n60365_, new_n60029_, new_n5606_ );
and  ( new_n60366_, new_n60365_, new_n60364_ );
nand ( new_n60367_, new_n60008_, new_n5915_ );
or   ( new_n60368_, new_n60142_, new_n6173_ );
and  ( new_n60369_, new_n60368_, new_n60367_ );
xor  ( new_n60370_, new_n60369_, new_n60366_ );
xor  ( new_n60371_, new_n60370_, new_n60363_ );
and  ( new_n60372_, new_n60371_, new_n60360_ );
xor  ( new_n60373_, new_n60371_, new_n60360_ );
not  ( new_n60374_, new_n60373_ );
or   ( new_n60375_, new_n60328_, new_n60321_ );
and  ( new_n60376_, new_n60328_, new_n60321_ );
or   ( new_n60377_, new_n60376_, new_n60317_ );
and  ( new_n60378_, new_n60377_, new_n60375_ );
nor  ( new_n60379_, new_n60378_, new_n60374_ );
nor  ( new_n60380_, new_n60379_, new_n60372_ );
and  ( new_n60381_, new_n60305_, new_n60304_ );
and  ( new_n60382_, new_n60306_, new_n60301_ );
or   ( new_n60383_, new_n60382_, new_n60381_ );
xor  ( new_n60384_, new_n59954_, new_n59953_ );
xor  ( new_n60385_, new_n59998_, new_n59997_ );
xor  ( new_n60386_, new_n60385_, new_n60384_ );
xor  ( new_n60387_, new_n60386_, new_n60383_ );
nor  ( new_n60388_, new_n60369_, new_n60366_ );
and  ( new_n60389_, new_n60370_, new_n60363_ );
or   ( new_n60390_, new_n60389_, new_n60388_ );
or   ( new_n60391_, new_n60296_, new_n60293_ );
nand ( new_n60392_, new_n60297_, new_n60290_ );
and  ( new_n60393_, new_n60392_, new_n60391_ );
or   ( new_n60394_, new_n60358_, new_n60355_ );
nand ( new_n60395_, new_n60359_, new_n60352_ );
and  ( new_n60396_, new_n60395_, new_n60394_ );
xor  ( new_n60397_, new_n60396_, new_n60393_ );
xor  ( new_n60398_, new_n60397_, new_n60390_ );
xor  ( new_n60399_, new_n60398_, new_n60387_ );
xor  ( new_n60400_, new_n60399_, new_n60380_ );
xor  ( new_n60401_, new_n60400_, new_n60348_ );
xor  ( new_n60402_, new_n60401_, new_n60248_ );
xor  ( new_n60403_, new_n60378_, new_n60374_ );
nand ( new_n60404_, new_n60342_, new_n60341_ );
nand ( new_n60405_, new_n60343_, new_n60337_ );
and  ( new_n60406_, new_n60405_, new_n60404_ );
xor  ( new_n60407_, new_n50788_, new_n3457_ );
or   ( new_n60408_, new_n60407_, new_n3896_ );
or   ( new_n60409_, new_n60202_, new_n3898_ );
and  ( new_n60410_, new_n60409_, new_n60408_ );
xor  ( new_n60411_, new_n51142_, new_n3113_ );
or   ( new_n60412_, new_n60411_, new_n3461_ );
or   ( new_n60413_, new_n60206_, new_n3463_ );
and  ( new_n60414_, new_n60413_, new_n60412_ );
nor  ( new_n60415_, new_n60414_, new_n60410_ );
nor  ( new_n60416_, new_n60315_, new_n8266_ );
xor  ( new_n60417_, new_n46789_, new_n7722_ );
nor  ( new_n60418_, new_n60417_, new_n8264_ );
or   ( new_n60419_, new_n60418_, new_n60416_ );
nand ( new_n60420_, new_n60414_, new_n60410_ );
and  ( new_n60421_, new_n60420_, new_n60419_ );
or   ( new_n60422_, new_n60421_, new_n60415_ );
xor  ( new_n60423_, new_n60211_, new_n60210_ );
nand ( new_n60424_, new_n60423_, new_n60422_ );
nor  ( new_n60425_, new_n60423_, new_n60422_ );
xor  ( new_n60426_, new_n50115_, new_n3892_ );
nor  ( new_n60427_, new_n60426_, new_n4302_ );
nor  ( new_n60428_, new_n60235_, new_n4304_ );
or   ( new_n60429_, new_n60428_, new_n60427_ );
xor  ( new_n60430_, new_n60229_, new_n60228_ );
and  ( new_n60431_, new_n60430_, new_n60429_ );
and  ( new_n60432_, new_n60124_, new_n4541_ );
xor  ( new_n60433_, new_n49488_, RIbb2e350_41 );
and  ( new_n60434_, new_n60433_, new_n4543_ );
nor  ( new_n60435_, new_n60434_, new_n60432_ );
xnor ( new_n60436_, new_n60430_, new_n60429_ );
nor  ( new_n60437_, new_n60436_, new_n60435_ );
nor  ( new_n60438_, new_n60437_, new_n60431_ );
or   ( new_n60439_, new_n60438_, new_n60425_ );
and  ( new_n60440_, new_n60439_, new_n60424_ );
xor  ( new_n60441_, new_n60440_, new_n60406_ );
xor  ( new_n60442_, new_n60182_, new_n60181_ );
xor  ( new_n60443_, new_n60442_, new_n60441_ );
xor  ( new_n60444_, new_n60443_, new_n60403_ );
xnor ( new_n60445_, new_n60436_, new_n60435_ );
and  ( new_n60446_, new_n53694_, new_n45578_ );
or   ( new_n60447_, new_n60446_, new_n2121_ );
xor  ( new_n60448_, new_n53306_, RIbb2e8f0_29 );
or   ( new_n60449_, new_n60448_, new_n2427_ );
or   ( new_n60450_, new_n60253_, new_n2425_ );
or   ( new_n60451_, new_n60450_, new_n60256_ );
and  ( new_n60452_, new_n60451_, new_n60449_ );
or   ( new_n60453_, new_n60452_, new_n60447_ );
xor  ( new_n60454_, new_n52280_, new_n2797_ );
or   ( new_n60455_, new_n60454_, new_n3117_ );
xor  ( new_n60456_, new_n51758_, new_n2797_ );
or   ( new_n60457_, new_n60456_, new_n3119_ );
and  ( new_n60458_, new_n60457_, new_n60455_ );
or   ( new_n60459_, new_n60458_, new_n60453_ );
xor  ( new_n60460_, new_n51446_, RIbb2e620_35 );
and  ( new_n60461_, new_n60460_, new_n3291_ );
xor  ( new_n60462_, new_n51477_, RIbb2e620_35 );
and  ( new_n60463_, new_n60462_, new_n3293_ );
nor  ( new_n60464_, new_n60463_, new_n60461_ );
xnor ( new_n60465_, new_n60458_, new_n60453_ );
or   ( new_n60466_, new_n60465_, new_n60464_ );
and  ( new_n60467_, new_n60466_, new_n60459_ );
xor  ( new_n60468_, new_n46427_, new_n8254_ );
or   ( new_n60469_, new_n60468_, new_n8876_ );
xor  ( new_n60470_, new_n46619_, new_n8254_ );
or   ( new_n60471_, new_n60470_, new_n8874_ );
and  ( new_n60472_, new_n60471_, new_n60469_ );
nor  ( new_n60473_, new_n60472_, new_n60467_ );
and  ( new_n60474_, new_n60472_, new_n60467_ );
xor  ( new_n60475_, new_n46958_, RIbb2ddb0_53 );
and  ( new_n60476_, new_n60475_, new_n7487_ );
xor  ( new_n60477_, new_n47303_, new_n7174_ );
nor  ( new_n60478_, new_n60477_, new_n7732_ );
nor  ( new_n60479_, new_n60478_, new_n60476_ );
nor  ( new_n60480_, new_n60479_, new_n60474_ );
nor  ( new_n60481_, new_n60480_, new_n60473_ );
or   ( new_n60482_, new_n60481_, new_n60445_ );
xor  ( new_n60483_, new_n49265_, new_n4705_ );
or   ( new_n60484_, new_n60483_, new_n5209_ );
xor  ( new_n60485_, new_n49427_, RIbb2e260_43 );
nand ( new_n60486_, new_n60485_, new_n4960_ );
and  ( new_n60487_, new_n60486_, new_n60484_ );
xor  ( new_n60488_, new_n48291_, new_n5594_ );
or   ( new_n60489_, new_n60488_, new_n6175_ );
xor  ( new_n60490_, new_n48518_, RIbb2e080_47 );
nand ( new_n60491_, new_n60490_, new_n5917_ );
and  ( new_n60492_, new_n60491_, new_n60489_ );
or   ( new_n60493_, new_n60492_, new_n60487_ );
xor  ( new_n60494_, new_n48756_, RIbb2e170_45 );
and  ( new_n60495_, new_n60494_, new_n5371_ );
xor  ( new_n60496_, new_n48908_, new_n5203_ );
nor  ( new_n60497_, new_n60496_, new_n5604_ );
or   ( new_n60498_, new_n60497_, new_n60495_ );
xor  ( new_n60499_, new_n60492_, new_n60487_ );
nand ( new_n60500_, new_n60499_, new_n60498_ );
and  ( new_n60501_, new_n60500_, new_n60493_ );
and  ( new_n60502_, new_n60481_, new_n60445_ );
or   ( new_n60503_, new_n60502_, new_n60501_ );
and  ( new_n60504_, new_n60503_, new_n60482_ );
xor  ( new_n60505_, new_n60414_, new_n60410_ );
xor  ( new_n60506_, new_n60505_, new_n60419_ );
and  ( new_n60507_, new_n60338_, new_n9738_ );
xor  ( new_n60508_, new_n45597_, RIbb2d9f0_61 );
and  ( new_n60509_, new_n60508_, new_n9740_ );
or   ( new_n60510_, new_n60509_, new_n60507_ );
nand ( new_n60511_, new_n60475_, new_n7489_ );
or   ( new_n60512_, new_n60134_, new_n7734_ );
and  ( new_n60513_, new_n60512_, new_n60511_ );
or   ( new_n60514_, new_n60128_, new_n7186_ );
xor  ( new_n60515_, new_n47046_, new_n6635_ );
or   ( new_n60516_, new_n60515_, new_n7184_ );
and  ( new_n60517_, new_n60516_, new_n60514_ );
xor  ( new_n60518_, new_n60517_, new_n60513_ );
xor  ( new_n60519_, new_n60518_, new_n60510_ );
nand ( new_n60520_, new_n60519_, new_n60506_ );
or   ( new_n60521_, new_n60519_, new_n60506_ );
and  ( new_n60522_, new_n60159_, new_n6508_ );
xor  ( new_n60523_, new_n47640_, new_n6163_ );
nor  ( new_n60524_, new_n60523_, new_n6645_ );
nor  ( new_n60525_, new_n60524_, new_n60522_ );
nand ( new_n60526_, new_n60140_, new_n5915_ );
or   ( new_n60527_, new_n60488_, new_n6173_ );
and  ( new_n60528_, new_n60527_, new_n60526_ );
nand ( new_n60529_, new_n60494_, new_n5373_ );
nand ( new_n60530_, new_n60279_, new_n5371_ );
and  ( new_n60531_, new_n60530_, new_n60529_ );
xor  ( new_n60532_, new_n60531_, new_n60528_ );
xnor ( new_n60533_, new_n60532_, new_n60525_ );
nand ( new_n60534_, new_n60533_, new_n60521_ );
and  ( new_n60535_, new_n60534_, new_n60520_ );
or   ( new_n60536_, new_n60535_, new_n60504_ );
and  ( new_n60537_, new_n60535_, new_n60504_ );
or   ( new_n60538_, new_n60262_, new_n2809_ );
xor  ( new_n60539_, new_n52293_, RIbb2e800_31 );
or   ( new_n60540_, new_n60539_, new_n2807_ );
and  ( new_n60541_, new_n60540_, new_n60538_ );
xor  ( new_n60542_, new_n52908_, RIbb2e8f0_29 );
nor  ( new_n60543_, new_n60542_, new_n2427_ );
nor  ( new_n60544_, new_n60448_, new_n2425_ );
or   ( new_n60545_, new_n60544_, new_n60543_ );
and  ( new_n60546_, new_n53694_, new_n2000_ );
nand ( new_n60547_, new_n60546_, new_n60545_ );
xor  ( new_n60548_, new_n52902_, RIbb2e800_31 );
nor  ( new_n60549_, new_n60548_, new_n2807_ );
nor  ( new_n60550_, new_n60539_, new_n2809_ );
or   ( new_n60551_, new_n60550_, new_n60549_ );
xor  ( new_n60552_, new_n60546_, new_n60545_ );
nand ( new_n60553_, new_n60552_, new_n60551_ );
and  ( new_n60554_, new_n60553_, new_n60547_ );
or   ( new_n60555_, new_n60554_, new_n60541_ );
and  ( new_n60556_, new_n60433_, new_n4541_ );
xor  ( new_n60557_, new_n49758_, new_n4292_ );
nor  ( new_n60558_, new_n60557_, new_n4709_ );
or   ( new_n60559_, new_n60558_, new_n60556_ );
xor  ( new_n60560_, new_n60554_, new_n60541_ );
nand ( new_n60561_, new_n60560_, new_n60559_ );
and  ( new_n60562_, new_n60561_, new_n60555_ );
or   ( new_n60563_, new_n60411_, new_n3463_ );
nand ( new_n60564_, new_n60460_, new_n3293_ );
and  ( new_n60565_, new_n60564_, new_n60563_ );
xor  ( new_n60566_, new_n50487_, new_n3892_ );
or   ( new_n60567_, new_n60566_, new_n4302_ );
or   ( new_n60568_, new_n60426_, new_n4304_ );
and  ( new_n60569_, new_n60568_, new_n60567_ );
or   ( new_n60570_, new_n60569_, new_n60565_ );
xor  ( new_n60571_, new_n50894_, new_n3457_ );
nor  ( new_n60572_, new_n60571_, new_n3896_ );
nor  ( new_n60573_, new_n60407_, new_n3898_ );
or   ( new_n60574_, new_n60573_, new_n60572_ );
xor  ( new_n60575_, new_n60569_, new_n60565_ );
nand ( new_n60576_, new_n60575_, new_n60574_ );
and  ( new_n60577_, new_n60576_, new_n60570_ );
nor  ( new_n60578_, new_n60577_, new_n60562_ );
xor  ( new_n60579_, new_n46962_, new_n7722_ );
nor  ( new_n60580_, new_n60579_, new_n8264_ );
nor  ( new_n60581_, new_n60417_, new_n8266_ );
or   ( new_n60582_, new_n60581_, new_n60580_ );
and  ( new_n60583_, new_n60267_, new_n2928_ );
nor  ( new_n60584_, new_n60456_, new_n3117_ );
or   ( new_n60585_, new_n60584_, new_n60583_ );
nor  ( new_n60586_, new_n60225_, new_n2427_ );
nor  ( new_n60587_, new_n60542_, new_n2425_ );
or   ( new_n60588_, new_n60587_, new_n60586_ );
xor  ( new_n60589_, new_n60259_, new_n60250_ );
xor  ( new_n60590_, new_n60589_, new_n60588_ );
xor  ( new_n60591_, new_n60590_, new_n60585_ );
and  ( new_n60592_, new_n60591_, new_n60582_ );
xor  ( new_n60593_, new_n48039_, RIbb2df90_49 );
and  ( new_n60594_, new_n60593_, new_n6510_ );
nor  ( new_n60595_, new_n60523_, new_n6647_ );
or   ( new_n60596_, new_n60595_, new_n60594_ );
xor  ( new_n60597_, new_n60591_, new_n60582_ );
and  ( new_n60598_, new_n60597_, new_n60596_ );
nor  ( new_n60599_, new_n60598_, new_n60592_ );
xnor ( new_n60600_, new_n60577_, new_n60562_ );
nor  ( new_n60601_, new_n60600_, new_n60599_ );
nor  ( new_n60602_, new_n60601_, new_n60578_ );
or   ( new_n60603_, new_n60602_, new_n60537_ );
nand ( new_n60604_, new_n60603_, new_n60536_ );
xnor ( new_n60605_, new_n60604_, new_n60444_ );
nor  ( new_n60606_, new_n60483_, new_n5207_ );
nor  ( new_n60607_, new_n60275_, new_n5209_ );
nor  ( new_n60608_, new_n60607_, new_n60606_ );
nand ( new_n60609_, new_n60589_, new_n60588_ );
nand ( new_n60610_, new_n60590_, new_n60585_ );
and  ( new_n60611_, new_n60610_, new_n60609_ );
or   ( new_n60612_, new_n60319_, new_n8876_ );
or   ( new_n60613_, new_n60468_, new_n8874_ );
and  ( new_n60614_, new_n60613_, new_n60612_ );
xor  ( new_n60615_, new_n60614_, new_n60611_ );
xor  ( new_n60616_, new_n60615_, new_n60608_ );
or   ( new_n60617_, new_n60515_, new_n7186_ );
xor  ( new_n60618_, new_n47296_, new_n6635_ );
or   ( new_n60619_, new_n60618_, new_n7184_ );
and  ( new_n60620_, new_n60619_, new_n60617_ );
or   ( new_n60621_, new_n45738_, new_n10052_ );
and  ( new_n60622_, new_n60621_, new_n10770_ );
and  ( new_n60623_, new_n45584_, RIbb2d888_64 );
or   ( new_n60624_, new_n60623_, new_n60622_ );
nand ( new_n60625_, new_n60623_, new_n10052_ );
and  ( new_n60626_, new_n60625_, new_n60624_ );
or   ( new_n60627_, new_n60626_, new_n60620_ );
and  ( new_n60628_, new_n60626_, new_n60620_ );
and  ( new_n60629_, new_n60508_, new_n9738_ );
xor  ( new_n60630_, new_n45928_, new_n9418_ );
nor  ( new_n60631_, new_n60630_, new_n10059_ );
nor  ( new_n60632_, new_n60631_, new_n60629_ );
or   ( new_n60633_, new_n60632_, new_n60628_ );
and  ( new_n60634_, new_n60633_, new_n60627_ );
or   ( new_n60635_, new_n60634_, new_n60616_ );
and  ( new_n60636_, new_n60634_, new_n60616_ );
xor  ( new_n60637_, new_n46037_, new_n8870_ );
nor  ( new_n60638_, new_n60637_, new_n9424_ );
xor  ( new_n60639_, new_n46137_, RIbb2dae0_59 );
and  ( new_n60640_, new_n60639_, new_n9187_ );
or   ( new_n60641_, new_n60640_, new_n60638_ );
xor  ( new_n60642_, new_n60560_, new_n60559_ );
and  ( new_n60643_, new_n60642_, new_n60641_ );
nor  ( new_n60644_, new_n60642_, new_n60641_ );
nor  ( new_n60645_, new_n60566_, new_n4304_ );
xor  ( new_n60646_, new_n50788_, new_n3892_ );
nor  ( new_n60647_, new_n60646_, new_n4302_ );
or   ( new_n60648_, new_n60647_, new_n60645_ );
xor  ( new_n60649_, new_n60552_, new_n60551_ );
and  ( new_n60650_, new_n60649_, new_n60648_ );
and  ( new_n60651_, new_n60485_, new_n4958_ );
xor  ( new_n60652_, new_n49488_, RIbb2e260_43 );
and  ( new_n60653_, new_n60652_, new_n4960_ );
or   ( new_n60654_, new_n60653_, new_n60651_ );
xor  ( new_n60655_, new_n60649_, new_n60648_ );
and  ( new_n60656_, new_n60655_, new_n60654_ );
nor  ( new_n60657_, new_n60656_, new_n60650_ );
nor  ( new_n60658_, new_n60657_, new_n60644_ );
nor  ( new_n60659_, new_n60658_, new_n60643_ );
or   ( new_n60660_, new_n60659_, new_n60636_ );
and  ( new_n60661_, new_n60660_, new_n60635_ );
xnor ( new_n60662_, new_n60330_, new_n60313_ );
xor  ( new_n60663_, new_n60662_, new_n60344_ );
or   ( new_n60664_, new_n60663_, new_n60661_ );
and  ( new_n60665_, new_n60663_, new_n60661_ );
xnor ( new_n60666_, new_n60600_, new_n60599_ );
nor  ( new_n60667_, new_n60637_, new_n9422_ );
nor  ( new_n60668_, new_n60334_, new_n9424_ );
nor  ( new_n60669_, new_n60668_, new_n60667_ );
xnor ( new_n60670_, new_n60270_, new_n60269_ );
or   ( new_n60671_, new_n60173_, new_n45584_ );
xor  ( new_n60672_, new_n45403_, new_n10052_ );
or   ( new_n60673_, new_n60672_, new_n21077_ );
and  ( new_n60674_, new_n60673_, new_n60671_ );
xor  ( new_n60675_, new_n60674_, new_n60670_ );
xor  ( new_n60676_, new_n60675_, new_n60669_ );
nor  ( new_n60677_, new_n60676_, new_n60666_ );
and  ( new_n60678_, new_n60676_, new_n60666_ );
or   ( new_n60679_, new_n60557_, new_n4711_ );
xor  ( new_n60680_, new_n50115_, new_n4292_ );
or   ( new_n60681_, new_n60680_, new_n4709_ );
and  ( new_n60682_, new_n60681_, new_n60679_ );
or   ( new_n60683_, new_n60571_, new_n3898_ );
xor  ( new_n60684_, new_n51142_, new_n3457_ );
or   ( new_n60685_, new_n60684_, new_n3896_ );
and  ( new_n60686_, new_n60685_, new_n60683_ );
nor  ( new_n60687_, new_n60686_, new_n60682_ );
xor  ( new_n60688_, new_n48291_, RIbb2df90_49 );
and  ( new_n60689_, new_n60688_, new_n6510_ );
and  ( new_n60690_, new_n60593_, new_n6508_ );
or   ( new_n60691_, new_n60690_, new_n60689_ );
xor  ( new_n60692_, new_n60686_, new_n60682_ );
and  ( new_n60693_, new_n60692_, new_n60691_ );
nor  ( new_n60694_, new_n60693_, new_n60687_ );
not  ( new_n60695_, new_n60694_ );
xor  ( new_n60696_, new_n46789_, new_n8254_ );
or   ( new_n60697_, new_n60696_, new_n8874_ );
or   ( new_n60698_, new_n60470_, new_n8876_ );
and  ( new_n60699_, new_n60698_, new_n60697_ );
nand ( new_n60700_, new_n60639_, new_n9185_ );
xor  ( new_n60701_, new_n46427_, new_n8870_ );
or   ( new_n60702_, new_n60701_, new_n9422_ );
and  ( new_n60703_, new_n60702_, new_n60700_ );
nor  ( new_n60704_, new_n60703_, new_n60699_ );
and  ( new_n60705_, new_n60490_, new_n5915_ );
xor  ( new_n60706_, new_n48756_, RIbb2e080_47 );
and  ( new_n60707_, new_n60706_, new_n5917_ );
or   ( new_n60708_, new_n60707_, new_n60705_ );
xor  ( new_n60709_, new_n60703_, new_n60699_ );
and  ( new_n60710_, new_n60709_, new_n60708_ );
nor  ( new_n60711_, new_n60710_, new_n60704_ );
not  ( new_n60712_, new_n60711_ );
and  ( new_n60713_, new_n60712_, new_n60695_ );
nor  ( new_n60714_, new_n60548_, new_n2809_ );
xor  ( new_n60715_, new_n52908_, RIbb2e800_31 );
nor  ( new_n60716_, new_n60715_, new_n2807_ );
or   ( new_n60717_, new_n60716_, new_n60714_ );
xor  ( new_n60718_, new_n60452_, new_n60447_ );
nand ( new_n60719_, new_n60718_, new_n60717_ );
and  ( new_n60720_, new_n60462_, new_n3291_ );
xor  ( new_n60721_, new_n51758_, new_n3113_ );
nor  ( new_n60722_, new_n60721_, new_n3461_ );
nor  ( new_n60723_, new_n60722_, new_n60720_ );
xnor ( new_n60724_, new_n60718_, new_n60717_ );
or   ( new_n60725_, new_n60724_, new_n60723_ );
and  ( new_n60726_, new_n60725_, new_n60719_ );
or   ( new_n60727_, new_n60579_, new_n8266_ );
xor  ( new_n60728_, new_n46958_, RIbb2dcc0_55 );
nand ( new_n60729_, new_n60728_, new_n8042_ );
and  ( new_n60730_, new_n60729_, new_n60727_ );
nor  ( new_n60731_, new_n60730_, new_n60726_ );
nor  ( new_n60732_, new_n60496_, new_n5606_ );
xor  ( new_n60733_, new_n49265_, new_n5203_ );
nor  ( new_n60734_, new_n60733_, new_n5604_ );
or   ( new_n60735_, new_n60734_, new_n60732_ );
xor  ( new_n60736_, new_n60730_, new_n60726_ );
and  ( new_n60737_, new_n60736_, new_n60735_ );
nor  ( new_n60738_, new_n60737_, new_n60731_ );
and  ( new_n60739_, new_n60711_, new_n60694_ );
nor  ( new_n60740_, new_n60739_, new_n60738_ );
nor  ( new_n60741_, new_n60740_, new_n60713_ );
nor  ( new_n60742_, new_n60741_, new_n60678_ );
nor  ( new_n60743_, new_n60742_, new_n60677_ );
or   ( new_n60744_, new_n60743_, new_n60665_ );
and  ( new_n60745_, new_n60744_, new_n60664_ );
or   ( new_n60746_, new_n60745_, new_n60605_ );
and  ( new_n60747_, new_n60745_, new_n60605_ );
xor  ( new_n60748_, new_n47046_, new_n7174_ );
or   ( new_n60749_, new_n60748_, new_n7732_ );
or   ( new_n60750_, new_n60477_, new_n7734_ );
and  ( new_n60751_, new_n60750_, new_n60749_ );
or   ( new_n60752_, new_n60618_, new_n7186_ );
xor  ( new_n60753_, new_n47640_, new_n6635_ );
or   ( new_n60754_, new_n60753_, new_n7184_ );
and  ( new_n60755_, new_n60754_, new_n60752_ );
nor  ( new_n60756_, new_n60755_, new_n60751_ );
nor  ( new_n60757_, new_n60630_, new_n10061_ );
xor  ( new_n60758_, new_n46037_, new_n9418_ );
nor  ( new_n60759_, new_n60758_, new_n10059_ );
nor  ( new_n60760_, new_n60759_, new_n60757_ );
and  ( new_n60761_, new_n60755_, new_n60751_ );
nor  ( new_n60762_, new_n60761_, new_n60760_ );
or   ( new_n60763_, new_n60762_, new_n60756_ );
xor  ( new_n60764_, new_n60575_, new_n60574_ );
and  ( new_n60765_, new_n60764_, new_n60763_ );
xor  ( new_n60766_, new_n60764_, new_n60763_ );
xor  ( new_n60767_, new_n60597_, new_n60596_ );
and  ( new_n60768_, new_n60767_, new_n60766_ );
nor  ( new_n60769_, new_n60768_, new_n60765_ );
xor  ( new_n60770_, new_n60481_, new_n60445_ );
xor  ( new_n60771_, new_n60770_, new_n60501_ );
nor  ( new_n60772_, new_n60771_, new_n60769_ );
xor  ( new_n60773_, new_n60771_, new_n60769_ );
xor  ( new_n60774_, new_n60519_, new_n60506_ );
xor  ( new_n60775_, new_n60774_, new_n60533_ );
and  ( new_n60776_, new_n60775_, new_n60773_ );
or   ( new_n60777_, new_n60776_, new_n60772_ );
xnor ( new_n60778_, new_n60535_, new_n60504_ );
xor  ( new_n60779_, new_n60778_, new_n60602_ );
nor  ( new_n60780_, new_n60779_, new_n60777_ );
nand ( new_n60781_, new_n60779_, new_n60777_ );
xor  ( new_n60782_, new_n60423_, new_n60422_ );
xor  ( new_n60783_, new_n60782_, new_n60438_ );
not  ( new_n60784_, new_n60783_ );
nor  ( new_n60785_, new_n60614_, new_n60611_ );
and  ( new_n60786_, new_n60614_, new_n60611_ );
nor  ( new_n60787_, new_n60786_, new_n60608_ );
nor  ( new_n60788_, new_n60787_, new_n60785_ );
xnor ( new_n60789_, new_n60137_, new_n60136_ );
or   ( new_n60790_, new_n60531_, new_n60528_ );
and  ( new_n60791_, new_n60531_, new_n60528_ );
or   ( new_n60792_, new_n60791_, new_n60525_ );
and  ( new_n60793_, new_n60792_, new_n60790_ );
xnor ( new_n60794_, new_n60793_, new_n60789_ );
xor  ( new_n60795_, new_n60794_, new_n60788_ );
xor  ( new_n60796_, new_n60795_, new_n60784_ );
nor  ( new_n60797_, new_n60517_, new_n60513_ );
and  ( new_n60798_, new_n60518_, new_n60510_ );
or   ( new_n60799_, new_n60798_, new_n60797_ );
xor  ( new_n60800_, new_n60162_, new_n60161_ );
xor  ( new_n60801_, new_n60800_, new_n60799_ );
nand ( new_n60802_, new_n60674_, new_n60670_ );
or   ( new_n60803_, new_n60674_, new_n60670_ );
nand ( new_n60804_, new_n60803_, new_n60669_ );
and  ( new_n60805_, new_n60804_, new_n60802_ );
xor  ( new_n60806_, new_n60805_, new_n60801_ );
xor  ( new_n60807_, new_n60806_, new_n60796_ );
not  ( new_n60808_, new_n60807_ );
and  ( new_n60809_, new_n60808_, new_n60781_ );
or   ( new_n60810_, new_n60809_, new_n60780_ );
or   ( new_n60811_, new_n60810_, new_n60747_ );
and  ( new_n60812_, new_n60811_, new_n60746_ );
and  ( new_n60813_, new_n60812_, new_n60402_ );
xor  ( new_n60814_, new_n60812_, new_n60402_ );
and  ( new_n60815_, new_n60443_, new_n60403_ );
and  ( new_n60816_, new_n60604_, new_n60444_ );
or   ( new_n60817_, new_n60816_, new_n60815_ );
and  ( new_n60818_, new_n60800_, new_n60799_ );
and  ( new_n60819_, new_n60805_, new_n60801_ );
or   ( new_n60820_, new_n60819_, new_n60818_ );
xnor ( new_n60821_, new_n60213_, new_n60194_ );
xor  ( new_n60822_, new_n60821_, new_n60240_ );
and  ( new_n60823_, new_n60822_, new_n60820_ );
nor  ( new_n60824_, new_n60822_, new_n60820_ );
nor  ( new_n60825_, new_n60793_, new_n60789_ );
and  ( new_n60826_, new_n60793_, new_n60789_ );
nor  ( new_n60827_, new_n60826_, new_n60788_ );
nor  ( new_n60828_, new_n60827_, new_n60825_ );
nor  ( new_n60829_, new_n60828_, new_n60824_ );
or   ( new_n60830_, new_n60829_, new_n60823_ );
or   ( new_n60831_, new_n60440_, new_n60406_ );
nand ( new_n60832_, new_n60442_, new_n60441_ );
and  ( new_n60833_, new_n60832_, new_n60831_ );
and  ( new_n60834_, new_n60307_, new_n60298_ );
and  ( new_n60835_, new_n60308_, new_n60287_ );
nor  ( new_n60836_, new_n60835_, new_n60834_ );
and  ( new_n60837_, new_n60192_, new_n9187_ );
and  ( new_n60838_, new_n59964_, new_n9185_ );
or   ( new_n60839_, new_n60838_, new_n60837_ );
nor  ( new_n60840_, new_n59911_, new_n8266_ );
and  ( new_n60841_, new_n60101_, new_n8042_ );
or   ( new_n60842_, new_n60841_, new_n60840_ );
nor  ( new_n60843_, new_n45119_, new_n10052_ );
or   ( new_n60844_, new_n44974_, RIbb2d900_63 );
and  ( new_n60845_, new_n60844_, RIbb2d888_64 );
or   ( new_n60846_, new_n60845_, new_n60843_ );
or   ( new_n60847_, new_n45209_, new_n10770_ );
and  ( new_n60848_, new_n60847_, new_n60846_ );
xor  ( new_n60849_, new_n60848_, new_n60842_ );
xor  ( new_n60850_, new_n60849_, new_n60839_ );
nor  ( new_n60851_, new_n60179_, new_n10059_ );
and  ( new_n60852_, new_n59917_, new_n9738_ );
nor  ( new_n60853_, new_n60852_, new_n60851_ );
or   ( new_n60854_, new_n60108_, new_n7184_ );
or   ( new_n60855_, new_n59895_, new_n7186_ );
and  ( new_n60856_, new_n60855_, new_n60854_ );
or   ( new_n60857_, new_n60114_, new_n8874_ );
nand ( new_n60858_, new_n59903_, new_n8649_ );
and  ( new_n60859_, new_n60858_, new_n60857_ );
xnor ( new_n60860_, new_n60859_, new_n60856_ );
nand ( new_n60861_, new_n60860_, new_n60853_ );
nor  ( new_n60862_, new_n60859_, new_n60856_ );
and  ( new_n60863_, new_n60859_, new_n60856_ );
nor  ( new_n60864_, new_n60863_, new_n60853_ );
not  ( new_n60865_, new_n60864_ );
or   ( new_n60866_, new_n60865_, new_n60862_ );
and  ( new_n60867_, new_n60866_, new_n60861_ );
xor  ( new_n60868_, new_n60867_, new_n60850_ );
xor  ( new_n60869_, new_n60868_, new_n60836_ );
xor  ( new_n60870_, new_n60869_, new_n60833_ );
xor  ( new_n60871_, new_n60870_, new_n60830_ );
xor  ( new_n60872_, new_n60871_, new_n60817_ );
xor  ( new_n60873_, new_n60822_, new_n60820_ );
xor  ( new_n60874_, new_n60873_, new_n60828_ );
nand ( new_n60875_, new_n60795_, new_n60784_ );
or   ( new_n60876_, new_n60795_, new_n60784_ );
nand ( new_n60877_, new_n60806_, new_n60876_ );
and  ( new_n60878_, new_n60877_, new_n60875_ );
or   ( new_n60879_, new_n60878_, new_n60874_ );
nand ( new_n60880_, new_n60878_, new_n60874_ );
xor  ( new_n60881_, new_n60346_, new_n60312_ );
nand ( new_n60882_, new_n60881_, new_n60880_ );
and  ( new_n60883_, new_n60882_, new_n60879_ );
xor  ( new_n60884_, new_n60883_, new_n60872_ );
and  ( new_n60885_, new_n60884_, new_n60814_ );
nor  ( new_n60886_, new_n60885_, new_n60813_ );
not  ( new_n60887_, new_n60886_ );
and  ( new_n60888_, new_n60848_, new_n60842_ );
and  ( new_n60889_, new_n60849_, new_n60839_ );
nor  ( new_n60890_, new_n60889_, new_n60888_ );
not  ( new_n60891_, new_n60890_ );
xor  ( new_n60892_, new_n59841_, new_n59840_ );
xor  ( new_n60893_, new_n60892_, new_n60891_ );
xor  ( new_n60894_, new_n59968_, new_n59967_ );
xor  ( new_n60895_, new_n60894_, new_n60893_ );
or   ( new_n60896_, new_n60243_, new_n60189_ );
and  ( new_n60897_, new_n60243_, new_n60189_ );
or   ( new_n60898_, new_n60897_, new_n60184_ );
and  ( new_n60899_, new_n60898_, new_n60896_ );
nor  ( new_n60900_, new_n60864_, new_n60862_ );
xnor ( new_n60901_, new_n59877_, new_n59873_ );
xor  ( new_n60902_, new_n60901_, new_n59882_ );
xnor ( new_n60903_, new_n59901_, new_n59897_ );
nand ( new_n60904_, new_n60903_, new_n59906_ );
not  ( new_n60905_, new_n59908_ );
or   ( new_n60906_, new_n60905_, new_n59902_ );
and  ( new_n60907_, new_n60906_, new_n60904_ );
xor  ( new_n60908_, new_n60907_, new_n60902_ );
xor  ( new_n60909_, new_n60908_, new_n60900_ );
xor  ( new_n60910_, new_n60909_, new_n60899_ );
xor  ( new_n60911_, new_n60910_, new_n60895_ );
nor  ( new_n60912_, new_n60245_, new_n60169_ );
nand ( new_n60913_, new_n60245_, new_n60169_ );
and  ( new_n60914_, new_n60913_, new_n60121_ );
or   ( new_n60915_, new_n60914_, new_n60912_ );
nor  ( new_n60916_, new_n60119_, new_n60100_ );
and  ( new_n60917_, new_n60119_, new_n60100_ );
not  ( new_n60918_, new_n60917_ );
and  ( new_n60919_, new_n60918_, new_n60099_ );
nor  ( new_n60920_, new_n60919_, new_n60916_ );
xnor ( new_n60921_, new_n60041_, new_n60040_ );
xor  ( new_n60922_, new_n60921_, new_n60075_ );
xnor ( new_n60923_, new_n60005_, new_n60000_ );
xor  ( new_n60924_, new_n60923_, new_n60020_ );
xnor ( new_n60925_, new_n60924_, new_n60922_ );
xor  ( new_n60926_, new_n60925_, new_n60920_ );
xnor ( new_n60927_, new_n60926_, new_n60915_ );
xor  ( new_n60928_, new_n60927_, new_n60911_ );
nand ( new_n60929_, new_n60871_, new_n60817_ );
nor  ( new_n60930_, new_n60871_, new_n60817_ );
or   ( new_n60931_, new_n60883_, new_n60930_ );
and  ( new_n60932_, new_n60931_, new_n60929_ );
xor  ( new_n60933_, new_n60932_, new_n60928_ );
nor  ( new_n60934_, new_n60400_, new_n60348_ );
and  ( new_n60935_, new_n60400_, new_n60348_ );
nor  ( new_n60936_, new_n60935_, new_n60248_ );
nor  ( new_n60937_, new_n60936_, new_n60934_ );
nor  ( new_n60938_, new_n60869_, new_n60833_ );
nand ( new_n60939_, new_n60869_, new_n60833_ );
and  ( new_n60940_, new_n60939_, new_n60830_ );
or   ( new_n60941_, new_n60940_, new_n60938_ );
and  ( new_n60942_, new_n60398_, new_n60387_ );
nor  ( new_n60943_, new_n60398_, new_n60387_ );
nor  ( new_n60944_, new_n60943_, new_n60380_ );
nor  ( new_n60945_, new_n60944_, new_n60942_ );
and  ( new_n60946_, new_n60867_, new_n60850_ );
nor  ( new_n60947_, new_n60867_, new_n60850_ );
nor  ( new_n60948_, new_n60947_, new_n60836_ );
or   ( new_n60949_, new_n60948_, new_n60946_ );
nor  ( new_n60950_, new_n60396_, new_n60393_ );
and  ( new_n60951_, new_n60397_, new_n60390_ );
or   ( new_n60952_, new_n60951_, new_n60950_ );
and  ( new_n60953_, new_n60385_, new_n60384_ );
and  ( new_n60954_, new_n60386_, new_n60383_ );
or   ( new_n60955_, new_n60954_, new_n60953_ );
xor  ( new_n60956_, new_n59921_, new_n59920_ );
xor  ( new_n60957_, new_n60956_, new_n60955_ );
xor  ( new_n60958_, new_n60957_, new_n60952_ );
xnor ( new_n60959_, new_n60958_, new_n60949_ );
xor  ( new_n60960_, new_n60959_, new_n60945_ );
xnor ( new_n60961_, new_n60960_, new_n60941_ );
xor  ( new_n60962_, new_n60961_, new_n60937_ );
xnor ( new_n60963_, new_n60962_, new_n60933_ );
and  ( new_n60964_, new_n60963_, new_n60887_ );
xor  ( new_n60965_, new_n59890_, new_n59889_ );
and  ( new_n60966_, new_n60892_, new_n60891_ );
and  ( new_n60967_, new_n60894_, new_n60893_ );
or   ( new_n60968_, new_n60967_, new_n60966_ );
xor  ( new_n60969_, new_n59971_, new_n59970_ );
xor  ( new_n60970_, new_n60969_, new_n60968_ );
xnor ( new_n60971_, new_n60970_, new_n60965_ );
nor  ( new_n60972_, new_n60909_, new_n60899_ );
nand ( new_n60973_, new_n60909_, new_n60899_ );
and  ( new_n60974_, new_n60973_, new_n60895_ );
or   ( new_n60975_, new_n60974_, new_n60972_ );
xor  ( new_n60976_, new_n59925_, new_n59924_ );
xnor ( new_n60977_, new_n59844_, new_n59843_ );
nand ( new_n60978_, new_n60907_, new_n60902_ );
nor  ( new_n60979_, new_n60907_, new_n60902_ );
or   ( new_n60980_, new_n60979_, new_n60900_ );
and  ( new_n60981_, new_n60980_, new_n60978_ );
xor  ( new_n60982_, new_n60981_, new_n60977_ );
xor  ( new_n60983_, new_n60982_, new_n60976_ );
xnor ( new_n60984_, new_n60983_, new_n60975_ );
xor  ( new_n60985_, new_n60984_, new_n60971_ );
not  ( new_n60986_, new_n60985_ );
nand ( new_n60987_, new_n60960_, new_n60941_ );
nor  ( new_n60988_, new_n60960_, new_n60941_ );
or   ( new_n60989_, new_n60988_, new_n60937_ );
and  ( new_n60990_, new_n60989_, new_n60987_ );
xor  ( new_n60991_, new_n60990_, new_n60986_ );
not  ( new_n60992_, new_n60991_ );
nor  ( new_n60993_, new_n60926_, new_n60915_ );
and  ( new_n60994_, new_n60926_, new_n60915_ );
nor  ( new_n60995_, new_n60994_, new_n60911_ );
nor  ( new_n60996_, new_n60995_, new_n60993_ );
and  ( new_n60997_, new_n60924_, new_n60922_ );
nor  ( new_n60998_, new_n60924_, new_n60922_ );
nor  ( new_n60999_, new_n60998_, new_n60920_ );
nor  ( new_n61000_, new_n60999_, new_n60997_ );
and  ( new_n61001_, new_n60956_, new_n60955_ );
or   ( new_n61002_, new_n60956_, new_n60955_ );
and  ( new_n61003_, new_n61002_, new_n60952_ );
or   ( new_n61004_, new_n61003_, new_n61001_ );
xnor ( new_n61005_, new_n60022_, new_n59984_ );
xor  ( new_n61006_, new_n61005_, new_n60077_ );
xor  ( new_n61007_, new_n61006_, new_n61004_ );
xor  ( new_n61008_, new_n61007_, new_n61000_ );
nand ( new_n61009_, new_n60958_, new_n60949_ );
nor  ( new_n61010_, new_n60958_, new_n60949_ );
or   ( new_n61011_, new_n61010_, new_n60945_ );
and  ( new_n61012_, new_n61011_, new_n61009_ );
xor  ( new_n61013_, new_n61012_, new_n61008_ );
xor  ( new_n61014_, new_n61013_, new_n60996_ );
xor  ( new_n61015_, new_n61014_, new_n60992_ );
or   ( new_n61016_, new_n60932_, new_n60928_ );
nand ( new_n61017_, new_n60932_, new_n60928_ );
nand ( new_n61018_, new_n60962_, new_n61017_ );
and  ( new_n61019_, new_n61018_, new_n61016_ );
and  ( new_n61020_, new_n61019_, new_n61015_ );
nor  ( new_n61021_, new_n61020_, new_n60964_ );
xor  ( new_n61022_, new_n60878_, new_n60874_ );
xor  ( new_n61023_, new_n61022_, new_n60881_ );
not  ( new_n61024_, new_n61023_ );
xor  ( new_n61025_, new_n60499_, new_n60498_ );
xnor ( new_n61026_, new_n60472_, new_n60467_ );
nand ( new_n61027_, new_n61026_, new_n60479_ );
not  ( new_n61028_, new_n60480_ );
or   ( new_n61029_, new_n61028_, new_n60473_ );
and  ( new_n61030_, new_n61029_, new_n61027_ );
and  ( new_n61031_, new_n61030_, new_n61025_ );
xor  ( new_n61032_, new_n61030_, new_n61025_ );
xnor ( new_n61033_, new_n60626_, new_n60620_ );
xor  ( new_n61034_, new_n61033_, new_n60632_ );
and  ( new_n61035_, new_n61034_, new_n61032_ );
or   ( new_n61036_, new_n61035_, new_n61031_ );
xnor ( new_n61037_, new_n60634_, new_n60616_ );
xor  ( new_n61038_, new_n61037_, new_n60659_ );
or   ( new_n61039_, new_n61038_, new_n61036_ );
nand ( new_n61040_, new_n61038_, new_n61036_ );
xnor ( new_n61041_, new_n60465_, new_n60464_ );
nand ( new_n61042_, new_n60652_, new_n4958_ );
xor  ( new_n61043_, new_n49758_, new_n4705_ );
or   ( new_n61044_, new_n61043_, new_n5207_ );
and  ( new_n61045_, new_n61044_, new_n61042_ );
or   ( new_n61046_, new_n60454_, new_n3119_ );
xor  ( new_n61047_, new_n52293_, RIbb2e710_33 );
or   ( new_n61048_, new_n61047_, new_n3117_ );
and  ( new_n61049_, new_n61048_, new_n61046_ );
or   ( new_n61050_, new_n61049_, new_n61045_ );
nor  ( new_n61051_, new_n60715_, new_n2809_ );
xor  ( new_n61052_, new_n53306_, RIbb2e800_31 );
nor  ( new_n61053_, new_n61052_, new_n2807_ );
or   ( new_n61054_, new_n61053_, new_n61051_ );
and  ( new_n61055_, new_n53694_, new_n2242_ );
and  ( new_n61056_, new_n61055_, new_n61054_ );
nor  ( new_n61057_, new_n61047_, new_n3119_ );
xor  ( new_n61058_, new_n52902_, RIbb2e710_33 );
nor  ( new_n61059_, new_n61058_, new_n3117_ );
or   ( new_n61060_, new_n61059_, new_n61057_ );
xor  ( new_n61061_, new_n61055_, new_n61054_ );
and  ( new_n61062_, new_n61061_, new_n61060_ );
nor  ( new_n61063_, new_n61062_, new_n61056_ );
and  ( new_n61064_, new_n61049_, new_n61045_ );
or   ( new_n61065_, new_n61064_, new_n61063_ );
and  ( new_n61066_, new_n61065_, new_n61050_ );
or   ( new_n61067_, new_n61066_, new_n61041_ );
xor  ( new_n61068_, new_n61066_, new_n61041_ );
and  ( new_n61069_, new_n45738_, RIbb2d888_64 );
nand ( new_n61070_, new_n61069_, RIbb2d900_63 );
or   ( new_n61071_, new_n46076_, RIbb2d888_64 );
or   ( new_n61072_, new_n61069_, RIbb2d900_63 );
and  ( new_n61073_, new_n61072_, new_n61071_ );
and  ( new_n61074_, new_n61073_, new_n61070_ );
nand ( new_n61075_, new_n61074_, new_n61068_ );
and  ( new_n61076_, new_n61075_, new_n61067_ );
xor  ( new_n61077_, new_n50487_, new_n4292_ );
or   ( new_n61078_, new_n61077_, new_n4709_ );
or   ( new_n61079_, new_n60680_, new_n4711_ );
and  ( new_n61080_, new_n61079_, new_n61078_ );
or   ( new_n61081_, new_n60646_, new_n4304_ );
xor  ( new_n61082_, new_n50894_, new_n3892_ );
or   ( new_n61083_, new_n61082_, new_n4302_ );
and  ( new_n61084_, new_n61083_, new_n61081_ );
or   ( new_n61085_, new_n61084_, new_n61080_ );
nor  ( new_n61086_, new_n60684_, new_n3898_ );
xor  ( new_n61087_, new_n51446_, RIbb2e530_37 );
and  ( new_n61088_, new_n61087_, new_n3733_ );
or   ( new_n61089_, new_n61088_, new_n61086_ );
xor  ( new_n61090_, new_n61084_, new_n61080_ );
nand ( new_n61091_, new_n61090_, new_n61089_ );
and  ( new_n61092_, new_n61091_, new_n61085_ );
xor  ( new_n61093_, new_n48908_, new_n5594_ );
or   ( new_n61094_, new_n61093_, new_n6173_ );
nand ( new_n61095_, new_n60706_, new_n5915_ );
and  ( new_n61096_, new_n61095_, new_n61094_ );
xor  ( new_n61097_, new_n46962_, new_n8254_ );
or   ( new_n61098_, new_n61097_, new_n8874_ );
or   ( new_n61099_, new_n60696_, new_n8876_ );
and  ( new_n61100_, new_n61099_, new_n61098_ );
or   ( new_n61101_, new_n61100_, new_n61096_ );
nor  ( new_n61102_, new_n60733_, new_n5606_ );
xor  ( new_n61103_, new_n49427_, RIbb2e170_45 );
and  ( new_n61104_, new_n61103_, new_n5373_ );
nor  ( new_n61105_, new_n61104_, new_n61102_ );
and  ( new_n61106_, new_n61100_, new_n61096_ );
or   ( new_n61107_, new_n61106_, new_n61105_ );
and  ( new_n61108_, new_n61107_, new_n61101_ );
or   ( new_n61109_, new_n61108_, new_n61092_ );
xor  ( new_n61110_, new_n61108_, new_n61092_ );
xnor ( new_n61111_, new_n60724_, new_n60723_ );
xor  ( new_n61112_, new_n46619_, new_n8870_ );
or   ( new_n61113_, new_n61112_, new_n9422_ );
or   ( new_n61114_, new_n60701_, new_n9424_ );
and  ( new_n61115_, new_n61114_, new_n61113_ );
nand ( new_n61116_, new_n61115_, new_n61111_ );
and  ( new_n61117_, new_n60688_, new_n6508_ );
xor  ( new_n61118_, new_n48518_, RIbb2df90_49 );
and  ( new_n61119_, new_n61118_, new_n6510_ );
nor  ( new_n61120_, new_n61119_, new_n61117_ );
or   ( new_n61121_, new_n61115_, new_n61111_ );
nand ( new_n61122_, new_n61121_, new_n61120_ );
and  ( new_n61123_, new_n61122_, new_n61116_ );
nand ( new_n61124_, new_n61123_, new_n61110_ );
and  ( new_n61125_, new_n61124_, new_n61109_ );
nor  ( new_n61126_, new_n61125_, new_n61076_ );
xor  ( new_n61127_, new_n60692_, new_n60691_ );
xor  ( new_n61128_, new_n60655_, new_n60654_ );
and  ( new_n61129_, new_n61128_, new_n61127_ );
and  ( new_n61130_, new_n53694_, new_n45845_ );
or   ( new_n61131_, new_n61130_, new_n2424_ );
or   ( new_n61132_, new_n61052_, new_n2809_ );
and  ( new_n61133_, new_n45843_, RIbb2e800_31 );
and  ( new_n61134_, new_n53694_, RIbb2e710_33 );
nor  ( new_n61135_, new_n61134_, new_n61133_ );
and  ( new_n61136_, RIbb2e788_32, new_n2421_ );
nor  ( new_n61137_, new_n53694_, RIbb2e710_33 );
nor  ( new_n61138_, new_n61137_, new_n61136_ );
or   ( new_n61139_, new_n61138_, new_n61135_ );
and  ( new_n61140_, new_n61139_, new_n61132_ );
or   ( new_n61141_, new_n61140_, new_n61131_ );
or   ( new_n61142_, new_n60721_, new_n3463_ );
xor  ( new_n61143_, new_n52280_, new_n3113_ );
or   ( new_n61144_, new_n61143_, new_n3461_ );
and  ( new_n61145_, new_n61144_, new_n61142_ );
or   ( new_n61146_, new_n61145_, new_n61141_ );
and  ( new_n61147_, new_n61087_, new_n3731_ );
xor  ( new_n61148_, new_n51477_, RIbb2e530_37 );
and  ( new_n61149_, new_n61148_, new_n3733_ );
or   ( new_n61150_, new_n61149_, new_n61147_ );
xor  ( new_n61151_, new_n61145_, new_n61141_ );
nand ( new_n61152_, new_n61151_, new_n61150_ );
and  ( new_n61153_, new_n61152_, new_n61146_ );
xor  ( new_n61154_, new_n47296_, RIbb2ddb0_53 );
nand ( new_n61155_, new_n61154_, new_n7489_ );
or   ( new_n61156_, new_n60748_, new_n7734_ );
and  ( new_n61157_, new_n61156_, new_n61155_ );
nor  ( new_n61158_, new_n61157_, new_n61153_ );
xor  ( new_n61159_, new_n47303_, new_n7722_ );
nor  ( new_n61160_, new_n61159_, new_n8264_ );
and  ( new_n61161_, new_n60728_, new_n8040_ );
nor  ( new_n61162_, new_n61161_, new_n61160_ );
xnor ( new_n61163_, new_n61157_, new_n61153_ );
nor  ( new_n61164_, new_n61163_, new_n61162_ );
or   ( new_n61165_, new_n61164_, new_n61158_ );
xor  ( new_n61166_, new_n61128_, new_n61127_ );
and  ( new_n61167_, new_n61166_, new_n61165_ );
nor  ( new_n61168_, new_n61167_, new_n61129_ );
xnor ( new_n61169_, new_n61125_, new_n61076_ );
nor  ( new_n61170_, new_n61169_, new_n61168_ );
nor  ( new_n61171_, new_n61170_, new_n61126_ );
nand ( new_n61172_, new_n61171_, new_n61040_ );
and  ( new_n61173_, new_n61172_, new_n61039_ );
xnor ( new_n61174_, new_n60663_, new_n60661_ );
xor  ( new_n61175_, new_n61174_, new_n60743_ );
nand ( new_n61176_, new_n61175_, new_n61173_ );
nor  ( new_n61177_, new_n61175_, new_n61173_ );
xor  ( new_n61178_, new_n60709_, new_n60708_ );
xnor ( new_n61179_, new_n60755_, new_n60751_ );
nand ( new_n61180_, new_n61179_, new_n60760_ );
not  ( new_n61181_, new_n60756_ );
nand ( new_n61182_, new_n60762_, new_n61181_ );
and  ( new_n61183_, new_n61182_, new_n61180_ );
and  ( new_n61184_, new_n61183_, new_n61178_ );
or   ( new_n61185_, new_n61183_, new_n61178_ );
xor  ( new_n61186_, new_n48039_, RIbb2dea0_51 );
and  ( new_n61187_, new_n61186_, new_n6910_ );
nor  ( new_n61188_, new_n60753_, new_n7186_ );
or   ( new_n61189_, new_n61188_, new_n61187_ );
xor  ( new_n61190_, new_n46137_, RIbb2d9f0_61 );
and  ( new_n61191_, new_n61190_, new_n9740_ );
nor  ( new_n61192_, new_n60758_, new_n10061_ );
nor  ( new_n61193_, new_n61192_, new_n61191_ );
not  ( new_n61194_, new_n61193_ );
and  ( new_n61195_, new_n61194_, new_n61189_ );
nor  ( new_n61196_, new_n61194_, new_n61189_ );
nor  ( new_n61197_, new_n45928_, new_n10052_ );
nor  ( new_n61198_, new_n61197_, new_n10769_ );
and  ( new_n61199_, new_n45597_, RIbb2d888_64 );
nor  ( new_n61200_, new_n61199_, new_n61198_ );
and  ( new_n61201_, new_n61199_, new_n10052_ );
nor  ( new_n61202_, new_n61201_, new_n61200_ );
nor  ( new_n61203_, new_n61202_, new_n61196_ );
or   ( new_n61204_, new_n61203_, new_n61195_ );
and  ( new_n61205_, new_n61204_, new_n61185_ );
or   ( new_n61206_, new_n61205_, new_n61184_ );
xnor ( new_n61207_, new_n60642_, new_n60641_ );
xor  ( new_n61208_, new_n61207_, new_n60657_ );
nand ( new_n61209_, new_n61208_, new_n61206_ );
xor  ( new_n61210_, new_n61208_, new_n61206_ );
xor  ( new_n61211_, new_n60711_, new_n60695_ );
nand ( new_n61212_, new_n61211_, new_n60738_ );
not  ( new_n61213_, new_n60740_ );
or   ( new_n61214_, new_n61213_, new_n60713_ );
and  ( new_n61215_, new_n61214_, new_n61212_ );
nand ( new_n61216_, new_n61215_, new_n61210_ );
and  ( new_n61217_, new_n61216_, new_n61209_ );
xor  ( new_n61218_, new_n60676_, new_n60666_ );
xor  ( new_n61219_, new_n61218_, new_n60741_ );
nor  ( new_n61220_, new_n61219_, new_n61217_ );
and  ( new_n61221_, new_n61219_, new_n61217_ );
xor  ( new_n61222_, new_n60775_, new_n60773_ );
not  ( new_n61223_, new_n61222_ );
nor  ( new_n61224_, new_n61223_, new_n61221_ );
nor  ( new_n61225_, new_n61224_, new_n61220_ );
or   ( new_n61226_, new_n61225_, new_n61177_ );
and  ( new_n61227_, new_n61226_, new_n61176_ );
and  ( new_n61228_, new_n61227_, new_n61024_ );
xor  ( new_n61229_, new_n61227_, new_n61024_ );
xor  ( new_n61230_, new_n60745_, new_n60605_ );
xor  ( new_n61231_, new_n61230_, new_n60810_ );
and  ( new_n61232_, new_n61231_, new_n61229_ );
nor  ( new_n61233_, new_n61232_, new_n61228_ );
not  ( new_n61234_, new_n61233_ );
xor  ( new_n61235_, new_n60884_, new_n60814_ );
and  ( new_n61236_, new_n61235_, new_n61234_ );
not  ( new_n61237_, new_n61236_ );
xor  ( new_n61238_, new_n60779_, new_n60777_ );
xor  ( new_n61239_, new_n61238_, new_n60808_ );
xor  ( new_n61240_, new_n60767_, new_n60766_ );
xor  ( new_n61241_, new_n61034_, new_n61032_ );
nand ( new_n61242_, new_n61241_, new_n61240_ );
nor  ( new_n61243_, new_n61241_, new_n61240_ );
xor  ( new_n61244_, new_n60736_, new_n60735_ );
xor  ( new_n61245_, new_n61074_, new_n61068_ );
and  ( new_n61246_, new_n61245_, new_n61244_ );
nor  ( new_n61247_, new_n61245_, new_n61244_ );
xor  ( new_n61248_, new_n51142_, new_n3892_ );
nor  ( new_n61249_, new_n61248_, new_n4302_ );
nor  ( new_n61250_, new_n61082_, new_n4304_ );
or   ( new_n61251_, new_n61250_, new_n61249_ );
xor  ( new_n61252_, new_n61061_, new_n61060_ );
and  ( new_n61253_, new_n61252_, new_n61251_ );
xor  ( new_n61254_, new_n50115_, new_n4705_ );
nor  ( new_n61255_, new_n61254_, new_n5207_ );
nor  ( new_n61256_, new_n61043_, new_n5209_ );
or   ( new_n61257_, new_n61256_, new_n61255_ );
xor  ( new_n61258_, new_n61252_, new_n61251_ );
and  ( new_n61259_, new_n61258_, new_n61257_ );
or   ( new_n61260_, new_n61259_, new_n61253_ );
xnor ( new_n61261_, new_n61049_, new_n61045_ );
xor  ( new_n61262_, new_n61261_, new_n61063_ );
and  ( new_n61263_, new_n61262_, new_n61260_ );
nor  ( new_n61264_, new_n61262_, new_n61260_ );
nor  ( new_n61265_, new_n61058_, new_n3119_ );
xor  ( new_n61266_, new_n52908_, RIbb2e710_33 );
nor  ( new_n61267_, new_n61266_, new_n3117_ );
or   ( new_n61268_, new_n61267_, new_n61265_ );
xor  ( new_n61269_, new_n61140_, new_n61131_ );
nand ( new_n61270_, new_n61269_, new_n61268_ );
xor  ( new_n61271_, new_n51758_, new_n3457_ );
nor  ( new_n61272_, new_n61271_, new_n3896_ );
and  ( new_n61273_, new_n61148_, new_n3731_ );
or   ( new_n61274_, new_n61273_, new_n61272_ );
xor  ( new_n61275_, new_n61269_, new_n61268_ );
nand ( new_n61276_, new_n61275_, new_n61274_ );
and  ( new_n61277_, new_n61276_, new_n61270_ );
xor  ( new_n61278_, new_n46958_, new_n8254_ );
or   ( new_n61279_, new_n61278_, new_n8874_ );
or   ( new_n61280_, new_n61097_, new_n8876_ );
and  ( new_n61281_, new_n61280_, new_n61279_ );
nor  ( new_n61282_, new_n61281_, new_n61277_ );
xor  ( new_n61283_, new_n47640_, new_n7174_ );
nor  ( new_n61284_, new_n61283_, new_n7732_ );
and  ( new_n61285_, new_n61154_, new_n7487_ );
or   ( new_n61286_, new_n61285_, new_n61284_ );
xor  ( new_n61287_, new_n61281_, new_n61277_ );
and  ( new_n61288_, new_n61287_, new_n61286_ );
nor  ( new_n61289_, new_n61288_, new_n61282_ );
nor  ( new_n61290_, new_n61289_, new_n61264_ );
nor  ( new_n61291_, new_n61290_, new_n61263_ );
nor  ( new_n61292_, new_n61291_, new_n61247_ );
nor  ( new_n61293_, new_n61292_, new_n61246_ );
or   ( new_n61294_, new_n61293_, new_n61243_ );
and  ( new_n61295_, new_n61294_, new_n61242_ );
xor  ( new_n61296_, new_n61038_, new_n61036_ );
xor  ( new_n61297_, new_n61296_, new_n61171_ );
or   ( new_n61298_, new_n61297_, new_n61295_ );
and  ( new_n61299_, new_n61297_, new_n61295_ );
xnor ( new_n61300_, new_n61169_, new_n61168_ );
xor  ( new_n61301_, new_n61123_, new_n61110_ );
xor  ( new_n61302_, new_n61183_, new_n61178_ );
xor  ( new_n61303_, new_n61302_, new_n61204_ );
nand ( new_n61304_, new_n61303_, new_n61301_ );
nor  ( new_n61305_, new_n61303_, new_n61301_ );
xor  ( new_n61306_, new_n46789_, new_n8870_ );
nor  ( new_n61307_, new_n61306_, new_n9422_ );
nor  ( new_n61308_, new_n61112_, new_n9424_ );
nor  ( new_n61309_, new_n61308_, new_n61307_ );
xor  ( new_n61310_, new_n48291_, new_n6635_ );
or   ( new_n61311_, new_n61310_, new_n7184_ );
nand ( new_n61312_, new_n61186_, new_n6908_ );
and  ( new_n61313_, new_n61312_, new_n61311_ );
or   ( new_n61314_, new_n61313_, new_n61309_ );
xnor ( new_n61315_, new_n61313_, new_n61309_ );
xor  ( new_n61316_, new_n45928_, new_n10052_ );
or   ( new_n61317_, new_n61316_, new_n21077_ );
or   ( new_n61318_, new_n46037_, new_n10052_ );
or   ( new_n61319_, new_n61318_, new_n10769_ );
and  ( new_n61320_, new_n61319_, new_n61317_ );
or   ( new_n61321_, new_n61320_, new_n61315_ );
and  ( new_n61322_, new_n61321_, new_n61314_ );
or   ( new_n61323_, new_n61248_, new_n4304_ );
xor  ( new_n61324_, new_n51446_, RIbb2e440_39 );
nand ( new_n61325_, new_n61324_, new_n4034_ );
and  ( new_n61326_, new_n61325_, new_n61323_ );
xor  ( new_n61327_, new_n49758_, new_n5203_ );
or   ( new_n61328_, new_n61327_, new_n5604_ );
xor  ( new_n61329_, new_n49488_, new_n5203_ );
or   ( new_n61330_, new_n61329_, new_n5606_ );
and  ( new_n61331_, new_n61330_, new_n61328_ );
nor  ( new_n61332_, new_n61331_, new_n61326_ );
xor  ( new_n61333_, new_n50894_, new_n4292_ );
nor  ( new_n61334_, new_n61333_, new_n4709_ );
xor  ( new_n61335_, new_n50788_, new_n4292_ );
nor  ( new_n61336_, new_n61335_, new_n4711_ );
nor  ( new_n61337_, new_n61336_, new_n61334_ );
xnor ( new_n61338_, new_n61331_, new_n61326_ );
nor  ( new_n61339_, new_n61338_, new_n61337_ );
or   ( new_n61340_, new_n61339_, new_n61332_ );
xor  ( new_n61341_, new_n61151_, new_n61150_ );
nand ( new_n61342_, new_n61341_, new_n61340_ );
nor  ( new_n61343_, new_n61341_, new_n61340_ );
or   ( new_n61344_, new_n61143_, new_n3463_ );
xor  ( new_n61345_, new_n52293_, RIbb2e620_35 );
or   ( new_n61346_, new_n61345_, new_n3461_ );
and  ( new_n61347_, new_n61346_, new_n61344_ );
nor  ( new_n61348_, new_n61266_, new_n3119_ );
xor  ( new_n61349_, new_n53306_, RIbb2e710_33 );
nor  ( new_n61350_, new_n61349_, new_n3117_ );
or   ( new_n61351_, new_n61350_, new_n61348_ );
and  ( new_n61352_, new_n53694_, new_n2613_ );
nand ( new_n61353_, new_n61352_, new_n61351_ );
xor  ( new_n61354_, new_n52902_, RIbb2e620_35 );
nor  ( new_n61355_, new_n61354_, new_n3461_ );
nor  ( new_n61356_, new_n61345_, new_n3463_ );
or   ( new_n61357_, new_n61356_, new_n61355_ );
xor  ( new_n61358_, new_n61352_, new_n61351_ );
nand ( new_n61359_, new_n61358_, new_n61357_ );
and  ( new_n61360_, new_n61359_, new_n61353_ );
nor  ( new_n61361_, new_n61360_, new_n61347_ );
xor  ( new_n61362_, new_n50487_, new_n4705_ );
nor  ( new_n61363_, new_n61362_, new_n5207_ );
nor  ( new_n61364_, new_n61254_, new_n5209_ );
or   ( new_n61365_, new_n61364_, new_n61363_ );
xor  ( new_n61366_, new_n61360_, new_n61347_ );
and  ( new_n61367_, new_n61366_, new_n61365_ );
nor  ( new_n61368_, new_n61367_, new_n61361_ );
or   ( new_n61369_, new_n61368_, new_n61343_ );
and  ( new_n61370_, new_n61369_, new_n61342_ );
nor  ( new_n61371_, new_n61370_, new_n61322_ );
xor  ( new_n61372_, new_n61370_, new_n61322_ );
xor  ( new_n61373_, new_n61193_, new_n61189_ );
xor  ( new_n61374_, new_n61373_, new_n61202_ );
and  ( new_n61375_, new_n61374_, new_n61372_ );
nor  ( new_n61376_, new_n61375_, new_n61371_ );
or   ( new_n61377_, new_n61376_, new_n61305_ );
and  ( new_n61378_, new_n61377_, new_n61304_ );
nor  ( new_n61379_, new_n61378_, new_n61300_ );
and  ( new_n61380_, new_n61378_, new_n61300_ );
or   ( new_n61381_, new_n61335_, new_n4709_ );
or   ( new_n61382_, new_n61077_, new_n4711_ );
and  ( new_n61383_, new_n61382_, new_n61381_ );
nand ( new_n61384_, new_n61103_, new_n5371_ );
or   ( new_n61385_, new_n61329_, new_n5604_ );
and  ( new_n61386_, new_n61385_, new_n61384_ );
nor  ( new_n61387_, new_n61386_, new_n61383_ );
xor  ( new_n61388_, new_n48756_, RIbb2df90_49 );
and  ( new_n61389_, new_n61388_, new_n6510_ );
and  ( new_n61390_, new_n61118_, new_n6508_ );
or   ( new_n61391_, new_n61390_, new_n61389_ );
xor  ( new_n61392_, new_n61386_, new_n61383_ );
and  ( new_n61393_, new_n61392_, new_n61391_ );
nor  ( new_n61394_, new_n61393_, new_n61387_ );
xnor ( new_n61395_, new_n61090_, new_n61089_ );
nor  ( new_n61396_, new_n61395_, new_n61394_ );
xnor ( new_n61397_, new_n61395_, new_n61394_ );
nand ( new_n61398_, new_n61190_, new_n9738_ );
xor  ( new_n61399_, new_n46427_, new_n9418_ );
or   ( new_n61400_, new_n61399_, new_n10059_ );
and  ( new_n61401_, new_n61400_, new_n61398_ );
xor  ( new_n61402_, new_n47046_, new_n7722_ );
or   ( new_n61403_, new_n61402_, new_n8264_ );
or   ( new_n61404_, new_n61159_, new_n8266_ );
and  ( new_n61405_, new_n61404_, new_n61403_ );
nor  ( new_n61406_, new_n61405_, new_n61401_ );
and  ( new_n61407_, new_n61405_, new_n61401_ );
nor  ( new_n61408_, new_n61093_, new_n6175_ );
xor  ( new_n61409_, new_n49265_, new_n5594_ );
nor  ( new_n61410_, new_n61409_, new_n6173_ );
nor  ( new_n61411_, new_n61410_, new_n61408_ );
nor  ( new_n61412_, new_n61411_, new_n61407_ );
nor  ( new_n61413_, new_n61412_, new_n61406_ );
nor  ( new_n61414_, new_n61413_, new_n61397_ );
or   ( new_n61415_, new_n61414_, new_n61396_ );
xnor ( new_n61416_, new_n61163_, new_n61162_ );
xor  ( new_n61417_, new_n61115_, new_n61111_ );
xor  ( new_n61418_, new_n61417_, new_n61120_ );
nand ( new_n61419_, new_n61418_, new_n61416_ );
nor  ( new_n61420_, new_n61418_, new_n61416_ );
xor  ( new_n61421_, new_n61100_, new_n61096_ );
xnor ( new_n61422_, new_n61421_, new_n61105_ );
or   ( new_n61423_, new_n61422_, new_n61420_ );
and  ( new_n61424_, new_n61423_, new_n61419_ );
and  ( new_n61425_, new_n61424_, new_n61415_ );
xor  ( new_n61426_, new_n61424_, new_n61415_ );
xor  ( new_n61427_, new_n61166_, new_n61165_ );
and  ( new_n61428_, new_n61427_, new_n61426_ );
nor  ( new_n61429_, new_n61428_, new_n61425_ );
nor  ( new_n61430_, new_n61429_, new_n61380_ );
nor  ( new_n61431_, new_n61430_, new_n61379_ );
or   ( new_n61432_, new_n61431_, new_n61299_ );
and  ( new_n61433_, new_n61432_, new_n61298_ );
and  ( new_n61434_, new_n61433_, new_n61239_ );
xnor ( new_n61435_, new_n61433_, new_n61239_ );
xnor ( new_n61436_, new_n61175_, new_n61173_ );
xor  ( new_n61437_, new_n61436_, new_n61225_ );
nor  ( new_n61438_, new_n61437_, new_n61435_ );
nor  ( new_n61439_, new_n61438_, new_n61434_ );
not  ( new_n61440_, new_n61439_ );
xor  ( new_n61441_, new_n61231_, new_n61229_ );
and  ( new_n61442_, new_n61441_, new_n61440_ );
xor  ( new_n61443_, new_n61219_, new_n61217_ );
xor  ( new_n61444_, new_n61443_, new_n61223_ );
xor  ( new_n61445_, new_n61215_, new_n61210_ );
xnor ( new_n61446_, new_n61241_, new_n61240_ );
xor  ( new_n61447_, new_n61446_, new_n61293_ );
nand ( new_n61448_, new_n61447_, new_n61445_ );
nor  ( new_n61449_, new_n61447_, new_n61445_ );
xor  ( new_n61450_, new_n61413_, new_n61397_ );
xnor ( new_n61451_, new_n61262_, new_n61260_ );
xor  ( new_n61452_, new_n61451_, new_n61289_ );
and  ( new_n61453_, new_n61452_, new_n61450_ );
or   ( new_n61454_, new_n61452_, new_n61450_ );
nor  ( new_n61455_, new_n61409_, new_n6175_ );
xor  ( new_n61456_, new_n49427_, RIbb2e080_47 );
and  ( new_n61457_, new_n61456_, new_n5917_ );
or   ( new_n61458_, new_n61457_, new_n61455_ );
xor  ( new_n61459_, new_n61275_, new_n61274_ );
and  ( new_n61460_, new_n61459_, new_n61458_ );
xor  ( new_n61461_, new_n48908_, new_n6163_ );
nor  ( new_n61462_, new_n61461_, new_n6645_ );
and  ( new_n61463_, new_n61388_, new_n6508_ );
or   ( new_n61464_, new_n61463_, new_n61462_ );
xor  ( new_n61465_, new_n61459_, new_n61458_ );
and  ( new_n61466_, new_n61465_, new_n61464_ );
or   ( new_n61467_, new_n61466_, new_n61460_ );
xor  ( new_n61468_, new_n61392_, new_n61391_ );
and  ( new_n61469_, new_n61468_, new_n61467_ );
nor  ( new_n61470_, new_n61468_, new_n61467_ );
and  ( new_n61471_, new_n53694_, new_n46355_ );
or   ( new_n61472_, new_n61471_, new_n2800_ );
or   ( new_n61473_, new_n61349_, new_n3119_ );
or   ( new_n61474_, new_n61134_, new_n3117_ );
or   ( new_n61475_, new_n61474_, new_n61137_ );
and  ( new_n61476_, new_n61475_, new_n61473_ );
or   ( new_n61477_, new_n61476_, new_n61472_ );
xor  ( new_n61478_, new_n52280_, new_n3457_ );
or   ( new_n61479_, new_n61478_, new_n3896_ );
or   ( new_n61480_, new_n61271_, new_n3898_ );
and  ( new_n61481_, new_n61480_, new_n61479_ );
or   ( new_n61482_, new_n61481_, new_n61477_ );
and  ( new_n61483_, new_n61324_, new_n4032_ );
xor  ( new_n61484_, new_n51477_, RIbb2e440_39 );
and  ( new_n61485_, new_n61484_, new_n4034_ );
nor  ( new_n61486_, new_n61485_, new_n61483_ );
not  ( new_n61487_, new_n61486_ );
xor  ( new_n61488_, new_n61481_, new_n61477_ );
nand ( new_n61489_, new_n61488_, new_n61487_ );
and  ( new_n61490_, new_n61489_, new_n61482_ );
or   ( new_n61491_, new_n61399_, new_n10061_ );
xor  ( new_n61492_, new_n46619_, new_n9418_ );
or   ( new_n61493_, new_n61492_, new_n10059_ );
and  ( new_n61494_, new_n61493_, new_n61491_ );
nor  ( new_n61495_, new_n61494_, new_n61490_ );
nor  ( new_n61496_, new_n61402_, new_n8266_ );
xor  ( new_n61497_, new_n47296_, RIbb2dcc0_55 );
and  ( new_n61498_, new_n61497_, new_n8042_ );
or   ( new_n61499_, new_n61498_, new_n61496_ );
xor  ( new_n61500_, new_n61494_, new_n61490_ );
and  ( new_n61501_, new_n61500_, new_n61499_ );
nor  ( new_n61502_, new_n61501_, new_n61495_ );
nor  ( new_n61503_, new_n61502_, new_n61470_ );
or   ( new_n61504_, new_n61503_, new_n61469_ );
and  ( new_n61505_, new_n61504_, new_n61454_ );
or   ( new_n61506_, new_n61505_, new_n61453_ );
xnor ( new_n61507_, new_n61245_, new_n61244_ );
xor  ( new_n61508_, new_n61507_, new_n61291_ );
and  ( new_n61509_, new_n61508_, new_n61506_ );
nor  ( new_n61510_, new_n61508_, new_n61506_ );
or   ( new_n61511_, new_n61283_, new_n7734_ );
xor  ( new_n61512_, new_n48039_, new_n7174_ );
or   ( new_n61513_, new_n61512_, new_n7732_ );
and  ( new_n61514_, new_n61513_, new_n61511_ );
or   ( new_n61515_, new_n61278_, new_n8876_ );
xor  ( new_n61516_, new_n47303_, new_n8254_ );
or   ( new_n61517_, new_n61516_, new_n8874_ );
and  ( new_n61518_, new_n61517_, new_n61515_ );
nor  ( new_n61519_, new_n61518_, new_n61514_ );
and  ( new_n61520_, new_n61518_, new_n61514_ );
nor  ( new_n61521_, new_n61306_, new_n9424_ );
xor  ( new_n61522_, new_n46962_, new_n8870_ );
nor  ( new_n61523_, new_n61522_, new_n9422_ );
nor  ( new_n61524_, new_n61523_, new_n61521_ );
nor  ( new_n61525_, new_n61524_, new_n61520_ );
nor  ( new_n61526_, new_n61525_, new_n61519_ );
not  ( new_n61527_, new_n61526_ );
xor  ( new_n61528_, new_n61258_, new_n61257_ );
and  ( new_n61529_, new_n61528_, new_n61527_ );
xor  ( new_n61530_, new_n61528_, new_n61527_ );
xnor ( new_n61531_, new_n61405_, new_n61401_ );
nand ( new_n61532_, new_n61531_, new_n61411_ );
not  ( new_n61533_, new_n61412_ );
or   ( new_n61534_, new_n61533_, new_n61406_ );
and  ( new_n61535_, new_n61534_, new_n61532_ );
and  ( new_n61536_, new_n61535_, new_n61530_ );
nor  ( new_n61537_, new_n61536_, new_n61529_ );
xnor ( new_n61538_, new_n61418_, new_n61416_ );
xor  ( new_n61539_, new_n61538_, new_n61422_ );
nor  ( new_n61540_, new_n61539_, new_n61537_ );
xor  ( new_n61541_, new_n61539_, new_n61537_ );
not  ( new_n61542_, new_n61541_ );
xor  ( new_n61543_, new_n61287_, new_n61286_ );
xor  ( new_n61544_, new_n61320_, new_n61315_ );
nand ( new_n61545_, new_n61544_, new_n61543_ );
nor  ( new_n61546_, new_n61544_, new_n61543_ );
or   ( new_n61547_, new_n61310_, new_n7186_ );
xor  ( new_n61548_, new_n48518_, new_n6635_ );
or   ( new_n61549_, new_n61548_, new_n7184_ );
and  ( new_n61550_, new_n61549_, new_n61547_ );
xor  ( new_n61551_, new_n46037_, new_n10052_ );
or   ( new_n61552_, new_n61551_, new_n21077_ );
or   ( new_n61553_, RIbb2d888_64, new_n10052_ );
or   ( new_n61554_, new_n61553_, new_n46137_ );
and  ( new_n61555_, new_n61554_, new_n61552_ );
nor  ( new_n61556_, new_n61555_, new_n61550_ );
and  ( new_n61557_, new_n61555_, new_n61550_ );
xor  ( new_n61558_, new_n50115_, new_n5203_ );
nor  ( new_n61559_, new_n61558_, new_n5604_ );
nor  ( new_n61560_, new_n61327_, new_n5606_ );
or   ( new_n61561_, new_n61560_, new_n61559_ );
xor  ( new_n61562_, new_n61358_, new_n61357_ );
and  ( new_n61563_, new_n61562_, new_n61561_ );
xor  ( new_n61564_, new_n50788_, new_n4705_ );
nor  ( new_n61565_, new_n61564_, new_n5207_ );
nor  ( new_n61566_, new_n61362_, new_n5209_ );
nor  ( new_n61567_, new_n61566_, new_n61565_ );
xnor ( new_n61568_, new_n61562_, new_n61561_ );
nor  ( new_n61569_, new_n61568_, new_n61567_ );
nor  ( new_n61570_, new_n61569_, new_n61563_ );
nor  ( new_n61571_, new_n61570_, new_n61557_ );
nor  ( new_n61572_, new_n61571_, new_n61556_ );
or   ( new_n61573_, new_n61572_, new_n61546_ );
and  ( new_n61574_, new_n61573_, new_n61545_ );
nor  ( new_n61575_, new_n61574_, new_n61542_ );
nor  ( new_n61576_, new_n61575_, new_n61540_ );
nor  ( new_n61577_, new_n61576_, new_n61510_ );
nor  ( new_n61578_, new_n61577_, new_n61509_ );
or   ( new_n61579_, new_n61578_, new_n61449_ );
and  ( new_n61580_, new_n61579_, new_n61448_ );
and  ( new_n61581_, new_n61580_, new_n61444_ );
xor  ( new_n61582_, new_n61580_, new_n61444_ );
not  ( new_n61583_, new_n61582_ );
xnor ( new_n61584_, new_n61297_, new_n61295_ );
xor  ( new_n61585_, new_n61584_, new_n61431_ );
nor  ( new_n61586_, new_n61585_, new_n61583_ );
nor  ( new_n61587_, new_n61586_, new_n61581_ );
not  ( new_n61588_, new_n61587_ );
xor  ( new_n61589_, new_n61437_, new_n61435_ );
and  ( new_n61590_, new_n61589_, new_n61588_ );
xor  ( new_n61591_, new_n61427_, new_n61426_ );
xnor ( new_n61592_, new_n61303_, new_n61301_ );
xor  ( new_n61593_, new_n61592_, new_n61376_ );
and  ( new_n61594_, new_n61593_, new_n61591_ );
nor  ( new_n61595_, new_n61593_, new_n61591_ );
xor  ( new_n61596_, new_n61374_, new_n61372_ );
xor  ( new_n61597_, new_n61452_, new_n61450_ );
xor  ( new_n61598_, new_n61597_, new_n61504_ );
and  ( new_n61599_, new_n61598_, new_n61596_ );
nor  ( new_n61600_, new_n61598_, new_n61596_ );
xnor ( new_n61601_, new_n61338_, new_n61337_ );
nand ( new_n61602_, new_n61497_, new_n8040_ );
xor  ( new_n61603_, new_n47640_, new_n7722_ );
or   ( new_n61604_, new_n61603_, new_n8264_ );
and  ( new_n61605_, new_n61604_, new_n61602_ );
xor  ( new_n61606_, new_n48291_, RIbb2ddb0_53 );
nand ( new_n61607_, new_n61606_, new_n7489_ );
or   ( new_n61608_, new_n61512_, new_n7734_ );
and  ( new_n61609_, new_n61608_, new_n61607_ );
or   ( new_n61610_, new_n61609_, new_n61605_ );
and  ( new_n61611_, new_n61609_, new_n61605_ );
and  ( new_n61612_, new_n46427_, new_n21077_ );
and  ( new_n61613_, new_n46137_, RIbb2d888_64 );
xor  ( new_n61614_, new_n61613_, new_n10052_ );
or   ( new_n61615_, new_n61614_, new_n61612_ );
or   ( new_n61616_, new_n61615_, new_n61611_ );
and  ( new_n61617_, new_n61616_, new_n61610_ );
or   ( new_n61618_, new_n61617_, new_n61601_ );
xor  ( new_n61619_, new_n61617_, new_n61601_ );
xor  ( new_n61620_, new_n61465_, new_n61464_ );
nand ( new_n61621_, new_n61620_, new_n61619_ );
and  ( new_n61622_, new_n61621_, new_n61618_ );
xor  ( new_n61623_, new_n61500_, new_n61499_ );
xnor ( new_n61624_, new_n61518_, new_n61514_ );
xor  ( new_n61625_, new_n61624_, new_n61524_ );
nand ( new_n61626_, new_n61625_, new_n61623_ );
nor  ( new_n61627_, new_n61625_, new_n61623_ );
xor  ( new_n61628_, new_n48756_, RIbb2dea0_51 );
nand ( new_n61629_, new_n61628_, new_n6910_ );
or   ( new_n61630_, new_n61548_, new_n7186_ );
and  ( new_n61631_, new_n61630_, new_n61629_ );
or   ( new_n61632_, new_n61522_, new_n9424_ );
xor  ( new_n61633_, new_n46958_, new_n8870_ );
or   ( new_n61634_, new_n61633_, new_n9422_ );
and  ( new_n61635_, new_n61634_, new_n61632_ );
nor  ( new_n61636_, new_n61635_, new_n61631_ );
and  ( new_n61637_, new_n61635_, new_n61631_ );
not  ( new_n61638_, new_n61637_ );
xor  ( new_n61639_, new_n61488_, new_n61487_ );
and  ( new_n61640_, new_n61639_, new_n61638_ );
nor  ( new_n61641_, new_n61640_, new_n61636_ );
or   ( new_n61642_, new_n61641_, new_n61627_ );
and  ( new_n61643_, new_n61642_, new_n61626_ );
nor  ( new_n61644_, new_n61643_, new_n61622_ );
and  ( new_n61645_, new_n61643_, new_n61622_ );
xor  ( new_n61646_, new_n61535_, new_n61530_ );
not  ( new_n61647_, new_n61646_ );
nor  ( new_n61648_, new_n61647_, new_n61645_ );
nor  ( new_n61649_, new_n61648_, new_n61644_ );
nor  ( new_n61650_, new_n61649_, new_n61600_ );
nor  ( new_n61651_, new_n61650_, new_n61599_ );
nor  ( new_n61652_, new_n61651_, new_n61595_ );
nor  ( new_n61653_, new_n61652_, new_n61594_ );
xor  ( new_n61654_, new_n61378_, new_n61300_ );
xor  ( new_n61655_, new_n61654_, new_n61429_ );
and  ( new_n61656_, new_n61655_, new_n61653_ );
xor  ( new_n61657_, new_n61655_, new_n61653_ );
not  ( new_n61658_, new_n61657_ );
xnor ( new_n61659_, new_n61447_, new_n61445_ );
xor  ( new_n61660_, new_n61659_, new_n61578_ );
nor  ( new_n61661_, new_n61660_, new_n61658_ );
nor  ( new_n61662_, new_n61661_, new_n61656_ );
not  ( new_n61663_, new_n61662_ );
xor  ( new_n61664_, new_n61585_, new_n61583_ );
and  ( new_n61665_, new_n61664_, new_n61663_ );
nor  ( new_n61666_, new_n61665_, new_n61590_ );
xor  ( new_n61667_, new_n49265_, new_n6163_ );
nor  ( new_n61668_, new_n61667_, new_n6645_ );
nor  ( new_n61669_, new_n61461_, new_n6647_ );
nor  ( new_n61670_, new_n61669_, new_n61668_ );
or   ( new_n61671_, new_n61333_, new_n4711_ );
xor  ( new_n61672_, new_n51142_, new_n4292_ );
or   ( new_n61673_, new_n61672_, new_n4709_ );
and  ( new_n61674_, new_n61673_, new_n61671_ );
nand ( new_n61675_, new_n61456_, new_n5915_ );
xor  ( new_n61676_, new_n49488_, new_n5594_ );
or   ( new_n61677_, new_n61676_, new_n6173_ );
and  ( new_n61678_, new_n61677_, new_n61675_ );
xor  ( new_n61679_, new_n61678_, new_n61674_ );
xor  ( new_n61680_, new_n61679_, new_n61670_ );
xor  ( new_n61681_, new_n49758_, new_n5594_ );
or   ( new_n61682_, new_n61681_, new_n6173_ );
or   ( new_n61683_, new_n61676_, new_n6175_ );
and  ( new_n61684_, new_n61683_, new_n61682_ );
or   ( new_n61685_, new_n61672_, new_n4711_ );
xor  ( new_n61686_, new_n51446_, RIbb2e350_41 );
nand ( new_n61687_, new_n61686_, new_n4543_ );
and  ( new_n61688_, new_n61687_, new_n61685_ );
or   ( new_n61689_, new_n61688_, new_n61684_ );
nor  ( new_n61690_, new_n61564_, new_n5209_ );
xor  ( new_n61691_, new_n50894_, new_n4705_ );
nor  ( new_n61692_, new_n61691_, new_n5207_ );
nor  ( new_n61693_, new_n61692_, new_n61690_ );
and  ( new_n61694_, new_n61688_, new_n61684_ );
or   ( new_n61695_, new_n61694_, new_n61693_ );
and  ( new_n61696_, new_n61695_, new_n61689_ );
nor  ( new_n61697_, new_n61696_, new_n61680_ );
nand ( new_n61698_, new_n61696_, new_n61680_ );
or   ( new_n61699_, new_n61478_, new_n3898_ );
xor  ( new_n61700_, new_n52293_, RIbb2e530_37 );
or   ( new_n61701_, new_n61700_, new_n3896_ );
and  ( new_n61702_, new_n61701_, new_n61699_ );
xor  ( new_n61703_, new_n52908_, RIbb2e620_35 );
nor  ( new_n61704_, new_n61703_, new_n3463_ );
xor  ( new_n61705_, new_n53306_, RIbb2e620_35 );
nor  ( new_n61706_, new_n61705_, new_n3461_ );
or   ( new_n61707_, new_n61706_, new_n61704_ );
and  ( new_n61708_, new_n53694_, new_n2928_ );
nand ( new_n61709_, new_n61708_, new_n61707_ );
xor  ( new_n61710_, new_n52902_, RIbb2e530_37 );
nor  ( new_n61711_, new_n61710_, new_n3896_ );
nor  ( new_n61712_, new_n61700_, new_n3898_ );
or   ( new_n61713_, new_n61712_, new_n61711_ );
xor  ( new_n61714_, new_n61708_, new_n61707_ );
nand ( new_n61715_, new_n61714_, new_n61713_ );
and  ( new_n61716_, new_n61715_, new_n61709_ );
nor  ( new_n61717_, new_n61716_, new_n61702_ );
nor  ( new_n61718_, new_n61558_, new_n5606_ );
xor  ( new_n61719_, new_n50487_, new_n5203_ );
nor  ( new_n61720_, new_n61719_, new_n5604_ );
or   ( new_n61721_, new_n61720_, new_n61718_ );
xor  ( new_n61722_, new_n61716_, new_n61702_ );
and  ( new_n61723_, new_n61722_, new_n61721_ );
or   ( new_n61724_, new_n61723_, new_n61717_ );
and  ( new_n61725_, new_n61724_, new_n61698_ );
or   ( new_n61726_, new_n61725_, new_n61697_ );
xnor ( new_n61727_, new_n61555_, new_n61550_ );
xor  ( new_n61728_, new_n61727_, new_n61570_ );
and  ( new_n61729_, new_n61728_, new_n61726_ );
or   ( new_n61730_, new_n61728_, new_n61726_ );
xnor ( new_n61731_, new_n61568_, new_n61567_ );
xor  ( new_n61732_, new_n48518_, RIbb2ddb0_53 );
and  ( new_n61733_, new_n61732_, new_n7489_ );
and  ( new_n61734_, new_n61606_, new_n7487_ );
nor  ( new_n61735_, new_n61734_, new_n61733_ );
xor  ( new_n61736_, new_n47303_, new_n8870_ );
or   ( new_n61737_, new_n61736_, new_n9422_ );
or   ( new_n61738_, new_n61633_, new_n9424_ );
and  ( new_n61739_, new_n61738_, new_n61737_ );
or   ( new_n61740_, new_n61739_, new_n61735_ );
and  ( new_n61741_, new_n61739_, new_n61735_ );
or   ( new_n61742_, new_n46619_, new_n10052_ );
and  ( new_n61743_, new_n61742_, new_n10770_ );
and  ( new_n61744_, new_n46427_, RIbb2d888_64 );
or   ( new_n61745_, new_n61744_, new_n61743_ );
nand ( new_n61746_, new_n61744_, new_n10052_ );
and  ( new_n61747_, new_n61746_, new_n61745_ );
or   ( new_n61748_, new_n61747_, new_n61741_ );
and  ( new_n61749_, new_n61748_, new_n61740_ );
nor  ( new_n61750_, new_n61749_, new_n61731_ );
and  ( new_n61751_, new_n61749_, new_n61731_ );
xor  ( new_n61752_, new_n48039_, RIbb2dcc0_55 );
and  ( new_n61753_, new_n61752_, new_n8042_ );
nor  ( new_n61754_, new_n61603_, new_n8266_ );
nor  ( new_n61755_, new_n61754_, new_n61753_ );
xor  ( new_n61756_, new_n47296_, RIbb2dbd0_57 );
nand ( new_n61757_, new_n61756_, new_n8651_ );
xor  ( new_n61758_, new_n47046_, new_n8254_ );
or   ( new_n61759_, new_n61758_, new_n8876_ );
and  ( new_n61760_, new_n61759_, new_n61757_ );
nor  ( new_n61761_, new_n61760_, new_n61755_ );
and  ( new_n61762_, new_n53694_, new_n46719_ );
or   ( new_n61763_, new_n61762_, new_n3116_ );
or   ( new_n61764_, new_n61705_, new_n3463_ );
and  ( new_n61765_, new_n53694_, RIbb2e620_35 );
nor  ( new_n61766_, new_n53694_, RIbb2e620_35 );
or   ( new_n61767_, new_n61766_, new_n3461_ );
or   ( new_n61768_, new_n61767_, new_n61765_ );
and  ( new_n61769_, new_n61768_, new_n61764_ );
or   ( new_n61770_, new_n61769_, new_n61763_ );
xor  ( new_n61771_, new_n51758_, new_n3892_ );
or   ( new_n61772_, new_n61771_, new_n4304_ );
xor  ( new_n61773_, new_n52280_, new_n3892_ );
or   ( new_n61774_, new_n61773_, new_n4302_ );
and  ( new_n61775_, new_n61774_, new_n61772_ );
nor  ( new_n61776_, new_n61775_, new_n61770_ );
and  ( new_n61777_, new_n61686_, new_n4541_ );
xor  ( new_n61778_, new_n51477_, RIbb2e350_41 );
and  ( new_n61779_, new_n61778_, new_n4543_ );
or   ( new_n61780_, new_n61779_, new_n61777_ );
xor  ( new_n61781_, new_n61775_, new_n61770_ );
and  ( new_n61782_, new_n61781_, new_n61780_ );
nor  ( new_n61783_, new_n61782_, new_n61776_ );
and  ( new_n61784_, new_n61760_, new_n61755_ );
nor  ( new_n61785_, new_n61784_, new_n61783_ );
nor  ( new_n61786_, new_n61785_, new_n61761_ );
nor  ( new_n61787_, new_n61786_, new_n61751_ );
nor  ( new_n61788_, new_n61787_, new_n61750_ );
not  ( new_n61789_, new_n61788_ );
and  ( new_n61790_, new_n61789_, new_n61730_ );
or   ( new_n61791_, new_n61790_, new_n61729_ );
xnor ( new_n61792_, new_n61544_, new_n61543_ );
xor  ( new_n61793_, new_n61792_, new_n61572_ );
nand ( new_n61794_, new_n61793_, new_n61791_ );
nor  ( new_n61795_, new_n61793_, new_n61791_ );
xor  ( new_n61796_, new_n61620_, new_n61619_ );
nor  ( new_n61797_, new_n61678_, new_n61674_ );
and  ( new_n61798_, new_n61678_, new_n61674_ );
nor  ( new_n61799_, new_n61798_, new_n61670_ );
nor  ( new_n61800_, new_n61799_, new_n61797_ );
xnor ( new_n61801_, new_n61366_, new_n61365_ );
xnor ( new_n61802_, new_n61801_, new_n61800_ );
or   ( new_n61803_, new_n61758_, new_n8874_ );
or   ( new_n61804_, new_n61516_, new_n8876_ );
and  ( new_n61805_, new_n61804_, new_n61803_ );
xor  ( new_n61806_, new_n46789_, new_n9418_ );
or   ( new_n61807_, new_n61806_, new_n10059_ );
or   ( new_n61808_, new_n61492_, new_n10061_ );
and  ( new_n61809_, new_n61808_, new_n61807_ );
or   ( new_n61810_, new_n61809_, new_n61805_ );
nor  ( new_n61811_, new_n61354_, new_n3463_ );
nor  ( new_n61812_, new_n61703_, new_n3461_ );
or   ( new_n61813_, new_n61812_, new_n61811_ );
xor  ( new_n61814_, new_n61476_, new_n61472_ );
nand ( new_n61815_, new_n61814_, new_n61813_ );
nor  ( new_n61816_, new_n61771_, new_n4302_ );
and  ( new_n61817_, new_n61484_, new_n4032_ );
or   ( new_n61818_, new_n61817_, new_n61816_ );
xor  ( new_n61819_, new_n61814_, new_n61813_ );
nand ( new_n61820_, new_n61819_, new_n61818_ );
and  ( new_n61821_, new_n61820_, new_n61815_ );
and  ( new_n61822_, new_n61809_, new_n61805_ );
or   ( new_n61823_, new_n61822_, new_n61821_ );
and  ( new_n61824_, new_n61823_, new_n61810_ );
xor  ( new_n61825_, new_n61824_, new_n61802_ );
nor  ( new_n61826_, new_n61825_, new_n61796_ );
nand ( new_n61827_, new_n61825_, new_n61796_ );
nor  ( new_n61828_, new_n61667_, new_n6647_ );
xor  ( new_n61829_, new_n49427_, RIbb2df90_49 );
and  ( new_n61830_, new_n61829_, new_n6510_ );
or   ( new_n61831_, new_n61830_, new_n61828_ );
xor  ( new_n61832_, new_n61819_, new_n61818_ );
and  ( new_n61833_, new_n61832_, new_n61831_ );
nor  ( new_n61834_, new_n61806_, new_n10061_ );
xor  ( new_n61835_, new_n46962_, new_n9418_ );
nor  ( new_n61836_, new_n61835_, new_n10059_ );
nor  ( new_n61837_, new_n61836_, new_n61834_ );
xnor ( new_n61838_, new_n61832_, new_n61831_ );
nor  ( new_n61839_, new_n61838_, new_n61837_ );
or   ( new_n61840_, new_n61839_, new_n61833_ );
xor  ( new_n61841_, new_n61635_, new_n61631_ );
xor  ( new_n61842_, new_n61841_, new_n61639_ );
nor  ( new_n61843_, new_n61842_, new_n61840_ );
nand ( new_n61844_, new_n61842_, new_n61840_ );
xor  ( new_n61845_, new_n61809_, new_n61805_ );
xor  ( new_n61846_, new_n61845_, new_n61821_ );
and  ( new_n61847_, new_n61846_, new_n61844_ );
or   ( new_n61848_, new_n61847_, new_n61843_ );
and  ( new_n61849_, new_n61848_, new_n61827_ );
or   ( new_n61850_, new_n61849_, new_n61826_ );
or   ( new_n61851_, new_n61850_, new_n61795_ );
and  ( new_n61852_, new_n61851_, new_n61794_ );
nor  ( new_n61853_, new_n61801_, new_n61800_ );
nor  ( new_n61854_, new_n61824_, new_n61802_ );
or   ( new_n61855_, new_n61854_, new_n61853_ );
xnor ( new_n61856_, new_n61341_, new_n61340_ );
xor  ( new_n61857_, new_n61856_, new_n61368_ );
nand ( new_n61858_, new_n61857_, new_n61855_ );
nor  ( new_n61859_, new_n61857_, new_n61855_ );
xor  ( new_n61860_, new_n61468_, new_n61467_ );
xor  ( new_n61861_, new_n61860_, new_n61502_ );
or   ( new_n61862_, new_n61861_, new_n61859_ );
and  ( new_n61863_, new_n61862_, new_n61858_ );
nor  ( new_n61864_, new_n61863_, new_n61852_ );
xor  ( new_n61865_, new_n61574_, new_n61542_ );
xor  ( new_n61866_, new_n61863_, new_n61852_ );
and  ( new_n61867_, new_n61866_, new_n61865_ );
nor  ( new_n61868_, new_n61867_, new_n61864_ );
not  ( new_n61869_, new_n61868_ );
xnor ( new_n61870_, new_n61508_, new_n61506_ );
xor  ( new_n61871_, new_n61870_, new_n61576_ );
nor  ( new_n61872_, new_n61871_, new_n61869_ );
xor  ( new_n61873_, new_n61871_, new_n61869_ );
not  ( new_n61874_, new_n61873_ );
xnor ( new_n61875_, new_n61593_, new_n61591_ );
xor  ( new_n61876_, new_n61875_, new_n61651_ );
nor  ( new_n61877_, new_n61876_, new_n61874_ );
nor  ( new_n61878_, new_n61877_, new_n61872_ );
not  ( new_n61879_, new_n61878_ );
xor  ( new_n61880_, new_n61660_, new_n61658_ );
and  ( new_n61881_, new_n61880_, new_n61879_ );
not  ( new_n61882_, new_n61881_ );
xor  ( new_n61883_, new_n61876_, new_n61874_ );
xor  ( new_n61884_, new_n61598_, new_n61596_ );
xor  ( new_n61885_, new_n61884_, new_n61649_ );
xor  ( new_n61886_, new_n61643_, new_n61622_ );
xor  ( new_n61887_, new_n61886_, new_n61647_ );
xor  ( new_n61888_, new_n61857_, new_n61855_ );
xor  ( new_n61889_, new_n61888_, new_n61861_ );
or   ( new_n61890_, new_n61889_, new_n61887_ );
and  ( new_n61891_, new_n61889_, new_n61887_ );
xor  ( new_n61892_, new_n61793_, new_n61791_ );
xor  ( new_n61893_, new_n61892_, new_n61850_ );
or   ( new_n61894_, new_n61893_, new_n61891_ );
and  ( new_n61895_, new_n61894_, new_n61890_ );
nor  ( new_n61896_, new_n61895_, new_n61885_ );
and  ( new_n61897_, new_n61895_, new_n61885_ );
not  ( new_n61898_, new_n61897_ );
xor  ( new_n61899_, new_n61866_, new_n61865_ );
and  ( new_n61900_, new_n61899_, new_n61898_ );
nor  ( new_n61901_, new_n61900_, new_n61896_ );
and  ( new_n61902_, new_n61901_, new_n61883_ );
not  ( new_n61903_, new_n61902_ );
and  ( new_n61904_, new_n61903_, new_n61882_ );
and  ( new_n61905_, new_n61904_, new_n61666_ );
xor  ( new_n61906_, new_n48908_, new_n6635_ );
nor  ( new_n61907_, new_n61906_, new_n7184_ );
and  ( new_n61908_, new_n61628_, new_n6908_ );
or   ( new_n61909_, new_n61908_, new_n61907_ );
xor  ( new_n61910_, new_n61722_, new_n61721_ );
and  ( new_n61911_, new_n61910_, new_n61909_ );
nor  ( new_n61912_, new_n61681_, new_n6175_ );
xor  ( new_n61913_, new_n50115_, new_n5594_ );
nor  ( new_n61914_, new_n61913_, new_n6173_ );
or   ( new_n61915_, new_n61914_, new_n61912_ );
xor  ( new_n61916_, new_n61714_, new_n61713_ );
and  ( new_n61917_, new_n61916_, new_n61915_ );
xor  ( new_n61918_, new_n50788_, new_n5203_ );
nor  ( new_n61919_, new_n61918_, new_n5604_ );
nor  ( new_n61920_, new_n61719_, new_n5606_ );
nor  ( new_n61921_, new_n61920_, new_n61919_ );
xnor ( new_n61922_, new_n61916_, new_n61915_ );
nor  ( new_n61923_, new_n61922_, new_n61921_ );
or   ( new_n61924_, new_n61923_, new_n61917_ );
xor  ( new_n61925_, new_n61910_, new_n61909_ );
and  ( new_n61926_, new_n61925_, new_n61924_ );
nor  ( new_n61927_, new_n61926_, new_n61911_ );
xor  ( new_n61928_, new_n61609_, new_n61605_ );
xor  ( new_n61929_, new_n61928_, new_n61615_ );
nor  ( new_n61930_, new_n61929_, new_n61927_ );
xor  ( new_n61931_, new_n61929_, new_n61927_ );
xor  ( new_n61932_, new_n61696_, new_n61680_ );
xor  ( new_n61933_, new_n61932_, new_n61724_ );
and  ( new_n61934_, new_n61933_, new_n61931_ );
or   ( new_n61935_, new_n61934_, new_n61930_ );
xnor ( new_n61936_, new_n61625_, new_n61623_ );
xor  ( new_n61937_, new_n61936_, new_n61641_ );
nor  ( new_n61938_, new_n61937_, new_n61935_ );
nand ( new_n61939_, new_n61937_, new_n61935_ );
or   ( new_n61940_, new_n61691_, new_n5209_ );
xor  ( new_n61941_, new_n51142_, new_n4705_ );
or   ( new_n61942_, new_n61941_, new_n5207_ );
and  ( new_n61943_, new_n61942_, new_n61940_ );
nand ( new_n61944_, new_n61829_, new_n6508_ );
xor  ( new_n61945_, new_n49488_, new_n6163_ );
or   ( new_n61946_, new_n61945_, new_n6645_ );
and  ( new_n61947_, new_n61946_, new_n61944_ );
or   ( new_n61948_, new_n61947_, new_n61943_ );
xor  ( new_n61949_, new_n47640_, new_n8254_ );
nor  ( new_n61950_, new_n61949_, new_n8874_ );
and  ( new_n61951_, new_n61756_, new_n8649_ );
or   ( new_n61952_, new_n61951_, new_n61950_ );
xor  ( new_n61953_, new_n61947_, new_n61943_ );
nand ( new_n61954_, new_n61953_, new_n61952_ );
and  ( new_n61955_, new_n61954_, new_n61948_ );
nor  ( new_n61956_, new_n61710_, new_n3898_ );
xor  ( new_n61957_, new_n52908_, RIbb2e530_37 );
nor  ( new_n61958_, new_n61957_, new_n3896_ );
or   ( new_n61959_, new_n61958_, new_n61956_ );
xor  ( new_n61960_, new_n61769_, new_n61763_ );
nand ( new_n61961_, new_n61960_, new_n61959_ );
xor  ( new_n61962_, new_n51758_, new_n4292_ );
nor  ( new_n61963_, new_n61962_, new_n4709_ );
and  ( new_n61964_, new_n61778_, new_n4541_ );
nor  ( new_n61965_, new_n61964_, new_n61963_ );
xnor ( new_n61966_, new_n61960_, new_n61959_ );
or   ( new_n61967_, new_n61966_, new_n61965_ );
and  ( new_n61968_, new_n61967_, new_n61961_ );
xor  ( new_n61969_, new_n46619_, new_n10052_ );
or   ( new_n61970_, new_n61969_, new_n21077_ );
or   ( new_n61971_, new_n46789_, new_n10052_ );
or   ( new_n61972_, new_n61971_, new_n10769_ );
and  ( new_n61973_, new_n61972_, new_n61970_ );
or   ( new_n61974_, new_n61973_, new_n61968_ );
xor  ( new_n61975_, new_n46958_, RIbb2d9f0_61 );
and  ( new_n61976_, new_n61975_, new_n9740_ );
nor  ( new_n61977_, new_n61835_, new_n10061_ );
or   ( new_n61978_, new_n61977_, new_n61976_ );
xor  ( new_n61979_, new_n61973_, new_n61968_ );
nand ( new_n61980_, new_n61979_, new_n61978_ );
and  ( new_n61981_, new_n61980_, new_n61974_ );
nor  ( new_n61982_, new_n61981_, new_n61955_ );
xor  ( new_n61983_, new_n48291_, new_n7722_ );
or   ( new_n61984_, new_n61983_, new_n8264_ );
nand ( new_n61985_, new_n61752_, new_n8040_ );
and  ( new_n61986_, new_n61985_, new_n61984_ );
xor  ( new_n61987_, new_n47046_, new_n8870_ );
or   ( new_n61988_, new_n61987_, new_n9422_ );
or   ( new_n61989_, new_n61736_, new_n9424_ );
and  ( new_n61990_, new_n61989_, new_n61988_ );
nor  ( new_n61991_, new_n61990_, new_n61986_ );
xor  ( new_n61992_, new_n48756_, RIbb2ddb0_53 );
and  ( new_n61993_, new_n61992_, new_n7489_ );
and  ( new_n61994_, new_n61732_, new_n7487_ );
or   ( new_n61995_, new_n61994_, new_n61993_ );
nand ( new_n61996_, new_n61990_, new_n61986_ );
and  ( new_n61997_, new_n61996_, new_n61995_ );
or   ( new_n61998_, new_n61997_, new_n61991_ );
xor  ( new_n61999_, new_n61981_, new_n61955_ );
and  ( new_n62000_, new_n61999_, new_n61998_ );
or   ( new_n62001_, new_n62000_, new_n61982_ );
xnor ( new_n62002_, new_n61749_, new_n61731_ );
xor  ( new_n62003_, new_n62002_, new_n61786_ );
nor  ( new_n62004_, new_n62003_, new_n62001_ );
nand ( new_n62005_, new_n62003_, new_n62001_ );
xor  ( new_n62006_, new_n61760_, new_n61755_ );
not  ( new_n62007_, new_n62006_ );
and  ( new_n62008_, new_n62007_, new_n61783_ );
not  ( new_n62009_, new_n61761_ );
and  ( new_n62010_, new_n61785_, new_n62009_ );
nor  ( new_n62011_, new_n62010_, new_n62008_ );
xnor ( new_n62012_, new_n61688_, new_n61684_ );
xor  ( new_n62013_, new_n62012_, new_n61693_ );
nand ( new_n62014_, new_n62013_, new_n62011_ );
xor  ( new_n62015_, new_n62013_, new_n62011_ );
xnor ( new_n62016_, new_n61739_, new_n61735_ );
xor  ( new_n62017_, new_n62016_, new_n61747_ );
nand ( new_n62018_, new_n62017_, new_n62015_ );
and  ( new_n62019_, new_n62018_, new_n62014_ );
and  ( new_n62020_, new_n62019_, new_n62005_ );
or   ( new_n62021_, new_n62020_, new_n62004_ );
and  ( new_n62022_, new_n62021_, new_n61939_ );
or   ( new_n62023_, new_n62022_, new_n61938_ );
xor  ( new_n62024_, new_n61889_, new_n61887_ );
xor  ( new_n62025_, new_n62024_, new_n61893_ );
nor  ( new_n62026_, new_n62025_, new_n62023_ );
and  ( new_n62027_, new_n62025_, new_n62023_ );
xor  ( new_n62028_, new_n61728_, new_n61726_ );
xor  ( new_n62029_, new_n62028_, new_n61789_ );
not  ( new_n62030_, new_n62029_ );
xor  ( new_n62031_, new_n61825_, new_n61796_ );
xor  ( new_n62032_, new_n62031_, new_n61848_ );
nor  ( new_n62033_, new_n62032_, new_n62030_ );
xor  ( new_n62034_, new_n62032_, new_n62030_ );
not  ( new_n62035_, new_n62034_ );
xnor ( new_n62036_, new_n61838_, new_n61837_ );
nor  ( new_n62037_, new_n61906_, new_n7186_ );
xor  ( new_n62038_, new_n49265_, new_n6635_ );
nor  ( new_n62039_, new_n62038_, new_n7184_ );
or   ( new_n62040_, new_n62039_, new_n62037_ );
xor  ( new_n62041_, new_n61781_, new_n61780_ );
nand ( new_n62042_, new_n62041_, new_n62040_ );
nor  ( new_n62043_, new_n62041_, new_n62040_ );
or   ( new_n62044_, new_n61773_, new_n4304_ );
xor  ( new_n62045_, new_n52293_, RIbb2e440_39 );
or   ( new_n62046_, new_n62045_, new_n4302_ );
and  ( new_n62047_, new_n62046_, new_n62044_ );
nor  ( new_n62048_, new_n61957_, new_n3898_ );
xor  ( new_n62049_, new_n53306_, RIbb2e530_37 );
nor  ( new_n62050_, new_n62049_, new_n3896_ );
or   ( new_n62051_, new_n62050_, new_n62048_ );
and  ( new_n62052_, new_n53694_, new_n3291_ );
nand ( new_n62053_, new_n62052_, new_n62051_ );
xor  ( new_n62054_, new_n52902_, RIbb2e440_39 );
nor  ( new_n62055_, new_n62054_, new_n4302_ );
nor  ( new_n62056_, new_n62045_, new_n4304_ );
or   ( new_n62057_, new_n62056_, new_n62055_ );
xor  ( new_n62058_, new_n62052_, new_n62051_ );
nand ( new_n62059_, new_n62058_, new_n62057_ );
and  ( new_n62060_, new_n62059_, new_n62053_ );
or   ( new_n62061_, new_n62060_, new_n62047_ );
xor  ( new_n62062_, new_n50487_, new_n5594_ );
nor  ( new_n62063_, new_n62062_, new_n6173_ );
nor  ( new_n62064_, new_n61913_, new_n6175_ );
or   ( new_n62065_, new_n62064_, new_n62063_ );
xor  ( new_n62066_, new_n62060_, new_n62047_ );
nand ( new_n62067_, new_n62066_, new_n62065_ );
and  ( new_n62068_, new_n62067_, new_n62061_ );
or   ( new_n62069_, new_n62068_, new_n62043_ );
and  ( new_n62070_, new_n62069_, new_n62042_ );
or   ( new_n62071_, new_n62070_, new_n62036_ );
and  ( new_n62072_, new_n62070_, new_n62036_ );
xnor ( new_n62073_, new_n61922_, new_n61921_ );
xor  ( new_n62074_, new_n47296_, new_n8870_ );
or   ( new_n62075_, new_n62074_, new_n9422_ );
or   ( new_n62076_, new_n61987_, new_n9424_ );
and  ( new_n62077_, new_n62076_, new_n62075_ );
or   ( new_n62078_, new_n62038_, new_n7186_ );
xor  ( new_n62079_, new_n49427_, RIbb2dea0_51 );
nand ( new_n62080_, new_n62079_, new_n6910_ );
and  ( new_n62081_, new_n62080_, new_n62078_ );
or   ( new_n62082_, new_n62081_, new_n62077_ );
xor  ( new_n62083_, new_n48908_, new_n7174_ );
nor  ( new_n62084_, new_n62083_, new_n7732_ );
and  ( new_n62085_, new_n61992_, new_n7487_ );
nor  ( new_n62086_, new_n62085_, new_n62084_ );
and  ( new_n62087_, new_n62081_, new_n62077_ );
or   ( new_n62088_, new_n62087_, new_n62086_ );
and  ( new_n62089_, new_n62088_, new_n62082_ );
nor  ( new_n62090_, new_n62089_, new_n62073_ );
and  ( new_n62091_, new_n53694_, new_n47102_ );
or   ( new_n62092_, new_n62091_, new_n3460_ );
or   ( new_n62093_, new_n62049_, new_n3898_ );
and  ( new_n62094_, new_n47100_, RIbb2e530_37 );
and  ( new_n62095_, new_n53694_, RIbb2e440_39 );
nor  ( new_n62096_, new_n62095_, new_n62094_ );
and  ( new_n62097_, RIbb2e4b8_38, new_n3457_ );
nor  ( new_n62098_, new_n53694_, RIbb2e440_39 );
nor  ( new_n62099_, new_n62098_, new_n62097_ );
or   ( new_n62100_, new_n62099_, new_n62096_ );
and  ( new_n62101_, new_n62100_, new_n62093_ );
or   ( new_n62102_, new_n62101_, new_n62092_ );
xor  ( new_n62103_, new_n52280_, new_n4292_ );
or   ( new_n62104_, new_n62103_, new_n4709_ );
or   ( new_n62105_, new_n61962_, new_n4711_ );
and  ( new_n62106_, new_n62105_, new_n62104_ );
or   ( new_n62107_, new_n62106_, new_n62102_ );
xor  ( new_n62108_, new_n51446_, RIbb2e260_43 );
and  ( new_n62109_, new_n62108_, new_n4958_ );
xor  ( new_n62110_, new_n51477_, RIbb2e260_43 );
and  ( new_n62111_, new_n62110_, new_n4960_ );
or   ( new_n62112_, new_n62111_, new_n62109_ );
xor  ( new_n62113_, new_n62106_, new_n62102_ );
nand ( new_n62114_, new_n62113_, new_n62112_ );
and  ( new_n62115_, new_n62114_, new_n62107_ );
xor  ( new_n62116_, new_n48518_, new_n7722_ );
or   ( new_n62117_, new_n62116_, new_n8264_ );
or   ( new_n62118_, new_n61983_, new_n8266_ );
and  ( new_n62119_, new_n62118_, new_n62117_ );
nor  ( new_n62120_, new_n62119_, new_n62115_ );
xor  ( new_n62121_, new_n47303_, new_n9418_ );
nor  ( new_n62122_, new_n62121_, new_n10059_ );
and  ( new_n62123_, new_n61975_, new_n9738_ );
nor  ( new_n62124_, new_n62123_, new_n62122_ );
xnor ( new_n62125_, new_n62119_, new_n62115_ );
nor  ( new_n62126_, new_n62125_, new_n62124_ );
or   ( new_n62127_, new_n62126_, new_n62120_ );
xor  ( new_n62128_, new_n62089_, new_n62073_ );
and  ( new_n62129_, new_n62128_, new_n62127_ );
nor  ( new_n62130_, new_n62129_, new_n62090_ );
or   ( new_n62131_, new_n62130_, new_n62072_ );
and  ( new_n62132_, new_n62131_, new_n62071_ );
xor  ( new_n62133_, new_n61842_, new_n61840_ );
xor  ( new_n62134_, new_n62133_, new_n61846_ );
or   ( new_n62135_, new_n62134_, new_n62132_ );
nand ( new_n62136_, new_n62134_, new_n62132_ );
xor  ( new_n62137_, new_n61933_, new_n61931_ );
nand ( new_n62138_, new_n62137_, new_n62136_ );
and  ( new_n62139_, new_n62138_, new_n62135_ );
nor  ( new_n62140_, new_n62139_, new_n62035_ );
nor  ( new_n62141_, new_n62140_, new_n62033_ );
nor  ( new_n62142_, new_n62141_, new_n62027_ );
nor  ( new_n62143_, new_n62142_, new_n62026_ );
not  ( new_n62144_, new_n62143_ );
xor  ( new_n62145_, new_n61895_, new_n61885_ );
xor  ( new_n62146_, new_n62145_, new_n61899_ );
nor  ( new_n62147_, new_n62146_, new_n62144_ );
xor  ( new_n62148_, new_n61937_, new_n61935_ );
xor  ( new_n62149_, new_n62148_, new_n62021_ );
or   ( new_n62150_, new_n61941_, new_n5209_ );
nand ( new_n62151_, new_n62108_, new_n4960_ );
and  ( new_n62152_, new_n62151_, new_n62150_ );
xor  ( new_n62153_, new_n49758_, new_n6163_ );
or   ( new_n62154_, new_n62153_, new_n6645_ );
or   ( new_n62155_, new_n61945_, new_n6647_ );
and  ( new_n62156_, new_n62155_, new_n62154_ );
or   ( new_n62157_, new_n62156_, new_n62152_ );
nor  ( new_n62158_, new_n61918_, new_n5606_ );
xor  ( new_n62159_, new_n50894_, new_n5203_ );
nor  ( new_n62160_, new_n62159_, new_n5604_ );
or   ( new_n62161_, new_n62160_, new_n62158_ );
xor  ( new_n62162_, new_n62156_, new_n62152_ );
nand ( new_n62163_, new_n62162_, new_n62161_ );
and  ( new_n62164_, new_n62163_, new_n62157_ );
xor  ( new_n62165_, new_n48039_, RIbb2dbd0_57 );
nand ( new_n62166_, new_n62165_, new_n8651_ );
or   ( new_n62167_, new_n61949_, new_n8876_ );
and  ( new_n62168_, new_n62167_, new_n62166_ );
xor  ( new_n62169_, new_n46789_, new_n10052_ );
or   ( new_n62170_, new_n62169_, new_n21077_ );
or   ( new_n62171_, new_n61553_, new_n46962_ );
and  ( new_n62172_, new_n62171_, new_n62170_ );
or   ( new_n62173_, new_n62172_, new_n62168_ );
and  ( new_n62174_, new_n62172_, new_n62168_ );
xnor ( new_n62175_, new_n61966_, new_n61965_ );
or   ( new_n62176_, new_n62175_, new_n62174_ );
and  ( new_n62177_, new_n62176_, new_n62173_ );
nor  ( new_n62178_, new_n62177_, new_n62164_ );
xor  ( new_n62179_, new_n61953_, new_n61952_ );
xor  ( new_n62180_, new_n62177_, new_n62164_ );
and  ( new_n62181_, new_n62180_, new_n62179_ );
or   ( new_n62182_, new_n62181_, new_n62178_ );
xor  ( new_n62183_, new_n61925_, new_n61924_ );
nand ( new_n62184_, new_n62183_, new_n62182_ );
xor  ( new_n62185_, new_n62183_, new_n62182_ );
xor  ( new_n62186_, new_n61999_, new_n61998_ );
nand ( new_n62187_, new_n62186_, new_n62185_ );
and  ( new_n62188_, new_n62187_, new_n62184_ );
xor  ( new_n62189_, new_n62003_, new_n62001_ );
xor  ( new_n62190_, new_n62189_, new_n62019_ );
or   ( new_n62191_, new_n62190_, new_n62188_ );
and  ( new_n62192_, new_n62190_, new_n62188_ );
xnor ( new_n62193_, new_n62017_, new_n62015_ );
xor  ( new_n62194_, new_n61990_, new_n61986_ );
xor  ( new_n62195_, new_n62194_, new_n61995_ );
xor  ( new_n62196_, new_n61979_, new_n61978_ );
nand ( new_n62197_, new_n62196_, new_n62195_ );
nor  ( new_n62198_, new_n62196_, new_n62195_ );
xor  ( new_n62199_, new_n62041_, new_n62040_ );
xor  ( new_n62200_, new_n62199_, new_n62068_ );
or   ( new_n62201_, new_n62200_, new_n62198_ );
and  ( new_n62202_, new_n62201_, new_n62197_ );
nor  ( new_n62203_, new_n62202_, new_n62193_ );
and  ( new_n62204_, new_n62202_, new_n62193_ );
xor  ( new_n62205_, new_n62070_, new_n62036_ );
xor  ( new_n62206_, new_n62205_, new_n62130_ );
nor  ( new_n62207_, new_n62206_, new_n62204_ );
nor  ( new_n62208_, new_n62207_, new_n62203_ );
or   ( new_n62209_, new_n62208_, new_n62192_ );
and  ( new_n62210_, new_n62209_, new_n62191_ );
nor  ( new_n62211_, new_n62210_, new_n62149_ );
xor  ( new_n62212_, new_n62139_, new_n62035_ );
xor  ( new_n62213_, new_n62210_, new_n62149_ );
and  ( new_n62214_, new_n62213_, new_n62212_ );
nor  ( new_n62215_, new_n62214_, new_n62211_ );
xor  ( new_n62216_, new_n62025_, new_n62023_ );
xor  ( new_n62217_, new_n62216_, new_n62141_ );
and  ( new_n62218_, new_n62217_, new_n62215_ );
nor  ( new_n62219_, new_n62218_, new_n62147_ );
xor  ( new_n62220_, new_n50788_, new_n5594_ );
nor  ( new_n62221_, new_n62220_, new_n6173_ );
nor  ( new_n62222_, new_n62062_, new_n6175_ );
or   ( new_n62223_, new_n62222_, new_n62221_ );
xor  ( new_n62224_, new_n62058_, new_n62057_ );
and  ( new_n62225_, new_n62224_, new_n62223_ );
and  ( new_n62226_, new_n62079_, new_n6908_ );
xor  ( new_n62227_, new_n49488_, RIbb2dea0_51 );
and  ( new_n62228_, new_n62227_, new_n6910_ );
nor  ( new_n62229_, new_n62228_, new_n62226_ );
xnor ( new_n62230_, new_n62224_, new_n62223_ );
nor  ( new_n62231_, new_n62230_, new_n62229_ );
or   ( new_n62232_, new_n62231_, new_n62225_ );
xor  ( new_n62233_, new_n62066_, new_n62065_ );
nand ( new_n62234_, new_n62233_, new_n62232_ );
nor  ( new_n62235_, new_n62121_, new_n10061_ );
xor  ( new_n62236_, new_n47046_, new_n9418_ );
nor  ( new_n62237_, new_n62236_, new_n10059_ );
nor  ( new_n62238_, new_n62237_, new_n62235_ );
xor  ( new_n62239_, new_n48756_, RIbb2dcc0_55 );
nand ( new_n62240_, new_n62239_, new_n8042_ );
or   ( new_n62241_, new_n62116_, new_n8266_ );
and  ( new_n62242_, new_n62241_, new_n62240_ );
nor  ( new_n62243_, new_n62242_, new_n62238_ );
nor  ( new_n62244_, new_n62054_, new_n4304_ );
xor  ( new_n62245_, new_n52908_, RIbb2e440_39 );
nor  ( new_n62246_, new_n62245_, new_n4302_ );
or   ( new_n62247_, new_n62246_, new_n62244_ );
xor  ( new_n62248_, new_n62101_, new_n62092_ );
and  ( new_n62249_, new_n62248_, new_n62247_ );
xor  ( new_n62250_, new_n52293_, RIbb2e350_41 );
nor  ( new_n62251_, new_n62250_, new_n4709_ );
nor  ( new_n62252_, new_n62103_, new_n4711_ );
or   ( new_n62253_, new_n62252_, new_n62251_ );
xor  ( new_n62254_, new_n62248_, new_n62247_ );
and  ( new_n62255_, new_n62254_, new_n62253_ );
nor  ( new_n62256_, new_n62255_, new_n62249_ );
and  ( new_n62257_, new_n62242_, new_n62238_ );
nor  ( new_n62258_, new_n62257_, new_n62256_ );
or   ( new_n62259_, new_n62258_, new_n62243_ );
xor  ( new_n62260_, new_n62233_, new_n62232_ );
nand ( new_n62261_, new_n62260_, new_n62259_ );
and  ( new_n62262_, new_n62261_, new_n62234_ );
xor  ( new_n62263_, new_n51142_, new_n5203_ );
or   ( new_n62264_, new_n62263_, new_n5604_ );
or   ( new_n62265_, new_n62159_, new_n5606_ );
and  ( new_n62266_, new_n62265_, new_n62264_ );
or   ( new_n62267_, new_n62153_, new_n6647_ );
xor  ( new_n62268_, new_n50115_, new_n6163_ );
or   ( new_n62269_, new_n62268_, new_n6645_ );
and  ( new_n62270_, new_n62269_, new_n62267_ );
nor  ( new_n62271_, new_n62270_, new_n62266_ );
and  ( new_n62272_, new_n62165_, new_n8649_ );
xor  ( new_n62273_, new_n48291_, RIbb2dbd0_57 );
and  ( new_n62274_, new_n62273_, new_n8651_ );
nor  ( new_n62275_, new_n62274_, new_n62272_ );
xnor ( new_n62276_, new_n62270_, new_n62266_ );
nor  ( new_n62277_, new_n62276_, new_n62275_ );
nor  ( new_n62278_, new_n62277_, new_n62271_ );
not  ( new_n62279_, new_n62278_ );
xor  ( new_n62280_, new_n62162_, new_n62161_ );
nand ( new_n62281_, new_n62280_, new_n62279_ );
xor  ( new_n62282_, new_n62280_, new_n62279_ );
not  ( new_n62283_, new_n62282_ );
xor  ( new_n62284_, new_n47640_, new_n8870_ );
or   ( new_n62285_, new_n62284_, new_n9422_ );
or   ( new_n62286_, new_n62074_, new_n9424_ );
and  ( new_n62287_, new_n62286_, new_n62285_ );
xor  ( new_n62288_, new_n49265_, new_n7174_ );
or   ( new_n62289_, new_n62288_, new_n7732_ );
or   ( new_n62290_, new_n62083_, new_n7734_ );
and  ( new_n62291_, new_n62290_, new_n62289_ );
or   ( new_n62292_, new_n62291_, new_n62287_ );
and  ( new_n62293_, new_n62291_, new_n62287_ );
and  ( new_n62294_, new_n46958_, new_n21077_ );
and  ( new_n62295_, new_n46962_, RIbb2d888_64 );
xor  ( new_n62296_, new_n62295_, new_n10052_ );
or   ( new_n62297_, new_n62296_, new_n62294_ );
or   ( new_n62298_, new_n62297_, new_n62293_ );
and  ( new_n62299_, new_n62298_, new_n62292_ );
or   ( new_n62300_, new_n62299_, new_n62283_ );
and  ( new_n62301_, new_n62300_, new_n62281_ );
nor  ( new_n62302_, new_n62301_, new_n62262_ );
xor  ( new_n62303_, new_n62128_, new_n62127_ );
xor  ( new_n62304_, new_n62301_, new_n62262_ );
and  ( new_n62305_, new_n62304_, new_n62303_ );
or   ( new_n62306_, new_n62305_, new_n62302_ );
xor  ( new_n62307_, new_n62186_, new_n62185_ );
and  ( new_n62308_, new_n62307_, new_n62306_ );
nor  ( new_n62309_, new_n62307_, new_n62306_ );
xnor ( new_n62310_, new_n62125_, new_n62124_ );
xor  ( new_n62311_, new_n62172_, new_n62168_ );
xor  ( new_n62312_, new_n62311_, new_n62175_ );
nor  ( new_n62313_, new_n62312_, new_n62310_ );
xor  ( new_n62314_, new_n62312_, new_n62310_ );
xnor ( new_n62315_, new_n62081_, new_n62077_ );
xor  ( new_n62316_, new_n62315_, new_n62086_ );
and  ( new_n62317_, new_n62316_, new_n62314_ );
nor  ( new_n62318_, new_n62317_, new_n62313_ );
xnor ( new_n62319_, new_n62180_, new_n62179_ );
nor  ( new_n62320_, new_n62319_, new_n62318_ );
xnor ( new_n62321_, new_n62319_, new_n62318_ );
xor  ( new_n62322_, new_n62196_, new_n62195_ );
xor  ( new_n62323_, new_n62322_, new_n62200_ );
nor  ( new_n62324_, new_n62323_, new_n62321_ );
nor  ( new_n62325_, new_n62324_, new_n62320_ );
nor  ( new_n62326_, new_n62325_, new_n62309_ );
nor  ( new_n62327_, new_n62326_, new_n62308_ );
not  ( new_n62328_, new_n62327_ );
xor  ( new_n62329_, new_n62134_, new_n62132_ );
xor  ( new_n62330_, new_n62329_, new_n62137_ );
and  ( new_n62331_, new_n62330_, new_n62328_ );
xor  ( new_n62332_, new_n62330_, new_n62328_ );
xnor ( new_n62333_, new_n62190_, new_n62188_ );
xor  ( new_n62334_, new_n62333_, new_n62208_ );
and  ( new_n62335_, new_n62334_, new_n62332_ );
nor  ( new_n62336_, new_n62335_, new_n62331_ );
xor  ( new_n62337_, new_n62213_, new_n62212_ );
not  ( new_n62338_, new_n62337_ );
and  ( new_n62339_, new_n62338_, new_n62336_ );
xor  ( new_n62340_, new_n62334_, new_n62332_ );
not  ( new_n62341_, new_n62340_ );
nor  ( new_n62342_, new_n62245_, new_n4304_ );
xor  ( new_n62343_, new_n53306_, RIbb2e440_39 );
nor  ( new_n62344_, new_n62343_, new_n4302_ );
or   ( new_n62345_, new_n62344_, new_n62342_ );
and  ( new_n62346_, new_n53694_, new_n3731_ );
nand ( new_n62347_, new_n62346_, new_n62345_ );
nor  ( new_n62348_, new_n62250_, new_n4711_ );
xor  ( new_n62349_, new_n52902_, RIbb2e350_41 );
nor  ( new_n62350_, new_n62349_, new_n4709_ );
or   ( new_n62351_, new_n62350_, new_n62348_ );
xor  ( new_n62352_, new_n62346_, new_n62345_ );
nand ( new_n62353_, new_n62352_, new_n62351_ );
and  ( new_n62354_, new_n62353_, new_n62347_ );
xor  ( new_n62355_, new_n51758_, new_n4705_ );
or   ( new_n62356_, new_n62355_, new_n5207_ );
nand ( new_n62357_, new_n62110_, new_n4958_ );
and  ( new_n62358_, new_n62357_, new_n62356_ );
nor  ( new_n62359_, new_n62358_, new_n62354_ );
xor  ( new_n62360_, new_n49758_, new_n6635_ );
nor  ( new_n62361_, new_n62360_, new_n7184_ );
and  ( new_n62362_, new_n62227_, new_n6908_ );
or   ( new_n62363_, new_n62362_, new_n62361_ );
xor  ( new_n62364_, new_n62358_, new_n62354_ );
and  ( new_n62365_, new_n62364_, new_n62363_ );
or   ( new_n62366_, new_n62365_, new_n62359_ );
xor  ( new_n62367_, new_n62113_, new_n62112_ );
and  ( new_n62368_, new_n62367_, new_n62366_ );
or   ( new_n62369_, new_n62263_, new_n5606_ );
xor  ( new_n62370_, new_n51446_, RIbb2e170_45 );
nand ( new_n62371_, new_n62370_, new_n5373_ );
and  ( new_n62372_, new_n62371_, new_n62369_ );
xor  ( new_n62373_, new_n50894_, new_n5594_ );
or   ( new_n62374_, new_n62373_, new_n6173_ );
or   ( new_n62375_, new_n62220_, new_n6175_ );
and  ( new_n62376_, new_n62375_, new_n62374_ );
nor  ( new_n62377_, new_n62376_, new_n62372_ );
xor  ( new_n62378_, new_n50487_, new_n6163_ );
nor  ( new_n62379_, new_n62378_, new_n6645_ );
nor  ( new_n62380_, new_n62268_, new_n6647_ );
or   ( new_n62381_, new_n62380_, new_n62379_ );
xor  ( new_n62382_, new_n62376_, new_n62372_ );
and  ( new_n62383_, new_n62382_, new_n62381_ );
nor  ( new_n62384_, new_n62383_, new_n62377_ );
xnor ( new_n62385_, new_n62367_, new_n62366_ );
nor  ( new_n62386_, new_n62385_, new_n62384_ );
nor  ( new_n62387_, new_n62386_, new_n62368_ );
not  ( new_n62388_, new_n62387_ );
xor  ( new_n62389_, new_n62260_, new_n62259_ );
and  ( new_n62390_, new_n62389_, new_n62388_ );
xor  ( new_n62391_, new_n62389_, new_n62388_ );
xnor ( new_n62392_, new_n62276_, new_n62275_ );
or   ( new_n62393_, new_n62288_, new_n7734_ );
xor  ( new_n62394_, new_n49427_, RIbb2ddb0_53 );
nand ( new_n62395_, new_n62394_, new_n7489_ );
and  ( new_n62396_, new_n62395_, new_n62393_ );
or   ( new_n62397_, new_n47303_, new_n10052_ );
and  ( new_n62398_, new_n62397_, new_n10770_ );
and  ( new_n62399_, new_n46958_, RIbb2d888_64 );
or   ( new_n62400_, new_n62399_, new_n62398_ );
nand ( new_n62401_, new_n62399_, new_n10052_ );
and  ( new_n62402_, new_n62401_, new_n62400_ );
or   ( new_n62403_, new_n62402_, new_n62396_ );
and  ( new_n62404_, new_n62402_, new_n62396_ );
xor  ( new_n62405_, new_n48908_, new_n7722_ );
nor  ( new_n62406_, new_n62405_, new_n8264_ );
and  ( new_n62407_, new_n62239_, new_n8040_ );
nor  ( new_n62408_, new_n62407_, new_n62406_ );
or   ( new_n62409_, new_n62408_, new_n62404_ );
and  ( new_n62410_, new_n62409_, new_n62403_ );
or   ( new_n62411_, new_n62410_, new_n62392_ );
and  ( new_n62412_, new_n62410_, new_n62392_ );
xor  ( new_n62413_, new_n48518_, RIbb2dbd0_57 );
and  ( new_n62414_, new_n62413_, new_n8651_ );
and  ( new_n62415_, new_n62273_, new_n8649_ );
or   ( new_n62416_, new_n62415_, new_n62414_ );
and  ( new_n62417_, new_n53694_, new_n47062_ );
or   ( new_n62418_, new_n62417_, new_n3895_ );
or   ( new_n62419_, new_n62343_, new_n4304_ );
or   ( new_n62420_, new_n62095_, new_n4302_ );
or   ( new_n62421_, new_n62420_, new_n62098_ );
and  ( new_n62422_, new_n62421_, new_n62419_ );
or   ( new_n62423_, new_n62422_, new_n62418_ );
or   ( new_n62424_, new_n62355_, new_n5209_ );
xor  ( new_n62425_, new_n52280_, new_n4705_ );
or   ( new_n62426_, new_n62425_, new_n5207_ );
and  ( new_n62427_, new_n62426_, new_n62424_ );
nand ( new_n62428_, new_n62427_, new_n62423_ );
or   ( new_n62429_, new_n62427_, new_n62423_ );
and  ( new_n62430_, new_n62370_, new_n5371_ );
xor  ( new_n62431_, new_n51477_, RIbb2e170_45 );
and  ( new_n62432_, new_n62431_, new_n5373_ );
nor  ( new_n62433_, new_n62432_, new_n62430_ );
nand ( new_n62434_, new_n62433_, new_n62429_ );
and  ( new_n62435_, new_n62434_, new_n62428_ );
and  ( new_n62436_, new_n62435_, new_n62416_ );
nor  ( new_n62437_, new_n62435_, new_n62416_ );
xor  ( new_n62438_, new_n47296_, RIbb2d9f0_61 );
and  ( new_n62439_, new_n62438_, new_n9740_ );
nor  ( new_n62440_, new_n62236_, new_n10061_ );
nor  ( new_n62441_, new_n62440_, new_n62439_ );
nor  ( new_n62442_, new_n62441_, new_n62437_ );
nor  ( new_n62443_, new_n62442_, new_n62436_ );
or   ( new_n62444_, new_n62443_, new_n62412_ );
nand ( new_n62445_, new_n62444_, new_n62411_ );
and  ( new_n62446_, new_n62445_, new_n62391_ );
or   ( new_n62447_, new_n62446_, new_n62390_ );
xor  ( new_n62448_, new_n62304_, new_n62303_ );
and  ( new_n62449_, new_n62448_, new_n62447_ );
or   ( new_n62450_, new_n62448_, new_n62447_ );
xor  ( new_n62451_, new_n62299_, new_n62283_ );
not  ( new_n62452_, new_n62451_ );
xnor ( new_n62453_, new_n62230_, new_n62229_ );
xor  ( new_n62454_, new_n62291_, new_n62287_ );
xor  ( new_n62455_, new_n62454_, new_n62297_ );
or   ( new_n62456_, new_n62455_, new_n62453_ );
nand ( new_n62457_, new_n62455_, new_n62453_ );
xor  ( new_n62458_, new_n62242_, new_n62238_ );
not  ( new_n62459_, new_n62458_ );
and  ( new_n62460_, new_n62459_, new_n62256_ );
not  ( new_n62461_, new_n62243_ );
and  ( new_n62462_, new_n62258_, new_n62461_ );
nor  ( new_n62463_, new_n62462_, new_n62460_ );
nand ( new_n62464_, new_n62463_, new_n62457_ );
and  ( new_n62465_, new_n62464_, new_n62456_ );
nor  ( new_n62466_, new_n62465_, new_n62452_ );
xor  ( new_n62467_, new_n62465_, new_n62452_ );
xor  ( new_n62468_, new_n62316_, new_n62314_ );
and  ( new_n62469_, new_n62468_, new_n62467_ );
or   ( new_n62470_, new_n62469_, new_n62466_ );
and  ( new_n62471_, new_n62470_, new_n62450_ );
or   ( new_n62472_, new_n62471_, new_n62449_ );
xnor ( new_n62473_, new_n62202_, new_n62193_ );
xor  ( new_n62474_, new_n62473_, new_n62206_ );
nor  ( new_n62475_, new_n62474_, new_n62472_ );
and  ( new_n62476_, new_n62474_, new_n62472_ );
xor  ( new_n62477_, new_n62307_, new_n62306_ );
xnor ( new_n62478_, new_n62477_, new_n62325_ );
nor  ( new_n62479_, new_n62478_, new_n62476_ );
nor  ( new_n62480_, new_n62479_, new_n62475_ );
not  ( new_n62481_, new_n62480_ );
and  ( new_n62482_, new_n62481_, new_n62341_ );
xor  ( new_n62483_, new_n62323_, new_n62321_ );
xor  ( new_n62484_, new_n62448_, new_n62447_ );
xor  ( new_n62485_, new_n62484_, new_n62470_ );
and  ( new_n62486_, new_n62485_, new_n62483_ );
nor  ( new_n62487_, new_n62485_, new_n62483_ );
xnor ( new_n62488_, new_n62445_, new_n62391_ );
xnor ( new_n62489_, new_n62385_, new_n62384_ );
xor  ( new_n62490_, new_n62382_, new_n62381_ );
xor  ( new_n62491_, new_n62364_, new_n62363_ );
nand ( new_n62492_, new_n62491_, new_n62490_ );
nor  ( new_n62493_, new_n62491_, new_n62490_ );
nor  ( new_n62494_, new_n62349_, new_n4711_ );
xor  ( new_n62495_, new_n52908_, RIbb2e350_41 );
nor  ( new_n62496_, new_n62495_, new_n4709_ );
or   ( new_n62497_, new_n62496_, new_n62494_ );
xor  ( new_n62498_, new_n62422_, new_n62418_ );
nand ( new_n62499_, new_n62498_, new_n62497_ );
nor  ( new_n62500_, new_n62425_, new_n5209_ );
xor  ( new_n62501_, new_n52293_, RIbb2e260_43 );
nor  ( new_n62502_, new_n62501_, new_n5207_ );
or   ( new_n62503_, new_n62502_, new_n62500_ );
xor  ( new_n62504_, new_n62498_, new_n62497_ );
nand ( new_n62505_, new_n62504_, new_n62503_ );
and  ( new_n62506_, new_n62505_, new_n62499_ );
xor  ( new_n62507_, new_n48756_, new_n8254_ );
or   ( new_n62508_, new_n62507_, new_n8874_ );
nand ( new_n62509_, new_n62413_, new_n8649_ );
and  ( new_n62510_, new_n62509_, new_n62508_ );
nor  ( new_n62511_, new_n62510_, new_n62506_ );
and  ( new_n62512_, new_n62438_, new_n9738_ );
xor  ( new_n62513_, new_n47640_, new_n9418_ );
nor  ( new_n62514_, new_n62513_, new_n10059_ );
nor  ( new_n62515_, new_n62514_, new_n62512_ );
and  ( new_n62516_, new_n62510_, new_n62506_ );
nor  ( new_n62517_, new_n62516_, new_n62515_ );
nor  ( new_n62518_, new_n62517_, new_n62511_ );
or   ( new_n62519_, new_n62518_, new_n62493_ );
and  ( new_n62520_, new_n62519_, new_n62492_ );
or   ( new_n62521_, new_n62520_, new_n62489_ );
and  ( new_n62522_, new_n62520_, new_n62489_ );
xor  ( new_n62523_, new_n48039_, RIbb2dae0_59 );
and  ( new_n62524_, new_n62523_, new_n9187_ );
nor  ( new_n62525_, new_n62284_, new_n9424_ );
or   ( new_n62526_, new_n62525_, new_n62524_ );
xor  ( new_n62527_, new_n62254_, new_n62253_ );
nand ( new_n62528_, new_n62527_, new_n62526_ );
nor  ( new_n62529_, new_n62373_, new_n6175_ );
xor  ( new_n62530_, new_n51142_, new_n5594_ );
nor  ( new_n62531_, new_n62530_, new_n6173_ );
or   ( new_n62532_, new_n62531_, new_n62529_ );
xor  ( new_n62533_, new_n62352_, new_n62351_ );
and  ( new_n62534_, new_n62533_, new_n62532_ );
and  ( new_n62535_, new_n62394_, new_n7487_ );
xor  ( new_n62536_, new_n49488_, RIbb2ddb0_53 );
and  ( new_n62537_, new_n62536_, new_n7489_ );
or   ( new_n62538_, new_n62537_, new_n62535_ );
xor  ( new_n62539_, new_n62533_, new_n62532_ );
and  ( new_n62540_, new_n62539_, new_n62538_ );
nor  ( new_n62541_, new_n62540_, new_n62534_ );
not  ( new_n62542_, new_n62541_ );
xor  ( new_n62543_, new_n62527_, new_n62526_ );
nand ( new_n62544_, new_n62543_, new_n62542_ );
and  ( new_n62545_, new_n62544_, new_n62528_ );
or   ( new_n62546_, new_n62545_, new_n62522_ );
and  ( new_n62547_, new_n62546_, new_n62521_ );
nor  ( new_n62548_, new_n62547_, new_n62488_ );
and  ( new_n62549_, new_n62547_, new_n62488_ );
not  ( new_n62550_, new_n62549_ );
xor  ( new_n62551_, new_n62468_, new_n62467_ );
and  ( new_n62552_, new_n62551_, new_n62550_ );
nor  ( new_n62553_, new_n62552_, new_n62548_ );
nor  ( new_n62554_, new_n62553_, new_n62487_ );
nor  ( new_n62555_, new_n62554_, new_n62486_ );
not  ( new_n62556_, new_n62555_ );
xor  ( new_n62557_, new_n62474_, new_n62472_ );
xnor ( new_n62558_, new_n62557_, new_n62478_ );
not  ( new_n62559_, new_n62558_ );
and  ( new_n62560_, new_n62559_, new_n62556_ );
xor  ( new_n62561_, new_n62435_, new_n62416_ );
xor  ( new_n62562_, new_n62561_, new_n62441_ );
xor  ( new_n62563_, new_n50788_, new_n6163_ );
or   ( new_n62564_, new_n62563_, new_n6645_ );
or   ( new_n62565_, new_n62378_, new_n6647_ );
and  ( new_n62566_, new_n62565_, new_n62564_ );
xor  ( new_n62567_, new_n50115_, new_n6635_ );
or   ( new_n62568_, new_n62567_, new_n7184_ );
or   ( new_n62569_, new_n62360_, new_n7186_ );
and  ( new_n62570_, new_n62569_, new_n62568_ );
or   ( new_n62571_, new_n62570_, new_n62566_ );
and  ( new_n62572_, new_n62523_, new_n9185_ );
xor  ( new_n62573_, new_n48291_, RIbb2dae0_59 );
and  ( new_n62574_, new_n62573_, new_n9187_ );
nor  ( new_n62575_, new_n62574_, new_n62572_ );
not  ( new_n62576_, new_n62575_ );
xor  ( new_n62577_, new_n62570_, new_n62566_ );
nand ( new_n62578_, new_n62577_, new_n62576_ );
and  ( new_n62579_, new_n62578_, new_n62571_ );
or   ( new_n62580_, new_n62405_, new_n8266_ );
xor  ( new_n62581_, new_n49265_, new_n7722_ );
or   ( new_n62582_, new_n62581_, new_n8264_ );
and  ( new_n62583_, new_n62582_, new_n62580_ );
xor  ( new_n62584_, new_n62427_, new_n62423_ );
xor  ( new_n62585_, new_n62584_, new_n62433_ );
and  ( new_n62586_, new_n62585_, new_n62583_ );
xor  ( new_n62587_, new_n47303_, new_n10052_ );
nor  ( new_n62588_, new_n62587_, new_n21077_ );
nor  ( new_n62589_, new_n47046_, new_n10052_ );
and  ( new_n62590_, new_n62589_, new_n10770_ );
nor  ( new_n62591_, new_n62590_, new_n62588_ );
or   ( new_n62592_, new_n62591_, new_n62586_ );
or   ( new_n62593_, new_n62585_, new_n62583_ );
and  ( new_n62594_, new_n62593_, new_n62592_ );
xnor ( new_n62595_, new_n62594_, new_n62579_ );
xor  ( new_n62596_, new_n62595_, new_n62562_ );
xor  ( new_n62597_, new_n62543_, new_n62542_ );
xor  ( new_n62598_, new_n51758_, new_n5203_ );
or   ( new_n62599_, new_n62598_, new_n5604_ );
nand ( new_n62600_, new_n62431_, new_n5371_ );
and  ( new_n62601_, new_n62600_, new_n62599_ );
nor  ( new_n62602_, new_n62495_, new_n4711_ );
xor  ( new_n62603_, new_n53306_, RIbb2e350_41 );
nor  ( new_n62604_, new_n62603_, new_n4709_ );
or   ( new_n62605_, new_n62604_, new_n62602_ );
and  ( new_n62606_, new_n53694_, new_n4032_ );
nand ( new_n62607_, new_n62606_, new_n62605_ );
nor  ( new_n62608_, new_n62501_, new_n5209_ );
xor  ( new_n62609_, new_n52902_, RIbb2e260_43 );
nor  ( new_n62610_, new_n62609_, new_n5207_ );
or   ( new_n62611_, new_n62610_, new_n62608_ );
xor  ( new_n62612_, new_n62606_, new_n62605_ );
nand ( new_n62613_, new_n62612_, new_n62611_ );
and  ( new_n62614_, new_n62613_, new_n62607_ );
or   ( new_n62615_, new_n62614_, new_n62601_ );
nor  ( new_n62616_, new_n62530_, new_n6175_ );
xor  ( new_n62617_, new_n51446_, RIbb2e080_47 );
and  ( new_n62618_, new_n62617_, new_n5917_ );
nor  ( new_n62619_, new_n62618_, new_n62616_ );
xnor ( new_n62620_, new_n62614_, new_n62601_ );
or   ( new_n62621_, new_n62620_, new_n62619_ );
and  ( new_n62622_, new_n62621_, new_n62615_ );
or   ( new_n62623_, new_n62567_, new_n7186_ );
xor  ( new_n62624_, new_n50487_, new_n6635_ );
or   ( new_n62625_, new_n62624_, new_n7184_ );
and  ( new_n62626_, new_n62625_, new_n62623_ );
or   ( new_n62627_, new_n62563_, new_n6647_ );
xor  ( new_n62628_, new_n50894_, new_n6163_ );
or   ( new_n62629_, new_n62628_, new_n6645_ );
and  ( new_n62630_, new_n62629_, new_n62627_ );
or   ( new_n62631_, new_n62630_, new_n62626_ );
and  ( new_n62632_, new_n62536_, new_n7487_ );
xor  ( new_n62633_, new_n49758_, new_n7174_ );
nor  ( new_n62634_, new_n62633_, new_n7732_ );
nor  ( new_n62635_, new_n62634_, new_n62632_ );
xnor ( new_n62636_, new_n62630_, new_n62626_ );
or   ( new_n62637_, new_n62636_, new_n62635_ );
and  ( new_n62638_, new_n62637_, new_n62631_ );
nor  ( new_n62639_, new_n62638_, new_n62622_ );
xor  ( new_n62640_, new_n62577_, new_n62576_ );
xor  ( new_n62641_, new_n62638_, new_n62622_ );
and  ( new_n62642_, new_n62641_, new_n62640_ );
or   ( new_n62643_, new_n62642_, new_n62639_ );
xnor ( new_n62644_, new_n62402_, new_n62396_ );
xor  ( new_n62645_, new_n62644_, new_n62408_ );
xor  ( new_n62646_, new_n62645_, new_n62643_ );
xor  ( new_n62647_, new_n62646_, new_n62597_ );
and  ( new_n62648_, new_n62647_, new_n62596_ );
nor  ( new_n62649_, new_n62647_, new_n62596_ );
xnor ( new_n62650_, new_n62641_, new_n62640_ );
xor  ( new_n62651_, new_n48291_, new_n9418_ );
or   ( new_n62652_, new_n62651_, new_n10059_ );
xor  ( new_n62653_, new_n48039_, RIbb2d9f0_61 );
nand ( new_n62654_, new_n62653_, new_n9738_ );
and  ( new_n62655_, new_n62654_, new_n62652_ );
xor  ( new_n62656_, new_n48756_, RIbb2dae0_59 );
nand ( new_n62657_, new_n62656_, new_n9187_ );
xor  ( new_n62658_, new_n48518_, RIbb2dae0_59 );
nand ( new_n62659_, new_n62658_, new_n9185_ );
and  ( new_n62660_, new_n62659_, new_n62657_ );
or   ( new_n62661_, new_n62660_, new_n62655_ );
xor  ( new_n62662_, new_n62660_, new_n62655_ );
nor  ( new_n62663_, new_n47640_, new_n10052_ );
or   ( new_n62664_, new_n62663_, RIbb2d888_64 );
and  ( new_n62665_, new_n47296_, new_n10052_ );
and  ( new_n62666_, new_n47986_, RIbb2d900_63 );
or   ( new_n62667_, new_n62666_, new_n21077_ );
or   ( new_n62668_, new_n62667_, new_n62665_ );
and  ( new_n62669_, new_n62668_, new_n62664_ );
nand ( new_n62670_, new_n62669_, new_n62662_ );
and  ( new_n62671_, new_n62670_, new_n62661_ );
or   ( new_n62672_, new_n62633_, new_n7734_ );
xor  ( new_n62673_, new_n50115_, new_n7174_ );
or   ( new_n62674_, new_n62673_, new_n7732_ );
and  ( new_n62675_, new_n62674_, new_n62672_ );
xor  ( new_n62676_, new_n50788_, new_n6635_ );
or   ( new_n62677_, new_n62676_, new_n7184_ );
or   ( new_n62678_, new_n62624_, new_n7186_ );
and  ( new_n62679_, new_n62678_, new_n62677_ );
or   ( new_n62680_, new_n62679_, new_n62675_ );
xor  ( new_n62681_, new_n48908_, new_n8254_ );
nor  ( new_n62682_, new_n62681_, new_n8876_ );
xor  ( new_n62683_, new_n49265_, new_n8254_ );
nor  ( new_n62684_, new_n62683_, new_n8874_ );
or   ( new_n62685_, new_n62684_, new_n62682_ );
xor  ( new_n62686_, new_n62679_, new_n62675_ );
nand ( new_n62687_, new_n62686_, new_n62685_ );
and  ( new_n62688_, new_n62687_, new_n62680_ );
or   ( new_n62689_, new_n62688_, new_n62671_ );
xnor ( new_n62690_, new_n62636_, new_n62635_ );
and  ( new_n62691_, new_n62688_, new_n62671_ );
or   ( new_n62692_, new_n62691_, new_n62690_ );
and  ( new_n62693_, new_n62692_, new_n62689_ );
nor  ( new_n62694_, new_n62693_, new_n62650_ );
and  ( new_n62695_, new_n62693_, new_n62650_ );
not  ( new_n62696_, new_n62695_ );
nor  ( new_n62697_, new_n62581_, new_n8266_ );
xor  ( new_n62698_, new_n49427_, RIbb2dcc0_55 );
and  ( new_n62699_, new_n62698_, new_n8042_ );
or   ( new_n62700_, new_n62699_, new_n62697_ );
xor  ( new_n62701_, new_n62504_, new_n62503_ );
and  ( new_n62702_, new_n62701_, new_n62700_ );
and  ( new_n62703_, new_n62573_, new_n9185_ );
and  ( new_n62704_, new_n62658_, new_n9187_ );
or   ( new_n62705_, new_n62704_, new_n62703_ );
xor  ( new_n62706_, new_n62701_, new_n62700_ );
and  ( new_n62707_, new_n62706_, new_n62705_ );
nor  ( new_n62708_, new_n62707_, new_n62702_ );
not  ( new_n62709_, new_n62708_ );
xor  ( new_n62710_, new_n62539_, new_n62538_ );
xor  ( new_n62711_, new_n62710_, new_n62709_ );
not  ( new_n62712_, new_n62711_ );
and  ( new_n62713_, new_n53694_, new_n47793_ );
or   ( new_n62714_, new_n62713_, new_n4295_ );
or   ( new_n62715_, new_n62603_, new_n4711_ );
and  ( new_n62716_, new_n53694_, RIbb2e350_41 );
nor  ( new_n62717_, new_n53694_, RIbb2e350_41 );
or   ( new_n62718_, new_n62717_, new_n4709_ );
or   ( new_n62719_, new_n62718_, new_n62716_ );
and  ( new_n62720_, new_n62719_, new_n62715_ );
or   ( new_n62721_, new_n62720_, new_n62714_ );
or   ( new_n62722_, new_n62598_, new_n5606_ );
xor  ( new_n62723_, new_n52280_, new_n5203_ );
or   ( new_n62724_, new_n62723_, new_n5604_ );
and  ( new_n62725_, new_n62724_, new_n62722_ );
or   ( new_n62726_, new_n62725_, new_n62721_ );
and  ( new_n62727_, new_n62617_, new_n5915_ );
xor  ( new_n62728_, new_n51477_, RIbb2e080_47 );
and  ( new_n62729_, new_n62728_, new_n5917_ );
or   ( new_n62730_, new_n62729_, new_n62727_ );
xor  ( new_n62731_, new_n62725_, new_n62721_ );
nand ( new_n62732_, new_n62731_, new_n62730_ );
and  ( new_n62733_, new_n62732_, new_n62726_ );
or   ( new_n62734_, new_n62681_, new_n8874_ );
or   ( new_n62735_, new_n62507_, new_n8876_ );
and  ( new_n62736_, new_n62735_, new_n62734_ );
or   ( new_n62737_, new_n62736_, new_n62733_ );
nor  ( new_n62738_, new_n62513_, new_n10061_ );
and  ( new_n62739_, new_n62653_, new_n9740_ );
nor  ( new_n62740_, new_n62739_, new_n62738_ );
and  ( new_n62741_, new_n62736_, new_n62733_ );
or   ( new_n62742_, new_n62741_, new_n62740_ );
and  ( new_n62743_, new_n62742_, new_n62737_ );
xor  ( new_n62744_, new_n62743_, new_n62712_ );
and  ( new_n62745_, new_n62744_, new_n62696_ );
nor  ( new_n62746_, new_n62745_, new_n62694_ );
nor  ( new_n62747_, new_n62746_, new_n62649_ );
nor  ( new_n62748_, new_n62747_, new_n62648_ );
not  ( new_n62749_, new_n62748_ );
nor  ( new_n62750_, new_n62594_, new_n62579_ );
and  ( new_n62751_, new_n62594_, new_n62579_ );
nor  ( new_n62752_, new_n62751_, new_n62562_ );
nor  ( new_n62753_, new_n62752_, new_n62750_ );
xor  ( new_n62754_, new_n62455_, new_n62453_ );
xor  ( new_n62755_, new_n62754_, new_n62463_ );
xnor ( new_n62756_, new_n62410_, new_n62392_ );
xor  ( new_n62757_, new_n62756_, new_n62443_ );
xnor ( new_n62758_, new_n62757_, new_n62755_ );
xor  ( new_n62759_, new_n62758_, new_n62753_ );
nor  ( new_n62760_, new_n62759_, new_n62749_ );
xor  ( new_n62761_, new_n62759_, new_n62749_ );
not  ( new_n62762_, new_n62761_ );
xnor ( new_n62763_, new_n62585_, new_n62583_ );
xor  ( new_n62764_, new_n62763_, new_n62591_ );
xnor ( new_n62765_, new_n62510_, new_n62506_ );
xor  ( new_n62766_, new_n62765_, new_n62515_ );
or   ( new_n62767_, new_n62766_, new_n62764_ );
and  ( new_n62768_, new_n62766_, new_n62764_ );
xnor ( new_n62769_, new_n62620_, new_n62619_ );
xor  ( new_n62770_, new_n47046_, new_n10052_ );
or   ( new_n62771_, new_n62770_, new_n21077_ );
nand ( new_n62772_, new_n62666_, new_n10770_ );
and  ( new_n62773_, new_n62772_, new_n62771_ );
nor  ( new_n62774_, new_n62773_, new_n62769_ );
nor  ( new_n62775_, new_n62628_, new_n6647_ );
xor  ( new_n62776_, new_n51142_, new_n6163_ );
nor  ( new_n62777_, new_n62776_, new_n6645_ );
or   ( new_n62778_, new_n62777_, new_n62775_ );
xor  ( new_n62779_, new_n62612_, new_n62611_ );
and  ( new_n62780_, new_n62779_, new_n62778_ );
and  ( new_n62781_, new_n62698_, new_n8040_ );
xor  ( new_n62782_, new_n49488_, RIbb2dcc0_55 );
and  ( new_n62783_, new_n62782_, new_n8042_ );
or   ( new_n62784_, new_n62783_, new_n62781_ );
xor  ( new_n62785_, new_n62779_, new_n62778_ );
and  ( new_n62786_, new_n62785_, new_n62784_ );
or   ( new_n62787_, new_n62786_, new_n62780_ );
xor  ( new_n62788_, new_n62773_, new_n62769_ );
and  ( new_n62789_, new_n62788_, new_n62787_ );
or   ( new_n62790_, new_n62789_, new_n62774_ );
or   ( new_n62791_, new_n62790_, new_n62768_ );
and  ( new_n62792_, new_n62791_, new_n62767_ );
xnor ( new_n62793_, new_n62491_, new_n62490_ );
xor  ( new_n62794_, new_n62793_, new_n62518_ );
and  ( new_n62795_, new_n62794_, new_n62792_ );
nor  ( new_n62796_, new_n62794_, new_n62792_ );
and  ( new_n62797_, new_n62710_, new_n62709_ );
nor  ( new_n62798_, new_n62743_, new_n62712_ );
nor  ( new_n62799_, new_n62798_, new_n62797_ );
nor  ( new_n62800_, new_n62799_, new_n62796_ );
nor  ( new_n62801_, new_n62800_, new_n62795_ );
nand ( new_n62802_, new_n62645_, new_n62643_ );
or   ( new_n62803_, new_n62645_, new_n62643_ );
nand ( new_n62804_, new_n62803_, new_n62597_ );
and  ( new_n62805_, new_n62804_, new_n62802_ );
xor  ( new_n62806_, new_n62520_, new_n62489_ );
xor  ( new_n62807_, new_n62806_, new_n62545_ );
xnor ( new_n62808_, new_n62807_, new_n62805_ );
xor  ( new_n62809_, new_n62808_, new_n62801_ );
nor  ( new_n62810_, new_n62809_, new_n62762_ );
nor  ( new_n62811_, new_n62810_, new_n62760_ );
not  ( new_n62812_, new_n62811_ );
and  ( new_n62813_, new_n62757_, new_n62755_ );
nor  ( new_n62814_, new_n62757_, new_n62755_ );
nor  ( new_n62815_, new_n62814_, new_n62753_ );
nor  ( new_n62816_, new_n62815_, new_n62813_ );
or   ( new_n62817_, new_n62807_, new_n62805_ );
and  ( new_n62818_, new_n62807_, new_n62805_ );
or   ( new_n62819_, new_n62818_, new_n62801_ );
and  ( new_n62820_, new_n62819_, new_n62817_ );
xor  ( new_n62821_, new_n62820_, new_n62816_ );
not  ( new_n62822_, new_n62821_ );
xor  ( new_n62823_, new_n62547_, new_n62488_ );
xor  ( new_n62824_, new_n62823_, new_n62551_ );
xor  ( new_n62825_, new_n62824_, new_n62822_ );
and  ( new_n62826_, new_n62825_, new_n62812_ );
not  ( new_n62827_, new_n62826_ );
xor  ( new_n62828_, new_n62809_, new_n62762_ );
xor  ( new_n62829_, new_n62794_, new_n62792_ );
xor  ( new_n62830_, new_n62829_, new_n62799_ );
xor  ( new_n62831_, new_n62706_, new_n62705_ );
xnor ( new_n62832_, new_n62736_, new_n62733_ );
xor  ( new_n62833_, new_n62832_, new_n62740_ );
and  ( new_n62834_, new_n62833_, new_n62831_ );
nor  ( new_n62835_, new_n62833_, new_n62831_ );
nor  ( new_n62836_, new_n62609_, new_n5209_ );
xor  ( new_n62837_, new_n52908_, RIbb2e260_43 );
nor  ( new_n62838_, new_n62837_, new_n5207_ );
or   ( new_n62839_, new_n62838_, new_n62836_ );
xor  ( new_n62840_, new_n62720_, new_n62714_ );
and  ( new_n62841_, new_n62840_, new_n62839_ );
and  ( new_n62842_, new_n62728_, new_n5915_ );
xor  ( new_n62843_, new_n51758_, new_n5594_ );
nor  ( new_n62844_, new_n62843_, new_n6173_ );
or   ( new_n62845_, new_n62844_, new_n62842_ );
xor  ( new_n62846_, new_n62840_, new_n62839_ );
and  ( new_n62847_, new_n62846_, new_n62845_ );
or   ( new_n62848_, new_n62847_, new_n62841_ );
xor  ( new_n62849_, new_n62731_, new_n62730_ );
and  ( new_n62850_, new_n62849_, new_n62848_ );
or   ( new_n62851_, new_n62673_, new_n7734_ );
xor  ( new_n62852_, new_n50487_, new_n7174_ );
or   ( new_n62853_, new_n62852_, new_n7732_ );
and  ( new_n62854_, new_n62853_, new_n62851_ );
or   ( new_n62855_, new_n62676_, new_n7186_ );
xor  ( new_n62856_, new_n50894_, new_n6635_ );
or   ( new_n62857_, new_n62856_, new_n7184_ );
and  ( new_n62858_, new_n62857_, new_n62855_ );
nor  ( new_n62859_, new_n62858_, new_n62854_ );
xor  ( new_n62860_, new_n49758_, new_n7722_ );
nor  ( new_n62861_, new_n62860_, new_n8264_ );
and  ( new_n62862_, new_n62782_, new_n8040_ );
or   ( new_n62863_, new_n62862_, new_n62861_ );
xor  ( new_n62864_, new_n62858_, new_n62854_ );
and  ( new_n62865_, new_n62864_, new_n62863_ );
or   ( new_n62866_, new_n62865_, new_n62859_ );
xor  ( new_n62867_, new_n62849_, new_n62848_ );
and  ( new_n62868_, new_n62867_, new_n62866_ );
nor  ( new_n62869_, new_n62868_, new_n62850_ );
nor  ( new_n62870_, new_n62869_, new_n62835_ );
or   ( new_n62871_, new_n62870_, new_n62834_ );
xor  ( new_n62872_, new_n62766_, new_n62764_ );
xor  ( new_n62873_, new_n62872_, new_n62790_ );
nand ( new_n62874_, new_n62873_, new_n62871_ );
nor  ( new_n62875_, new_n62873_, new_n62871_ );
or   ( new_n62876_, new_n62723_, new_n5606_ );
xor  ( new_n62877_, new_n52293_, RIbb2e170_45 );
or   ( new_n62878_, new_n62877_, new_n5604_ );
and  ( new_n62879_, new_n62878_, new_n62876_ );
nor  ( new_n62880_, new_n62837_, new_n5209_ );
xor  ( new_n62881_, new_n53306_, RIbb2e260_43 );
nor  ( new_n62882_, new_n62881_, new_n5207_ );
or   ( new_n62883_, new_n62882_, new_n62880_ );
and  ( new_n62884_, new_n53694_, new_n4541_ );
nand ( new_n62885_, new_n62884_, new_n62883_ );
nor  ( new_n62886_, new_n62877_, new_n5606_ );
xor  ( new_n62887_, new_n52902_, RIbb2e170_45 );
nor  ( new_n62888_, new_n62887_, new_n5604_ );
or   ( new_n62889_, new_n62888_, new_n62886_ );
xor  ( new_n62890_, new_n62884_, new_n62883_ );
nand ( new_n62891_, new_n62890_, new_n62889_ );
and  ( new_n62892_, new_n62891_, new_n62885_ );
nor  ( new_n62893_, new_n62892_, new_n62879_ );
nor  ( new_n62894_, new_n62776_, new_n6647_ );
xor  ( new_n62895_, new_n51446_, RIbb2df90_49 );
and  ( new_n62896_, new_n62895_, new_n6510_ );
or   ( new_n62897_, new_n62896_, new_n62894_ );
xor  ( new_n62898_, new_n62892_, new_n62879_ );
and  ( new_n62899_, new_n62898_, new_n62897_ );
or   ( new_n62900_, new_n62899_, new_n62893_ );
xor  ( new_n62901_, new_n62686_, new_n62685_ );
and  ( new_n62902_, new_n62901_, new_n62900_ );
nor  ( new_n62903_, new_n53695_, new_n48294_ );
or   ( new_n62904_, new_n62903_, new_n4708_ );
or   ( new_n62905_, new_n62881_, new_n5209_ );
and  ( new_n62906_, new_n53694_, RIbb2e260_43 );
nor  ( new_n62907_, new_n53694_, RIbb2e260_43 );
or   ( new_n62908_, new_n62907_, new_n5207_ );
or   ( new_n62909_, new_n62908_, new_n62906_ );
and  ( new_n62910_, new_n62909_, new_n62905_ );
or   ( new_n62911_, new_n62910_, new_n62904_ );
or   ( new_n62912_, new_n62843_, new_n6175_ );
xor  ( new_n62913_, new_n52280_, new_n5594_ );
or   ( new_n62914_, new_n62913_, new_n6173_ );
and  ( new_n62915_, new_n62914_, new_n62912_ );
nor  ( new_n62916_, new_n62915_, new_n62911_ );
and  ( new_n62917_, new_n62895_, new_n6508_ );
xor  ( new_n62918_, new_n51477_, RIbb2df90_49 );
and  ( new_n62919_, new_n62918_, new_n6510_ );
or   ( new_n62920_, new_n62919_, new_n62917_ );
xor  ( new_n62921_, new_n62915_, new_n62911_ );
and  ( new_n62922_, new_n62921_, new_n62920_ );
or   ( new_n62923_, new_n62922_, new_n62916_ );
xor  ( new_n62924_, new_n62846_, new_n62845_ );
and  ( new_n62925_, new_n62924_, new_n62923_ );
xor  ( new_n62926_, new_n48908_, new_n8870_ );
nor  ( new_n62927_, new_n62926_, new_n9422_ );
and  ( new_n62928_, new_n62656_, new_n9185_ );
or   ( new_n62929_, new_n62928_, new_n62927_ );
xor  ( new_n62930_, new_n62924_, new_n62923_ );
and  ( new_n62931_, new_n62930_, new_n62929_ );
nor  ( new_n62932_, new_n62931_, new_n62925_ );
xnor ( new_n62933_, new_n62901_, new_n62900_ );
nor  ( new_n62934_, new_n62933_, new_n62932_ );
or   ( new_n62935_, new_n62934_, new_n62902_ );
xor  ( new_n62936_, new_n62788_, new_n62787_ );
and  ( new_n62937_, new_n62936_, new_n62935_ );
or   ( new_n62938_, new_n62683_, new_n8876_ );
xor  ( new_n62939_, new_n49427_, RIbb2dbd0_57 );
nand ( new_n62940_, new_n62939_, new_n8651_ );
and  ( new_n62941_, new_n62940_, new_n62938_ );
or   ( new_n62942_, new_n62651_, new_n10061_ );
xor  ( new_n62943_, new_n48518_, RIbb2d9f0_61 );
nand ( new_n62944_, new_n62943_, new_n9740_ );
and  ( new_n62945_, new_n62944_, new_n62942_ );
nor  ( new_n62946_, new_n62945_, new_n62941_ );
and  ( new_n62947_, new_n57100_, new_n48040_ );
xor  ( new_n62948_, new_n47640_, new_n10052_ );
nor  ( new_n62949_, new_n62948_, new_n21077_ );
nor  ( new_n62950_, new_n62949_, new_n62947_ );
and  ( new_n62951_, new_n62945_, new_n62941_ );
nor  ( new_n62952_, new_n62951_, new_n62950_ );
or   ( new_n62953_, new_n62952_, new_n62946_ );
xor  ( new_n62954_, new_n62785_, new_n62784_ );
and  ( new_n62955_, new_n62954_, new_n62953_ );
xor  ( new_n62956_, new_n62669_, new_n62662_ );
xor  ( new_n62957_, new_n62954_, new_n62953_ );
and  ( new_n62958_, new_n62957_, new_n62956_ );
nor  ( new_n62959_, new_n62958_, new_n62955_ );
not  ( new_n62960_, new_n62959_ );
xor  ( new_n62961_, new_n62936_, new_n62935_ );
and  ( new_n62962_, new_n62961_, new_n62960_ );
nor  ( new_n62963_, new_n62962_, new_n62937_ );
or   ( new_n62964_, new_n62963_, new_n62875_ );
and  ( new_n62965_, new_n62964_, new_n62874_ );
nor  ( new_n62966_, new_n62965_, new_n62830_ );
and  ( new_n62967_, new_n62965_, new_n62830_ );
not  ( new_n62968_, new_n62967_ );
xor  ( new_n62969_, new_n62647_, new_n62596_ );
xnor ( new_n62970_, new_n62969_, new_n62746_ );
and  ( new_n62971_, new_n62970_, new_n62968_ );
nor  ( new_n62972_, new_n62971_, new_n62966_ );
and  ( new_n62973_, new_n62972_, new_n62828_ );
xor  ( new_n62974_, new_n62693_, new_n62650_ );
xor  ( new_n62975_, new_n62974_, new_n62744_ );
xnor ( new_n62976_, new_n62873_, new_n62871_ );
xor  ( new_n62977_, new_n62976_, new_n62963_ );
or   ( new_n62978_, new_n62977_, new_n62975_ );
xor  ( new_n62979_, new_n62977_, new_n62975_ );
xor  ( new_n62980_, new_n62688_, new_n62671_ );
xor  ( new_n62981_, new_n62980_, new_n62690_ );
xor  ( new_n62982_, new_n62833_, new_n62831_ );
xor  ( new_n62983_, new_n62982_, new_n62869_ );
or   ( new_n62984_, new_n62983_, new_n62981_ );
nand ( new_n62985_, new_n62983_, new_n62981_ );
xor  ( new_n62986_, new_n62961_, new_n62960_ );
nand ( new_n62987_, new_n62986_, new_n62985_ );
and  ( new_n62988_, new_n62987_, new_n62984_ );
nand ( new_n62989_, new_n62988_, new_n62979_ );
and  ( new_n62990_, new_n62989_, new_n62978_ );
xor  ( new_n62991_, new_n62965_, new_n62830_ );
xor  ( new_n62992_, new_n62991_, new_n62970_ );
and  ( new_n62993_, new_n62992_, new_n62990_ );
nor  ( new_n62994_, new_n62992_, new_n62990_ );
xor  ( new_n62995_, new_n62988_, new_n62979_ );
nor  ( new_n62996_, new_n62860_, new_n8266_ );
xor  ( new_n62997_, new_n50115_, new_n7722_ );
nor  ( new_n62998_, new_n62997_, new_n8264_ );
or   ( new_n62999_, new_n62998_, new_n62996_ );
xor  ( new_n63000_, new_n62890_, new_n62889_ );
and  ( new_n63001_, new_n63000_, new_n62999_ );
and  ( new_n63002_, new_n62939_, new_n8649_ );
xor  ( new_n63003_, new_n49488_, RIbb2dbd0_57 );
and  ( new_n63004_, new_n63003_, new_n8651_ );
or   ( new_n63005_, new_n63004_, new_n63002_ );
xor  ( new_n63006_, new_n63000_, new_n62999_ );
and  ( new_n63007_, new_n63006_, new_n63005_ );
or   ( new_n63008_, new_n63007_, new_n63001_ );
xor  ( new_n63009_, new_n62898_, new_n62897_ );
and  ( new_n63010_, new_n63009_, new_n63008_ );
xor  ( new_n63011_, new_n63009_, new_n63008_ );
xor  ( new_n63012_, new_n62864_, new_n62863_ );
and  ( new_n63013_, new_n63012_, new_n63011_ );
nor  ( new_n63014_, new_n63013_, new_n63010_ );
not  ( new_n63015_, new_n63014_ );
xor  ( new_n63016_, new_n62867_, new_n62866_ );
and  ( new_n63017_, new_n63016_, new_n63015_ );
xor  ( new_n63018_, new_n63016_, new_n63015_ );
xor  ( new_n63019_, new_n62957_, new_n62956_ );
and  ( new_n63020_, new_n63019_, new_n63018_ );
or   ( new_n63021_, new_n63020_, new_n63017_ );
xor  ( new_n63022_, new_n62983_, new_n62981_ );
xor  ( new_n63023_, new_n63022_, new_n62986_ );
nand ( new_n63024_, new_n63023_, new_n63021_ );
nor  ( new_n63025_, new_n63023_, new_n63021_ );
xnor ( new_n63026_, new_n62933_, new_n62932_ );
or   ( new_n63027_, new_n62997_, new_n8266_ );
xor  ( new_n63028_, new_n50487_, new_n7722_ );
or   ( new_n63029_, new_n63028_, new_n8264_ );
and  ( new_n63030_, new_n63029_, new_n63027_ );
xor  ( new_n63031_, new_n50788_, new_n7174_ );
or   ( new_n63032_, new_n63031_, new_n7734_ );
xor  ( new_n63033_, new_n50894_, new_n7174_ );
or   ( new_n63034_, new_n63033_, new_n7732_ );
and  ( new_n63035_, new_n63034_, new_n63032_ );
nor  ( new_n63036_, new_n63035_, new_n63030_ );
xor  ( new_n63037_, new_n51142_, new_n6635_ );
nor  ( new_n63038_, new_n63037_, new_n7186_ );
xor  ( new_n63039_, new_n51446_, RIbb2dea0_51 );
and  ( new_n63040_, new_n63039_, new_n6910_ );
nor  ( new_n63041_, new_n63040_, new_n63038_ );
and  ( new_n63042_, new_n63035_, new_n63030_ );
nor  ( new_n63043_, new_n63042_, new_n63041_ );
or   ( new_n63044_, new_n63043_, new_n63036_ );
xor  ( new_n63045_, new_n62921_, new_n62920_ );
and  ( new_n63046_, new_n63045_, new_n63044_ );
or   ( new_n63047_, new_n62913_, new_n6175_ );
xor  ( new_n63048_, new_n52293_, RIbb2e080_47 );
or   ( new_n63049_, new_n63048_, new_n6173_ );
and  ( new_n63050_, new_n63049_, new_n63047_ );
xor  ( new_n63051_, new_n52908_, RIbb2e170_45 );
nor  ( new_n63052_, new_n63051_, new_n5606_ );
xor  ( new_n63053_, new_n53306_, RIbb2e170_45 );
nor  ( new_n63054_, new_n63053_, new_n5604_ );
or   ( new_n63055_, new_n63054_, new_n63052_ );
and  ( new_n63056_, new_n53694_, new_n4958_ );
nand ( new_n63057_, new_n63056_, new_n63055_ );
xor  ( new_n63058_, new_n52902_, RIbb2e080_47 );
nor  ( new_n63059_, new_n63058_, new_n6173_ );
nor  ( new_n63060_, new_n63048_, new_n6175_ );
nor  ( new_n63061_, new_n63060_, new_n63059_ );
xnor ( new_n63062_, new_n63056_, new_n63055_ );
or   ( new_n63063_, new_n63062_, new_n63061_ );
and  ( new_n63064_, new_n63063_, new_n63057_ );
nor  ( new_n63065_, new_n63064_, new_n63050_ );
and  ( new_n63066_, new_n63003_, new_n8649_ );
xor  ( new_n63067_, new_n49758_, new_n8254_ );
nor  ( new_n63068_, new_n63067_, new_n8874_ );
nor  ( new_n63069_, new_n63068_, new_n63066_ );
not  ( new_n63070_, new_n63069_ );
xor  ( new_n63071_, new_n63064_, new_n63050_ );
and  ( new_n63072_, new_n63071_, new_n63070_ );
or   ( new_n63073_, new_n63072_, new_n63065_ );
xor  ( new_n63074_, new_n63045_, new_n63044_ );
and  ( new_n63075_, new_n63074_, new_n63073_ );
or   ( new_n63076_, new_n63075_, new_n63046_ );
xnor ( new_n63077_, new_n62945_, new_n62941_ );
nand ( new_n63078_, new_n63077_, new_n62950_ );
not  ( new_n63079_, new_n62946_ );
nand ( new_n63080_, new_n62952_, new_n63079_ );
and  ( new_n63081_, new_n63080_, new_n63078_ );
nand ( new_n63082_, new_n63081_, new_n63076_ );
nor  ( new_n63083_, new_n63081_, new_n63076_ );
xor  ( new_n63084_, new_n48756_, RIbb2d9f0_61 );
and  ( new_n63085_, new_n63084_, new_n9738_ );
xor  ( new_n63086_, new_n48908_, new_n9418_ );
nor  ( new_n63087_, new_n63086_, new_n10059_ );
nor  ( new_n63088_, new_n63087_, new_n63085_ );
not  ( new_n63089_, new_n63088_ );
and  ( new_n63090_, new_n62918_, new_n6508_ );
xor  ( new_n63091_, new_n51758_, new_n6163_ );
nor  ( new_n63092_, new_n63091_, new_n6645_ );
or   ( new_n63093_, new_n63092_, new_n63090_ );
nor  ( new_n63094_, new_n62887_, new_n5606_ );
nor  ( new_n63095_, new_n63051_, new_n5604_ );
or   ( new_n63096_, new_n63095_, new_n63094_ );
xor  ( new_n63097_, new_n62910_, new_n62904_ );
xor  ( new_n63098_, new_n63097_, new_n63096_ );
xor  ( new_n63099_, new_n63098_, new_n63093_ );
and  ( new_n63100_, new_n63099_, new_n63089_ );
xor  ( new_n63101_, new_n63099_, new_n63089_ );
and  ( new_n63102_, new_n48291_, RIbb2d888_64 );
nand ( new_n63103_, new_n63102_, RIbb2d900_63 );
or   ( new_n63104_, new_n63102_, RIbb2d900_63 );
or   ( new_n63105_, new_n48519_, RIbb2d888_64 );
and  ( new_n63106_, new_n63105_, new_n63104_ );
and  ( new_n63107_, new_n63106_, new_n63103_ );
and  ( new_n63108_, new_n63107_, new_n63101_ );
or   ( new_n63109_, new_n63108_, new_n63100_ );
xor  ( new_n63110_, new_n63006_, new_n63005_ );
and  ( new_n63111_, new_n63110_, new_n63109_ );
xor  ( new_n63112_, new_n63110_, new_n63109_ );
nor  ( new_n63113_, new_n62852_, new_n7734_ );
nor  ( new_n63114_, new_n63031_, new_n7732_ );
nor  ( new_n63115_, new_n63114_, new_n63113_ );
or   ( new_n63116_, new_n62856_, new_n7186_ );
or   ( new_n63117_, new_n63037_, new_n7184_ );
and  ( new_n63118_, new_n63117_, new_n63116_ );
xnor ( new_n63119_, new_n63118_, new_n63115_ );
and  ( new_n63120_, new_n62943_, new_n9738_ );
and  ( new_n63121_, new_n63084_, new_n9740_ );
nor  ( new_n63122_, new_n63121_, new_n63120_ );
xor  ( new_n63123_, new_n63122_, new_n63119_ );
and  ( new_n63124_, new_n63123_, new_n63112_ );
nor  ( new_n63125_, new_n63124_, new_n63111_ );
or   ( new_n63126_, new_n63125_, new_n63083_ );
and  ( new_n63127_, new_n63126_, new_n63082_ );
nor  ( new_n63128_, new_n63127_, new_n63026_ );
and  ( new_n63129_, new_n63127_, new_n63026_ );
nor  ( new_n63130_, new_n63118_, new_n63115_ );
and  ( new_n63131_, new_n63118_, new_n63115_ );
nor  ( new_n63132_, new_n63122_, new_n63131_ );
nor  ( new_n63133_, new_n63132_, new_n63130_ );
xnor ( new_n63134_, new_n62930_, new_n62929_ );
nor  ( new_n63135_, new_n63134_, new_n63133_ );
xnor ( new_n63136_, new_n63134_, new_n63133_ );
nor  ( new_n63137_, new_n62926_, new_n9424_ );
xor  ( new_n63138_, new_n49265_, new_n8870_ );
nor  ( new_n63139_, new_n63138_, new_n9422_ );
nor  ( new_n63140_, new_n63139_, new_n63137_ );
nand ( new_n63141_, new_n63097_, new_n63096_ );
nand ( new_n63142_, new_n63098_, new_n63093_ );
and  ( new_n63143_, new_n63142_, new_n63141_ );
or   ( new_n63144_, new_n63143_, new_n63140_ );
and  ( new_n63145_, new_n63143_, new_n63140_ );
or   ( new_n63146_, new_n48291_, new_n10052_ );
and  ( new_n63147_, new_n63146_, new_n10770_ );
and  ( new_n63148_, new_n48039_, RIbb2d888_64 );
or   ( new_n63149_, new_n63148_, new_n63147_ );
nand ( new_n63150_, new_n63148_, new_n10052_ );
and  ( new_n63151_, new_n63150_, new_n63149_ );
or   ( new_n63152_, new_n63151_, new_n63145_ );
and  ( new_n63153_, new_n63152_, new_n63144_ );
nor  ( new_n63154_, new_n63153_, new_n63136_ );
nor  ( new_n63155_, new_n63154_, new_n63135_ );
nor  ( new_n63156_, new_n63155_, new_n63129_ );
nor  ( new_n63157_, new_n63156_, new_n63128_ );
or   ( new_n63158_, new_n63157_, new_n63025_ );
and  ( new_n63159_, new_n63158_, new_n63024_ );
nor  ( new_n63160_, new_n63159_, new_n62995_ );
and  ( new_n63161_, new_n63159_, new_n62995_ );
xnor ( new_n63162_, new_n63019_, new_n63018_ );
xor  ( new_n63163_, new_n63012_, new_n63011_ );
xor  ( new_n63164_, new_n63153_, new_n63136_ );
nand ( new_n63165_, new_n63164_, new_n63163_ );
xor  ( new_n63166_, new_n63164_, new_n63163_ );
nor  ( new_n63167_, new_n53695_, new_n48671_ );
or   ( new_n63168_, new_n63167_, new_n5206_ );
or   ( new_n63169_, new_n63053_, new_n5606_ );
and  ( new_n63170_, new_n53694_, RIbb2e170_45 );
nor  ( new_n63171_, new_n53694_, RIbb2e170_45 );
or   ( new_n63172_, new_n63171_, new_n5604_ );
or   ( new_n63173_, new_n63172_, new_n63170_ );
and  ( new_n63174_, new_n63173_, new_n63169_ );
or   ( new_n63175_, new_n63174_, new_n63168_ );
or   ( new_n63176_, new_n63091_, new_n6647_ );
xor  ( new_n63177_, new_n52280_, new_n6163_ );
or   ( new_n63178_, new_n63177_, new_n6645_ );
and  ( new_n63179_, new_n63178_, new_n63176_ );
or   ( new_n63180_, new_n63179_, new_n63175_ );
and  ( new_n63181_, new_n63039_, new_n6908_ );
xor  ( new_n63182_, new_n51477_, RIbb2dea0_51 );
and  ( new_n63183_, new_n63182_, new_n6910_ );
or   ( new_n63184_, new_n63183_, new_n63181_ );
xor  ( new_n63185_, new_n63179_, new_n63175_ );
nand ( new_n63186_, new_n63185_, new_n63184_ );
and  ( new_n63187_, new_n63186_, new_n63180_ );
or   ( new_n63188_, new_n63138_, new_n9424_ );
xor  ( new_n63189_, new_n49427_, new_n8870_ );
or   ( new_n63190_, new_n63189_, new_n9422_ );
and  ( new_n63191_, new_n63190_, new_n63188_ );
nor  ( new_n63192_, new_n63191_, new_n63187_ );
xor  ( new_n63193_, new_n63071_, new_n63070_ );
xor  ( new_n63194_, new_n63191_, new_n63187_ );
and  ( new_n63195_, new_n63194_, new_n63193_ );
or   ( new_n63196_, new_n63195_, new_n63192_ );
xnor ( new_n63197_, new_n63143_, new_n63140_ );
xor  ( new_n63198_, new_n63197_, new_n63151_ );
or   ( new_n63199_, new_n63198_, new_n63196_ );
nand ( new_n63200_, new_n63198_, new_n63196_ );
xnor ( new_n63201_, new_n63035_, new_n63030_ );
nand ( new_n63202_, new_n63201_, new_n63041_ );
not  ( new_n63203_, new_n63036_ );
nand ( new_n63204_, new_n63043_, new_n63203_ );
and  ( new_n63205_, new_n63204_, new_n63202_ );
xnor ( new_n63206_, new_n63062_, new_n63061_ );
or   ( new_n63207_, new_n63067_, new_n8876_ );
xor  ( new_n63208_, new_n50115_, new_n8254_ );
or   ( new_n63209_, new_n63208_, new_n8874_ );
and  ( new_n63210_, new_n63209_, new_n63207_ );
nand ( new_n63211_, new_n63210_, new_n63206_ );
xor  ( new_n63212_, new_n50788_, new_n7722_ );
nor  ( new_n63213_, new_n63212_, new_n8264_ );
nor  ( new_n63214_, new_n63028_, new_n8266_ );
nor  ( new_n63215_, new_n63214_, new_n63213_ );
or   ( new_n63216_, new_n63210_, new_n63206_ );
nand ( new_n63217_, new_n63216_, new_n63215_ );
and  ( new_n63218_, new_n63217_, new_n63211_ );
and  ( new_n63219_, new_n63218_, new_n63205_ );
or   ( new_n63220_, new_n63189_, new_n9424_ );
xor  ( new_n63221_, new_n49488_, new_n8870_ );
or   ( new_n63222_, new_n63221_, new_n9422_ );
and  ( new_n63223_, new_n63222_, new_n63220_ );
or   ( new_n63224_, new_n63033_, new_n7734_ );
xor  ( new_n63225_, new_n51142_, new_n7174_ );
or   ( new_n63226_, new_n63225_, new_n7732_ );
and  ( new_n63227_, new_n63226_, new_n63224_ );
nor  ( new_n63228_, new_n63227_, new_n63223_ );
xor  ( new_n63229_, new_n49265_, new_n9418_ );
nor  ( new_n63230_, new_n63229_, new_n10059_ );
nor  ( new_n63231_, new_n63086_, new_n10061_ );
nor  ( new_n63232_, new_n63231_, new_n63230_ );
and  ( new_n63233_, new_n63227_, new_n63223_ );
nor  ( new_n63234_, new_n63233_, new_n63232_ );
nor  ( new_n63235_, new_n63234_, new_n63228_ );
not  ( new_n63236_, new_n63235_ );
xor  ( new_n63237_, new_n63218_, new_n63205_ );
and  ( new_n63238_, new_n63237_, new_n63236_ );
nor  ( new_n63239_, new_n63238_, new_n63219_ );
nand ( new_n63240_, new_n63239_, new_n63200_ );
and  ( new_n63241_, new_n63240_, new_n63199_ );
nand ( new_n63242_, new_n63241_, new_n63166_ );
and  ( new_n63243_, new_n63242_, new_n63165_ );
nor  ( new_n63244_, new_n63243_, new_n63162_ );
and  ( new_n63245_, new_n63243_, new_n63162_ );
xor  ( new_n63246_, new_n63127_, new_n63026_ );
xor  ( new_n63247_, new_n63246_, new_n63155_ );
nor  ( new_n63248_, new_n63247_, new_n63245_ );
nor  ( new_n63249_, new_n63248_, new_n63244_ );
not  ( new_n63250_, new_n63249_ );
xnor ( new_n63251_, new_n63023_, new_n63021_ );
xor  ( new_n63252_, new_n63251_, new_n63157_ );
and  ( new_n63253_, new_n63252_, new_n63250_ );
nor  ( new_n63254_, new_n63252_, new_n63250_ );
xor  ( new_n63255_, new_n63241_, new_n63166_ );
xnor ( new_n63256_, new_n63081_, new_n63076_ );
xor  ( new_n63257_, new_n63256_, new_n63125_ );
nor  ( new_n63258_, new_n63257_, new_n63255_ );
and  ( new_n63259_, new_n63257_, new_n63255_ );
xor  ( new_n63260_, new_n63074_, new_n63073_ );
xor  ( new_n63261_, new_n63123_, new_n63112_ );
nor  ( new_n63262_, new_n63261_, new_n63260_ );
and  ( new_n63263_, new_n63261_, new_n63260_ );
xnor ( new_n63264_, new_n63107_, new_n63101_ );
nor  ( new_n63265_, new_n63058_, new_n6175_ );
xor  ( new_n63266_, new_n52908_, RIbb2e080_47 );
nor  ( new_n63267_, new_n63266_, new_n6173_ );
or   ( new_n63268_, new_n63267_, new_n63265_ );
xor  ( new_n63269_, new_n63174_, new_n63168_ );
and  ( new_n63270_, new_n63269_, new_n63268_ );
nor  ( new_n63271_, new_n63177_, new_n6647_ );
xor  ( new_n63272_, new_n52293_, RIbb2df90_49 );
nor  ( new_n63273_, new_n63272_, new_n6645_ );
or   ( new_n63274_, new_n63273_, new_n63271_ );
xor  ( new_n63275_, new_n63269_, new_n63268_ );
and  ( new_n63276_, new_n63275_, new_n63274_ );
or   ( new_n63277_, new_n63276_, new_n63270_ );
xor  ( new_n63278_, new_n63185_, new_n63184_ );
nand ( new_n63279_, new_n63278_, new_n63277_ );
xor  ( new_n63280_, new_n63278_, new_n63277_ );
or   ( new_n63281_, new_n49271_, RIbb2d888_64 );
or   ( new_n63282_, new_n48519_, new_n10770_ );
and  ( new_n63283_, new_n48518_, RIbb2d888_64 );
or   ( new_n63284_, new_n63283_, RIbb2d900_63 );
and  ( new_n63285_, new_n63284_, new_n63282_ );
and  ( new_n63286_, new_n63285_, new_n63281_ );
nand ( new_n63287_, new_n63286_, new_n63280_ );
and  ( new_n63288_, new_n63287_, new_n63279_ );
and  ( new_n63289_, new_n63288_, new_n63264_ );
xor  ( new_n63290_, new_n63194_, new_n63193_ );
nor  ( new_n63291_, new_n63288_, new_n63264_ );
nor  ( new_n63292_, new_n63291_, new_n63290_ );
nor  ( new_n63293_, new_n63292_, new_n63289_ );
nor  ( new_n63294_, new_n63293_, new_n63263_ );
nor  ( new_n63295_, new_n63294_, new_n63262_ );
nor  ( new_n63296_, new_n63295_, new_n63259_ );
nor  ( new_n63297_, new_n63296_, new_n63258_ );
xnor ( new_n63298_, new_n63243_, new_n63162_ );
xor  ( new_n63299_, new_n63298_, new_n63247_ );
and  ( new_n63300_, new_n63299_, new_n63297_ );
nor  ( new_n63301_, new_n63299_, new_n63297_ );
xor  ( new_n63302_, new_n63257_, new_n63255_ );
xnor ( new_n63303_, new_n63302_, new_n63295_ );
xor  ( new_n63304_, new_n63237_, new_n63236_ );
not  ( new_n63305_, new_n63304_ );
nor  ( new_n63306_, new_n63266_, new_n6175_ );
xor  ( new_n63307_, new_n53306_, RIbb2e080_47 );
nor  ( new_n63308_, new_n63307_, new_n6173_ );
or   ( new_n63309_, new_n63308_, new_n63306_ );
and  ( new_n63310_, new_n53694_, new_n5371_ );
nand ( new_n63311_, new_n63310_, new_n63309_ );
nor  ( new_n63312_, new_n63272_, new_n6647_ );
xor  ( new_n63313_, new_n52902_, RIbb2df90_49 );
nor  ( new_n63314_, new_n63313_, new_n6645_ );
nor  ( new_n63315_, new_n63314_, new_n63312_ );
not  ( new_n63316_, new_n63315_ );
xor  ( new_n63317_, new_n63310_, new_n63309_ );
nand ( new_n63318_, new_n63317_, new_n63316_ );
and  ( new_n63319_, new_n63318_, new_n63311_ );
xor  ( new_n63320_, new_n51758_, new_n6635_ );
or   ( new_n63321_, new_n63320_, new_n7184_ );
nand ( new_n63322_, new_n63182_, new_n6908_ );
and  ( new_n63323_, new_n63322_, new_n63321_ );
or   ( new_n63324_, new_n63323_, new_n63319_ );
xor  ( new_n63325_, new_n50487_, new_n8254_ );
nor  ( new_n63326_, new_n63325_, new_n8874_ );
nor  ( new_n63327_, new_n63208_, new_n8876_ );
nor  ( new_n63328_, new_n63327_, new_n63326_ );
not  ( new_n63329_, new_n63328_ );
xor  ( new_n63330_, new_n63323_, new_n63319_ );
nand ( new_n63331_, new_n63330_, new_n63329_ );
and  ( new_n63332_, new_n63331_, new_n63324_ );
xor  ( new_n63333_, new_n49758_, new_n8870_ );
or   ( new_n63334_, new_n63333_, new_n9422_ );
or   ( new_n63335_, new_n63221_, new_n9424_ );
and  ( new_n63336_, new_n63335_, new_n63334_ );
or   ( new_n63337_, new_n63212_, new_n8266_ );
xor  ( new_n63338_, new_n50894_, new_n7722_ );
or   ( new_n63339_, new_n63338_, new_n8264_ );
and  ( new_n63340_, new_n63339_, new_n63337_ );
or   ( new_n63341_, new_n63340_, new_n63336_ );
nor  ( new_n63342_, new_n63225_, new_n7734_ );
xor  ( new_n63343_, new_n51446_, RIbb2ddb0_53 );
and  ( new_n63344_, new_n63343_, new_n7489_ );
nor  ( new_n63345_, new_n63344_, new_n63342_ );
and  ( new_n63346_, new_n63340_, new_n63336_ );
or   ( new_n63347_, new_n63346_, new_n63345_ );
and  ( new_n63348_, new_n63347_, new_n63341_ );
or   ( new_n63349_, new_n63348_, new_n63332_ );
and  ( new_n63350_, new_n63348_, new_n63332_ );
xor  ( new_n63351_, new_n63210_, new_n63206_ );
xor  ( new_n63352_, new_n63351_, new_n63215_ );
or   ( new_n63353_, new_n63352_, new_n63350_ );
and  ( new_n63354_, new_n63353_, new_n63349_ );
or   ( new_n63355_, new_n63354_, new_n63305_ );
xor  ( new_n63356_, new_n63354_, new_n63305_ );
nor  ( new_n63357_, new_n53695_, new_n49294_ );
or   ( new_n63358_, new_n63357_, new_n5597_ );
or   ( new_n63359_, new_n63307_, new_n6175_ );
and  ( new_n63360_, new_n53694_, RIbb2e080_47 );
nor  ( new_n63361_, new_n53694_, RIbb2e080_47 );
or   ( new_n63362_, new_n63361_, new_n6173_ );
or   ( new_n63363_, new_n63362_, new_n63360_ );
and  ( new_n63364_, new_n63363_, new_n63359_ );
or   ( new_n63365_, new_n63364_, new_n63358_ );
or   ( new_n63366_, new_n63320_, new_n7186_ );
xor  ( new_n63367_, new_n52280_, new_n6635_ );
or   ( new_n63368_, new_n63367_, new_n7184_ );
and  ( new_n63369_, new_n63368_, new_n63366_ );
nor  ( new_n63370_, new_n63369_, new_n63365_ );
xor  ( new_n63371_, new_n51477_, RIbb2ddb0_53 );
and  ( new_n63372_, new_n63371_, new_n7489_ );
and  ( new_n63373_, new_n63343_, new_n7487_ );
or   ( new_n63374_, new_n63373_, new_n63372_ );
xor  ( new_n63375_, new_n63369_, new_n63365_ );
and  ( new_n63376_, new_n63375_, new_n63374_ );
or   ( new_n63377_, new_n63376_, new_n63370_ );
xor  ( new_n63378_, new_n63275_, new_n63274_ );
and  ( new_n63379_, new_n63378_, new_n63377_ );
nor  ( new_n63380_, new_n63229_, new_n10061_ );
xor  ( new_n63381_, new_n49427_, RIbb2d9f0_61 );
and  ( new_n63382_, new_n63381_, new_n9740_ );
nor  ( new_n63383_, new_n63382_, new_n63380_ );
not  ( new_n63384_, new_n63383_ );
xor  ( new_n63385_, new_n63378_, new_n63377_ );
and  ( new_n63386_, new_n63385_, new_n63384_ );
or   ( new_n63387_, new_n63386_, new_n63379_ );
xnor ( new_n63388_, new_n63227_, new_n63223_ );
nand ( new_n63389_, new_n63388_, new_n63232_ );
not  ( new_n63390_, new_n63234_ );
or   ( new_n63391_, new_n63390_, new_n63228_ );
and  ( new_n63392_, new_n63391_, new_n63389_ );
or   ( new_n63393_, new_n63392_, new_n63387_ );
and  ( new_n63394_, new_n63392_, new_n63387_ );
xor  ( new_n63395_, new_n63286_, new_n63280_ );
or   ( new_n63396_, new_n63395_, new_n63394_ );
and  ( new_n63397_, new_n63396_, new_n63393_ );
nand ( new_n63398_, new_n63397_, new_n63356_ );
and  ( new_n63399_, new_n63398_, new_n63355_ );
xor  ( new_n63400_, new_n63198_, new_n63196_ );
xor  ( new_n63401_, new_n63400_, new_n63239_ );
or   ( new_n63402_, new_n63401_, new_n63399_ );
and  ( new_n63403_, new_n63401_, new_n63399_ );
xor  ( new_n63404_, new_n63261_, new_n63260_ );
xnor ( new_n63405_, new_n63404_, new_n63293_ );
or   ( new_n63406_, new_n63405_, new_n63403_ );
and  ( new_n63407_, new_n63406_, new_n63402_ );
nor  ( new_n63408_, new_n63407_, new_n63303_ );
and  ( new_n63409_, new_n63407_, new_n63303_ );
xnor ( new_n63410_, new_n63288_, new_n63264_ );
xor  ( new_n63411_, new_n63410_, new_n63290_ );
xor  ( new_n63412_, new_n63330_, new_n63329_ );
not  ( new_n63413_, new_n63412_ );
xor  ( new_n63414_, new_n50788_, new_n8254_ );
or   ( new_n63415_, new_n63414_, new_n8874_ );
or   ( new_n63416_, new_n63325_, new_n8876_ );
and  ( new_n63417_, new_n63416_, new_n63415_ );
xor  ( new_n63418_, new_n51142_, new_n7722_ );
or   ( new_n63419_, new_n63418_, new_n8264_ );
or   ( new_n63420_, new_n63338_, new_n8266_ );
and  ( new_n63421_, new_n63420_, new_n63419_ );
or   ( new_n63422_, new_n63421_, new_n63417_ );
nand ( new_n63423_, new_n63421_, new_n63417_ );
xor  ( new_n63424_, new_n63317_, new_n63316_ );
nand ( new_n63425_, new_n63424_, new_n63423_ );
and  ( new_n63426_, new_n63425_, new_n63422_ );
nor  ( new_n63427_, new_n63426_, new_n63413_ );
xor  ( new_n63428_, new_n63426_, new_n63413_ );
not  ( new_n63429_, new_n63428_ );
or   ( new_n63430_, new_n48908_, new_n10052_ );
and  ( new_n63431_, new_n63430_, new_n10770_ );
and  ( new_n63432_, new_n48756_, RIbb2d888_64 );
or   ( new_n63433_, new_n63432_, new_n63431_ );
nand ( new_n63434_, new_n63432_, new_n10052_ );
and  ( new_n63435_, new_n63434_, new_n63433_ );
nor  ( new_n63436_, new_n63435_, new_n63429_ );
or   ( new_n63437_, new_n63436_, new_n63427_ );
xnor ( new_n63438_, new_n63348_, new_n63332_ );
xor  ( new_n63439_, new_n63438_, new_n63352_ );
nand ( new_n63440_, new_n63439_, new_n63437_ );
nor  ( new_n63441_, new_n63439_, new_n63437_ );
nor  ( new_n63442_, new_n63333_, new_n9424_ );
xor  ( new_n63443_, new_n50115_, new_n8870_ );
nor  ( new_n63444_, new_n63443_, new_n9422_ );
nor  ( new_n63445_, new_n63444_, new_n63442_ );
nand ( new_n63446_, new_n63381_, new_n9738_ );
xor  ( new_n63447_, new_n49488_, new_n9418_ );
or   ( new_n63448_, new_n63447_, new_n10059_ );
and  ( new_n63449_, new_n63448_, new_n63446_ );
nor  ( new_n63450_, new_n63449_, new_n63445_ );
xor  ( new_n63451_, new_n63449_, new_n63445_ );
xor  ( new_n63452_, new_n48908_, new_n10052_ );
or   ( new_n63453_, new_n63452_, new_n21077_ );
or   ( new_n63454_, new_n49265_, new_n10052_ );
or   ( new_n63455_, new_n63454_, new_n10769_ );
nand ( new_n63456_, new_n63455_, new_n63453_ );
and  ( new_n63457_, new_n63456_, new_n63451_ );
or   ( new_n63458_, new_n63457_, new_n63450_ );
xnor ( new_n63459_, new_n63340_, new_n63336_ );
xor  ( new_n63460_, new_n63459_, new_n63345_ );
and  ( new_n63461_, new_n63460_, new_n63458_ );
nor  ( new_n63462_, new_n63460_, new_n63458_ );
not  ( new_n63463_, new_n63462_ );
xor  ( new_n63464_, new_n63385_, new_n63384_ );
and  ( new_n63465_, new_n63464_, new_n63463_ );
nor  ( new_n63466_, new_n63465_, new_n63461_ );
or   ( new_n63467_, new_n63466_, new_n63441_ );
and  ( new_n63468_, new_n63467_, new_n63440_ );
and  ( new_n63469_, new_n63468_, new_n63411_ );
nor  ( new_n63470_, new_n63468_, new_n63411_ );
xor  ( new_n63471_, new_n63397_, new_n63356_ );
nor  ( new_n63472_, new_n63471_, new_n63470_ );
nor  ( new_n63473_, new_n63472_, new_n63469_ );
xnor ( new_n63474_, new_n63401_, new_n63399_ );
xor  ( new_n63475_, new_n63474_, new_n63405_ );
nor  ( new_n63476_, new_n63475_, new_n63473_ );
and  ( new_n63477_, new_n63475_, new_n63473_ );
xnor ( new_n63478_, new_n63439_, new_n63437_ );
xor  ( new_n63479_, new_n63478_, new_n63466_ );
xor  ( new_n63480_, new_n63392_, new_n63387_ );
xor  ( new_n63481_, new_n63480_, new_n63395_ );
nor  ( new_n63482_, new_n63481_, new_n63479_ );
and  ( new_n63483_, new_n63481_, new_n63479_ );
xnor ( new_n63484_, new_n63456_, new_n63451_ );
xor  ( new_n63485_, new_n50487_, new_n8870_ );
or   ( new_n63486_, new_n63485_, new_n9422_ );
or   ( new_n63487_, new_n63443_, new_n9424_ );
and  ( new_n63488_, new_n63487_, new_n63486_ );
xor  ( new_n63489_, new_n49758_, new_n9418_ );
or   ( new_n63490_, new_n63489_, new_n10059_ );
or   ( new_n63491_, new_n63447_, new_n10061_ );
and  ( new_n63492_, new_n63491_, new_n63490_ );
or   ( new_n63493_, new_n63492_, new_n63488_ );
nor  ( new_n63494_, new_n63418_, new_n8266_ );
xor  ( new_n63495_, new_n51446_, RIbb2dcc0_55 );
and  ( new_n63496_, new_n63495_, new_n8042_ );
nor  ( new_n63497_, new_n63496_, new_n63494_ );
and  ( new_n63498_, new_n63492_, new_n63488_ );
or   ( new_n63499_, new_n63498_, new_n63497_ );
and  ( new_n63500_, new_n63499_, new_n63493_ );
or   ( new_n63501_, new_n63500_, new_n63484_ );
nor  ( new_n63502_, new_n53695_, new_n49685_ );
or   ( new_n63503_, new_n63502_, new_n6166_ );
xor  ( new_n63504_, new_n53306_, RIbb2df90_49 );
or   ( new_n63505_, new_n63504_, new_n6647_ );
and  ( new_n63506_, new_n49684_, RIbb2df90_49 );
and  ( new_n63507_, new_n53694_, RIbb2dea0_51 );
nor  ( new_n63508_, new_n63507_, new_n63506_ );
and  ( new_n63509_, RIbb2df18_50, new_n6163_ );
nor  ( new_n63510_, new_n53694_, RIbb2dea0_51 );
nor  ( new_n63511_, new_n63510_, new_n63509_ );
or   ( new_n63512_, new_n63511_, new_n63508_ );
and  ( new_n63513_, new_n63512_, new_n63505_ );
or   ( new_n63514_, new_n63513_, new_n63503_ );
xor  ( new_n63515_, new_n52280_, new_n7174_ );
or   ( new_n63516_, new_n63515_, new_n7732_ );
xor  ( new_n63517_, new_n51758_, new_n7174_ );
or   ( new_n63518_, new_n63517_, new_n7734_ );
and  ( new_n63519_, new_n63518_, new_n63516_ );
nor  ( new_n63520_, new_n63519_, new_n63514_ );
and  ( new_n63521_, new_n63495_, new_n8040_ );
xor  ( new_n63522_, new_n51477_, RIbb2dcc0_55 );
and  ( new_n63523_, new_n63522_, new_n8042_ );
nor  ( new_n63524_, new_n63523_, new_n63521_ );
xnor ( new_n63525_, new_n63519_, new_n63514_ );
nor  ( new_n63526_, new_n63525_, new_n63524_ );
nor  ( new_n63527_, new_n63526_, new_n63520_ );
and  ( new_n63528_, new_n63371_, new_n7487_ );
nor  ( new_n63529_, new_n63517_, new_n7732_ );
or   ( new_n63530_, new_n63529_, new_n63528_ );
nor  ( new_n63531_, new_n63313_, new_n6647_ );
xor  ( new_n63532_, new_n52908_, RIbb2df90_49 );
nor  ( new_n63533_, new_n63532_, new_n6645_ );
or   ( new_n63534_, new_n63533_, new_n63531_ );
xor  ( new_n63535_, new_n63364_, new_n63358_ );
xor  ( new_n63536_, new_n63535_, new_n63534_ );
xnor ( new_n63537_, new_n63536_, new_n63530_ );
or   ( new_n63538_, new_n63537_, new_n63527_ );
xnor ( new_n63539_, new_n63537_, new_n63527_ );
xor  ( new_n63540_, new_n49265_, new_n10052_ );
or   ( new_n63541_, new_n63540_, new_n21077_ );
or   ( new_n63542_, new_n61553_, new_n49427_ );
and  ( new_n63543_, new_n63542_, new_n63541_ );
or   ( new_n63544_, new_n63543_, new_n63539_ );
and  ( new_n63545_, new_n63544_, new_n63538_ );
and  ( new_n63546_, new_n63500_, new_n63484_ );
or   ( new_n63547_, new_n63546_, new_n63545_ );
and  ( new_n63548_, new_n63547_, new_n63501_ );
and  ( new_n63549_, new_n63535_, new_n63534_ );
and  ( new_n63550_, new_n63536_, new_n63530_ );
or   ( new_n63551_, new_n63550_, new_n63549_ );
xor  ( new_n63552_, new_n63375_, new_n63374_ );
nand ( new_n63553_, new_n63552_, new_n63551_ );
or   ( new_n63554_, new_n63367_, new_n7186_ );
xor  ( new_n63555_, new_n52293_, RIbb2dea0_51 );
or   ( new_n63556_, new_n63555_, new_n7184_ );
and  ( new_n63557_, new_n63556_, new_n63554_ );
nor  ( new_n63558_, new_n63504_, new_n6645_ );
nor  ( new_n63559_, new_n63532_, new_n6647_ );
or   ( new_n63560_, new_n63559_, new_n63558_ );
and  ( new_n63561_, new_n53694_, new_n5915_ );
nand ( new_n63562_, new_n63561_, new_n63560_ );
xor  ( new_n63563_, new_n52902_, RIbb2dea0_51 );
nor  ( new_n63564_, new_n63563_, new_n7184_ );
nor  ( new_n63565_, new_n63555_, new_n7186_ );
or   ( new_n63566_, new_n63565_, new_n63564_ );
xor  ( new_n63567_, new_n63561_, new_n63560_ );
nand ( new_n63568_, new_n63567_, new_n63566_ );
and  ( new_n63569_, new_n63568_, new_n63562_ );
nor  ( new_n63570_, new_n63569_, new_n63557_ );
nor  ( new_n63571_, new_n63414_, new_n8876_ );
xor  ( new_n63572_, new_n50894_, new_n8254_ );
nor  ( new_n63573_, new_n63572_, new_n8874_ );
or   ( new_n63574_, new_n63573_, new_n63571_ );
xor  ( new_n63575_, new_n63569_, new_n63557_ );
and  ( new_n63576_, new_n63575_, new_n63574_ );
or   ( new_n63577_, new_n63576_, new_n63570_ );
xor  ( new_n63578_, new_n63552_, new_n63551_ );
nand ( new_n63579_, new_n63578_, new_n63577_ );
and  ( new_n63580_, new_n63579_, new_n63553_ );
and  ( new_n63581_, new_n63580_, new_n63548_ );
nor  ( new_n63582_, new_n63580_, new_n63548_ );
xor  ( new_n63583_, new_n63435_, new_n63429_ );
nor  ( new_n63584_, new_n63583_, new_n63582_ );
nor  ( new_n63585_, new_n63584_, new_n63581_ );
nor  ( new_n63586_, new_n63585_, new_n63483_ );
nor  ( new_n63587_, new_n63586_, new_n63482_ );
xor  ( new_n63588_, new_n63468_, new_n63411_ );
xor  ( new_n63589_, new_n63588_, new_n63471_ );
nor  ( new_n63590_, new_n63589_, new_n63587_ );
and  ( new_n63591_, new_n63589_, new_n63587_ );
xor  ( new_n63592_, new_n63578_, new_n63577_ );
xor  ( new_n63593_, new_n63421_, new_n63417_ );
xor  ( new_n63594_, new_n63593_, new_n63424_ );
nor  ( new_n63595_, new_n63594_, new_n63592_ );
and  ( new_n63596_, new_n63594_, new_n63592_ );
not  ( new_n63597_, new_n63596_ );
nor  ( new_n63598_, new_n63563_, new_n7186_ );
xor  ( new_n63599_, new_n52908_, RIbb2dea0_51 );
nor  ( new_n63600_, new_n63599_, new_n7184_ );
or   ( new_n63601_, new_n63600_, new_n63598_ );
xor  ( new_n63602_, new_n63513_, new_n63503_ );
nand ( new_n63603_, new_n63602_, new_n63601_ );
nor  ( new_n63604_, new_n63515_, new_n7734_ );
xor  ( new_n63605_, new_n52293_, RIbb2ddb0_53 );
nor  ( new_n63606_, new_n63605_, new_n7732_ );
or   ( new_n63607_, new_n63606_, new_n63604_ );
xor  ( new_n63608_, new_n63602_, new_n63601_ );
nand ( new_n63609_, new_n63608_, new_n63607_ );
and  ( new_n63610_, new_n63609_, new_n63603_ );
xor  ( new_n63611_, new_n50788_, new_n8870_ );
or   ( new_n63612_, new_n63611_, new_n9422_ );
or   ( new_n63613_, new_n63485_, new_n9424_ );
and  ( new_n63614_, new_n63613_, new_n63612_ );
nor  ( new_n63615_, new_n63614_, new_n63610_ );
nor  ( new_n63616_, new_n63489_, new_n10061_ );
xor  ( new_n63617_, new_n50115_, new_n9418_ );
nor  ( new_n63618_, new_n63617_, new_n10059_ );
or   ( new_n63619_, new_n63618_, new_n63616_ );
xor  ( new_n63620_, new_n63614_, new_n63610_ );
and  ( new_n63621_, new_n63620_, new_n63619_ );
or   ( new_n63622_, new_n63621_, new_n63615_ );
xor  ( new_n63623_, new_n63575_, new_n63574_ );
and  ( new_n63624_, new_n63623_, new_n63622_ );
xor  ( new_n63625_, new_n51142_, new_n8254_ );
nor  ( new_n63626_, new_n63625_, new_n8874_ );
nor  ( new_n63627_, new_n63572_, new_n8876_ );
or   ( new_n63628_, new_n63627_, new_n63626_ );
xor  ( new_n63629_, new_n63567_, new_n63566_ );
and  ( new_n63630_, new_n63629_, new_n63628_ );
xor  ( new_n63631_, new_n63629_, new_n63628_ );
or   ( new_n63632_, new_n49979_, RIbb2d888_64 );
and  ( new_n63633_, new_n49427_, RIbb2d888_64 );
xor  ( new_n63634_, new_n63633_, RIbb2d900_63 );
and  ( new_n63635_, new_n63634_, new_n63632_ );
and  ( new_n63636_, new_n63635_, new_n63631_ );
nor  ( new_n63637_, new_n63636_, new_n63630_ );
xnor ( new_n63638_, new_n63623_, new_n63622_ );
nor  ( new_n63639_, new_n63638_, new_n63637_ );
nor  ( new_n63640_, new_n63639_, new_n63624_ );
and  ( new_n63641_, new_n63640_, new_n63597_ );
nor  ( new_n63642_, new_n63641_, new_n63595_ );
xor  ( new_n63643_, new_n63460_, new_n63458_ );
xor  ( new_n63644_, new_n63643_, new_n63464_ );
nor  ( new_n63645_, new_n63644_, new_n63642_ );
xnor ( new_n63646_, new_n63644_, new_n63642_ );
xor  ( new_n63647_, new_n63580_, new_n63548_ );
xor  ( new_n63648_, new_n63647_, new_n63583_ );
nor  ( new_n63649_, new_n63648_, new_n63646_ );
nor  ( new_n63650_, new_n63649_, new_n63645_ );
not  ( new_n63651_, new_n63650_ );
xnor ( new_n63652_, new_n63481_, new_n63479_ );
xor  ( new_n63653_, new_n63652_, new_n63585_ );
and  ( new_n63654_, new_n63653_, new_n63651_ );
nor  ( new_n63655_, new_n63653_, new_n63651_ );
xnor ( new_n63656_, new_n63492_, new_n63488_ );
xor  ( new_n63657_, new_n63656_, new_n63497_ );
xor  ( new_n63658_, new_n63543_, new_n63539_ );
and  ( new_n63659_, new_n63658_, new_n63657_ );
xnor ( new_n63660_, new_n63525_, new_n63524_ );
or   ( new_n63661_, new_n63617_, new_n10061_ );
xor  ( new_n63662_, new_n50487_, new_n9418_ );
or   ( new_n63663_, new_n63662_, new_n10059_ );
and  ( new_n63664_, new_n63663_, new_n63661_ );
xor  ( new_n63665_, new_n50894_, new_n8870_ );
or   ( new_n63666_, new_n63665_, new_n9422_ );
or   ( new_n63667_, new_n63611_, new_n9424_ );
and  ( new_n63668_, new_n63667_, new_n63666_ );
or   ( new_n63669_, new_n63668_, new_n63664_ );
and  ( new_n63670_, new_n63668_, new_n63664_ );
nor  ( new_n63671_, new_n49758_, new_n10052_ );
nor  ( new_n63672_, new_n63671_, new_n10769_ );
and  ( new_n63673_, new_n49488_, RIbb2d888_64 );
nor  ( new_n63674_, new_n63673_, new_n63672_ );
and  ( new_n63675_, new_n63673_, new_n10052_ );
nor  ( new_n63676_, new_n63675_, new_n63674_ );
or   ( new_n63677_, new_n63676_, new_n63670_ );
and  ( new_n63678_, new_n63677_, new_n63669_ );
and  ( new_n63679_, new_n63678_, new_n63660_ );
or   ( new_n63680_, new_n63625_, new_n8876_ );
xor  ( new_n63681_, new_n51446_, RIbb2dbd0_57 );
nand ( new_n63682_, new_n63681_, new_n8651_ );
and  ( new_n63683_, new_n63682_, new_n63680_ );
xor  ( new_n63684_, new_n51758_, new_n7722_ );
or   ( new_n63685_, new_n63684_, new_n8264_ );
nand ( new_n63686_, new_n63522_, new_n8040_ );
and  ( new_n63687_, new_n63686_, new_n63685_ );
nor  ( new_n63688_, new_n63687_, new_n63683_ );
xor  ( new_n63689_, new_n53306_, RIbb2dea0_51 );
nor  ( new_n63690_, new_n63689_, new_n7184_ );
nor  ( new_n63691_, new_n63599_, new_n7186_ );
or   ( new_n63692_, new_n63691_, new_n63690_ );
and  ( new_n63693_, new_n53694_, new_n6508_ );
and  ( new_n63694_, new_n63693_, new_n63692_ );
nor  ( new_n63695_, new_n63605_, new_n7734_ );
xor  ( new_n63696_, new_n52902_, RIbb2ddb0_53 );
nor  ( new_n63697_, new_n63696_, new_n7732_ );
or   ( new_n63698_, new_n63697_, new_n63695_ );
xor  ( new_n63699_, new_n63693_, new_n63692_ );
and  ( new_n63700_, new_n63699_, new_n63698_ );
nor  ( new_n63701_, new_n63700_, new_n63694_ );
and  ( new_n63702_, new_n63687_, new_n63683_ );
nor  ( new_n63703_, new_n63702_, new_n63701_ );
nor  ( new_n63704_, new_n63703_, new_n63688_ );
nor  ( new_n63705_, new_n63704_, new_n63679_ );
nor  ( new_n63706_, new_n63678_, new_n63660_ );
nor  ( new_n63707_, new_n63706_, new_n63705_ );
not  ( new_n63708_, new_n63707_ );
xor  ( new_n63709_, new_n63658_, new_n63657_ );
and  ( new_n63710_, new_n63709_, new_n63708_ );
nor  ( new_n63711_, new_n63710_, new_n63659_ );
xor  ( new_n63712_, new_n63500_, new_n63484_ );
xor  ( new_n63713_, new_n63712_, new_n63545_ );
and  ( new_n63714_, new_n63713_, new_n63711_ );
xor  ( new_n63715_, new_n63713_, new_n63711_ );
xor  ( new_n63716_, new_n63594_, new_n63592_ );
xor  ( new_n63717_, new_n63716_, new_n63640_ );
and  ( new_n63718_, new_n63717_, new_n63715_ );
nor  ( new_n63719_, new_n63718_, new_n63714_ );
not  ( new_n63720_, new_n63719_ );
xor  ( new_n63721_, new_n63648_, new_n63646_ );
and  ( new_n63722_, new_n63721_, new_n63720_ );
nor  ( new_n63723_, new_n63721_, new_n63720_ );
xor  ( new_n63724_, new_n63717_, new_n63715_ );
xnor ( new_n63725_, new_n63638_, new_n63637_ );
xor  ( new_n63726_, new_n63620_, new_n63619_ );
xor  ( new_n63727_, new_n63635_, new_n63631_ );
nand ( new_n63728_, new_n63727_, new_n63726_ );
nor  ( new_n63729_, new_n63727_, new_n63726_ );
and  ( new_n63730_, new_n53694_, new_n50306_ );
or   ( new_n63731_, new_n63730_, new_n6638_ );
or   ( new_n63732_, new_n63689_, new_n7186_ );
or   ( new_n63733_, new_n63507_, new_n7184_ );
or   ( new_n63734_, new_n63733_, new_n63510_ );
and  ( new_n63735_, new_n63734_, new_n63732_ );
or   ( new_n63736_, new_n63735_, new_n63731_ );
or   ( new_n63737_, new_n63684_, new_n8266_ );
xor  ( new_n63738_, new_n52280_, new_n7722_ );
or   ( new_n63739_, new_n63738_, new_n8264_ );
and  ( new_n63740_, new_n63739_, new_n63737_ );
nor  ( new_n63741_, new_n63740_, new_n63736_ );
and  ( new_n63742_, new_n63681_, new_n8649_ );
xor  ( new_n63743_, new_n51477_, RIbb2dbd0_57 );
and  ( new_n63744_, new_n63743_, new_n8651_ );
or   ( new_n63745_, new_n63744_, new_n63742_ );
xor  ( new_n63746_, new_n63740_, new_n63736_ );
and  ( new_n63747_, new_n63746_, new_n63745_ );
or   ( new_n63748_, new_n63747_, new_n63741_ );
xor  ( new_n63749_, new_n63608_, new_n63607_ );
and  ( new_n63750_, new_n63749_, new_n63748_ );
nor  ( new_n63751_, new_n63749_, new_n63748_ );
xor  ( new_n63752_, new_n50788_, new_n9418_ );
nor  ( new_n63753_, new_n63752_, new_n10059_ );
nor  ( new_n63754_, new_n63662_, new_n10061_ );
or   ( new_n63755_, new_n63754_, new_n63753_ );
xor  ( new_n63756_, new_n63699_, new_n63698_ );
and  ( new_n63757_, new_n63756_, new_n63755_ );
nor  ( new_n63758_, new_n63665_, new_n9424_ );
xor  ( new_n63759_, new_n51142_, new_n8870_ );
nor  ( new_n63760_, new_n63759_, new_n9422_ );
or   ( new_n63761_, new_n63760_, new_n63758_ );
xor  ( new_n63762_, new_n63756_, new_n63755_ );
and  ( new_n63763_, new_n63762_, new_n63761_ );
nor  ( new_n63764_, new_n63763_, new_n63757_ );
nor  ( new_n63765_, new_n63764_, new_n63751_ );
nor  ( new_n63766_, new_n63765_, new_n63750_ );
or   ( new_n63767_, new_n63766_, new_n63729_ );
and  ( new_n63768_, new_n63767_, new_n63728_ );
or   ( new_n63769_, new_n63768_, new_n63725_ );
xor  ( new_n63770_, new_n63709_, new_n63708_ );
nand ( new_n63771_, new_n63768_, new_n63725_ );
nand ( new_n63772_, new_n63771_, new_n63770_ );
and  ( new_n63773_, new_n63772_, new_n63769_ );
and  ( new_n63774_, new_n63773_, new_n63724_ );
nor  ( new_n63775_, new_n63773_, new_n63724_ );
nor  ( new_n63776_, new_n63696_, new_n7734_ );
xor  ( new_n63777_, new_n52908_, RIbb2ddb0_53 );
nor  ( new_n63778_, new_n63777_, new_n7732_ );
or   ( new_n63779_, new_n63778_, new_n63776_ );
xor  ( new_n63780_, new_n63735_, new_n63731_ );
nand ( new_n63781_, new_n63780_, new_n63779_ );
nor  ( new_n63782_, new_n63738_, new_n8266_ );
xor  ( new_n63783_, new_n52293_, RIbb2dcc0_55 );
nor  ( new_n63784_, new_n63783_, new_n8264_ );
nor  ( new_n63785_, new_n63784_, new_n63782_ );
xnor ( new_n63786_, new_n63780_, new_n63779_ );
or   ( new_n63787_, new_n63786_, new_n63785_ );
and  ( new_n63788_, new_n63787_, new_n63781_ );
xor  ( new_n63789_, new_n49758_, new_n10052_ );
or   ( new_n63790_, new_n63789_, new_n21077_ );
or   ( new_n63791_, new_n50115_, new_n10052_ );
or   ( new_n63792_, new_n63791_, new_n10769_ );
and  ( new_n63793_, new_n63792_, new_n63790_ );
nor  ( new_n63794_, new_n63793_, new_n63788_ );
xor  ( new_n63795_, new_n63793_, new_n63788_ );
xor  ( new_n63796_, new_n63746_, new_n63745_ );
and  ( new_n63797_, new_n63796_, new_n63795_ );
nor  ( new_n63798_, new_n63797_, new_n63794_ );
not  ( new_n63799_, new_n63798_ );
xnor ( new_n63800_, new_n63687_, new_n63683_ );
xor  ( new_n63801_, new_n63800_, new_n63701_ );
nor  ( new_n63802_, new_n63801_, new_n63799_ );
xor  ( new_n63803_, new_n63801_, new_n63799_ );
xnor ( new_n63804_, new_n63668_, new_n63664_ );
xnor ( new_n63805_, new_n63804_, new_n63676_ );
and  ( new_n63806_, new_n63805_, new_n63803_ );
nor  ( new_n63807_, new_n63806_, new_n63802_ );
xnor ( new_n63808_, new_n63678_, new_n63660_ );
xor  ( new_n63809_, new_n63808_, new_n63704_ );
nor  ( new_n63810_, new_n63809_, new_n63807_ );
xor  ( new_n63811_, new_n63809_, new_n63807_ );
not  ( new_n63812_, new_n63811_ );
xnor ( new_n63813_, new_n63727_, new_n63726_ );
xor  ( new_n63814_, new_n63813_, new_n63766_ );
nor  ( new_n63815_, new_n63814_, new_n63812_ );
nor  ( new_n63816_, new_n63815_, new_n63810_ );
xor  ( new_n63817_, new_n63768_, new_n63725_ );
xor  ( new_n63818_, new_n63817_, new_n63770_ );
nor  ( new_n63819_, new_n63818_, new_n63816_ );
and  ( new_n63820_, new_n63818_, new_n63816_ );
xor  ( new_n63821_, new_n63814_, new_n63812_ );
not  ( new_n63822_, new_n63821_ );
xnor ( new_n63823_, new_n63805_, new_n63803_ );
xnor ( new_n63824_, new_n63749_, new_n63748_ );
xor  ( new_n63825_, new_n63824_, new_n63764_ );
or   ( new_n63826_, new_n63825_, new_n63823_ );
nand ( new_n63827_, new_n63825_, new_n63823_ );
nand ( new_n63828_, new_n63743_, new_n8649_ );
xor  ( new_n63829_, new_n51758_, new_n8254_ );
or   ( new_n63830_, new_n63829_, new_n8874_ );
and  ( new_n63831_, new_n63830_, new_n63828_ );
nor  ( new_n63832_, new_n63777_, new_n7734_ );
xor  ( new_n63833_, new_n53306_, RIbb2ddb0_53 );
nor  ( new_n63834_, new_n63833_, new_n7732_ );
or   ( new_n63835_, new_n63834_, new_n63832_ );
and  ( new_n63836_, new_n53694_, new_n6908_ );
nand ( new_n63837_, new_n63836_, new_n63835_ );
nor  ( new_n63838_, new_n63783_, new_n8266_ );
xor  ( new_n63839_, new_n52902_, RIbb2dcc0_55 );
nor  ( new_n63840_, new_n63839_, new_n8264_ );
nor  ( new_n63841_, new_n63840_, new_n63838_ );
xnor ( new_n63842_, new_n63836_, new_n63835_ );
or   ( new_n63843_, new_n63842_, new_n63841_ );
and  ( new_n63844_, new_n63843_, new_n63837_ );
nor  ( new_n63845_, new_n63844_, new_n63831_ );
nor  ( new_n63846_, new_n63752_, new_n10061_ );
xor  ( new_n63847_, new_n50894_, new_n9418_ );
nor  ( new_n63848_, new_n63847_, new_n10059_ );
or   ( new_n63849_, new_n63848_, new_n63846_ );
xor  ( new_n63850_, new_n63844_, new_n63831_ );
and  ( new_n63851_, new_n63850_, new_n63849_ );
or   ( new_n63852_, new_n63851_, new_n63845_ );
xor  ( new_n63853_, new_n63762_, new_n63761_ );
and  ( new_n63854_, new_n63853_, new_n63852_ );
xnor ( new_n63855_, new_n63786_, new_n63785_ );
xor  ( new_n63856_, new_n50115_, new_n10052_ );
or   ( new_n63857_, new_n63856_, new_n21077_ );
or   ( new_n63858_, new_n50487_, new_n10052_ );
or   ( new_n63859_, new_n63858_, new_n10769_ );
and  ( new_n63860_, new_n63859_, new_n63857_ );
nor  ( new_n63861_, new_n63860_, new_n63855_ );
nor  ( new_n63862_, new_n63759_, new_n9424_ );
xor  ( new_n63863_, new_n51446_, RIbb2dae0_59 );
and  ( new_n63864_, new_n63863_, new_n9187_ );
or   ( new_n63865_, new_n63864_, new_n63862_ );
xor  ( new_n63866_, new_n63860_, new_n63855_ );
and  ( new_n63867_, new_n63866_, new_n63865_ );
nor  ( new_n63868_, new_n63867_, new_n63861_ );
not  ( new_n63869_, new_n63868_ );
xor  ( new_n63870_, new_n63853_, new_n63852_ );
and  ( new_n63871_, new_n63870_, new_n63869_ );
nor  ( new_n63872_, new_n63871_, new_n63854_ );
nand ( new_n63873_, new_n63872_, new_n63827_ );
and  ( new_n63874_, new_n63873_, new_n63826_ );
nor  ( new_n63875_, new_n63874_, new_n63822_ );
and  ( new_n63876_, new_n63874_, new_n63822_ );
xor  ( new_n63877_, new_n63850_, new_n63849_ );
and  ( new_n63878_, new_n63863_, new_n9185_ );
xor  ( new_n63879_, new_n51477_, RIbb2dae0_59 );
and  ( new_n63880_, new_n63879_, new_n9187_ );
or   ( new_n63881_, new_n63880_, new_n63878_ );
nor  ( new_n63882_, new_n63829_, new_n8876_ );
xor  ( new_n63883_, new_n52280_, new_n8254_ );
nor  ( new_n63884_, new_n63883_, new_n8874_ );
nor  ( new_n63885_, new_n63884_, new_n63882_ );
not  ( new_n63886_, new_n63885_ );
or   ( new_n63887_, new_n63886_, new_n63881_ );
and  ( new_n63888_, new_n63886_, new_n63881_ );
nor  ( new_n63889_, new_n53695_, new_n50765_ );
or   ( new_n63890_, new_n63889_, new_n7177_ );
or   ( new_n63891_, new_n63833_, new_n7734_ );
and  ( new_n63892_, new_n50764_, RIbb2ddb0_53 );
and  ( new_n63893_, new_n53694_, RIbb2dcc0_55 );
nor  ( new_n63894_, new_n63893_, new_n63892_ );
and  ( new_n63895_, RIbb2dd38_54, new_n7174_ );
nor  ( new_n63896_, new_n53694_, RIbb2dcc0_55 );
nor  ( new_n63897_, new_n63896_, new_n63895_ );
or   ( new_n63898_, new_n63897_, new_n63894_ );
and  ( new_n63899_, new_n63898_, new_n63891_ );
nor  ( new_n63900_, new_n63899_, new_n63890_ );
or   ( new_n63901_, new_n63900_, new_n63888_ );
and  ( new_n63902_, new_n63901_, new_n63887_ );
and  ( new_n63903_, new_n63902_, new_n63877_ );
xnor ( new_n63904_, new_n63842_, new_n63841_ );
xor  ( new_n63905_, new_n50487_, new_n10052_ );
or   ( new_n63906_, new_n63905_, new_n21077_ );
or   ( new_n63907_, new_n50788_, new_n10052_ );
or   ( new_n63908_, new_n63907_, new_n10769_ );
and  ( new_n63909_, new_n63908_, new_n63906_ );
nor  ( new_n63910_, new_n63909_, new_n63904_ );
nor  ( new_n63911_, new_n63847_, new_n10061_ );
xor  ( new_n63912_, new_n51142_, new_n9418_ );
nor  ( new_n63913_, new_n63912_, new_n10059_ );
or   ( new_n63914_, new_n63913_, new_n63911_ );
xor  ( new_n63915_, new_n63909_, new_n63904_ );
and  ( new_n63916_, new_n63915_, new_n63914_ );
nor  ( new_n63917_, new_n63916_, new_n63910_ );
not  ( new_n63918_, new_n63917_ );
xor  ( new_n63919_, new_n63902_, new_n63877_ );
and  ( new_n63920_, new_n63919_, new_n63918_ );
or   ( new_n63921_, new_n63920_, new_n63903_ );
xor  ( new_n63922_, new_n63796_, new_n63795_ );
and  ( new_n63923_, new_n63922_, new_n63921_ );
nor  ( new_n63924_, new_n63922_, new_n63921_ );
not  ( new_n63925_, new_n63924_ );
xor  ( new_n63926_, new_n63870_, new_n63869_ );
and  ( new_n63927_, new_n63926_, new_n63925_ );
nor  ( new_n63928_, new_n63927_, new_n63923_ );
xor  ( new_n63929_, new_n63825_, new_n63823_ );
xor  ( new_n63930_, new_n63929_, new_n63872_ );
nor  ( new_n63931_, new_n63930_, new_n63928_ );
and  ( new_n63932_, new_n63930_, new_n63928_ );
nor  ( new_n63933_, new_n63839_, new_n8266_ );
xor  ( new_n63934_, new_n52908_, RIbb2dcc0_55 );
nor  ( new_n63935_, new_n63934_, new_n8264_ );
or   ( new_n63936_, new_n63935_, new_n63933_ );
xor  ( new_n63937_, new_n63899_, new_n63890_ );
nand ( new_n63938_, new_n63937_, new_n63936_ );
nor  ( new_n63939_, new_n63883_, new_n8876_ );
xor  ( new_n63940_, new_n52293_, RIbb2dbd0_57 );
nor  ( new_n63941_, new_n63940_, new_n8874_ );
nor  ( new_n63942_, new_n63941_, new_n63939_ );
xnor ( new_n63943_, new_n63937_, new_n63936_ );
or   ( new_n63944_, new_n63943_, new_n63942_ );
and  ( new_n63945_, new_n63944_, new_n63938_ );
xor  ( new_n63946_, new_n63885_, new_n63881_ );
xor  ( new_n63947_, new_n63946_, new_n63900_ );
nor  ( new_n63948_, new_n63947_, new_n63945_ );
nand ( new_n63949_, new_n63947_, new_n63945_ );
xor  ( new_n63950_, new_n53306_, RIbb2dcc0_55 );
nor  ( new_n63951_, new_n63950_, new_n8264_ );
nor  ( new_n63952_, new_n63934_, new_n8266_ );
or   ( new_n63953_, new_n63952_, new_n63951_ );
and  ( new_n63954_, new_n53694_, new_n7487_ );
and  ( new_n63955_, new_n63954_, new_n63953_ );
xor  ( new_n63956_, new_n52902_, RIbb2dbd0_57 );
nor  ( new_n63957_, new_n63956_, new_n8874_ );
nor  ( new_n63958_, new_n63940_, new_n8876_ );
nor  ( new_n63959_, new_n63958_, new_n63957_ );
xnor ( new_n63960_, new_n63954_, new_n63953_ );
nor  ( new_n63961_, new_n63960_, new_n63959_ );
nor  ( new_n63962_, new_n63961_, new_n63955_ );
or   ( new_n63963_, new_n63912_, new_n10061_ );
xor  ( new_n63964_, new_n51446_, RIbb2d9f0_61 );
nand ( new_n63965_, new_n63964_, new_n9740_ );
and  ( new_n63966_, new_n63965_, new_n63963_ );
nor  ( new_n63967_, new_n63966_, new_n63962_ );
and  ( new_n63968_, new_n63966_, new_n63962_ );
and  ( new_n63969_, new_n63879_, new_n9185_ );
xor  ( new_n63970_, new_n51758_, new_n8870_ );
nor  ( new_n63971_, new_n63970_, new_n9422_ );
nor  ( new_n63972_, new_n63971_, new_n63969_ );
nor  ( new_n63973_, new_n63972_, new_n63968_ );
or   ( new_n63974_, new_n63973_, new_n63967_ );
and  ( new_n63975_, new_n63974_, new_n63949_ );
or   ( new_n63976_, new_n63975_, new_n63948_ );
xor  ( new_n63977_, new_n63866_, new_n63865_ );
and  ( new_n63978_, new_n63977_, new_n63976_ );
nor  ( new_n63979_, new_n63977_, new_n63976_ );
not  ( new_n63980_, new_n63979_ );
xor  ( new_n63981_, new_n63919_, new_n63918_ );
and  ( new_n63982_, new_n63981_, new_n63980_ );
nor  ( new_n63983_, new_n63982_, new_n63978_ );
not  ( new_n63984_, new_n63983_ );
xor  ( new_n63985_, new_n63922_, new_n63921_ );
xor  ( new_n63986_, new_n63985_, new_n63926_ );
and  ( new_n63987_, new_n63986_, new_n63984_ );
nor  ( new_n63988_, new_n63986_, new_n63984_ );
xor  ( new_n63989_, new_n63915_, new_n63914_ );
xor  ( new_n63990_, new_n63947_, new_n63945_ );
xor  ( new_n63991_, new_n63990_, new_n63974_ );
and  ( new_n63992_, new_n63991_, new_n63989_ );
nor  ( new_n63993_, new_n63991_, new_n63989_ );
xnor ( new_n63994_, new_n63943_, new_n63942_ );
xor  ( new_n63995_, new_n50788_, new_n10052_ );
or   ( new_n63996_, new_n63995_, new_n21077_ );
or   ( new_n63997_, new_n50894_, new_n10052_ );
or   ( new_n63998_, new_n63997_, new_n10769_ );
and  ( new_n63999_, new_n63998_, new_n63996_ );
nor  ( new_n64000_, new_n63999_, new_n63994_ );
and  ( new_n64001_, new_n63999_, new_n63994_ );
not  ( new_n64002_, new_n64001_ );
nor  ( new_n64003_, new_n63970_, new_n9424_ );
xor  ( new_n64004_, new_n52280_, new_n8870_ );
nor  ( new_n64005_, new_n64004_, new_n9422_ );
nor  ( new_n64006_, new_n64005_, new_n64003_ );
and  ( new_n64007_, new_n63964_, new_n9738_ );
xor  ( new_n64008_, new_n51477_, RIbb2d9f0_61 );
and  ( new_n64009_, new_n64008_, new_n9740_ );
nor  ( new_n64010_, new_n64009_, new_n64007_ );
and  ( new_n64011_, new_n64010_, new_n64006_ );
nor  ( new_n64012_, new_n64010_, new_n64006_ );
nor  ( new_n64013_, new_n53695_, new_n51217_ );
or   ( new_n64014_, new_n64013_, new_n7725_ );
or   ( new_n64015_, new_n63950_, new_n8266_ );
or   ( new_n64016_, new_n63893_, new_n8264_ );
or   ( new_n64017_, new_n64016_, new_n63896_ );
and  ( new_n64018_, new_n64017_, new_n64015_ );
nor  ( new_n64019_, new_n64018_, new_n64014_ );
nor  ( new_n64020_, new_n64019_, new_n64012_ );
nor  ( new_n64021_, new_n64020_, new_n64011_ );
and  ( new_n64022_, new_n64021_, new_n64002_ );
nor  ( new_n64023_, new_n64022_, new_n64000_ );
nor  ( new_n64024_, new_n64023_, new_n63993_ );
nor  ( new_n64025_, new_n64024_, new_n63992_ );
not  ( new_n64026_, new_n64025_ );
xor  ( new_n64027_, new_n63977_, new_n63976_ );
xor  ( new_n64028_, new_n64027_, new_n63981_ );
and  ( new_n64029_, new_n64028_, new_n64026_ );
nor  ( new_n64030_, new_n64028_, new_n64026_ );
xor  ( new_n64031_, new_n63966_, new_n63962_ );
not  ( new_n64032_, new_n64031_ );
and  ( new_n64033_, new_n64032_, new_n63972_ );
not  ( new_n64034_, new_n63967_ );
and  ( new_n64035_, new_n63973_, new_n64034_ );
nor  ( new_n64036_, new_n64035_, new_n64033_ );
not  ( new_n64037_, new_n64036_ );
xnor ( new_n64038_, new_n63960_, new_n63959_ );
xor  ( new_n64039_, new_n50894_, new_n10052_ );
or   ( new_n64040_, new_n64039_, new_n21077_ );
or   ( new_n64041_, new_n51142_, new_n10052_ );
or   ( new_n64042_, new_n64041_, new_n10769_ );
and  ( new_n64043_, new_n64042_, new_n64040_ );
or   ( new_n64044_, new_n64043_, new_n64038_ );
and  ( new_n64045_, new_n64043_, new_n64038_ );
nor  ( new_n64046_, new_n63956_, new_n8876_ );
xor  ( new_n64047_, new_n52908_, RIbb2dbd0_57 );
nor  ( new_n64048_, new_n64047_, new_n8874_ );
or   ( new_n64049_, new_n64048_, new_n64046_ );
xor  ( new_n64050_, new_n64018_, new_n64014_ );
and  ( new_n64051_, new_n64050_, new_n64049_ );
nor  ( new_n64052_, new_n64050_, new_n64049_ );
and  ( new_n64053_, new_n64008_, new_n9738_ );
xor  ( new_n64054_, new_n51758_, new_n9418_ );
nor  ( new_n64055_, new_n64054_, new_n10059_ );
nor  ( new_n64056_, new_n64055_, new_n64053_ );
nor  ( new_n64057_, new_n64056_, new_n64052_ );
nor  ( new_n64058_, new_n64057_, new_n64051_ );
or   ( new_n64059_, new_n64058_, new_n64045_ );
and  ( new_n64060_, new_n64059_, new_n64044_ );
and  ( new_n64061_, new_n64060_, new_n64037_ );
xor  ( new_n64062_, new_n64060_, new_n64037_ );
xor  ( new_n64063_, new_n63999_, new_n63994_ );
xnor ( new_n64064_, new_n64063_, new_n64021_ );
and  ( new_n64065_, new_n64064_, new_n64062_ );
nor  ( new_n64066_, new_n64065_, new_n64061_ );
xnor ( new_n64067_, new_n63991_, new_n63989_ );
xor  ( new_n64068_, new_n64067_, new_n64023_ );
and  ( new_n64069_, new_n64068_, new_n64066_ );
nor  ( new_n64070_, new_n64068_, new_n64066_ );
xnor ( new_n64071_, new_n64064_, new_n64062_ );
xnor ( new_n64072_, new_n64010_, new_n64006_ );
xor  ( new_n64073_, new_n64072_, new_n64019_ );
nor  ( new_n64074_, new_n64004_, new_n9424_ );
xor  ( new_n64075_, new_n52293_, RIbb2dae0_59 );
nor  ( new_n64076_, new_n64075_, new_n9422_ );
nor  ( new_n64077_, new_n64076_, new_n64074_ );
nor  ( new_n64078_, new_n64047_, new_n8876_ );
xor  ( new_n64079_, new_n53306_, RIbb2dbd0_57 );
nor  ( new_n64080_, new_n64079_, new_n8874_ );
or   ( new_n64081_, new_n64080_, new_n64078_ );
and  ( new_n64082_, new_n53694_, new_n8040_ );
nand ( new_n64083_, new_n64082_, new_n64081_ );
nor  ( new_n64084_, new_n64075_, new_n9424_ );
xor  ( new_n64085_, new_n52902_, RIbb2dae0_59 );
nor  ( new_n64086_, new_n64085_, new_n9422_ );
or   ( new_n64087_, new_n64086_, new_n64084_ );
xor  ( new_n64088_, new_n64082_, new_n64081_ );
nand ( new_n64089_, new_n64088_, new_n64087_ );
and  ( new_n64090_, new_n64089_, new_n64083_ );
or   ( new_n64091_, new_n64090_, new_n64077_ );
and  ( new_n64092_, new_n64090_, new_n64077_ );
xor  ( new_n64093_, new_n51142_, new_n10052_ );
or   ( new_n64094_, new_n64093_, new_n21077_ );
or   ( new_n64095_, new_n61553_, new_n51446_ );
and  ( new_n64096_, new_n64095_, new_n64094_ );
or   ( new_n64097_, new_n64096_, new_n64092_ );
and  ( new_n64098_, new_n64097_, new_n64091_ );
nand ( new_n64099_, new_n64098_, new_n64073_ );
nor  ( new_n64100_, new_n64098_, new_n64073_ );
xor  ( new_n64101_, new_n64043_, new_n64038_ );
xnor ( new_n64102_, new_n64101_, new_n64058_ );
or   ( new_n64103_, new_n64102_, new_n64100_ );
and  ( new_n64104_, new_n64103_, new_n64099_ );
and  ( new_n64105_, new_n64104_, new_n64071_ );
nor  ( new_n64106_, new_n64104_, new_n64071_ );
xor  ( new_n64107_, new_n64050_, new_n64049_ );
xnor ( new_n64108_, new_n64107_, new_n64056_ );
nor  ( new_n64109_, new_n53695_, new_n51962_ );
or   ( new_n64110_, new_n64109_, new_n8257_ );
or   ( new_n64111_, new_n64079_, new_n8876_ );
and  ( new_n64112_, new_n51961_, RIbb2dbd0_57 );
and  ( new_n64113_, new_n53694_, RIbb2dae0_59 );
nor  ( new_n64114_, new_n64113_, new_n64112_ );
and  ( new_n64115_, RIbb2db58_58, new_n8254_ );
nor  ( new_n64116_, new_n53694_, RIbb2dae0_59 );
nor  ( new_n64117_, new_n64116_, new_n64115_ );
or   ( new_n64118_, new_n64117_, new_n64114_ );
and  ( new_n64119_, new_n64118_, new_n64111_ );
or   ( new_n64120_, new_n64119_, new_n64110_ );
xor  ( new_n64121_, new_n52280_, new_n9418_ );
or   ( new_n64122_, new_n64121_, new_n10059_ );
or   ( new_n64123_, new_n64054_, new_n10061_ );
and  ( new_n64124_, new_n64123_, new_n64122_ );
nand ( new_n64125_, new_n64124_, new_n64120_ );
nor  ( new_n64126_, new_n64124_, new_n64120_ );
and  ( new_n64127_, new_n51446_, RIbb2d888_64 );
and  ( new_n64128_, new_n64127_, RIbb2d900_63 );
not  ( new_n64129_, new_n64128_ );
and  ( new_n64130_, new_n51477_, new_n21077_ );
nor  ( new_n64131_, new_n64127_, RIbb2d900_63 );
nor  ( new_n64132_, new_n64131_, new_n64130_ );
and  ( new_n64133_, new_n64132_, new_n64129_ );
or   ( new_n64134_, new_n64133_, new_n64126_ );
and  ( new_n64135_, new_n64134_, new_n64125_ );
nor  ( new_n64136_, new_n64135_, new_n64108_ );
xor  ( new_n64137_, new_n64135_, new_n64108_ );
not  ( new_n64138_, new_n64137_ );
xnor ( new_n64139_, new_n64090_, new_n64077_ );
xor  ( new_n64140_, new_n64139_, new_n64096_ );
nor  ( new_n64141_, new_n64140_, new_n64138_ );
or   ( new_n64142_, new_n64141_, new_n64136_ );
xnor ( new_n64143_, new_n64098_, new_n64073_ );
xor  ( new_n64144_, new_n64143_, new_n64102_ );
nor  ( new_n64145_, new_n64144_, new_n64142_ );
and  ( new_n64146_, new_n64144_, new_n64142_ );
nor  ( new_n64147_, new_n64085_, new_n9424_ );
xor  ( new_n64148_, new_n52908_, RIbb2dae0_59 );
nor  ( new_n64149_, new_n64148_, new_n9422_ );
or   ( new_n64150_, new_n64149_, new_n64147_ );
xor  ( new_n64151_, new_n64119_, new_n64110_ );
and  ( new_n64152_, new_n64151_, new_n64150_ );
nor  ( new_n64153_, new_n64121_, new_n10061_ );
xor  ( new_n64154_, new_n52293_, RIbb2d9f0_61 );
nor  ( new_n64155_, new_n64154_, new_n10059_ );
nor  ( new_n64156_, new_n64155_, new_n64153_ );
not  ( new_n64157_, new_n64156_ );
xor  ( new_n64158_, new_n64151_, new_n64150_ );
and  ( new_n64159_, new_n64158_, new_n64157_ );
nor  ( new_n64160_, new_n64159_, new_n64152_ );
not  ( new_n64161_, new_n64160_ );
xor  ( new_n64162_, new_n64088_, new_n64087_ );
and  ( new_n64163_, new_n64162_, new_n64161_ );
xor  ( new_n64164_, new_n64162_, new_n64161_ );
not  ( new_n64165_, new_n64164_ );
xnor ( new_n64166_, new_n64124_, new_n64120_ );
xor  ( new_n64167_, new_n64166_, new_n64133_ );
nor  ( new_n64168_, new_n64167_, new_n64165_ );
nor  ( new_n64169_, new_n64168_, new_n64163_ );
xor  ( new_n64170_, new_n64140_, new_n64138_ );
nor  ( new_n64171_, new_n64170_, new_n64169_ );
and  ( new_n64172_, new_n64170_, new_n64169_ );
nor  ( new_n64173_, new_n64148_, new_n9424_ );
xor  ( new_n64174_, new_n53306_, RIbb2dae0_59 );
nor  ( new_n64175_, new_n64174_, new_n9422_ );
or   ( new_n64176_, new_n64175_, new_n64173_ );
and  ( new_n64177_, new_n53694_, new_n8649_ );
nand ( new_n64178_, new_n64177_, new_n64176_ );
xor  ( new_n64179_, new_n52902_, RIbb2d9f0_61 );
nor  ( new_n64180_, new_n64179_, new_n10059_ );
nor  ( new_n64181_, new_n64154_, new_n10061_ );
nor  ( new_n64182_, new_n64181_, new_n64180_ );
not  ( new_n64183_, new_n64182_ );
xor  ( new_n64184_, new_n64177_, new_n64176_ );
nand ( new_n64185_, new_n64184_, new_n64183_ );
and  ( new_n64186_, new_n64185_, new_n64178_ );
or   ( new_n64187_, new_n51758_, new_n10052_ );
and  ( new_n64188_, new_n64187_, new_n10770_ );
and  ( new_n64189_, new_n51477_, RIbb2d888_64 );
or   ( new_n64190_, new_n64189_, new_n64188_ );
nand ( new_n64191_, new_n64189_, new_n10052_ );
and  ( new_n64192_, new_n64191_, new_n64190_ );
nor  ( new_n64193_, new_n64192_, new_n64186_ );
and  ( new_n64194_, new_n64192_, new_n64186_ );
xor  ( new_n64195_, new_n64158_, new_n64157_ );
not  ( new_n64196_, new_n64195_ );
nor  ( new_n64197_, new_n64196_, new_n64194_ );
nor  ( new_n64198_, new_n64197_, new_n64193_ );
and  ( new_n64199_, new_n53694_, new_n52349_ );
or   ( new_n64200_, new_n64199_, new_n8873_ );
or   ( new_n64201_, new_n64174_, new_n9424_ );
or   ( new_n64202_, new_n64113_, new_n9422_ );
or   ( new_n64203_, new_n64202_, new_n64116_ );
and  ( new_n64204_, new_n64203_, new_n64201_ );
or   ( new_n64205_, new_n64204_, new_n64200_ );
xor  ( new_n64206_, new_n51758_, new_n10052_ );
or   ( new_n64207_, new_n64206_, new_n21077_ );
or   ( new_n64208_, new_n52280_, new_n10052_ );
or   ( new_n64209_, new_n64208_, new_n10769_ );
and  ( new_n64210_, new_n64209_, new_n64207_ );
nor  ( new_n64211_, new_n64210_, new_n64205_ );
and  ( new_n64212_, new_n64210_, new_n64205_ );
xor  ( new_n64213_, new_n64184_, new_n64183_ );
not  ( new_n64214_, new_n64213_ );
nor  ( new_n64215_, new_n64214_, new_n64212_ );
nor  ( new_n64216_, new_n64215_, new_n64211_ );
xor  ( new_n64217_, new_n64192_, new_n64186_ );
xor  ( new_n64218_, new_n64217_, new_n64195_ );
not  ( new_n64219_, new_n64218_ );
and  ( new_n64220_, new_n64219_, new_n64216_ );
nor  ( new_n64221_, new_n64179_, new_n10061_ );
xor  ( new_n64222_, new_n52908_, RIbb2d9f0_61 );
nor  ( new_n64223_, new_n64222_, new_n10059_ );
nor  ( new_n64224_, new_n64223_, new_n64221_ );
not  ( new_n64225_, new_n64224_ );
xor  ( new_n64226_, new_n64204_, new_n64200_ );
and  ( new_n64227_, new_n64226_, new_n64225_ );
xor  ( new_n64228_, new_n64226_, new_n64225_ );
not  ( new_n64229_, new_n64228_ );
xor  ( new_n64230_, new_n52280_, new_n10052_ );
or   ( new_n64231_, new_n64230_, new_n21077_ );
nand ( new_n64232_, new_n52293_, RIbb2d900_63 );
or   ( new_n64233_, new_n64232_, RIbb2d888_64 );
and  ( new_n64234_, new_n64233_, new_n64231_ );
nor  ( new_n64235_, new_n64234_, new_n64229_ );
nor  ( new_n64236_, new_n64235_, new_n64227_ );
xor  ( new_n64237_, new_n64210_, new_n64205_ );
xor  ( new_n64238_, new_n64237_, new_n64213_ );
not  ( new_n64239_, new_n64238_ );
and  ( new_n64240_, new_n64239_, new_n64236_ );
xor  ( new_n64241_, new_n64234_, new_n64229_ );
or   ( new_n64242_, new_n53695_, new_n9424_ );
xor  ( new_n64243_, new_n52293_, RIbb2d900_63 );
or   ( new_n64244_, new_n64243_, new_n21077_ );
nand ( new_n64245_, new_n52902_, RIbb2d900_63 );
or   ( new_n64246_, new_n64245_, RIbb2d888_64 );
and  ( new_n64247_, new_n64246_, new_n64244_ );
nor  ( new_n64248_, new_n64247_, new_n64242_ );
and  ( new_n64249_, new_n64247_, new_n64242_ );
nor  ( new_n64250_, new_n64222_, new_n10061_ );
xor  ( new_n64251_, new_n53306_, RIbb2d9f0_61 );
nor  ( new_n64252_, new_n64251_, new_n10059_ );
nor  ( new_n64253_, new_n64252_, new_n64250_ );
nor  ( new_n64254_, new_n64253_, new_n64249_ );
nor  ( new_n64255_, new_n64254_, new_n64248_ );
not  ( new_n64256_, new_n64255_ );
and  ( new_n64257_, new_n64256_, new_n64241_ );
nor  ( new_n64258_, new_n64256_, new_n64241_ );
nor  ( new_n64259_, new_n53695_, new_n52849_ );
nor  ( new_n64260_, new_n64259_, new_n9421_ );
not  ( new_n64261_, new_n64260_ );
or   ( new_n64262_, new_n64251_, new_n10061_ );
and  ( new_n64263_, new_n53694_, RIbb2d9f0_61 );
nor  ( new_n64264_, new_n53694_, RIbb2d9f0_61 );
or   ( new_n64265_, new_n64264_, new_n10059_ );
or   ( new_n64266_, new_n64265_, new_n64263_ );
and  ( new_n64267_, new_n64266_, new_n64262_ );
nor  ( new_n64268_, new_n64267_, new_n64261_ );
xor  ( new_n64269_, new_n64247_, new_n64242_ );
xor  ( new_n64270_, new_n64269_, new_n64253_ );
not  ( new_n64271_, new_n64270_ );
and  ( new_n64272_, new_n64271_, new_n64268_ );
nor  ( new_n64273_, new_n64271_, new_n64268_ );
xor  ( new_n64274_, new_n52908_, RIbb2d900_63 );
nor  ( new_n64275_, new_n64274_, new_n21077_ );
and  ( new_n64276_, new_n57100_, new_n53306_ );
nor  ( new_n64277_, new_n64276_, new_n64275_ );
and  ( new_n64278_, new_n53694_, new_n9738_ );
nor  ( new_n64279_, new_n53306_, new_n21077_ );
not  ( new_n64280_, new_n64279_ );
nor  ( new_n64281_, new_n53694_, new_n10052_ );
and  ( new_n64282_, new_n64281_, new_n64280_ );
nor  ( new_n64283_, new_n64282_, new_n64278_ );
nor  ( new_n64284_, new_n64283_, new_n64277_ );
xor  ( new_n64285_, new_n64267_, new_n64261_ );
and  ( new_n64286_, new_n64285_, new_n64284_ );
nor  ( new_n64287_, new_n64285_, new_n64284_ );
xor  ( new_n64288_, new_n52902_, RIbb2d900_63 );
nor  ( new_n64289_, new_n64288_, new_n21077_ );
and  ( new_n64290_, new_n52908_, RIbb2d900_63 );
and  ( new_n64291_, new_n64290_, new_n21077_ );
nor  ( new_n64292_, new_n64291_, new_n64289_ );
nor  ( new_n64293_, new_n64292_, new_n64287_ );
nor  ( new_n64294_, new_n64293_, new_n64286_ );
nor  ( new_n64295_, new_n64294_, new_n64273_ );
nor  ( new_n64296_, new_n64295_, new_n64272_ );
nor  ( new_n64297_, new_n64296_, new_n64258_ );
nor  ( new_n64298_, new_n64297_, new_n64257_ );
nor  ( new_n64299_, new_n64298_, new_n64240_ );
not  ( new_n64300_, new_n64299_ );
nor  ( new_n64301_, new_n64239_, new_n64236_ );
nor  ( new_n64302_, new_n64219_, new_n64216_ );
nor  ( new_n64303_, new_n64302_, new_n64301_ );
and  ( new_n64304_, new_n64303_, new_n64300_ );
nor  ( new_n64305_, new_n64304_, new_n64220_ );
not  ( new_n64306_, new_n64305_ );
and  ( new_n64307_, new_n64306_, new_n64198_ );
not  ( new_n64308_, new_n64307_ );
xor  ( new_n64309_, new_n64167_, new_n64165_ );
and  ( new_n64310_, new_n64309_, new_n64308_ );
nor  ( new_n64311_, new_n64306_, new_n64198_ );
nor  ( new_n64312_, new_n64311_, new_n64310_ );
nor  ( new_n64313_, new_n64312_, new_n64172_ );
nor  ( new_n64314_, new_n64313_, new_n64171_ );
nor  ( new_n64315_, new_n64314_, new_n64146_ );
nor  ( new_n64316_, new_n64315_, new_n64145_ );
nor  ( new_n64317_, new_n64316_, new_n64106_ );
nor  ( new_n64318_, new_n64317_, new_n64105_ );
nor  ( new_n64319_, new_n64318_, new_n64070_ );
nor  ( new_n64320_, new_n64319_, new_n64069_ );
nor  ( new_n64321_, new_n64320_, new_n64030_ );
nor  ( new_n64322_, new_n64321_, new_n64029_ );
nor  ( new_n64323_, new_n64322_, new_n63988_ );
nor  ( new_n64324_, new_n64323_, new_n63987_ );
nor  ( new_n64325_, new_n64324_, new_n63932_ );
nor  ( new_n64326_, new_n64325_, new_n63931_ );
not  ( new_n64327_, new_n64326_ );
nor  ( new_n64328_, new_n64327_, new_n63876_ );
nor  ( new_n64329_, new_n64328_, new_n63875_ );
nor  ( new_n64330_, new_n64329_, new_n63820_ );
nor  ( new_n64331_, new_n64330_, new_n63819_ );
nor  ( new_n64332_, new_n64331_, new_n63775_ );
nor  ( new_n64333_, new_n64332_, new_n63774_ );
nor  ( new_n64334_, new_n64333_, new_n63723_ );
nor  ( new_n64335_, new_n64334_, new_n63722_ );
nor  ( new_n64336_, new_n64335_, new_n63655_ );
nor  ( new_n64337_, new_n64336_, new_n63654_ );
nor  ( new_n64338_, new_n64337_, new_n63591_ );
nor  ( new_n64339_, new_n64338_, new_n63590_ );
nor  ( new_n64340_, new_n64339_, new_n63477_ );
nor  ( new_n64341_, new_n64340_, new_n63476_ );
not  ( new_n64342_, new_n64341_ );
nor  ( new_n64343_, new_n64342_, new_n63409_ );
nor  ( new_n64344_, new_n64343_, new_n63408_ );
nor  ( new_n64345_, new_n64344_, new_n63301_ );
nor  ( new_n64346_, new_n64345_, new_n63300_ );
nor  ( new_n64347_, new_n64346_, new_n63254_ );
nor  ( new_n64348_, new_n64347_, new_n63253_ );
nor  ( new_n64349_, new_n64348_, new_n63161_ );
nor  ( new_n64350_, new_n64349_, new_n63160_ );
nor  ( new_n64351_, new_n64350_, new_n62994_ );
nor  ( new_n64352_, new_n64351_, new_n62993_ );
nor  ( new_n64353_, new_n64352_, new_n62973_ );
and  ( new_n64354_, new_n64353_, new_n62827_ );
not  ( new_n64355_, new_n64354_ );
and  ( new_n64356_, new_n62820_, new_n62816_ );
nor  ( new_n64357_, new_n62824_, new_n62822_ );
nor  ( new_n64358_, new_n64357_, new_n64356_ );
xor  ( new_n64359_, new_n62485_, new_n62483_ );
xnor ( new_n64360_, new_n64359_, new_n62553_ );
and  ( new_n64361_, new_n64360_, new_n64358_ );
not  ( new_n64362_, new_n64361_ );
nor  ( new_n64363_, new_n62825_, new_n62812_ );
nor  ( new_n64364_, new_n62972_, new_n62828_ );
and  ( new_n64365_, new_n64364_, new_n62827_ );
nor  ( new_n64366_, new_n64365_, new_n64363_ );
and  ( new_n64367_, new_n64366_, new_n64362_ );
and  ( new_n64368_, new_n64367_, new_n64355_ );
not  ( new_n64369_, new_n64368_ );
nor  ( new_n64370_, new_n64360_, new_n64358_ );
and  ( new_n64371_, new_n62558_, new_n62555_ );
nor  ( new_n64372_, new_n64371_, new_n64370_ );
and  ( new_n64373_, new_n64372_, new_n64369_ );
nor  ( new_n64374_, new_n64373_, new_n62560_ );
nor  ( new_n64375_, new_n64374_, new_n62482_ );
not  ( new_n64376_, new_n64375_ );
nor  ( new_n64377_, new_n64376_, new_n62339_ );
and  ( new_n64378_, new_n64377_, new_n62219_ );
and  ( new_n64379_, new_n64378_, new_n61905_ );
not  ( new_n64380_, new_n64379_ );
and  ( new_n64381_, new_n62146_, new_n62144_ );
nor  ( new_n64382_, new_n62217_, new_n62215_ );
and  ( new_n64383_, new_n62480_, new_n62340_ );
nor  ( new_n64384_, new_n62338_, new_n62336_ );
nor  ( new_n64385_, new_n64384_, new_n64383_ );
nor  ( new_n64386_, new_n64385_, new_n62339_ );
nor  ( new_n64387_, new_n64386_, new_n64382_ );
not  ( new_n64388_, new_n64387_ );
and  ( new_n64389_, new_n64388_, new_n62219_ );
nor  ( new_n64390_, new_n64389_, new_n64381_ );
not  ( new_n64391_, new_n64390_ );
and  ( new_n64392_, new_n64391_, new_n61905_ );
not  ( new_n64393_, new_n64392_ );
nor  ( new_n64394_, new_n61589_, new_n61588_ );
nor  ( new_n64395_, new_n61664_, new_n61663_ );
not  ( new_n64396_, new_n64395_ );
nor  ( new_n64397_, new_n61880_, new_n61879_ );
nor  ( new_n64398_, new_n61901_, new_n61883_ );
and  ( new_n64399_, new_n64398_, new_n61882_ );
nor  ( new_n64400_, new_n64399_, new_n64397_ );
and  ( new_n64401_, new_n64400_, new_n64396_ );
not  ( new_n64402_, new_n64401_ );
and  ( new_n64403_, new_n64402_, new_n61666_ );
nor  ( new_n64404_, new_n64403_, new_n64394_ );
and  ( new_n64405_, new_n64404_, new_n64393_ );
and  ( new_n64406_, new_n64405_, new_n64380_ );
nor  ( new_n64407_, new_n64406_, new_n61442_ );
and  ( new_n64408_, new_n64407_, new_n61237_ );
and  ( new_n64409_, new_n64408_, new_n61021_ );
xor  ( new_n64410_, new_n60081_, new_n59976_ );
xor  ( new_n64411_, new_n64410_, new_n60084_ );
not  ( new_n64412_, new_n64411_ );
and  ( new_n64413_, new_n61006_, new_n61004_ );
nor  ( new_n64414_, new_n61006_, new_n61004_ );
nor  ( new_n64415_, new_n64414_, new_n61000_ );
or   ( new_n64416_, new_n64415_, new_n64413_ );
xor  ( new_n64417_, new_n59851_, new_n59846_ );
xnor ( new_n64418_, new_n64417_, new_n59855_ );
or   ( new_n64419_, new_n60981_, new_n60977_ );
nand ( new_n64420_, new_n60981_, new_n60977_ );
nand ( new_n64421_, new_n64420_, new_n60976_ );
and  ( new_n64422_, new_n64421_, new_n64419_ );
xor  ( new_n64423_, new_n59736_, new_n59734_ );
xor  ( new_n64424_, new_n64423_, new_n59760_ );
xnor ( new_n64425_, new_n64424_, new_n64422_ );
xor  ( new_n64426_, new_n64425_, new_n64418_ );
nand ( new_n64427_, new_n64426_, new_n64416_ );
nor  ( new_n64428_, new_n64426_, new_n64416_ );
and  ( new_n64429_, new_n60983_, new_n60975_ );
nor  ( new_n64430_, new_n60983_, new_n60975_ );
nor  ( new_n64431_, new_n64430_, new_n60971_ );
nor  ( new_n64432_, new_n64431_, new_n64429_ );
or   ( new_n64433_, new_n64432_, new_n64428_ );
and  ( new_n64434_, new_n64433_, new_n64427_ );
and  ( new_n64435_, new_n64434_, new_n64412_ );
xor  ( new_n64436_, new_n64434_, new_n64412_ );
not  ( new_n64437_, new_n64436_ );
xor  ( new_n64438_, new_n59974_, new_n59973_ );
or   ( new_n64439_, new_n60969_, new_n60968_ );
and  ( new_n64440_, new_n60969_, new_n60968_ );
or   ( new_n64441_, new_n64440_, new_n60965_ );
and  ( new_n64442_, new_n64441_, new_n64439_ );
and  ( new_n64443_, new_n64442_, new_n64438_ );
nor  ( new_n64444_, new_n64442_, new_n64438_ );
xor  ( new_n64445_, new_n60079_, new_n59983_ );
not  ( new_n64446_, new_n64445_ );
nor  ( new_n64447_, new_n64446_, new_n64444_ );
nor  ( new_n64448_, new_n64447_, new_n64443_ );
xnor ( new_n64449_, new_n59860_, new_n59859_ );
or   ( new_n64450_, new_n64424_, new_n64422_ );
and  ( new_n64451_, new_n64424_, new_n64422_ );
or   ( new_n64452_, new_n64451_, new_n64418_ );
and  ( new_n64453_, new_n64452_, new_n64450_ );
xnor ( new_n64454_, new_n64453_, new_n64449_ );
xor  ( new_n64455_, new_n64454_, new_n64448_ );
nor  ( new_n64456_, new_n64455_, new_n64437_ );
nor  ( new_n64457_, new_n64456_, new_n64435_ );
not  ( new_n64458_, new_n64457_ );
xor  ( new_n64459_, new_n59867_, new_n59862_ );
xnor ( new_n64460_, new_n64459_, new_n60087_ );
not  ( new_n64461_, new_n64460_ );
or   ( new_n64462_, new_n64453_, new_n64449_ );
and  ( new_n64463_, new_n64453_, new_n64449_ );
or   ( new_n64464_, new_n64463_, new_n64448_ );
and  ( new_n64465_, new_n64464_, new_n64462_ );
xor  ( new_n64466_, new_n59778_, new_n59776_ );
xor  ( new_n64467_, new_n64466_, new_n59783_ );
xor  ( new_n64468_, new_n64467_, new_n64465_ );
xor  ( new_n64469_, new_n64468_, new_n64461_ );
and  ( new_n64470_, new_n64469_, new_n64458_ );
xor  ( new_n64471_, new_n60089_, new_n59799_ );
xor  ( new_n64472_, new_n64471_, new_n60094_ );
or   ( new_n64473_, new_n64467_, new_n64465_ );
and  ( new_n64474_, new_n64467_, new_n64465_ );
or   ( new_n64475_, new_n64474_, new_n64461_ );
and  ( new_n64476_, new_n64475_, new_n64473_ );
and  ( new_n64477_, new_n64476_, new_n64472_ );
nor  ( new_n64478_, new_n64477_, new_n64470_ );
nor  ( new_n64479_, new_n61012_, new_n61008_ );
and  ( new_n64480_, new_n61012_, new_n61008_ );
not  ( new_n64481_, new_n64480_ );
and  ( new_n64482_, new_n64481_, new_n60996_ );
nor  ( new_n64483_, new_n64482_, new_n64479_ );
xor  ( new_n64484_, new_n64442_, new_n64438_ );
xor  ( new_n64485_, new_n64484_, new_n64446_ );
and  ( new_n64486_, new_n64485_, new_n64483_ );
xor  ( new_n64487_, new_n64485_, new_n64483_ );
not  ( new_n64488_, new_n64487_ );
xnor ( new_n64489_, new_n64426_, new_n64416_ );
xor  ( new_n64490_, new_n64489_, new_n64432_ );
nor  ( new_n64491_, new_n64490_, new_n64488_ );
nor  ( new_n64492_, new_n64491_, new_n64486_ );
not  ( new_n64493_, new_n64492_ );
xor  ( new_n64494_, new_n64455_, new_n64437_ );
and  ( new_n64495_, new_n64494_, new_n64493_ );
not  ( new_n64496_, new_n64495_ );
and  ( new_n64497_, new_n60990_, new_n60986_ );
nor  ( new_n64498_, new_n61014_, new_n60992_ );
nor  ( new_n64499_, new_n64498_, new_n64497_ );
not  ( new_n64500_, new_n64499_ );
xor  ( new_n64501_, new_n64490_, new_n64488_ );
and  ( new_n64502_, new_n64501_, new_n64500_ );
not  ( new_n64503_, new_n64502_ );
and  ( new_n64504_, new_n64503_, new_n64496_ );
and  ( new_n64505_, new_n64504_, new_n64478_ );
and  ( new_n64506_, new_n64505_, new_n64409_ );
not  ( new_n64507_, new_n64506_ );
nor  ( new_n64508_, new_n64476_, new_n64472_ );
nor  ( new_n64509_, new_n60963_, new_n60887_ );
not  ( new_n64510_, new_n64509_ );
nor  ( new_n64511_, new_n61235_, new_n61234_ );
nor  ( new_n64512_, new_n61441_, new_n61440_ );
and  ( new_n64513_, new_n64512_, new_n61237_ );
nor  ( new_n64514_, new_n64513_, new_n64511_ );
and  ( new_n64515_, new_n64514_, new_n64510_ );
not  ( new_n64516_, new_n64515_ );
and  ( new_n64517_, new_n64516_, new_n61021_ );
nor  ( new_n64518_, new_n61019_, new_n61015_ );
nor  ( new_n64519_, new_n64518_, new_n64517_ );
not  ( new_n64520_, new_n64519_ );
and  ( new_n64521_, new_n64520_, new_n64504_ );
not  ( new_n64522_, new_n64521_ );
nor  ( new_n64523_, new_n64469_, new_n64458_ );
not  ( new_n64524_, new_n64523_ );
nor  ( new_n64525_, new_n64494_, new_n64493_ );
nor  ( new_n64526_, new_n64501_, new_n64500_ );
and  ( new_n64527_, new_n64526_, new_n64496_ );
nor  ( new_n64528_, new_n64527_, new_n64525_ );
and  ( new_n64529_, new_n64528_, new_n64524_ );
and  ( new_n64530_, new_n64529_, new_n64522_ );
not  ( new_n64531_, new_n64530_ );
and  ( new_n64532_, new_n64531_, new_n64478_ );
nor  ( new_n64533_, new_n64532_, new_n64508_ );
and  ( new_n64534_, new_n64533_, new_n64507_ );
nor  ( new_n64535_, new_n64534_, new_n60098_ );
nor  ( new_n64536_, new_n64535_, new_n60097_ );
nor  ( new_n64537_, new_n64536_, new_n59796_ );
nor  ( new_n64538_, new_n64537_, new_n59795_ );
nor  ( new_n64539_, new_n64538_, new_n59602_ );
nor  ( new_n64540_, new_n64539_, new_n59601_ );
nor  ( new_n64541_, new_n64540_, new_n59478_ );
nor  ( new_n64542_, new_n64541_, new_n59477_ );
not  ( new_n64543_, new_n64542_ );
and  ( new_n64544_, new_n59459_, new_n59450_ );
and  ( new_n64545_, new_n59460_, new_n59447_ );
nor  ( new_n64546_, new_n64545_, new_n64544_ );
xor  ( new_n64547_, new_n58638_, new_n58636_ );
xor  ( new_n64548_, new_n64547_, new_n58642_ );
nor  ( new_n64549_, new_n64548_, new_n64546_ );
xor  ( new_n64550_, new_n64548_, new_n64546_ );
xnor ( new_n64551_, new_n58492_, new_n58490_ );
or   ( new_n64552_, new_n59457_, new_n59455_ );
nand ( new_n64553_, new_n59457_, new_n59455_ );
nand ( new_n64554_, new_n64553_, new_n59454_ );
and  ( new_n64555_, new_n64554_, new_n64552_ );
xor  ( new_n64556_, new_n64555_, new_n64551_ );
or   ( new_n64557_, new_n59468_, new_n59464_ );
nand ( new_n64558_, new_n59468_, new_n59464_ );
nand ( new_n64559_, new_n64558_, new_n59463_ );
and  ( new_n64560_, new_n64559_, new_n64557_ );
xor  ( new_n64561_, new_n64560_, new_n64556_ );
and  ( new_n64562_, new_n64561_, new_n64550_ );
nor  ( new_n64563_, new_n64562_, new_n64549_ );
nor  ( new_n64564_, new_n64555_, new_n64551_ );
and  ( new_n64565_, new_n64560_, new_n64556_ );
nor  ( new_n64566_, new_n64565_, new_n64564_ );
not  ( new_n64567_, new_n64566_ );
xor  ( new_n64568_, new_n58349_, new_n58348_ );
xor  ( new_n64569_, new_n64568_, new_n64567_ );
not  ( new_n64570_, new_n64569_ );
xor  ( new_n64571_, new_n58496_, new_n58494_ );
xor  ( new_n64572_, new_n64571_, new_n58644_ );
xor  ( new_n64573_, new_n64572_, new_n64570_ );
not  ( new_n64574_, new_n64573_ );
and  ( new_n64575_, new_n64574_, new_n64563_ );
and  ( new_n64576_, new_n59470_, new_n59461_ );
nor  ( new_n64577_, new_n59475_, new_n59471_ );
nor  ( new_n64578_, new_n64577_, new_n64576_ );
xor  ( new_n64579_, new_n64561_, new_n64550_ );
not  ( new_n64580_, new_n64579_ );
and  ( new_n64581_, new_n64580_, new_n64578_ );
nor  ( new_n64582_, new_n64581_, new_n64575_ );
and  ( new_n64583_, new_n64582_, new_n64543_ );
not  ( new_n64584_, new_n64583_ );
and  ( new_n64585_, new_n64568_, new_n64567_ );
nor  ( new_n64586_, new_n64572_, new_n64570_ );
nor  ( new_n64587_, new_n64586_, new_n64585_ );
not  ( new_n64588_, new_n64587_ );
xor  ( new_n64589_, new_n58646_, new_n58370_ );
and  ( new_n64590_, new_n64589_, new_n64588_ );
nor  ( new_n64591_, new_n64574_, new_n64563_ );
nor  ( new_n64592_, new_n64580_, new_n64578_ );
nor  ( new_n64593_, new_n64592_, new_n64591_ );
nor  ( new_n64594_, new_n64593_, new_n64575_ );
nor  ( new_n64595_, new_n64594_, new_n64590_ );
and  ( new_n64596_, new_n64595_, new_n64584_ );
not  ( new_n64597_, new_n64596_ );
nor  ( new_n64598_, new_n64589_, new_n64588_ );
nor  ( new_n64599_, new_n58651_, new_n58649_ );
nor  ( new_n64600_, new_n64599_, new_n64598_ );
and  ( new_n64601_, new_n64600_, new_n64597_ );
nor  ( new_n64602_, new_n64601_, new_n58652_ );
nor  ( new_n64603_, new_n64602_, new_n58364_ );
nor  ( new_n64604_, new_n58363_, new_n58265_ );
nor  ( new_n64605_, new_n64604_, new_n64603_ );
not  ( new_n64606_, new_n64605_ );
nor  ( new_n64607_, new_n64606_, new_n58264_ );
nor  ( new_n64608_, new_n64607_, new_n58263_ );
nor  ( new_n64609_, new_n64608_, new_n57798_ );
nor  ( new_n64610_, new_n64609_, new_n57797_ );
not  ( new_n64611_, new_n64610_ );
nor  ( new_n64612_, new_n64611_, new_n57686_ );
nor  ( new_n64613_, new_n64612_, new_n57685_ );
not  ( new_n64614_, new_n64613_ );
nor  ( new_n64615_, new_n64614_, new_n57377_ );
nor  ( new_n64616_, new_n64615_, new_n57376_ );
not  ( new_n64617_, new_n64616_ );
nor  ( new_n64618_, new_n64617_, new_n57125_ );
nor  ( new_n64619_, new_n64618_, new_n57124_ );
nor  ( new_n64620_, new_n64619_, new_n56880_ );
nor  ( new_n64621_, new_n64620_, new_n56879_ );
nor  ( new_n64622_, new_n64621_, new_n56573_ );
nor  ( new_n64623_, new_n64622_, new_n56572_ );
not  ( new_n64624_, new_n64623_ );
and  ( new_n64625_, new_n64624_, new_n56361_ );
not  ( new_n64626_, new_n64625_ );
nor  ( new_n64627_, new_n56359_, new_n56356_ );
nor  ( new_n64628_, new_n55961_, new_n55730_ );
nor  ( new_n64629_, new_n64628_, new_n64627_ );
and  ( new_n64630_, new_n64629_, new_n64626_ );
nor  ( new_n64631_, new_n64630_, new_n55962_ );
nor  ( new_n64632_, new_n64631_, new_n55729_ );
nor  ( new_n64633_, new_n64632_, new_n55728_ );
nor  ( new_n64634_, new_n64633_, new_n55454_ );
not  ( new_n64635_, new_n64634_ );
nor  ( new_n64636_, new_n55336_, new_n55327_ );
and  ( new_n64637_, new_n55336_, new_n55327_ );
nor  ( new_n64638_, new_n64637_, new_n54863_ );
nor  ( new_n64639_, new_n64638_, new_n64636_ );
nor  ( new_n64640_, new_n54860_, new_n54714_ );
and  ( new_n64641_, new_n54862_, new_n54861_ );
nor  ( new_n64642_, new_n64641_, new_n64640_ );
nor  ( new_n64643_, new_n55333_, new_n55330_ );
and  ( new_n64644_, new_n55335_, new_n55334_ );
or   ( new_n64645_, new_n64644_, new_n64643_ );
xor  ( new_n64646_, new_n54500_, new_n54499_ );
xor  ( new_n64647_, new_n64646_, new_n64645_ );
xnor ( new_n64648_, new_n64647_, new_n64642_ );
nor  ( new_n64649_, new_n64648_, new_n64639_ );
and  ( new_n64650_, new_n55453_, new_n55338_ );
nor  ( new_n64651_, new_n64650_, new_n64649_ );
and  ( new_n64652_, new_n64651_, new_n64635_ );
not  ( new_n64653_, new_n64652_ );
xor  ( new_n64654_, new_n54261_, new_n54259_ );
xor  ( new_n64655_, new_n64654_, new_n54502_ );
nand ( new_n64656_, new_n64646_, new_n64645_ );
nor  ( new_n64657_, new_n64646_, new_n64645_ );
or   ( new_n64658_, new_n64657_, new_n64642_ );
and  ( new_n64659_, new_n64658_, new_n64656_ );
nor  ( new_n64660_, new_n64659_, new_n64655_ );
and  ( new_n64661_, new_n64648_, new_n64639_ );
nor  ( new_n64662_, new_n64661_, new_n64660_ );
and  ( new_n64663_, new_n64662_, new_n64653_ );
not  ( new_n64664_, new_n64663_ );
and  ( new_n64665_, new_n64659_, new_n64655_ );
nor  ( new_n64666_, new_n54506_, new_n54258_ );
nor  ( new_n64667_, new_n64666_, new_n64665_ );
and  ( new_n64668_, new_n64667_, new_n64664_ );
nor  ( new_n64669_, new_n64668_, new_n54507_ );
not  ( new_n64670_, new_n64669_ );
nor  ( new_n64671_, new_n64670_, new_n54257_ );
nor  ( new_n64672_, new_n64671_, new_n54256_ );
nor  ( new_n64673_, new_n64672_, new_n53989_ );
nor  ( new_n64674_, new_n64673_, new_n53988_ );
nor  ( new_n64675_, new_n64674_, new_n53559_ );
nor  ( new_n64676_, new_n64675_, new_n53558_ );
and  ( new_n64677_, new_n64676_, new_n53267_ );
nor  ( new_n64678_, new_n64677_, new_n53265_ );
not  ( new_n64679_, new_n64678_ );
nor  ( new_n64680_, new_n64679_, new_n52836_ );
not  ( new_n64681_, new_n64680_ );
nor  ( new_n64682_, new_n52821_, new_n52817_ );
and  ( new_n64683_, new_n52826_, new_n52822_ );
nor  ( new_n64684_, new_n64683_, new_n64682_ );
not  ( new_n64685_, new_n64684_ );
xor  ( new_n64686_, new_n51811_, new_n51809_ );
xor  ( new_n64687_, new_n64686_, new_n51814_ );
xor  ( new_n64688_, new_n64687_, new_n64685_ );
xor  ( new_n64689_, new_n52125_, new_n52017_ );
xor  ( new_n64690_, new_n64689_, new_n64688_ );
not  ( new_n64691_, new_n64690_ );
nor  ( new_n64692_, new_n52829_, new_n52827_ );
and  ( new_n64693_, new_n52829_, new_n52827_ );
nor  ( new_n64694_, new_n52834_, new_n64693_ );
nor  ( new_n64695_, new_n64694_, new_n64692_ );
and  ( new_n64696_, new_n64695_, new_n64691_ );
not  ( new_n64697_, new_n64696_ );
and  ( new_n64698_, new_n52835_, new_n52815_ );
and  ( new_n64699_, new_n64687_, new_n64685_ );
and  ( new_n64700_, new_n64689_, new_n64688_ );
nor  ( new_n64701_, new_n64700_, new_n64699_ );
xor  ( new_n64702_, new_n51835_, new_n51834_ );
xor  ( new_n64703_, new_n64702_, new_n52127_ );
and  ( new_n64704_, new_n64703_, new_n64701_ );
nor  ( new_n64705_, new_n64704_, new_n64698_ );
and  ( new_n64706_, new_n64705_, new_n64697_ );
and  ( new_n64707_, new_n64706_, new_n64681_ );
not  ( new_n64708_, new_n64707_ );
not  ( new_n64709_, new_n64704_ );
nor  ( new_n64710_, new_n64695_, new_n64691_ );
and  ( new_n64711_, new_n64710_, new_n64709_ );
not  ( new_n64712_, new_n64711_ );
nor  ( new_n64713_, new_n64703_, new_n64701_ );
nor  ( new_n64714_, new_n52132_, new_n51833_ );
nor  ( new_n64715_, new_n64714_, new_n64713_ );
and  ( new_n64716_, new_n64715_, new_n64712_ );
and  ( new_n64717_, new_n64716_, new_n64708_ );
nor  ( new_n64718_, new_n64717_, new_n52133_ );
nor  ( new_n64719_, new_n64718_, new_n51832_ );
nor  ( new_n64720_, new_n64719_, new_n51831_ );
nor  ( new_n64721_, new_n64720_, new_n51522_ );
nor  ( new_n64722_, new_n64721_, new_n51521_ );
nor  ( new_n64723_, new_n64722_, new_n51261_ );
nor  ( new_n64724_, new_n64723_, new_n51260_ );
nor  ( new_n64725_, new_n64724_, new_n50868_ );
nor  ( new_n64726_, new_n64725_, new_n50867_ );
nor  ( new_n64727_, new_n64726_, new_n50623_ );
nor  ( new_n64728_, new_n64727_, new_n50622_ );
nor  ( new_n64729_, new_n64728_, new_n50294_ );
nor  ( new_n64730_, new_n64729_, new_n50293_ );
nor  ( new_n64731_, new_n64730_, new_n50155_ );
nor  ( new_n64732_, new_n64731_, new_n50154_ );
nor  ( new_n64733_, new_n64732_, new_n49888_ );
nor  ( new_n64734_, new_n64733_, new_n49887_ );
nor  ( new_n64735_, new_n64734_, new_n49619_ );
nor  ( new_n64736_, new_n64735_, new_n49618_ );
not  ( new_n64737_, new_n64736_ );
nor  ( new_n64738_, new_n64737_, new_n49361_ );
nor  ( new_n64739_, new_n64738_, new_n49360_ );
nor  ( new_n64740_, new_n64739_, new_n49115_ );
nor  ( new_n64741_, new_n64740_, new_n49114_ );
nor  ( new_n64742_, new_n64741_, new_n48794_ );
nor  ( new_n64743_, new_n64742_, new_n48793_ );
nor  ( new_n64744_, new_n64743_, new_n48632_ );
nor  ( new_n64745_, new_n64744_, new_n48631_ );
nor  ( new_n64746_, new_n64745_, new_n48209_ );
nor  ( new_n64747_, new_n64746_, new_n48208_ );
nor  ( new_n64748_, new_n64747_, new_n48156_ );
nor  ( new_n64749_, new_n64748_, new_n48155_ );
nor  ( new_n64750_, new_n64749_, new_n47915_ );
not  ( new_n64751_, new_n64750_ );
and  ( new_n64752_, new_n47912_, new_n47874_ );
nor  ( new_n64753_, new_n47912_, new_n47874_ );
nor  ( new_n64754_, new_n64753_, new_n47840_ );
nor  ( new_n64755_, new_n64754_, new_n64752_ );
xor  ( new_n64756_, new_n46862_, new_n46861_ );
not  ( new_n64757_, new_n64756_ );
or   ( new_n64758_, new_n47862_, new_n47858_ );
and  ( new_n64759_, new_n47862_, new_n47858_ );
or   ( new_n64760_, new_n64759_, new_n47857_ );
and  ( new_n64761_, new_n64760_, new_n64758_ );
xor  ( new_n64762_, new_n64761_, new_n64757_ );
xnor ( new_n64763_, new_n46542_, new_n46541_ );
nand ( new_n64764_, new_n47855_, new_n47850_ );
nor  ( new_n64765_, new_n47855_, new_n47850_ );
or   ( new_n64766_, new_n64765_, new_n47845_ );
and  ( new_n64767_, new_n64766_, new_n64764_ );
xor  ( new_n64768_, new_n64767_, new_n64763_ );
xor  ( new_n64769_, new_n46680_, new_n46679_ );
xor  ( new_n64770_, new_n64769_, new_n46686_ );
xor  ( new_n64771_, new_n64770_, new_n64768_ );
xor  ( new_n64772_, new_n64771_, new_n64762_ );
nand ( new_n64773_, new_n47908_, new_n47888_ );
nor  ( new_n64774_, new_n47908_, new_n47888_ );
or   ( new_n64775_, new_n64774_, new_n47885_ );
and  ( new_n64776_, new_n64775_, new_n64773_ );
xnor ( new_n64777_, new_n46843_, new_n46842_ );
nor  ( new_n64778_, new_n47905_, new_n47903_ );
nand ( new_n64779_, new_n47870_, new_n47866_ );
or   ( new_n64780_, new_n47870_, new_n47866_ );
nand ( new_n64781_, new_n64780_, new_n47865_ );
and  ( new_n64782_, new_n64781_, new_n64779_ );
xor  ( new_n64783_, new_n64782_, new_n64778_ );
xor  ( new_n64784_, new_n64783_, new_n64777_ );
xor  ( new_n64785_, new_n64784_, new_n64776_ );
xor  ( new_n64786_, new_n64785_, new_n64772_ );
not  ( new_n64787_, new_n64786_ );
nand ( new_n64788_, new_n47872_, new_n47864_ );
nand ( new_n64789_, new_n47873_, new_n47843_ );
and  ( new_n64790_, new_n64789_, new_n64788_ );
nand ( new_n64791_, new_n47910_, new_n47881_ );
nor  ( new_n64792_, new_n47910_, new_n47881_ );
or   ( new_n64793_, new_n64792_, new_n47878_ );
and  ( new_n64794_, new_n64793_, new_n64791_ );
xor  ( new_n64795_, new_n64794_, new_n64790_ );
xor  ( new_n64796_, new_n64795_, new_n64787_ );
nor  ( new_n64797_, new_n64796_, new_n64755_ );
and  ( new_n64798_, new_n47914_, new_n47836_ );
nor  ( new_n64799_, new_n64798_, new_n64797_ );
and  ( new_n64800_, new_n64799_, new_n64751_ );
not  ( new_n64801_, new_n64800_ );
nor  ( new_n64802_, new_n64761_, new_n64757_ );
and  ( new_n64803_, new_n64771_, new_n64762_ );
nor  ( new_n64804_, new_n64803_, new_n64802_ );
not  ( new_n64805_, new_n64804_ );
xnor ( new_n64806_, new_n46865_, new_n46864_ );
or   ( new_n64807_, new_n64782_, new_n64778_ );
and  ( new_n64808_, new_n64782_, new_n64778_ );
or   ( new_n64809_, new_n64808_, new_n64777_ );
and  ( new_n64810_, new_n64809_, new_n64807_ );
xor  ( new_n64811_, new_n64810_, new_n64806_ );
xor  ( new_n64812_, new_n64811_, new_n64805_ );
nor  ( new_n64813_, new_n64767_, new_n64763_ );
and  ( new_n64814_, new_n64770_, new_n64768_ );
nor  ( new_n64815_, new_n64814_, new_n64813_ );
xor  ( new_n64816_, new_n46696_, new_n46691_ );
xor  ( new_n64817_, new_n46545_, new_n46544_ );
xor  ( new_n64818_, new_n64817_, new_n46547_ );
xnor ( new_n64819_, new_n64818_, new_n64816_ );
xnor ( new_n64820_, new_n64819_, new_n64815_ );
or   ( new_n64821_, new_n64784_, new_n64776_ );
nand ( new_n64822_, new_n64784_, new_n64776_ );
nand ( new_n64823_, new_n64822_, new_n64772_ );
and  ( new_n64824_, new_n64823_, new_n64821_ );
xor  ( new_n64825_, new_n64824_, new_n64820_ );
xor  ( new_n64826_, new_n64825_, new_n64812_ );
not  ( new_n64827_, new_n64826_ );
nor  ( new_n64828_, new_n64794_, new_n64790_ );
and  ( new_n64829_, new_n64794_, new_n64790_ );
nor  ( new_n64830_, new_n64829_, new_n64787_ );
nor  ( new_n64831_, new_n64830_, new_n64828_ );
and  ( new_n64832_, new_n64831_, new_n64827_ );
and  ( new_n64833_, new_n64796_, new_n64755_ );
nor  ( new_n64834_, new_n64833_, new_n64832_ );
and  ( new_n64835_, new_n64834_, new_n64801_ );
nand ( new_n64836_, new_n64818_, new_n64816_ );
or   ( new_n64837_, new_n64819_, new_n64815_ );
and  ( new_n64838_, new_n64837_, new_n64836_ );
or   ( new_n64839_, new_n64810_, new_n64806_ );
nand ( new_n64840_, new_n64811_, new_n64805_ );
and  ( new_n64841_, new_n64840_, new_n64839_ );
nor  ( new_n64842_, new_n64841_, new_n64838_ );
xor  ( new_n64843_, new_n46872_, new_n46871_ );
xor  ( new_n64844_, new_n64841_, new_n64838_ );
and  ( new_n64845_, new_n64844_, new_n64843_ );
nor  ( new_n64846_, new_n64845_, new_n64842_ );
xor  ( new_n64847_, new_n46715_, new_n46713_ );
xor  ( new_n64848_, new_n64847_, new_n46874_ );
and  ( new_n64849_, new_n64848_, new_n64846_ );
not  ( new_n64850_, new_n64849_ );
nor  ( new_n64851_, new_n64824_, new_n64820_ );
and  ( new_n64852_, new_n64825_, new_n64812_ );
nor  ( new_n64853_, new_n64852_, new_n64851_ );
xor  ( new_n64854_, new_n64844_, new_n64843_ );
not  ( new_n64855_, new_n64854_ );
nand ( new_n64856_, new_n64855_, new_n64853_ );
and  ( new_n64857_, new_n64856_, new_n64850_ );
and  ( new_n64858_, new_n64857_, new_n64835_ );
and  ( new_n64859_, new_n64858_, new_n46877_ );
nand ( new_n64860_, new_n64859_, new_n46709_ );
nor  ( new_n64861_, new_n64860_, new_n46030_ );
not  ( new_n64862_, new_n64861_ );
or   ( new_n64863_, new_n45515_, new_n45397_ );
or   ( new_n64864_, new_n46021_, new_n46012_ );
or   ( new_n64865_, new_n64864_, new_n46027_ );
or   ( new_n64866_, new_n46026_, new_n46025_ );
or   ( new_n64867_, new_n45574_, new_n45572_ );
and  ( new_n64868_, new_n64867_, new_n64866_ );
and  ( new_n64869_, new_n64868_, new_n64865_ );
or   ( new_n64870_, new_n64869_, new_n45576_ );
and  ( new_n64871_, new_n64870_, new_n64863_ );
or   ( new_n64872_, new_n46876_, new_n46711_ );
nor  ( new_n64873_, new_n64848_, new_n64846_ );
nor  ( new_n64874_, new_n64855_, new_n64853_ );
nor  ( new_n64875_, new_n64831_, new_n64827_ );
or   ( new_n64876_, new_n64875_, new_n64874_ );
and  ( new_n64877_, new_n64876_, new_n64856_ );
and  ( new_n64878_, new_n64877_, new_n64850_ );
nor  ( new_n64879_, new_n64878_, new_n64873_ );
not  ( new_n64880_, new_n64879_ );
nand ( new_n64881_, new_n64880_, new_n46877_ );
and  ( new_n64882_, new_n64881_, new_n64872_ );
not  ( new_n64883_, new_n64882_ );
nand ( new_n64884_, new_n64883_, new_n46709_ );
or   ( new_n64885_, new_n46336_, new_n46331_ );
and  ( new_n64886_, new_n46329_, new_n46320_ );
and  ( new_n64887_, new_n46529_, new_n46528_ );
and  ( new_n64888_, new_n46706_, new_n46705_ );
and  ( new_n64889_, new_n64888_, new_n46530_ );
or   ( new_n64890_, new_n64889_, new_n64887_ );
or   ( new_n64891_, new_n64890_, new_n64886_ );
nand ( new_n64892_, new_n64891_, new_n46338_ );
and  ( new_n64893_, new_n64892_, new_n64885_ );
and  ( new_n64894_, new_n64893_, new_n64884_ );
or   ( new_n64895_, new_n64894_, new_n46029_ );
and  ( new_n64896_, new_n64895_, new_n64871_ );
nor  ( new_n64897_, new_n64896_, new_n45396_ );
not  ( new_n64898_, new_n64897_ );
or   ( new_n64899_, new_n45296_, new_n45281_ );
or   ( new_n64900_, new_n45394_, new_n45393_ );
or   ( new_n64901_, new_n45277_, new_n45248_ );
and  ( new_n64902_, new_n64901_, new_n64900_ );
or   ( new_n64903_, new_n64902_, new_n45298_ );
and  ( new_n64904_, new_n64903_, new_n64899_ );
and  ( new_n64905_, new_n45294_, new_n45287_ );
nor  ( new_n64906_, new_n45295_, new_n45284_ );
nor  ( new_n64907_, new_n64906_, new_n64905_ );
not  ( new_n64908_, new_n64907_ );
and  ( new_n64909_, new_n45291_, new_n45290_ );
and  ( new_n64910_, new_n45293_, new_n45292_ );
or   ( new_n64911_, new_n64910_, new_n64909_ );
xor  ( new_n64912_, new_n44555_, new_n44554_ );
xor  ( new_n64913_, new_n44735_, new_n44734_ );
xor  ( new_n64914_, new_n64913_, new_n64912_ );
xor  ( new_n64915_, new_n64914_, new_n64911_ );
nand ( new_n64916_, new_n64915_, new_n64908_ );
and  ( new_n64917_, new_n64916_, new_n64904_ );
and  ( new_n64918_, new_n64917_, new_n64898_ );
and  ( new_n64919_, new_n64918_, new_n64862_ );
not  ( new_n64920_, new_n64919_ );
nor  ( new_n64921_, new_n64915_, new_n64908_ );
and  ( new_n64922_, new_n64913_, new_n64912_ );
and  ( new_n64923_, new_n64914_, new_n64911_ );
nor  ( new_n64924_, new_n64923_, new_n64922_ );
xor  ( new_n64925_, new_n44739_, new_n44738_ );
not  ( new_n64926_, new_n64925_ );
and  ( new_n64927_, new_n64926_, new_n64924_ );
nor  ( new_n64928_, new_n64927_, new_n64921_ );
and  ( new_n64929_, new_n64928_, new_n64920_ );
and  ( new_n64930_, new_n64929_, new_n44757_ );
not  ( new_n64931_, new_n64930_ );
nor  ( new_n64932_, new_n64926_, new_n64924_ );
and  ( new_n64933_, new_n44749_, new_n44741_ );
nor  ( new_n64934_, new_n64933_, new_n64932_ );
not  ( new_n64935_, new_n64934_ );
and  ( new_n64936_, new_n64935_, new_n44757_ );
nor  ( new_n64937_, new_n44755_, new_n44753_ );
nor  ( new_n64938_, new_n64937_, new_n64936_ );
and  ( new_n64939_, new_n64938_, new_n64931_ );
nor  ( new_n64940_, new_n64939_, new_n44544_ );
nor  ( new_n64941_, new_n64940_, new_n44543_ );
nor  ( new_n64942_, new_n64941_, new_n44456_ );
and  ( new_n64943_, new_n44455_, new_n44454_ );
nor  ( new_n64944_, new_n64943_, new_n64942_ );
nor  ( new_n64945_, new_n64944_, new_n44303_ );
nor  ( new_n64946_, new_n64945_, new_n44302_ );
or   ( new_n64947_, new_n64946_, new_n44267_ );
and  ( new_n64948_, new_n64947_, new_n44266_ );
xnor ( new_n64949_, new_n64948_, new_n44133_ );
or   ( new_n64950_, new_n64949_, new_n44129_ );
xor  ( new_n64951_, RIbb33f30_217, RIbb33d50_213 );
not  ( new_n64952_, RIbb345c0_231 );
xor  ( new_n64953_, RIbb34bd8_244, new_n64952_ );
xor  ( new_n64954_, RIbb34db8_248, RIbb338a0_203 );
xor  ( new_n64955_, new_n64954_, new_n64953_ );
xnor ( new_n64956_, new_n64955_, new_n64951_ );
xor  ( new_n64957_, RIbb34cc8_246, RIbb347a0_235 );
xnor ( new_n64958_, RIbb34110_221, RIbb33990_205 );
xor  ( new_n64959_, RIbb34d40_247, RIbb33c60_211 );
xor  ( new_n64960_, new_n64959_, new_n64958_ );
xor  ( new_n64961_, new_n64960_, new_n64957_ );
xnor ( new_n64962_, RIbb34098_220, RIbb33a08_206 );
not  ( new_n64963_, RIbb336c0_199 );
xor  ( new_n64964_, RIbb34278_224, new_n64963_ );
xor  ( new_n64965_, new_n64964_, new_n64962_ );
xor  ( new_n64966_, new_n64965_, new_n64961_ );
xor  ( new_n64967_, new_n64966_, new_n64956_ );
xnor ( new_n64968_, RIbb34188_222, RIbb33828_202 );
xnor ( new_n64969_, new_n64968_, new_n64967_ );
xor  ( new_n64970_, RIbb349f8_240, RIbb33738_200 );
not  ( new_n64971_, RIbb33a80_207 );
xor  ( new_n64972_, RIbb34908_238, new_n64971_ );
xor  ( new_n64973_, new_n64972_, new_n64970_ );
not  ( new_n64974_, RIbb346b0_233 );
xor  ( new_n64975_, new_n64974_, RIbb34638_232 );
xnor ( new_n64976_, RIbb34ea8_250, RIbb34548_230 );
xor  ( new_n64977_, RIbb35010_253, RIbb334e0_195 );
xor  ( new_n64978_, new_n64977_, new_n64976_ );
xor  ( new_n64979_, new_n64978_, new_n64975_ );
xor  ( new_n64980_, new_n64979_, new_n64973_ );
xnor ( new_n64981_, RIbb34980_239, RIbb33918_204 );
xor  ( new_n64982_, RIbb35088_254, RIbb34728_234 );
xor  ( new_n64983_, new_n64982_, new_n64981_ );
xor  ( new_n64984_, new_n64983_, new_n64980_ );
xor  ( new_n64985_, new_n64984_, new_n64969_ );
not  ( new_n64986_, RIbb342f0_225 );
xor  ( new_n64987_, new_n64986_, RIbb33648_198 );
xor  ( new_n64988_, new_n64987_, RIbb34c50_245 );
xnor ( new_n64989_, RIbb34890_237, RIbb33cd8_212 );
xor  ( new_n64990_, new_n64989_, new_n64988_ );
xnor ( new_n64991_, new_n64990_, new_n64985_ );
xor  ( new_n64992_, RIbb35100_255, RIbb33468_194 );
xnor ( new_n64993_, RIbb34818_236, RIbb33eb8_216 );
xor  ( new_n64994_, new_n64993_, new_n64992_ );
xor  ( new_n64995_, RIbb34b60_243, RIbb344d0_229 );
xnor ( new_n64996_, RIbb34ae8_242, RIbb34458_228 );
xor  ( new_n64997_, RIbb34e30_249, RIbb33558_196 );
xor  ( new_n64998_, new_n64997_, new_n64996_ );
xor  ( new_n64999_, new_n64998_, new_n64995_ );
xor  ( new_n65000_, RIbb343e0_227, RIbb34368_226 );
not  ( new_n65001_, RIbb333f0_193 );
xor  ( new_n65002_, RIbb35178_256, new_n65001_ );
xor  ( new_n65003_, RIbb34a70_241, RIbb335d0_197 );
xor  ( new_n65004_, new_n65003_, new_n65002_ );
xor  ( new_n65005_, new_n65004_, new_n65000_ );
not  ( new_n65006_, RIbb34020_219 );
xor  ( new_n65007_, new_n65006_, RIbb33af8_208 );
not  ( new_n65008_, RIbb33b70_209 );
xor  ( new_n65009_, RIbb33fa8_218, new_n65008_ );
xor  ( new_n65010_, new_n65009_, new_n65007_ );
xor  ( new_n65011_, new_n65010_, new_n65005_ );
xor  ( new_n65012_, new_n65011_, new_n64999_ );
not  ( new_n65013_, RIbb337b0_201 );
xor  ( new_n65014_, RIbb34200_223, new_n65013_ );
xor  ( new_n65015_, new_n65014_, new_n65012_ );
xor  ( new_n65016_, new_n65015_, new_n64994_ );
xnor ( new_n65017_, RIbb33e40_215, RIbb33dc8_214 );
not  ( new_n65018_, RIbb34f20_251 );
xor  ( new_n65019_, RIbb34f98_252, RIbb33be8_210 );
xor  ( new_n65020_, new_n65019_, new_n65018_ );
xor  ( new_n65021_, new_n65020_, new_n65017_ );
xor  ( new_n65022_, new_n65021_, new_n65016_ );
xor  ( new_n65023_, new_n65022_, new_n64991_ );
nand ( new_n65024_, new_n64949_, new_n44129_ );
and  ( new_n65025_, new_n65024_, new_n65023_ );
and  ( new_n65026_, new_n65025_, new_n64950_ );
xnor ( new_n65027_, new_n65026_, new_n43446_ );
or   ( new_n65028_, new_n42726_, new_n42724_ );
and  ( new_n65029_, new_n42726_, new_n42724_ );
or   ( new_n65030_, new_n42731_, new_n65029_ );
and  ( new_n65031_, new_n65030_, new_n65028_ );
not  ( new_n65032_, new_n21693_ );
nand ( new_n65033_, new_n21710_, new_n65032_ );
or   ( new_n65034_, new_n283_, new_n21701_ );
or   ( new_n65035_, new_n286_, new_n21703_ );
and  ( new_n65036_, new_n65035_, new_n65034_ );
or   ( new_n65037_, new_n317_, new_n21694_ );
or   ( new_n65038_, new_n320_, new_n21696_ );
and  ( new_n65039_, new_n65038_, new_n65037_ );
xor  ( new_n65040_, new_n65039_, new_n278_ );
xor  ( new_n65041_, new_n65040_, new_n65036_ );
xor  ( new_n65042_, new_n65041_, new_n65033_ );
xor  ( new_n65043_, new_n65042_, new_n65031_ );
and  ( new_n65044_, new_n42733_, new_n42719_ );
and  ( new_n65045_, new_n42734_, new_n42718_ );
or   ( new_n65046_, new_n65045_, new_n65044_ );
and  ( new_n65047_, new_n267_, RIbb31938_136 );
and  ( new_n65048_, new_n265_, RIbb318c0_135 );
or   ( new_n65049_, new_n65048_, new_n65047_ );
and  ( new_n65050_, RIbb319b0_137, RIbb2f610_1 );
xnor ( new_n65051_, new_n65050_, new_n65049_ );
xor  ( new_n65052_, new_n65051_, new_n21626_ );
xor  ( new_n65053_, new_n65052_, new_n65046_ );
xor  ( new_n65054_, new_n65053_, new_n65043_ );
or   ( new_n65055_, new_n42732_, new_n42723_ );
and  ( new_n65056_, new_n298_, RIbb31848_134 );
and  ( new_n65057_, new_n295_, RIbb317d0_133 );
or   ( new_n65058_, new_n65057_, new_n65056_ );
not  ( new_n65059_, new_n21780_ );
not  ( new_n65060_, new_n21784_ );
and  ( new_n65061_, new_n65060_, new_n65059_ );
or   ( new_n65062_, new_n65060_, new_n65059_ );
and  ( new_n65063_, new_n65062_, new_n21776_ );
or   ( new_n65064_, new_n65063_, new_n65061_ );
or   ( new_n65065_, new_n21722_, new_n21719_ );
and  ( new_n65066_, new_n21722_, new_n21719_ );
or   ( new_n65067_, new_n65066_, new_n21715_ );
and  ( new_n65068_, new_n65067_, new_n65065_ );
xor  ( new_n65069_, new_n65068_, new_n65064_ );
xor  ( new_n65070_, new_n65069_, new_n65058_ );
xor  ( new_n65071_, new_n65070_, new_n65055_ );
xor  ( new_n65072_, new_n65071_, new_n65054_ );
xnor ( new_n65073_, new_n65072_, new_n65027_ );
nor  ( new_n65074_, new_n65073_, new_n21791_ );
and  ( new_n65075_, new_n65073_, new_n21791_ );
xor  ( new_n65076_, new_n43441_, new_n42735_ );
xnor ( new_n65077_, new_n44265_, new_n44264_ );
xor  ( new_n65078_, new_n65077_, new_n64946_ );
and  ( new_n65079_, new_n65078_, new_n65023_ );
xnor ( new_n65080_, new_n65079_, new_n43444_ );
nor  ( new_n65081_, new_n65080_, new_n65076_ );
and  ( new_n65082_, new_n65080_, new_n65076_ );
xor  ( new_n65083_, new_n42738_, new_n42737_ );
xnor ( new_n65084_, new_n65083_, new_n43434_ );
not  ( new_n65085_, new_n65023_ );
xor  ( new_n65086_, new_n44455_, new_n44454_ );
xor  ( new_n65087_, new_n65086_, new_n64941_ );
nor  ( new_n65088_, new_n65087_, new_n65085_ );
nor  ( new_n65089_, new_n65088_, new_n65084_ );
and  ( new_n65090_, new_n65088_, new_n65084_ );
xor  ( new_n65091_, new_n42743_, new_n42742_ );
xnor ( new_n65092_, new_n65091_, new_n43421_ );
nor  ( new_n65093_, new_n64932_, new_n64929_ );
xor  ( new_n65094_, new_n44749_, new_n44741_ );
xor  ( new_n65095_, new_n65094_, new_n65093_ );
nor  ( new_n65096_, new_n65095_, new_n65085_ );
nor  ( new_n65097_, new_n65096_, new_n65092_ );
and  ( new_n65098_, new_n65096_, new_n65092_ );
xor  ( new_n65099_, new_n42748_, new_n42747_ );
xnor ( new_n65100_, new_n65099_, new_n43414_ );
xor  ( new_n65101_, new_n64915_, new_n64907_ );
and  ( new_n65102_, new_n64894_, new_n64860_ );
or   ( new_n65103_, new_n65102_, new_n46030_ );
or   ( new_n65104_, new_n64871_, new_n45396_ );
and  ( new_n65105_, new_n65104_, new_n64904_ );
and  ( new_n65106_, new_n65105_, new_n65103_ );
xor  ( new_n65107_, new_n65106_, new_n65101_ );
and  ( new_n65108_, new_n65107_, new_n65023_ );
nor  ( new_n65109_, new_n65108_, new_n65100_ );
and  ( new_n65110_, new_n65108_, new_n65100_ );
xor  ( new_n65111_, new_n42753_, new_n42752_ );
xnor ( new_n65112_, new_n65111_, new_n43371_ );
xor  ( new_n65113_, new_n46336_, new_n46331_ );
or   ( new_n65114_, new_n64883_, new_n64859_ );
and  ( new_n65115_, new_n65114_, new_n46708_ );
or   ( new_n65116_, new_n65115_, new_n64891_ );
and  ( new_n65117_, new_n65116_, new_n46330_ );
xor  ( new_n65118_, new_n65117_, new_n65113_ );
and  ( new_n65119_, new_n65118_, new_n65023_ );
nor  ( new_n65120_, new_n65119_, new_n65112_ );
and  ( new_n65121_, new_n65119_, new_n65112_ );
xor  ( new_n65122_, new_n42758_, new_n42757_ );
xnor ( new_n65123_, new_n65122_, new_n43357_ );
xor  ( new_n65124_, new_n46706_, new_n46705_ );
xor  ( new_n65125_, new_n65124_, new_n65114_ );
and  ( new_n65126_, new_n65125_, new_n65023_ );
nor  ( new_n65127_, new_n65126_, new_n65123_ );
and  ( new_n65128_, new_n65126_, new_n65123_ );
xor  ( new_n65129_, new_n42761_, new_n42760_ );
xnor ( new_n65130_, new_n65129_, new_n43355_ );
nor  ( new_n65131_, new_n64880_, new_n64858_ );
xor  ( new_n65132_, new_n46876_, new_n46711_ );
xor  ( new_n65133_, new_n65132_, new_n65131_ );
nor  ( new_n65134_, new_n65133_, new_n65085_ );
nor  ( new_n65135_, new_n65134_, new_n65130_ );
and  ( new_n65136_, new_n65134_, new_n65130_ );
xor  ( new_n65137_, new_n42766_, new_n42765_ );
xnor ( new_n65138_, new_n65137_, new_n43348_ );
nor  ( new_n65139_, new_n64875_, new_n64835_ );
xor  ( new_n65140_, new_n64855_, new_n64853_ );
xor  ( new_n65141_, new_n65140_, new_n65139_ );
nor  ( new_n65142_, new_n65141_, new_n65085_ );
nor  ( new_n65143_, new_n65142_, new_n65138_ );
and  ( new_n65144_, new_n65142_, new_n65138_ );
xor  ( new_n65145_, new_n42771_, new_n42770_ );
xnor ( new_n65146_, new_n65145_, new_n43334_ );
xnor ( new_n65147_, new_n47914_, new_n47836_ );
xor  ( new_n65148_, new_n65147_, new_n64749_ );
and  ( new_n65149_, new_n65148_, new_n65023_ );
nor  ( new_n65150_, new_n65149_, new_n65146_ );
and  ( new_n65151_, new_n65149_, new_n65146_ );
xnor ( new_n65152_, new_n42774_, new_n42773_ );
xnor ( new_n65153_, new_n48154_, new_n48152_ );
xor  ( new_n65154_, new_n65153_, new_n64747_ );
nand ( new_n65155_, new_n65154_, new_n65023_ );
xor  ( new_n65156_, new_n65155_, new_n43332_ );
xor  ( new_n65157_, new_n65156_, new_n65152_ );
xor  ( new_n65158_, new_n48207_, new_n48205_ );
xor  ( new_n65159_, new_n65158_, new_n64745_ );
nor  ( new_n65160_, new_n65159_, new_n65085_ );
xor  ( new_n65161_, new_n43327_, new_n42777_ );
xor  ( new_n65162_, new_n65161_, new_n43330_ );
not  ( new_n65163_, new_n65162_ );
nor  ( new_n65164_, new_n65163_, new_n65160_ );
and  ( new_n65165_, new_n65163_, new_n65160_ );
xor  ( new_n65166_, new_n42779_, new_n42778_ );
xnor ( new_n65167_, new_n65166_, new_n43325_ );
xor  ( new_n65168_, new_n48630_, new_n48210_ );
xor  ( new_n65169_, new_n65168_, new_n64743_ );
nor  ( new_n65170_, new_n65169_, new_n65085_ );
nor  ( new_n65171_, new_n65170_, new_n65167_ );
and  ( new_n65172_, new_n65170_, new_n65167_ );
xor  ( new_n65173_, new_n42784_, new_n42783_ );
xnor ( new_n65174_, new_n65173_, new_n43317_ );
xnor ( new_n65175_, new_n49113_, new_n49112_ );
xor  ( new_n65176_, new_n65175_, new_n64739_ );
and  ( new_n65177_, new_n65176_, new_n65023_ );
nor  ( new_n65178_, new_n65177_, new_n65174_ );
and  ( new_n65179_, new_n65177_, new_n65174_ );
xor  ( new_n65180_, new_n42787_, new_n42786_ );
xnor ( new_n65181_, new_n65180_, new_n43314_ );
xor  ( new_n65182_, new_n49359_, new_n49116_ );
and  ( new_n65183_, new_n65182_, new_n64736_ );
not  ( new_n65184_, new_n65183_ );
or   ( new_n65185_, new_n65182_, new_n64736_ );
and  ( new_n65186_, new_n65185_, new_n65023_ );
and  ( new_n65187_, new_n65186_, new_n65184_ );
nor  ( new_n65188_, new_n65187_, new_n65181_ );
and  ( new_n65189_, new_n65187_, new_n65181_ );
xor  ( new_n65190_, new_n42790_, new_n42789_ );
xnor ( new_n65191_, new_n65190_, new_n43312_ );
xor  ( new_n65192_, new_n49617_, new_n49615_ );
and  ( new_n65193_, new_n65192_, new_n64734_ );
not  ( new_n65194_, new_n65193_ );
or   ( new_n65195_, new_n65192_, new_n64734_ );
and  ( new_n65196_, new_n65195_, new_n65023_ );
and  ( new_n65197_, new_n65196_, new_n65194_ );
nor  ( new_n65198_, new_n65197_, new_n65191_ );
and  ( new_n65199_, new_n65197_, new_n65191_ );
xor  ( new_n65200_, new_n42795_, new_n42794_ );
xnor ( new_n65201_, new_n65200_, new_n43304_ );
xor  ( new_n65202_, new_n50153_, new_n50152_ );
and  ( new_n65203_, new_n65202_, new_n64730_ );
not  ( new_n65204_, new_n65203_ );
or   ( new_n65205_, new_n65202_, new_n64730_ );
and  ( new_n65206_, new_n65205_, new_n65023_ );
and  ( new_n65207_, new_n65206_, new_n65204_ );
nor  ( new_n65208_, new_n65207_, new_n65201_ );
and  ( new_n65209_, new_n65207_, new_n65201_ );
xor  ( new_n65210_, new_n42798_, new_n42797_ );
xnor ( new_n65211_, new_n65210_, new_n43302_ );
xor  ( new_n65212_, new_n50292_, new_n50157_ );
and  ( new_n65213_, new_n65212_, new_n64728_ );
not  ( new_n65214_, new_n65213_ );
or   ( new_n65215_, new_n65212_, new_n64728_ );
and  ( new_n65216_, new_n65215_, new_n65023_ );
and  ( new_n65217_, new_n65216_, new_n65214_ );
nor  ( new_n65218_, new_n65217_, new_n65211_ );
and  ( new_n65219_, new_n65217_, new_n65211_ );
xor  ( new_n65220_, new_n42803_, new_n42802_ );
xnor ( new_n65221_, new_n65220_, new_n43294_ );
xor  ( new_n65222_, new_n50866_, new_n50865_ );
xor  ( new_n65223_, new_n65222_, new_n64724_ );
and  ( new_n65224_, new_n65223_, new_n65023_ );
nor  ( new_n65225_, new_n65224_, new_n65221_ );
and  ( new_n65226_, new_n65224_, new_n65221_ );
xor  ( new_n65227_, new_n42806_, new_n42805_ );
xnor ( new_n65228_, new_n65227_, new_n43291_ );
xor  ( new_n65229_, new_n51259_, new_n51258_ );
and  ( new_n65230_, new_n65229_, new_n64722_ );
not  ( new_n65231_, new_n65230_ );
or   ( new_n65232_, new_n65229_, new_n64722_ );
and  ( new_n65233_, new_n65232_, new_n65023_ );
and  ( new_n65234_, new_n65233_, new_n65231_ );
nor  ( new_n65235_, new_n65234_, new_n65228_ );
and  ( new_n65236_, new_n65234_, new_n65228_ );
xor  ( new_n65237_, new_n42809_, new_n42808_ );
xnor ( new_n65238_, new_n65237_, new_n43288_ );
xor  ( new_n65239_, new_n51520_, new_n51263_ );
and  ( new_n65240_, new_n65239_, new_n64720_ );
not  ( new_n65241_, new_n65240_ );
or   ( new_n65242_, new_n65239_, new_n64720_ );
and  ( new_n65243_, new_n65242_, new_n65023_ );
and  ( new_n65244_, new_n65243_, new_n65241_ );
nor  ( new_n65245_, new_n65244_, new_n65238_ );
and  ( new_n65246_, new_n65244_, new_n65238_ );
xor  ( new_n65247_, new_n42812_, new_n42811_ );
xnor ( new_n65248_, new_n65247_, new_n43286_ );
xor  ( new_n65249_, new_n51830_, new_n51828_ );
and  ( new_n65250_, new_n65249_, new_n64718_ );
not  ( new_n65251_, new_n65250_ );
or   ( new_n65252_, new_n65249_, new_n64718_ );
and  ( new_n65253_, new_n65252_, new_n65023_ );
and  ( new_n65254_, new_n65253_, new_n65251_ );
nor  ( new_n65255_, new_n65254_, new_n65248_ );
and  ( new_n65256_, new_n65254_, new_n65248_ );
xor  ( new_n65257_, new_n42817_, new_n42816_ );
xnor ( new_n65258_, new_n65257_, new_n43266_ );
xor  ( new_n65259_, new_n52835_, new_n52815_ );
xor  ( new_n65260_, new_n65259_, new_n64679_ );
and  ( new_n65261_, new_n65260_, new_n65023_ );
nor  ( new_n65262_, new_n65261_, new_n65258_ );
and  ( new_n65263_, new_n65261_, new_n65258_ );
xor  ( new_n65264_, new_n42820_, new_n42819_ );
xnor ( new_n65265_, new_n65264_, new_n43263_ );
xor  ( new_n65266_, new_n53264_, new_n53262_ );
xor  ( new_n65267_, new_n65266_, new_n64676_ );
and  ( new_n65268_, new_n65267_, new_n65023_ );
nor  ( new_n65269_, new_n65268_, new_n65265_ );
and  ( new_n65270_, new_n65268_, new_n65265_ );
xor  ( new_n65271_, new_n42823_, new_n42822_ );
xnor ( new_n65272_, new_n65271_, new_n43260_ );
xor  ( new_n65273_, new_n53557_, new_n53555_ );
and  ( new_n65274_, new_n65273_, new_n64674_ );
not  ( new_n65275_, new_n65274_ );
or   ( new_n65276_, new_n65273_, new_n64674_ );
and  ( new_n65277_, new_n65276_, new_n65023_ );
and  ( new_n65278_, new_n65277_, new_n65275_ );
nor  ( new_n65279_, new_n65278_, new_n65272_ );
and  ( new_n65280_, new_n65278_, new_n65272_ );
xor  ( new_n65281_, new_n42826_, new_n42825_ );
xnor ( new_n65282_, new_n65281_, new_n43257_ );
xor  ( new_n65283_, new_n53987_, new_n53986_ );
xnor ( new_n65284_, new_n65283_, new_n64672_ );
nor  ( new_n65285_, new_n65284_, new_n65085_ );
nor  ( new_n65286_, new_n65285_, new_n65282_ );
and  ( new_n65287_, new_n65285_, new_n65282_ );
xor  ( new_n65288_, new_n42829_, new_n42828_ );
xnor ( new_n65289_, new_n65288_, new_n43255_ );
xor  ( new_n65290_, new_n54255_, new_n54254_ );
xor  ( new_n65291_, new_n65290_, new_n64669_ );
nor  ( new_n65292_, new_n65291_, new_n65085_ );
nor  ( new_n65293_, new_n65292_, new_n65289_ );
and  ( new_n65294_, new_n65292_, new_n65289_ );
xor  ( new_n65295_, new_n42834_, new_n42833_ );
xnor ( new_n65296_, new_n65295_, new_n43248_ );
nor  ( new_n65297_, new_n64661_, new_n64652_ );
xor  ( new_n65298_, new_n64659_, new_n64655_ );
xor  ( new_n65299_, new_n65298_, new_n65297_ );
nor  ( new_n65300_, new_n65299_, new_n65085_ );
nor  ( new_n65301_, new_n65300_, new_n65296_ );
and  ( new_n65302_, new_n65300_, new_n65296_ );
xor  ( new_n65303_, new_n42839_, new_n42838_ );
xnor ( new_n65304_, new_n65303_, new_n43240_ );
xor  ( new_n65305_, new_n55453_, new_n55338_ );
and  ( new_n65306_, new_n65305_, new_n64633_ );
not  ( new_n65307_, new_n65306_ );
or   ( new_n65308_, new_n65305_, new_n64633_ );
and  ( new_n65309_, new_n65308_, new_n65023_ );
and  ( new_n65310_, new_n65309_, new_n65307_ );
nor  ( new_n65311_, new_n65310_, new_n65304_ );
and  ( new_n65312_, new_n65310_, new_n65304_ );
xor  ( new_n65313_, new_n42842_, new_n42841_ );
xnor ( new_n65314_, new_n65313_, new_n43237_ );
xor  ( new_n65315_, new_n55727_, new_n55725_ );
and  ( new_n65316_, new_n65315_, new_n64631_ );
not  ( new_n65317_, new_n65316_ );
or   ( new_n65318_, new_n65315_, new_n64631_ );
and  ( new_n65319_, new_n65318_, new_n65023_ );
and  ( new_n65320_, new_n65319_, new_n65317_ );
nor  ( new_n65321_, new_n65320_, new_n65314_ );
and  ( new_n65322_, new_n65320_, new_n65314_ );
xor  ( new_n65323_, new_n42845_, new_n42844_ );
xnor ( new_n65324_, new_n65323_, new_n43234_ );
or   ( new_n65325_, new_n64627_, new_n64625_ );
xor  ( new_n65326_, new_n55961_, new_n55730_ );
xor  ( new_n65327_, new_n65326_, new_n65325_ );
and  ( new_n65328_, new_n65327_, new_n65023_ );
nor  ( new_n65329_, new_n65328_, new_n65324_ );
and  ( new_n65330_, new_n65328_, new_n65324_ );
xor  ( new_n65331_, new_n42848_, new_n42847_ );
xnor ( new_n65332_, new_n65331_, new_n43231_ );
xor  ( new_n65333_, new_n56359_, new_n56356_ );
and  ( new_n65334_, new_n65333_, new_n64624_ );
not  ( new_n65335_, new_n65334_ );
or   ( new_n65336_, new_n65333_, new_n64624_ );
and  ( new_n65337_, new_n65336_, new_n65023_ );
and  ( new_n65338_, new_n65337_, new_n65335_ );
nor  ( new_n65339_, new_n65338_, new_n65332_ );
and  ( new_n65340_, new_n65338_, new_n65332_ );
xor  ( new_n65341_, new_n42851_, new_n42850_ );
xnor ( new_n65342_, new_n65341_, new_n43229_ );
and  ( new_n65343_, new_n65085_, RIbb2f610_1 );
not  ( new_n65344_, new_n64621_ );
xor  ( new_n65345_, new_n56571_, new_n56363_ );
and  ( new_n65346_, new_n65345_, new_n65344_ );
not  ( new_n65347_, new_n65346_ );
or   ( new_n65348_, new_n65345_, new_n65344_ );
and  ( new_n65349_, new_n65348_, new_n65023_ );
and  ( new_n65350_, new_n65349_, new_n65347_ );
nor  ( new_n65351_, new_n65350_, new_n65343_ );
not  ( new_n65352_, new_n65351_ );
nor  ( new_n65353_, new_n65352_, new_n65342_ );
and  ( new_n65354_, new_n65352_, new_n65342_ );
xor  ( new_n65355_, new_n42856_, new_n42855_ );
xnor ( new_n65356_, new_n65355_, new_n43221_ );
and  ( new_n65357_, new_n65085_, RIbb2f520_3 );
xor  ( new_n65358_, new_n57123_, new_n56881_ );
and  ( new_n65359_, new_n65358_, new_n64616_ );
not  ( new_n65360_, new_n65359_ );
or   ( new_n65361_, new_n65358_, new_n64616_ );
and  ( new_n65362_, new_n65361_, new_n65023_ );
and  ( new_n65363_, new_n65362_, new_n65360_ );
nor  ( new_n65364_, new_n65363_, new_n65357_ );
not  ( new_n65365_, new_n65364_ );
nor  ( new_n65366_, new_n65365_, new_n65356_ );
and  ( new_n65367_, new_n65365_, new_n65356_ );
xor  ( new_n65368_, new_n42859_, new_n42858_ );
xnor ( new_n65369_, new_n65368_, new_n43218_ );
and  ( new_n65370_, new_n65085_, RIbb2f4a8_4 );
xor  ( new_n65371_, new_n57375_, new_n57128_ );
and  ( new_n65372_, new_n65371_, new_n64614_ );
not  ( new_n65373_, new_n65372_ );
or   ( new_n65374_, new_n65371_, new_n64614_ );
and  ( new_n65375_, new_n65374_, new_n65023_ );
and  ( new_n65376_, new_n65375_, new_n65373_ );
nor  ( new_n65377_, new_n65376_, new_n65370_ );
not  ( new_n65378_, new_n65377_ );
nor  ( new_n65379_, new_n65378_, new_n65369_ );
and  ( new_n65380_, new_n65378_, new_n65369_ );
xor  ( new_n65381_, new_n42862_, new_n42861_ );
xnor ( new_n65382_, new_n65381_, new_n43215_ );
and  ( new_n65383_, new_n65085_, RIbb2f430_5 );
xor  ( new_n65384_, new_n57684_, new_n57379_ );
and  ( new_n65385_, new_n65384_, new_n64610_ );
not  ( new_n65386_, new_n65385_ );
or   ( new_n65387_, new_n65384_, new_n64610_ );
and  ( new_n65388_, new_n65387_, new_n65023_ );
and  ( new_n65389_, new_n65388_, new_n65386_ );
nor  ( new_n65390_, new_n65389_, new_n65383_ );
not  ( new_n65391_, new_n65390_ );
nor  ( new_n65392_, new_n65391_, new_n65382_ );
and  ( new_n65393_, new_n65391_, new_n65382_ );
xor  ( new_n65394_, new_n42865_, new_n42864_ );
xnor ( new_n65395_, new_n65394_, new_n43212_ );
and  ( new_n65396_, new_n65085_, RIbb2f3b8_6 );
xor  ( new_n65397_, new_n57796_, new_n57794_ );
and  ( new_n65398_, new_n65397_, new_n64608_ );
not  ( new_n65399_, new_n65398_ );
or   ( new_n65400_, new_n65397_, new_n64608_ );
and  ( new_n65401_, new_n65400_, new_n65023_ );
and  ( new_n65402_, new_n65401_, new_n65399_ );
nor  ( new_n65403_, new_n65402_, new_n65396_ );
not  ( new_n65404_, new_n65403_ );
nor  ( new_n65405_, new_n65404_, new_n65395_ );
and  ( new_n65406_, new_n65404_, new_n65395_ );
xor  ( new_n65407_, new_n42868_, new_n42867_ );
xnor ( new_n65408_, new_n65407_, new_n43209_ );
and  ( new_n65409_, new_n65085_, RIbb2f340_7 );
xor  ( new_n65410_, new_n58262_, new_n58260_ );
not  ( new_n65411_, new_n65410_ );
and  ( new_n65412_, new_n65411_, new_n64605_ );
not  ( new_n65413_, new_n65412_ );
or   ( new_n65414_, new_n65411_, new_n64605_ );
and  ( new_n65415_, new_n65414_, new_n65023_ );
and  ( new_n65416_, new_n65415_, new_n65413_ );
nor  ( new_n65417_, new_n65416_, new_n65409_ );
not  ( new_n65418_, new_n65417_ );
nor  ( new_n65419_, new_n65418_, new_n65408_ );
and  ( new_n65420_, new_n65418_, new_n65408_ );
xor  ( new_n65421_, new_n42871_, new_n42870_ );
xnor ( new_n65422_, new_n65421_, new_n43206_ );
and  ( new_n65423_, new_n65085_, RIbb2f2c8_8 );
not  ( new_n65424_, new_n64602_ );
xor  ( new_n65425_, new_n58363_, new_n58265_ );
and  ( new_n65426_, new_n65425_, new_n65424_ );
not  ( new_n65427_, new_n65426_ );
or   ( new_n65428_, new_n65425_, new_n65424_ );
and  ( new_n65429_, new_n65428_, new_n65023_ );
and  ( new_n65430_, new_n65429_, new_n65427_ );
nor  ( new_n65431_, new_n65430_, new_n65423_ );
not  ( new_n65432_, new_n65431_ );
nor  ( new_n65433_, new_n65432_, new_n65422_ );
and  ( new_n65434_, new_n65432_, new_n65422_ );
xor  ( new_n65435_, new_n42874_, new_n42873_ );
xnor ( new_n65436_, new_n65435_, new_n43203_ );
xor  ( new_n65437_, new_n58651_, new_n58648_ );
or   ( new_n65438_, new_n64598_, new_n64596_ );
and  ( new_n65439_, new_n65438_, new_n65437_ );
not  ( new_n65440_, new_n58652_ );
and  ( new_n65441_, new_n64601_, new_n65440_ );
or   ( new_n65442_, new_n65441_, new_n65439_ );
and  ( new_n65443_, new_n65442_, new_n65023_ );
and  ( new_n65444_, new_n65085_, new_n329_ );
nor  ( new_n65445_, new_n65444_, new_n65443_ );
nor  ( new_n65446_, new_n65445_, new_n65436_ );
and  ( new_n65447_, new_n65445_, new_n65436_ );
xor  ( new_n65448_, new_n42877_, new_n42876_ );
xnor ( new_n65449_, new_n65448_, new_n43200_ );
and  ( new_n65450_, new_n65085_, RIbb2f1d8_10 );
nor  ( new_n65451_, new_n64594_, new_n64583_ );
not  ( new_n65452_, new_n65451_ );
xor  ( new_n65453_, new_n64589_, new_n64588_ );
and  ( new_n65454_, new_n65453_, new_n65452_ );
not  ( new_n65455_, new_n65454_ );
or   ( new_n65456_, new_n65453_, new_n65452_ );
and  ( new_n65457_, new_n65456_, new_n65023_ );
and  ( new_n65458_, new_n65457_, new_n65455_ );
nor  ( new_n65459_, new_n65458_, new_n65450_ );
not  ( new_n65460_, new_n65459_ );
nor  ( new_n65461_, new_n65460_, new_n65449_ );
and  ( new_n65462_, new_n65460_, new_n65449_ );
xor  ( new_n65463_, new_n42880_, new_n42879_ );
xnor ( new_n65464_, new_n65463_, new_n43197_ );
and  ( new_n65465_, new_n65085_, RIbb2f160_11 );
xor  ( new_n65466_, new_n64574_, new_n64563_ );
nor  ( new_n65467_, new_n64581_, new_n64542_ );
nor  ( new_n65468_, new_n65467_, new_n64592_ );
not  ( new_n65469_, new_n65468_ );
and  ( new_n65470_, new_n65469_, new_n65466_ );
not  ( new_n65471_, new_n65470_ );
or   ( new_n65472_, new_n65469_, new_n65466_ );
and  ( new_n65473_, new_n65472_, new_n65023_ );
and  ( new_n65474_, new_n65473_, new_n65471_ );
nor  ( new_n65475_, new_n65474_, new_n65465_ );
not  ( new_n65476_, new_n65475_ );
nor  ( new_n65477_, new_n65476_, new_n65464_ );
and  ( new_n65478_, new_n65476_, new_n65464_ );
xor  ( new_n65479_, new_n42883_, new_n42882_ );
xnor ( new_n65480_, new_n65479_, new_n43194_ );
xor  ( new_n65481_, new_n64580_, new_n64578_ );
xor  ( new_n65482_, new_n65481_, new_n64543_ );
and  ( new_n65483_, new_n65482_, new_n65023_ );
and  ( new_n65484_, new_n65085_, RIbb2f0e8_12 );
nor  ( new_n65485_, new_n65484_, new_n65483_ );
not  ( new_n65486_, new_n65485_ );
nor  ( new_n65487_, new_n65486_, new_n65480_ );
and  ( new_n65488_, new_n65486_, new_n65480_ );
xor  ( new_n65489_, new_n42886_, new_n42885_ );
xnor ( new_n65490_, new_n65489_, new_n43191_ );
and  ( new_n65491_, new_n65085_, RIbb2f070_13 );
not  ( new_n65492_, new_n64540_ );
xor  ( new_n65493_, new_n59476_, new_n59443_ );
and  ( new_n65494_, new_n65493_, new_n65492_ );
not  ( new_n65495_, new_n65494_ );
or   ( new_n65496_, new_n65493_, new_n65492_ );
and  ( new_n65497_, new_n65496_, new_n65023_ );
and  ( new_n65498_, new_n65497_, new_n65495_ );
nor  ( new_n65499_, new_n65498_, new_n65491_ );
not  ( new_n65500_, new_n65499_ );
nor  ( new_n65501_, new_n65500_, new_n65490_ );
and  ( new_n65502_, new_n65500_, new_n65490_ );
xor  ( new_n65503_, new_n42889_, new_n42888_ );
xnor ( new_n65504_, new_n65503_, new_n43188_ );
and  ( new_n65505_, new_n65085_, RIbb2eff8_14 );
not  ( new_n65506_, new_n64538_ );
xor  ( new_n65507_, new_n59600_, new_n59599_ );
and  ( new_n65508_, new_n65507_, new_n65506_ );
not  ( new_n65509_, new_n65508_ );
or   ( new_n65510_, new_n65507_, new_n65506_ );
and  ( new_n65511_, new_n65510_, new_n65023_ );
and  ( new_n65512_, new_n65511_, new_n65509_ );
nor  ( new_n65513_, new_n65512_, new_n65505_ );
not  ( new_n65514_, new_n65513_ );
nor  ( new_n65515_, new_n65514_, new_n65504_ );
and  ( new_n65516_, new_n65514_, new_n65504_ );
xor  ( new_n65517_, new_n42892_, new_n42891_ );
xnor ( new_n65518_, new_n65517_, new_n43185_ );
and  ( new_n65519_, new_n65085_, new_n520_ );
xor  ( new_n65520_, new_n59794_, new_n59793_ );
and  ( new_n65521_, new_n65520_, new_n64536_ );
not  ( new_n65522_, new_n65521_ );
or   ( new_n65523_, new_n65520_, new_n64536_ );
and  ( new_n65524_, new_n65523_, new_n65023_ );
and  ( new_n65525_, new_n65524_, new_n65522_ );
nor  ( new_n65526_, new_n65525_, new_n65519_ );
nor  ( new_n65527_, new_n65526_, new_n65518_ );
and  ( new_n65528_, new_n65526_, new_n65518_ );
xor  ( new_n65529_, new_n42895_, new_n42894_ );
xnor ( new_n65530_, new_n65529_, new_n43182_ );
and  ( new_n65531_, new_n65085_, RIbb2ef08_16 );
not  ( new_n65532_, new_n64534_ );
xor  ( new_n65533_, new_n60096_, new_n59798_ );
and  ( new_n65534_, new_n65533_, new_n65532_ );
not  ( new_n65535_, new_n65534_ );
or   ( new_n65536_, new_n65533_, new_n65532_ );
and  ( new_n65537_, new_n65536_, new_n65023_ );
and  ( new_n65538_, new_n65537_, new_n65535_ );
nor  ( new_n65539_, new_n65538_, new_n65531_ );
not  ( new_n65540_, new_n65539_ );
nor  ( new_n65541_, new_n65540_, new_n65530_ );
and  ( new_n65542_, new_n65540_, new_n65530_ );
xor  ( new_n65543_, new_n42898_, new_n42897_ );
xnor ( new_n65544_, new_n65543_, new_n43179_ );
and  ( new_n65545_, new_n65085_, RIbb2ee90_17 );
xor  ( new_n65546_, new_n64476_, new_n64472_ );
nor  ( new_n65547_, new_n64520_, new_n64409_ );
not  ( new_n65548_, new_n65547_ );
and  ( new_n65549_, new_n65548_, new_n64504_ );
not  ( new_n65550_, new_n65549_ );
and  ( new_n65551_, new_n65550_, new_n64528_ );
nor  ( new_n65552_, new_n65551_, new_n64470_ );
nor  ( new_n65553_, new_n65552_, new_n64523_ );
not  ( new_n65554_, new_n65553_ );
and  ( new_n65555_, new_n65554_, new_n65546_ );
not  ( new_n65556_, new_n65555_ );
or   ( new_n65557_, new_n65554_, new_n65546_ );
and  ( new_n65558_, new_n65557_, new_n65023_ );
and  ( new_n65559_, new_n65558_, new_n65556_ );
nor  ( new_n65560_, new_n65559_, new_n65545_ );
not  ( new_n65561_, new_n65560_ );
nor  ( new_n65562_, new_n65561_, new_n65544_ );
and  ( new_n65563_, new_n65561_, new_n65544_ );
xor  ( new_n65564_, new_n42901_, new_n42900_ );
xnor ( new_n65565_, new_n65564_, new_n43176_ );
and  ( new_n65566_, new_n65085_, RIbb2ee18_18 );
not  ( new_n65567_, new_n65551_ );
xor  ( new_n65568_, new_n64469_, new_n64458_ );
and  ( new_n65569_, new_n65568_, new_n65567_ );
not  ( new_n65570_, new_n65569_ );
or   ( new_n65571_, new_n65568_, new_n65567_ );
and  ( new_n65572_, new_n65571_, new_n65023_ );
and  ( new_n65573_, new_n65572_, new_n65570_ );
nor  ( new_n65574_, new_n65573_, new_n65566_ );
not  ( new_n65575_, new_n65574_ );
nor  ( new_n65576_, new_n65575_, new_n65565_ );
and  ( new_n65577_, new_n65575_, new_n65565_ );
xor  ( new_n65578_, new_n42904_, new_n42903_ );
xnor ( new_n65579_, new_n65578_, new_n43173_ );
and  ( new_n65580_, new_n65085_, RIbb2eda0_19 );
and  ( new_n65581_, new_n65548_, new_n64503_ );
nor  ( new_n65582_, new_n65581_, new_n64526_ );
xor  ( new_n65583_, new_n64494_, new_n64493_ );
not  ( new_n65584_, new_n65583_ );
and  ( new_n65585_, new_n65584_, new_n65582_ );
not  ( new_n65586_, new_n65585_ );
or   ( new_n65587_, new_n65584_, new_n65582_ );
and  ( new_n65588_, new_n65587_, new_n65023_ );
and  ( new_n65589_, new_n65588_, new_n65586_ );
nor  ( new_n65590_, new_n65589_, new_n65580_ );
not  ( new_n65591_, new_n65590_ );
nor  ( new_n65592_, new_n65591_, new_n65579_ );
and  ( new_n65593_, new_n65591_, new_n65579_ );
xor  ( new_n65594_, new_n42907_, new_n42906_ );
xnor ( new_n65595_, new_n65594_, new_n43170_ );
and  ( new_n65596_, new_n65085_, RIbb2ed28_20 );
xor  ( new_n65597_, new_n64501_, new_n64500_ );
and  ( new_n65598_, new_n65597_, new_n65548_ );
not  ( new_n65599_, new_n65598_ );
or   ( new_n65600_, new_n65597_, new_n65548_ );
and  ( new_n65601_, new_n65600_, new_n65023_ );
and  ( new_n65602_, new_n65601_, new_n65599_ );
nor  ( new_n65603_, new_n65602_, new_n65596_ );
not  ( new_n65604_, new_n65603_ );
nor  ( new_n65605_, new_n65604_, new_n65595_ );
and  ( new_n65606_, new_n65604_, new_n65595_ );
xor  ( new_n65607_, new_n42910_, new_n42909_ );
xnor ( new_n65608_, new_n65607_, new_n43167_ );
and  ( new_n65609_, new_n65085_, RIbb2ecb0_21 );
xor  ( new_n65610_, new_n61019_, new_n61015_ );
not  ( new_n65611_, new_n64408_ );
and  ( new_n65612_, new_n64514_, new_n65611_ );
and  ( new_n65613_, new_n65612_, new_n64510_ );
nor  ( new_n65614_, new_n65613_, new_n60964_ );
and  ( new_n65615_, new_n65614_, new_n65610_ );
not  ( new_n65616_, new_n65615_ );
or   ( new_n65617_, new_n65614_, new_n65610_ );
and  ( new_n65618_, new_n65617_, new_n65023_ );
and  ( new_n65619_, new_n65618_, new_n65616_ );
nor  ( new_n65620_, new_n65619_, new_n65609_ );
not  ( new_n65621_, new_n65620_ );
nor  ( new_n65622_, new_n65621_, new_n65608_ );
and  ( new_n65623_, new_n65621_, new_n65608_ );
xor  ( new_n65624_, new_n42913_, new_n42912_ );
xnor ( new_n65625_, new_n65624_, new_n43164_ );
and  ( new_n65626_, new_n65085_, RIbb2ec38_22 );
not  ( new_n65627_, new_n65612_ );
xor  ( new_n65628_, new_n60963_, new_n60887_ );
and  ( new_n65629_, new_n65628_, new_n65627_ );
not  ( new_n65630_, new_n65629_ );
or   ( new_n65631_, new_n65628_, new_n65627_ );
and  ( new_n65632_, new_n65631_, new_n65023_ );
and  ( new_n65633_, new_n65632_, new_n65630_ );
nor  ( new_n65634_, new_n65633_, new_n65626_ );
not  ( new_n65635_, new_n65634_ );
nor  ( new_n65636_, new_n65635_, new_n65625_ );
and  ( new_n65637_, new_n65635_, new_n65625_ );
xor  ( new_n65638_, new_n42916_, new_n42915_ );
xnor ( new_n65639_, new_n65638_, new_n43161_ );
and  ( new_n65640_, new_n65085_, RIbb2ebc0_23 );
nor  ( new_n65641_, new_n64512_, new_n64407_ );
xor  ( new_n65642_, new_n61235_, new_n61234_ );
not  ( new_n65643_, new_n65642_ );
and  ( new_n65644_, new_n65643_, new_n65641_ );
not  ( new_n65645_, new_n65644_ );
or   ( new_n65646_, new_n65643_, new_n65641_ );
and  ( new_n65647_, new_n65646_, new_n65023_ );
and  ( new_n65648_, new_n65647_, new_n65645_ );
nor  ( new_n65649_, new_n65648_, new_n65640_ );
not  ( new_n65650_, new_n65649_ );
nor  ( new_n65651_, new_n65650_, new_n65639_ );
and  ( new_n65652_, new_n65650_, new_n65639_ );
xor  ( new_n65653_, new_n42919_, new_n42918_ );
xnor ( new_n65654_, new_n65653_, new_n43158_ );
and  ( new_n65655_, new_n65085_, RIbb2eb48_24 );
not  ( new_n65656_, new_n64406_ );
xor  ( new_n65657_, new_n61441_, new_n61440_ );
and  ( new_n65658_, new_n65657_, new_n65656_ );
not  ( new_n65659_, new_n65658_ );
or   ( new_n65660_, new_n65657_, new_n65656_ );
and  ( new_n65661_, new_n65660_, new_n65023_ );
and  ( new_n65662_, new_n65661_, new_n65659_ );
nor  ( new_n65663_, new_n65662_, new_n65655_ );
not  ( new_n65664_, new_n65663_ );
nor  ( new_n65665_, new_n65664_, new_n65654_ );
and  ( new_n65666_, new_n65664_, new_n65654_ );
xor  ( new_n65667_, new_n42922_, new_n42921_ );
xnor ( new_n65668_, new_n65667_, new_n43155_ );
and  ( new_n65669_, new_n65085_, RIbb2ead0_25 );
xor  ( new_n65670_, new_n61589_, new_n61588_ );
nor  ( new_n65671_, new_n64391_, new_n64378_ );
not  ( new_n65672_, new_n65671_ );
and  ( new_n65673_, new_n65672_, new_n61904_ );
not  ( new_n65674_, new_n65673_ );
and  ( new_n65675_, new_n65674_, new_n64400_ );
nor  ( new_n65676_, new_n65675_, new_n61665_ );
nor  ( new_n65677_, new_n65676_, new_n64395_ );
not  ( new_n65678_, new_n65677_ );
and  ( new_n65679_, new_n65678_, new_n65670_ );
not  ( new_n65680_, new_n65679_ );
or   ( new_n65681_, new_n65678_, new_n65670_ );
and  ( new_n65682_, new_n65681_, new_n65023_ );
and  ( new_n65683_, new_n65682_, new_n65680_ );
nor  ( new_n65684_, new_n65683_, new_n65669_ );
not  ( new_n65685_, new_n65684_ );
nor  ( new_n65686_, new_n65685_, new_n65668_ );
and  ( new_n65687_, new_n65685_, new_n65668_ );
xor  ( new_n65688_, new_n42925_, new_n42924_ );
xnor ( new_n65689_, new_n65688_, new_n43152_ );
and  ( new_n65690_, new_n65085_, RIbb2ea58_26 );
not  ( new_n65691_, new_n65675_ );
xor  ( new_n65692_, new_n61664_, new_n61663_ );
and  ( new_n65693_, new_n65692_, new_n65691_ );
not  ( new_n65694_, new_n65693_ );
or   ( new_n65695_, new_n65692_, new_n65691_ );
and  ( new_n65696_, new_n65695_, new_n65023_ );
and  ( new_n65697_, new_n65696_, new_n65694_ );
nor  ( new_n65698_, new_n65697_, new_n65690_ );
not  ( new_n65699_, new_n65698_ );
nor  ( new_n65700_, new_n65699_, new_n65689_ );
and  ( new_n65701_, new_n65699_, new_n65689_ );
xor  ( new_n65702_, new_n42928_, new_n42927_ );
xnor ( new_n65703_, new_n65702_, new_n43149_ );
and  ( new_n65704_, new_n65085_, RIbb2e9e0_27 );
xor  ( new_n65705_, new_n61880_, new_n61879_ );
and  ( new_n65706_, new_n65672_, new_n61903_ );
nor  ( new_n65707_, new_n65706_, new_n64398_ );
not  ( new_n65708_, new_n65707_ );
and  ( new_n65709_, new_n65708_, new_n65705_ );
not  ( new_n65710_, new_n65709_ );
or   ( new_n65711_, new_n65708_, new_n65705_ );
and  ( new_n65712_, new_n65711_, new_n65023_ );
and  ( new_n65713_, new_n65712_, new_n65710_ );
nor  ( new_n65714_, new_n65713_, new_n65704_ );
not  ( new_n65715_, new_n65714_ );
nor  ( new_n65716_, new_n65715_, new_n65703_ );
and  ( new_n65717_, new_n65715_, new_n65703_ );
xor  ( new_n65718_, new_n42931_, new_n42930_ );
xnor ( new_n65719_, new_n65718_, new_n43146_ );
and  ( new_n65720_, new_n65085_, RIbb2e968_28 );
xor  ( new_n65721_, new_n61901_, new_n61883_ );
and  ( new_n65722_, new_n65721_, new_n65672_ );
not  ( new_n65723_, new_n65722_ );
or   ( new_n65724_, new_n65721_, new_n65672_ );
and  ( new_n65725_, new_n65724_, new_n65023_ );
and  ( new_n65726_, new_n65725_, new_n65723_ );
nor  ( new_n65727_, new_n65726_, new_n65720_ );
not  ( new_n65728_, new_n65727_ );
nor  ( new_n65729_, new_n65728_, new_n65719_ );
and  ( new_n65730_, new_n65728_, new_n65719_ );
xor  ( new_n65731_, new_n42934_, new_n42933_ );
xnor ( new_n65732_, new_n65731_, new_n43143_ );
and  ( new_n65733_, new_n65085_, RIbb2e8f0_29 );
xor  ( new_n65734_, new_n62146_, new_n62144_ );
nor  ( new_n65735_, new_n64386_, new_n64377_ );
nor  ( new_n65736_, new_n65735_, new_n62218_ );
nor  ( new_n65737_, new_n65736_, new_n64382_ );
not  ( new_n65738_, new_n65737_ );
and  ( new_n65739_, new_n65738_, new_n65734_ );
not  ( new_n65740_, new_n65739_ );
or   ( new_n65741_, new_n65738_, new_n65734_ );
and  ( new_n65742_, new_n65741_, new_n65023_ );
and  ( new_n65743_, new_n65742_, new_n65740_ );
nor  ( new_n65744_, new_n65743_, new_n65733_ );
not  ( new_n65745_, new_n65744_ );
nor  ( new_n65746_, new_n65745_, new_n65732_ );
and  ( new_n65747_, new_n65745_, new_n65732_ );
xor  ( new_n65748_, new_n42937_, new_n42936_ );
xnor ( new_n65749_, new_n65748_, new_n43140_ );
and  ( new_n65750_, new_n65085_, RIbb2e878_30 );
not  ( new_n65751_, new_n65735_ );
xor  ( new_n65752_, new_n62217_, new_n62215_ );
and  ( new_n65753_, new_n65752_, new_n65751_ );
not  ( new_n65754_, new_n65753_ );
or   ( new_n65755_, new_n65752_, new_n65751_ );
and  ( new_n65756_, new_n65755_, new_n65023_ );
and  ( new_n65757_, new_n65756_, new_n65754_ );
nor  ( new_n65758_, new_n65757_, new_n65750_ );
not  ( new_n65759_, new_n65758_ );
nor  ( new_n65760_, new_n65759_, new_n65749_ );
and  ( new_n65761_, new_n65759_, new_n65749_ );
xor  ( new_n65762_, new_n42940_, new_n42939_ );
xnor ( new_n65763_, new_n65762_, new_n43137_ );
and  ( new_n65764_, new_n65085_, RIbb2e800_31 );
xor  ( new_n65765_, new_n62338_, new_n62336_ );
nor  ( new_n65766_, new_n64383_, new_n64375_ );
not  ( new_n65767_, new_n65766_ );
and  ( new_n65768_, new_n65767_, new_n65765_ );
not  ( new_n65769_, new_n65768_ );
or   ( new_n65770_, new_n65767_, new_n65765_ );
and  ( new_n65771_, new_n65770_, new_n65023_ );
and  ( new_n65772_, new_n65771_, new_n65769_ );
nor  ( new_n65773_, new_n65772_, new_n65764_ );
not  ( new_n65774_, new_n65773_ );
nor  ( new_n65775_, new_n65774_, new_n65763_ );
and  ( new_n65776_, new_n65774_, new_n65763_ );
xor  ( new_n65777_, new_n62480_, new_n62340_ );
xor  ( new_n65778_, new_n65777_, new_n64374_ );
and  ( new_n65779_, new_n65778_, new_n65023_ );
and  ( new_n65780_, new_n65085_, new_n45843_ );
or   ( new_n65781_, new_n65780_, new_n65779_ );
xnor ( new_n65782_, new_n42943_, new_n42942_ );
xor  ( new_n65783_, new_n65782_, new_n43135_ );
xor  ( new_n65784_, new_n65783_, new_n65781_ );
xor  ( new_n65785_, new_n62558_, new_n62556_ );
or   ( new_n65786_, new_n64370_, new_n64368_ );
and  ( new_n65787_, new_n65786_, new_n65785_ );
not  ( new_n65788_, new_n62560_ );
and  ( new_n65789_, new_n64373_, new_n65788_ );
or   ( new_n65790_, new_n65789_, new_n65787_ );
and  ( new_n65791_, new_n65790_, new_n65023_ );
and  ( new_n65792_, new_n65085_, new_n2797_ );
nor  ( new_n65793_, new_n65792_, new_n65791_ );
xor  ( new_n65794_, new_n43130_, new_n42946_ );
xor  ( new_n65795_, new_n65794_, new_n43133_ );
not  ( new_n65796_, new_n65795_ );
nor  ( new_n65797_, new_n65796_, new_n65793_ );
and  ( new_n65798_, new_n65796_, new_n65793_ );
xor  ( new_n65799_, new_n42952_, new_n42951_ );
xnor ( new_n65800_, new_n65799_, new_n43125_ );
and  ( new_n65801_, new_n65085_, RIbb2e620_35 );
nor  ( new_n65802_, new_n64364_, new_n64353_ );
xor  ( new_n65803_, new_n62825_, new_n62812_ );
not  ( new_n65804_, new_n65803_ );
and  ( new_n65805_, new_n65804_, new_n65802_ );
not  ( new_n65806_, new_n65805_ );
or   ( new_n65807_, new_n65804_, new_n65802_ );
and  ( new_n65808_, new_n65807_, new_n65023_ );
and  ( new_n65809_, new_n65808_, new_n65806_ );
nor  ( new_n65810_, new_n65809_, new_n65801_ );
not  ( new_n65811_, new_n65810_ );
nor  ( new_n65812_, new_n65811_, new_n65800_ );
and  ( new_n65813_, new_n65811_, new_n65800_ );
xor  ( new_n65814_, new_n42955_, new_n42954_ );
xnor ( new_n65815_, new_n65814_, new_n43122_ );
and  ( new_n65816_, new_n65085_, RIbb2e5a8_36 );
not  ( new_n65817_, new_n64352_ );
xor  ( new_n65818_, new_n62972_, new_n62828_ );
and  ( new_n65819_, new_n65818_, new_n65817_ );
not  ( new_n65820_, new_n65819_ );
or   ( new_n65821_, new_n65818_, new_n65817_ );
and  ( new_n65822_, new_n65821_, new_n65023_ );
and  ( new_n65823_, new_n65822_, new_n65820_ );
nor  ( new_n65824_, new_n65823_, new_n65816_ );
not  ( new_n65825_, new_n65824_ );
nor  ( new_n65826_, new_n65825_, new_n65815_ );
and  ( new_n65827_, new_n65825_, new_n65815_ );
xor  ( new_n65828_, new_n42958_, new_n42957_ );
xnor ( new_n65829_, new_n65828_, new_n43119_ );
xor  ( new_n65830_, new_n62992_, new_n62990_ );
xor  ( new_n65831_, new_n65830_, new_n64350_ );
nor  ( new_n65832_, new_n65831_, new_n65085_ );
and  ( new_n65833_, new_n65085_, RIbb2e530_37 );
nor  ( new_n65834_, new_n65833_, new_n65832_ );
not  ( new_n65835_, new_n65834_ );
nor  ( new_n65836_, new_n65835_, new_n65829_ );
and  ( new_n65837_, new_n65835_, new_n65829_ );
xor  ( new_n65838_, new_n42961_, new_n42960_ );
xnor ( new_n65839_, new_n65838_, new_n43116_ );
xnor ( new_n65840_, new_n63159_, new_n62995_ );
xor  ( new_n65841_, new_n65840_, new_n64348_ );
and  ( new_n65842_, new_n65841_, new_n65023_ );
and  ( new_n65843_, new_n65085_, RIbb2e4b8_38 );
nor  ( new_n65844_, new_n65843_, new_n65842_ );
not  ( new_n65845_, new_n65844_ );
nor  ( new_n65846_, new_n65845_, new_n65839_ );
and  ( new_n65847_, new_n65845_, new_n65839_ );
xor  ( new_n65848_, new_n42964_, new_n42963_ );
xnor ( new_n65849_, new_n65848_, new_n43113_ );
and  ( new_n65850_, new_n65085_, RIbb2e440_39 );
not  ( new_n65851_, new_n64346_ );
xor  ( new_n65852_, new_n63252_, new_n63250_ );
and  ( new_n65853_, new_n65852_, new_n65851_ );
not  ( new_n65854_, new_n65853_ );
or   ( new_n65855_, new_n65852_, new_n65851_ );
and  ( new_n65856_, new_n65855_, new_n65023_ );
and  ( new_n65857_, new_n65856_, new_n65854_ );
nor  ( new_n65858_, new_n65857_, new_n65850_ );
not  ( new_n65859_, new_n65858_ );
nor  ( new_n65860_, new_n65859_, new_n65849_ );
and  ( new_n65861_, new_n65859_, new_n65849_ );
xor  ( new_n65862_, new_n42967_, new_n42966_ );
xnor ( new_n65863_, new_n65862_, new_n43110_ );
and  ( new_n65864_, new_n65085_, RIbb2e3c8_40 );
not  ( new_n65865_, new_n64344_ );
xor  ( new_n65866_, new_n63299_, new_n63297_ );
and  ( new_n65867_, new_n65866_, new_n65865_ );
not  ( new_n65868_, new_n65867_ );
or   ( new_n65869_, new_n65866_, new_n65865_ );
and  ( new_n65870_, new_n65869_, new_n65023_ );
and  ( new_n65871_, new_n65870_, new_n65868_ );
nor  ( new_n65872_, new_n65871_, new_n65864_ );
not  ( new_n65873_, new_n65872_ );
nor  ( new_n65874_, new_n65873_, new_n65863_ );
and  ( new_n65875_, new_n65873_, new_n65863_ );
xor  ( new_n65876_, new_n42970_, new_n42969_ );
xnor ( new_n65877_, new_n65876_, new_n43107_ );
and  ( new_n65878_, new_n65085_, RIbb2e350_41 );
xor  ( new_n65879_, new_n63407_, new_n63303_ );
and  ( new_n65880_, new_n65879_, new_n64341_ );
not  ( new_n65881_, new_n65880_ );
or   ( new_n65882_, new_n65879_, new_n64341_ );
and  ( new_n65883_, new_n65882_, new_n65023_ );
and  ( new_n65884_, new_n65883_, new_n65881_ );
nor  ( new_n65885_, new_n65884_, new_n65878_ );
not  ( new_n65886_, new_n65885_ );
nor  ( new_n65887_, new_n65886_, new_n65877_ );
and  ( new_n65888_, new_n65886_, new_n65877_ );
xor  ( new_n65889_, new_n42973_, new_n42972_ );
xnor ( new_n65890_, new_n65889_, new_n43104_ );
and  ( new_n65891_, new_n65085_, RIbb2e2d8_42 );
xor  ( new_n65892_, new_n63475_, new_n63473_ );
and  ( new_n65893_, new_n65892_, new_n64339_ );
not  ( new_n65894_, new_n65893_ );
or   ( new_n65895_, new_n65892_, new_n64339_ );
and  ( new_n65896_, new_n65895_, new_n65023_ );
and  ( new_n65897_, new_n65896_, new_n65894_ );
nor  ( new_n65898_, new_n65897_, new_n65891_ );
not  ( new_n65899_, new_n65898_ );
nor  ( new_n65900_, new_n65899_, new_n65890_ );
and  ( new_n65901_, new_n65899_, new_n65890_ );
xor  ( new_n65902_, new_n42976_, new_n42975_ );
xnor ( new_n65903_, new_n65902_, new_n43101_ );
and  ( new_n65904_, new_n65085_, RIbb2e260_43 );
xor  ( new_n65905_, new_n63589_, new_n63587_ );
and  ( new_n65906_, new_n65905_, new_n64337_ );
not  ( new_n65907_, new_n65906_ );
or   ( new_n65908_, new_n65905_, new_n64337_ );
and  ( new_n65909_, new_n65908_, new_n65023_ );
and  ( new_n65910_, new_n65909_, new_n65907_ );
nor  ( new_n65911_, new_n65910_, new_n65904_ );
not  ( new_n65912_, new_n65911_ );
nor  ( new_n65913_, new_n65912_, new_n65903_ );
and  ( new_n65914_, new_n65912_, new_n65903_ );
xor  ( new_n65915_, new_n42979_, new_n42978_ );
xnor ( new_n65916_, new_n65915_, new_n43098_ );
and  ( new_n65917_, new_n65085_, RIbb2e1e8_44 );
xor  ( new_n65918_, new_n63653_, new_n63651_ );
and  ( new_n65919_, new_n65918_, new_n64335_ );
not  ( new_n65920_, new_n65919_ );
or   ( new_n65921_, new_n65918_, new_n64335_ );
and  ( new_n65922_, new_n65921_, new_n65023_ );
and  ( new_n65923_, new_n65922_, new_n65920_ );
nor  ( new_n65924_, new_n65923_, new_n65917_ );
not  ( new_n65925_, new_n65924_ );
nor  ( new_n65926_, new_n65925_, new_n65916_ );
and  ( new_n65927_, new_n65925_, new_n65916_ );
xor  ( new_n65928_, new_n42982_, new_n42981_ );
xnor ( new_n65929_, new_n65928_, new_n43095_ );
and  ( new_n65930_, new_n65085_, RIbb2e170_45 );
xor  ( new_n65931_, new_n63721_, new_n63720_ );
and  ( new_n65932_, new_n65931_, new_n64333_ );
not  ( new_n65933_, new_n65932_ );
or   ( new_n65934_, new_n65931_, new_n64333_ );
and  ( new_n65935_, new_n65934_, new_n65023_ );
and  ( new_n65936_, new_n65935_, new_n65933_ );
nor  ( new_n65937_, new_n65936_, new_n65930_ );
not  ( new_n65938_, new_n65937_ );
nor  ( new_n65939_, new_n65938_, new_n65929_ );
and  ( new_n65940_, new_n65938_, new_n65929_ );
xor  ( new_n65941_, new_n42985_, new_n42984_ );
xnor ( new_n65942_, new_n65941_, new_n43092_ );
and  ( new_n65943_, new_n65085_, RIbb2e0f8_46 );
xor  ( new_n65944_, new_n63773_, new_n63724_ );
and  ( new_n65945_, new_n65944_, new_n64331_ );
not  ( new_n65946_, new_n65945_ );
or   ( new_n65947_, new_n65944_, new_n64331_ );
and  ( new_n65948_, new_n65947_, new_n65023_ );
and  ( new_n65949_, new_n65948_, new_n65946_ );
nor  ( new_n65950_, new_n65949_, new_n65943_ );
not  ( new_n65951_, new_n65950_ );
nor  ( new_n65952_, new_n65951_, new_n65942_ );
and  ( new_n65953_, new_n65951_, new_n65942_ );
xor  ( new_n65954_, new_n42988_, new_n42987_ );
xor  ( new_n65955_, new_n65954_, new_n43090_ );
and  ( new_n65956_, new_n65085_, RIbb2e080_47 );
xor  ( new_n65957_, new_n63818_, new_n63816_ );
and  ( new_n65958_, new_n65957_, new_n64329_ );
not  ( new_n65959_, new_n65958_ );
or   ( new_n65960_, new_n65957_, new_n64329_ );
and  ( new_n65961_, new_n65960_, new_n65023_ );
and  ( new_n65962_, new_n65961_, new_n65959_ );
nor  ( new_n65963_, new_n65962_, new_n65956_ );
and  ( new_n65964_, new_n65963_, new_n65955_ );
nor  ( new_n65965_, new_n65963_, new_n65955_ );
xor  ( new_n65966_, new_n42992_, new_n42991_ );
xor  ( new_n65967_, new_n65966_, new_n43088_ );
and  ( new_n65968_, new_n65085_, RIbb2e008_48 );
xor  ( new_n65969_, new_n63874_, new_n63822_ );
and  ( new_n65970_, new_n65969_, new_n64327_ );
not  ( new_n65971_, new_n65970_ );
or   ( new_n65972_, new_n65969_, new_n64327_ );
and  ( new_n65973_, new_n65972_, new_n65023_ );
and  ( new_n65974_, new_n65973_, new_n65971_ );
nor  ( new_n65975_, new_n65974_, new_n65968_ );
and  ( new_n65976_, new_n65975_, new_n65967_ );
nor  ( new_n65977_, new_n65975_, new_n65967_ );
xor  ( new_n65978_, new_n42996_, new_n42995_ );
xnor ( new_n65979_, new_n65978_, new_n43086_ );
and  ( new_n65980_, new_n65085_, RIbb2df90_49 );
not  ( new_n65981_, new_n64324_ );
xor  ( new_n65982_, new_n63930_, new_n63928_ );
and  ( new_n65983_, new_n65982_, new_n65981_ );
not  ( new_n65984_, new_n65983_ );
or   ( new_n65985_, new_n65982_, new_n65981_ );
and  ( new_n65986_, new_n65985_, new_n65023_ );
and  ( new_n65987_, new_n65986_, new_n65984_ );
nor  ( new_n65988_, new_n65987_, new_n65980_ );
not  ( new_n65989_, new_n65988_ );
nor  ( new_n65990_, new_n65989_, new_n65979_ );
and  ( new_n65991_, new_n65989_, new_n65979_ );
xor  ( new_n65992_, new_n43000_, new_n42999_ );
xnor ( new_n65993_, new_n65992_, new_n43083_ );
and  ( new_n65994_, new_n65085_, RIbb2df18_50 );
not  ( new_n65995_, new_n64322_ );
xor  ( new_n65996_, new_n63986_, new_n63984_ );
and  ( new_n65997_, new_n65996_, new_n65995_ );
not  ( new_n65998_, new_n65997_ );
or   ( new_n65999_, new_n65996_, new_n65995_ );
and  ( new_n66000_, new_n65999_, new_n65023_ );
and  ( new_n66001_, new_n66000_, new_n65998_ );
nor  ( new_n66002_, new_n66001_, new_n65994_ );
not  ( new_n66003_, new_n66002_ );
nor  ( new_n66004_, new_n66003_, new_n65993_ );
and  ( new_n66005_, new_n66003_, new_n65993_ );
xor  ( new_n66006_, new_n43003_, new_n43002_ );
xnor ( new_n66007_, new_n66006_, new_n43080_ );
and  ( new_n66008_, new_n65085_, RIbb2dea0_51 );
not  ( new_n66009_, new_n64320_ );
xor  ( new_n66010_, new_n64028_, new_n64026_ );
and  ( new_n66011_, new_n66010_, new_n66009_ );
not  ( new_n66012_, new_n66011_ );
or   ( new_n66013_, new_n66010_, new_n66009_ );
and  ( new_n66014_, new_n66013_, new_n65023_ );
and  ( new_n66015_, new_n66014_, new_n66012_ );
nor  ( new_n66016_, new_n66015_, new_n66008_ );
not  ( new_n66017_, new_n66016_ );
nor  ( new_n66018_, new_n66017_, new_n66007_ );
and  ( new_n66019_, new_n66017_, new_n66007_ );
xor  ( new_n66020_, new_n43006_, new_n43005_ );
xnor ( new_n66021_, new_n66020_, new_n43077_ );
and  ( new_n66022_, new_n65085_, RIbb2de28_52 );
not  ( new_n66023_, new_n64318_ );
xor  ( new_n66024_, new_n64068_, new_n64066_ );
and  ( new_n66025_, new_n66024_, new_n66023_ );
not  ( new_n66026_, new_n66025_ );
or   ( new_n66027_, new_n66024_, new_n66023_ );
and  ( new_n66028_, new_n66027_, new_n65023_ );
and  ( new_n66029_, new_n66028_, new_n66026_ );
nor  ( new_n66030_, new_n66029_, new_n66022_ );
not  ( new_n66031_, new_n66030_ );
nor  ( new_n66032_, new_n66031_, new_n66021_ );
and  ( new_n66033_, new_n66031_, new_n66021_ );
xor  ( new_n66034_, new_n43012_, new_n43011_ );
xor  ( new_n66035_, new_n64144_, new_n64142_ );
xor  ( new_n66036_, new_n66035_, new_n64314_ );
or   ( new_n66037_, new_n66036_, new_n65085_ );
or   ( new_n66038_, new_n65023_, new_n50764_ );
and  ( new_n66039_, new_n66038_, new_n66037_ );
xnor ( new_n66040_, new_n66039_, new_n66034_ );
xor  ( new_n66041_, new_n66040_, new_n43072_ );
xnor ( new_n66042_, new_n43009_, new_n43008_ );
xor  ( new_n66043_, new_n66042_, new_n43074_ );
xor  ( new_n66044_, new_n64104_, new_n64071_ );
xor  ( new_n66045_, new_n66044_, new_n64316_ );
or   ( new_n66046_, new_n66045_, new_n65085_ );
or   ( new_n66047_, new_n65023_, new_n7174_ );
and  ( new_n66048_, new_n66047_, new_n66046_ );
xor  ( new_n66049_, new_n66048_, new_n66043_ );
or   ( new_n66050_, new_n66049_, new_n66041_ );
or   ( new_n66051_, new_n66050_, new_n66033_ );
or   ( new_n66052_, new_n66051_, new_n66032_ );
or   ( new_n66053_, new_n66052_, new_n66019_ );
or   ( new_n66054_, new_n66053_, new_n66018_ );
or   ( new_n66055_, new_n66054_, new_n66005_ );
or   ( new_n66056_, new_n66055_, new_n66004_ );
or   ( new_n66057_, new_n66056_, new_n65991_ );
or   ( new_n66058_, new_n66057_, new_n65990_ );
or   ( new_n66059_, new_n66058_, new_n65977_ );
or   ( new_n66060_, new_n66059_, new_n65976_ );
or   ( new_n66061_, new_n66060_, new_n65965_ );
or   ( new_n66062_, new_n66061_, new_n65964_ );
or   ( new_n66063_, new_n66062_, new_n65953_ );
or   ( new_n66064_, new_n66063_, new_n65952_ );
or   ( new_n66065_, new_n66064_, new_n65940_ );
or   ( new_n66066_, new_n66065_, new_n65939_ );
or   ( new_n66067_, new_n66066_, new_n65927_ );
or   ( new_n66068_, new_n66067_, new_n65926_ );
or   ( new_n66069_, new_n66068_, new_n65914_ );
or   ( new_n66070_, new_n66069_, new_n65913_ );
or   ( new_n66071_, new_n66070_, new_n65901_ );
or   ( new_n66072_, new_n66071_, new_n65900_ );
or   ( new_n66073_, new_n66072_, new_n65888_ );
or   ( new_n66074_, new_n66073_, new_n65887_ );
or   ( new_n66075_, new_n66074_, new_n65875_ );
or   ( new_n66076_, new_n66075_, new_n65874_ );
or   ( new_n66077_, new_n66076_, new_n65861_ );
or   ( new_n66078_, new_n66077_, new_n65860_ );
or   ( new_n66079_, new_n66078_, new_n65847_ );
or   ( new_n66080_, new_n66079_, new_n65846_ );
or   ( new_n66081_, new_n66080_, new_n65837_ );
or   ( new_n66082_, new_n66081_, new_n65836_ );
or   ( new_n66083_, new_n66082_, new_n65827_ );
or   ( new_n66084_, new_n66083_, new_n65826_ );
or   ( new_n66085_, new_n66084_, new_n65813_ );
or   ( new_n66086_, new_n66085_, new_n65812_ );
xnor ( new_n66087_, new_n42948_, new_n42947_ );
xor  ( new_n66088_, new_n66087_, new_n43128_ );
or   ( new_n66089_, new_n65023_, new_n46353_ );
and  ( new_n66090_, new_n64366_, new_n64355_ );
xor  ( new_n66091_, new_n64360_, new_n64358_ );
not  ( new_n66092_, new_n66091_ );
nor  ( new_n66093_, new_n66092_, new_n66090_ );
and  ( new_n66094_, new_n66092_, new_n66090_ );
or   ( new_n66095_, new_n66094_, new_n65085_ );
or   ( new_n66096_, new_n66095_, new_n66093_ );
and  ( new_n66097_, new_n66096_, new_n66089_ );
xor  ( new_n66098_, new_n66097_, new_n66088_ );
or   ( new_n66099_, new_n66098_, new_n66086_ );
or   ( new_n66100_, new_n66099_, new_n65798_ );
or   ( new_n66101_, new_n66100_, new_n65797_ );
or   ( new_n66102_, new_n66101_, new_n65784_ );
or   ( new_n66103_, new_n66102_, new_n65776_ );
or   ( new_n66104_, new_n66103_, new_n65775_ );
or   ( new_n66105_, new_n66104_, new_n65761_ );
or   ( new_n66106_, new_n66105_, new_n65760_ );
or   ( new_n66107_, new_n66106_, new_n65747_ );
or   ( new_n66108_, new_n66107_, new_n65746_ );
or   ( new_n66109_, new_n66108_, new_n65730_ );
or   ( new_n66110_, new_n66109_, new_n65729_ );
or   ( new_n66111_, new_n66110_, new_n65717_ );
or   ( new_n66112_, new_n66111_, new_n65716_ );
or   ( new_n66113_, new_n66112_, new_n65701_ );
or   ( new_n66114_, new_n66113_, new_n65700_ );
or   ( new_n66115_, new_n66114_, new_n65687_ );
or   ( new_n66116_, new_n66115_, new_n65686_ );
or   ( new_n66117_, new_n66116_, new_n65666_ );
or   ( new_n66118_, new_n66117_, new_n65665_ );
or   ( new_n66119_, new_n66118_, new_n65652_ );
or   ( new_n66120_, new_n66119_, new_n65651_ );
or   ( new_n66121_, new_n66120_, new_n65637_ );
or   ( new_n66122_, new_n66121_, new_n65636_ );
or   ( new_n66123_, new_n66122_, new_n65623_ );
or   ( new_n66124_, new_n66123_, new_n65622_ );
or   ( new_n66125_, new_n66124_, new_n65606_ );
or   ( new_n66126_, new_n66125_, new_n65605_ );
or   ( new_n66127_, new_n66126_, new_n65593_ );
or   ( new_n66128_, new_n66127_, new_n65592_ );
or   ( new_n66129_, new_n66128_, new_n65577_ );
or   ( new_n66130_, new_n66129_, new_n65576_ );
or   ( new_n66131_, new_n66130_, new_n65563_ );
or   ( new_n66132_, new_n66131_, new_n65562_ );
or   ( new_n66133_, new_n66132_, new_n65542_ );
or   ( new_n66134_, new_n66133_, new_n65541_ );
or   ( new_n66135_, new_n66134_, new_n65528_ );
or   ( new_n66136_, new_n66135_, new_n65527_ );
or   ( new_n66137_, new_n66136_, new_n65516_ );
or   ( new_n66138_, new_n66137_, new_n65515_ );
or   ( new_n66139_, new_n66138_, new_n65502_ );
or   ( new_n66140_, new_n66139_, new_n65501_ );
or   ( new_n66141_, new_n66140_, new_n65488_ );
or   ( new_n66142_, new_n66141_, new_n65487_ );
or   ( new_n66143_, new_n66142_, new_n65478_ );
or   ( new_n66144_, new_n66143_, new_n65477_ );
or   ( new_n66145_, new_n66144_, new_n65462_ );
or   ( new_n66146_, new_n66145_, new_n65461_ );
or   ( new_n66147_, new_n66146_, new_n65447_ );
or   ( new_n66148_, new_n66147_, new_n65446_ );
or   ( new_n66149_, new_n66148_, new_n65434_ );
or   ( new_n66150_, new_n66149_, new_n65433_ );
or   ( new_n66151_, new_n66150_, new_n65420_ );
or   ( new_n66152_, new_n66151_, new_n65419_ );
or   ( new_n66153_, new_n66152_, new_n65406_ );
or   ( new_n66154_, new_n66153_, new_n65405_ );
or   ( new_n66155_, new_n66154_, new_n65393_ );
or   ( new_n66156_, new_n66155_, new_n65392_ );
or   ( new_n66157_, new_n66156_, new_n65380_ );
or   ( new_n66158_, new_n66157_, new_n65379_ );
or   ( new_n66159_, new_n66158_, new_n65367_ );
or   ( new_n66160_, new_n66159_, new_n65366_ );
or   ( new_n66161_, new_n66160_, new_n65354_ );
or   ( new_n66162_, new_n66161_, new_n65353_ );
or   ( new_n66163_, new_n66162_, new_n65340_ );
or   ( new_n66164_, new_n66163_, new_n65339_ );
or   ( new_n66165_, new_n66164_, new_n65330_ );
or   ( new_n66166_, new_n66165_, new_n65329_ );
or   ( new_n66167_, new_n66166_, new_n65322_ );
or   ( new_n66168_, new_n66167_, new_n65321_ );
or   ( new_n66169_, new_n66168_, new_n65312_ );
or   ( new_n66170_, new_n66169_, new_n65311_ );
or   ( new_n66171_, new_n66170_, new_n65302_ );
or   ( new_n66172_, new_n66171_, new_n65301_ );
or   ( new_n66173_, new_n66172_, new_n65294_ );
or   ( new_n66174_, new_n66173_, new_n65293_ );
or   ( new_n66175_, new_n66174_, new_n65287_ );
or   ( new_n66176_, new_n66175_, new_n65286_ );
or   ( new_n66177_, new_n66176_, new_n65280_ );
or   ( new_n66178_, new_n66177_, new_n65279_ );
or   ( new_n66179_, new_n66178_, new_n65270_ );
or   ( new_n66180_, new_n66179_, new_n65269_ );
or   ( new_n66181_, new_n66180_, new_n65263_ );
or   ( new_n66182_, new_n66181_, new_n65262_ );
or   ( new_n66183_, new_n66182_, new_n65256_ );
or   ( new_n66184_, new_n66183_, new_n65255_ );
or   ( new_n66185_, new_n66184_, new_n65246_ );
or   ( new_n66186_, new_n66185_, new_n65245_ );
or   ( new_n66187_, new_n66186_, new_n65236_ );
or   ( new_n66188_, new_n66187_, new_n65235_ );
or   ( new_n66189_, new_n66188_, new_n65226_ );
or   ( new_n66190_, new_n66189_, new_n65225_ );
or   ( new_n66191_, new_n66190_, new_n65219_ );
or   ( new_n66192_, new_n66191_, new_n65218_ );
or   ( new_n66193_, new_n66192_, new_n65209_ );
or   ( new_n66194_, new_n66193_, new_n65208_ );
or   ( new_n66195_, new_n66194_, new_n65199_ );
or   ( new_n66196_, new_n66195_, new_n65198_ );
or   ( new_n66197_, new_n66196_, new_n65189_ );
or   ( new_n66198_, new_n66197_, new_n65188_ );
or   ( new_n66199_, new_n66198_, new_n65179_ );
or   ( new_n66200_, new_n66199_, new_n65178_ );
or   ( new_n66201_, new_n66200_, new_n65172_ );
or   ( new_n66202_, new_n66201_, new_n65171_ );
or   ( new_n66203_, new_n66202_, new_n65165_ );
or   ( new_n66204_, new_n66203_, new_n65164_ );
or   ( new_n66205_, new_n66204_, new_n65157_ );
or   ( new_n66206_, new_n66205_, new_n65151_ );
or   ( new_n66207_, new_n66206_, new_n65150_ );
or   ( new_n66208_, new_n66207_, new_n65144_ );
or   ( new_n66209_, new_n66208_, new_n65143_ );
or   ( new_n66210_, new_n66209_, new_n65136_ );
or   ( new_n66211_, new_n66210_, new_n65135_ );
or   ( new_n66212_, new_n66211_, new_n65128_ );
or   ( new_n66213_, new_n66212_, new_n65127_ );
or   ( new_n66214_, new_n66213_, new_n65121_ );
or   ( new_n66215_, new_n66214_, new_n65120_ );
or   ( new_n66216_, new_n66215_, new_n65110_ );
or   ( new_n66217_, new_n66216_, new_n65109_ );
or   ( new_n66218_, new_n66217_, new_n65098_ );
or   ( new_n66219_, new_n66218_, new_n65097_ );
or   ( new_n66220_, new_n66219_, new_n65090_ );
or   ( new_n66221_, new_n66220_, new_n65089_ );
or   ( new_n66222_, new_n66221_, new_n65082_ );
or   ( new_n66223_, new_n66222_, new_n65081_ );
or   ( new_n66224_, new_n66223_, new_n65075_ );
or   ( new_n66225_, new_n66224_, new_n65074_ );
xnor ( new_n66226_, RIbb35178_256, RIbb35100_255 );
xnor ( new_n66227_, RIbb34ae8_242, RIbb34a70_241 );
xor  ( new_n66228_, RIbb34cc8_246, RIbb34c50_245 );
xor  ( new_n66229_, new_n66228_, new_n66227_ );
xor  ( new_n66230_, new_n66229_, new_n66226_ );
xor  ( new_n66231_, RIbb34ea8_250, RIbb34e30_249 );
xor  ( new_n66232_, RIbb35088_254, RIbb35010_253 );
xor  ( new_n66233_, new_n66232_, new_n66231_ );
xor  ( new_n66234_, RIbb349f8_240, RIbb34980_239 );
xor  ( new_n66235_, RIbb34548_230, RIbb344d0_229 );
xor  ( new_n66236_, new_n66235_, new_n65000_ );
xor  ( new_n66237_, new_n66236_, new_n66234_ );
xor  ( new_n66238_, RIbb34818_236, RIbb347a0_235 );
xor  ( new_n66239_, RIbb34728_234, new_n64974_ );
xor  ( new_n66240_, RIbb34908_238, RIbb34890_237 );
xor  ( new_n66241_, new_n66240_, new_n66239_ );
xor  ( new_n66242_, new_n66241_, new_n66238_ );
xor  ( new_n66243_, RIbb34638_232, new_n64952_ );
xor  ( new_n66244_, RIbb34458_228, new_n64986_ );
xor  ( new_n66245_, new_n66244_, new_n66243_ );
xor  ( new_n66246_, new_n66245_, new_n66242_ );
xor  ( new_n66247_, new_n66246_, new_n66237_ );
xor  ( new_n66248_, RIbb34f98_252, new_n65018_ );
xor  ( new_n66249_, new_n66248_, new_n66247_ );
xor  ( new_n66250_, new_n66249_, new_n66233_ );
xor  ( new_n66251_, RIbb33af8_208, new_n64971_ );
xor  ( new_n66252_, RIbb33468_194, new_n65001_ );
xor  ( new_n66253_, RIbb33648_198, RIbb335d0_197 );
xor  ( new_n66254_, new_n66253_, new_n66252_ );
xor  ( new_n66255_, new_n66254_, new_n66251_ );
xor  ( new_n66256_, RIbb33918_204, RIbb338a0_203 );
xor  ( new_n66257_, RIbb33828_202, new_n65013_ );
xor  ( new_n66258_, RIbb33a08_206, RIbb33990_205 );
xor  ( new_n66259_, new_n66258_, new_n66257_ );
xor  ( new_n66260_, new_n66259_, new_n66256_ );
xor  ( new_n66261_, RIbb33738_200, new_n64963_ );
xnor ( new_n66262_, RIbb33558_196, RIbb334e0_195 );
xor  ( new_n66263_, new_n66262_, new_n66261_ );
xor  ( new_n66264_, new_n66263_, new_n66260_ );
xor  ( new_n66265_, new_n66264_, new_n66255_ );
xor  ( new_n66266_, RIbb34098_220, new_n65006_ );
xor  ( new_n66267_, new_n66266_, new_n66265_ );
xor  ( new_n66268_, RIbb33eb8_216, RIbb33e40_215 );
xnor ( new_n66269_, RIbb33cd8_212, RIbb33c60_211 );
xor  ( new_n66270_, new_n66269_, new_n66268_ );
xnor ( new_n66271_, RIbb34278_224, RIbb34200_223 );
xor  ( new_n66272_, RIbb33be8_210, new_n65008_ );
xor  ( new_n66273_, RIbb33dc8_214, RIbb33d50_213 );
xor  ( new_n66274_, new_n66273_, new_n66272_ );
xor  ( new_n66275_, new_n66274_, new_n66271_ );
xor  ( new_n66276_, new_n66275_, new_n66270_ );
xnor ( new_n66277_, RIbb33fa8_218, RIbb33f30_217 );
xor  ( new_n66278_, RIbb34188_222, RIbb34110_221 );
xor  ( new_n66279_, new_n66278_, new_n66277_ );
xor  ( new_n66280_, new_n66279_, new_n66276_ );
xor  ( new_n66281_, new_n66280_, new_n66267_ );
xnor ( new_n66282_, RIbb34db8_248, RIbb34d40_247 );
xnor ( new_n66283_, RIbb34bd8_244, RIbb34b60_243 );
xor  ( new_n66284_, new_n66283_, new_n66282_ );
xor  ( new_n66285_, new_n66284_, new_n66281_ );
xor  ( new_n66286_, new_n66285_, new_n66250_ );
xor  ( new_n66287_, new_n66286_, new_n66230_ );
and  ( eq, new_n66287_, new_n66225_ );
endmodule


