module miter ( 
    RI2af433cd5b80_17, RI2af433cd5b08_16, RI2af433cd5a90_15,
    RI2af433cd5a18_14, RI2af433cd59a0_13, RI2af433cd5928_12,
    RI2af433cd58b0_11, RI2af433cd5838_10, RI2af433cd57c0_9,
    RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6, RI2af433cd55e0_5,
    RI2af433cd5568_4, RI2af433cd54f0_3, RI2af433cd5478_2, RI2af433cc8a70_1,
    RI2af433cd5bf8_18, RI2af433cd5c70_19, RI2af433cd5ce8_20,
    RI2af433cd5d60_21, RI2af433cd5dd8_22, RI2af433cd5e50_23,
    RI2af433cd5ec8_24, RI2af433cd5f40_25, RI2af433cd5fb8_26,
    RI2af433cd6030_27, RI2af433cd60a8_28, RI2af433cd6120_29,
    RI2af433cd6198_30, RI2af433cd6210_31, RI2af433cd6288_32,
    RI2af433cd6300_33, RI2af433cd6378_34, RI2af433cd63f0_35,
    RI2af433cd6468_36, RI2af433cd64e0_37, RI2af433cd6558_38,
    RI2af433cd65d0_39, RI2af433cd6648_40, RI2af433cd66c0_41,
    RI2af433cd6738_42, RI2af433cd67b0_43, RI2af433cd6828_44,
    RI2af433cd68a0_45, RI2af433cd6918_46, RI2af433cd6990_47,
    RI2af433cd6a08_48, RI2af433cd6a80_49, RI2af433cd6af8_50,
    RI2af433cd6b70_51, RI2af433cd6be8_52, RI2af433cd6c60_53,
    RI2af433cd6cd8_54, RI2af433cd6d50_55, RI2af433cd6dc8_56,
    RI2af433cd6e40_57, RI2af433cd6eb8_58, RI2af433cd6f30_59,
    RI2af433cd6fa8_60, RI2af433cd7020_61, RI2af433cd7098_62,
    RI2af433cd7110_63, RI2af433cd7188_64, RI2af433cd7200_65,
    RI2af433cd7278_66, RI2af433cd72f0_67, RI2af433cd7368_68,
    RI2af433cd73e0_69, RI2af433cd7458_70, RI2af433cd74d0_71,
    RI2af433cd7548_72, RI2af433cd75c0_73, RI2af433cd7638_74,
    RI2af433cd76b0_75, RI2af433cd7728_76, RI2af433cd77a0_77,
    RI2af433cd7818_78, RI2af433cd7890_79, RI2af433cd7908_80,
    RI2af433cd7980_81, RI2af433cd79f8_82, RI2af433cd7a70_83,
    RI2af433cd7ae8_84, RI2af433cd7b60_85, RI2af433cd7bd8_86,
    RI2af433cd7c50_87, RI2af433cd7cc8_88, RI2af433cd7d40_89,
    RI2af433cd7db8_90, RI2af433cd7e30_91, RI2af433cd7ea8_92,
    RI2af433cd7f20_93, RI2af433cd7f98_94, RI2af433cd8010_95,
    RI2af433cd8088_96, RI2af433cd8100_97, RI2af433cd8178_98,
    RI2af433cd81f0_99, RI2af433cd8268_100, RI2af433cd82e0_101,
    RI2af433cd8358_102, RI2af433cd83d0_103, RI2af433cd8448_104,
    RI2af433cd84c0_105, RI2af433cd8538_106, RI2af433cd85b0_107,
    RI2af433cd8628_108, RI2af433cd86a0_109, RI2af433cd8718_110,
    RI2af433cd8790_111, RI2af433cd8808_112, RI2af433cd8880_113,
    RI2af433cd88f8_114, RI2af433cd8970_115, RI2af433cd89e8_116,
    RI2af433cd8a60_117, RI2af433cd8ad8_118, RI2af433cd8b50_119,
    RI2af433cd8bc8_120, RI2af433cd8c40_121, RI2af433cd8cb8_122,
    RI2af433cd8d30_123, RI2af433cd8da8_124, RI2af433cd8e20_125,
    RI2af433cd8e98_126, RI2af433cd8f10_127, RI2af433cd8f88_128,
    RI2af433cd9000_129, RI2af433cd9078_130, RI2af433cd90f0_131,
    RI2af433cd9168_132, RI2af433cd91e0_133, RI2af433cd9258_134,
    RI2af433cd92d0_135, RI2af433cd9348_136, RI2af433cd93c0_137,
    RI2af433cd9438_138, RI2af433cd94b0_139, RI2af433cd9528_140,
    RI2af433cd95a0_141, RI2af433cd9618_142, RI2af433cd9690_143,
    RI2af433cd9708_144, RI2af433cd9780_145, RI2af433cd97f8_146,
    RI2af433cd9870_147, RI2af433cd98e8_148, RI2af433cd9960_149,
    RI2af433cd99d8_150, RI2af433cd9a50_151, RI2af433cd9ac8_152,
    RI2af433cd9b40_153, RI2af433cd9bb8_154, RI2af433cd9c30_155,
    RI2af433cd9ca8_156, RI2af433cd9d20_157, RI2af433cd9d98_158,
    RI2af433cd9e10_159, RI2af433cd9e88_160, RI2af433cd9f00_161,
    RI2af433cd9f78_162, RI2af433cd9ff0_163, RI2af433cda068_164,
    RI2af433cda0e0_165, RI2af433cda158_166, RI2af433cda1d0_167,
    RI2af433cda248_168, RI2af433cda2c0_169, RI2af433cda338_170,
    RI2af433cda3b0_171, RI2af433cda428_172, RI2af433cda4a0_173,
    RI2af433cda518_174, RI2af433cda590_175, RI2af433cda608_176,
    RI2af433cda680_177, RI2af433cda6f8_178, RI2af433cda770_179,
    RI2af433cda7e8_180, RI2af433cda860_181, RI2af433cda8d8_182,
    RI2af433cda950_183, RI2af433cda9c8_184, RI2af433cdaa40_185,
    RI2af433cdaab8_186, RI2af433cdab30_187, RI2af433cdaba8_188,
    RI2af433cdac20_189, RI2af433cdac98_190, RI2af433cdad10_191,
    RI2af433cdad88_192, RI2af433cdae00_193, RI2af433cdae78_194,
    RI2af433cdaef0_195, RI2af433cdaf68_196, RI2af433cdafe0_197,
    RI2af433cdb058_198, RI2af433cdb0d0_199, RI2af433cdb148_200,
    RI2af433cdb1c0_201, RI2af433cdb238_202, RI2af433cdb2b0_203,
    RI2af433cdb328_204, RI2af433cdb3a0_205, RI2af433cdb418_206,
    RI2af433cdb490_207, RI2af433cdb508_208, RI2af433cdb580_209,
    RI2af433cdb5f8_210, RI2af433cdb670_211, RI2af433cdb6e8_212,
    RI2af433cdb760_213, RI2af433cdb7d8_214, RI2af433cdb850_215,
    RI2af433cdb8c8_216, RI2af433cdb940_217,
    eq  );
  input  RI2af433cd5b80_17, RI2af433cd5b08_16, RI2af433cd5a90_15,
    RI2af433cd5a18_14, RI2af433cd59a0_13, RI2af433cd5928_12,
    RI2af433cd58b0_11, RI2af433cd5838_10, RI2af433cd57c0_9,
    RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6, RI2af433cd55e0_5,
    RI2af433cd5568_4, RI2af433cd54f0_3, RI2af433cd5478_2, RI2af433cc8a70_1,
    RI2af433cd5bf8_18, RI2af433cd5c70_19, RI2af433cd5ce8_20,
    RI2af433cd5d60_21, RI2af433cd5dd8_22, RI2af433cd5e50_23,
    RI2af433cd5ec8_24, RI2af433cd5f40_25, RI2af433cd5fb8_26,
    RI2af433cd6030_27, RI2af433cd60a8_28, RI2af433cd6120_29,
    RI2af433cd6198_30, RI2af433cd6210_31, RI2af433cd6288_32,
    RI2af433cd6300_33, RI2af433cd6378_34, RI2af433cd63f0_35,
    RI2af433cd6468_36, RI2af433cd64e0_37, RI2af433cd6558_38,
    RI2af433cd65d0_39, RI2af433cd6648_40, RI2af433cd66c0_41,
    RI2af433cd6738_42, RI2af433cd67b0_43, RI2af433cd6828_44,
    RI2af433cd68a0_45, RI2af433cd6918_46, RI2af433cd6990_47,
    RI2af433cd6a08_48, RI2af433cd6a80_49, RI2af433cd6af8_50,
    RI2af433cd6b70_51, RI2af433cd6be8_52, RI2af433cd6c60_53,
    RI2af433cd6cd8_54, RI2af433cd6d50_55, RI2af433cd6dc8_56,
    RI2af433cd6e40_57, RI2af433cd6eb8_58, RI2af433cd6f30_59,
    RI2af433cd6fa8_60, RI2af433cd7020_61, RI2af433cd7098_62,
    RI2af433cd7110_63, RI2af433cd7188_64, RI2af433cd7200_65,
    RI2af433cd7278_66, RI2af433cd72f0_67, RI2af433cd7368_68,
    RI2af433cd73e0_69, RI2af433cd7458_70, RI2af433cd74d0_71,
    RI2af433cd7548_72, RI2af433cd75c0_73, RI2af433cd7638_74,
    RI2af433cd76b0_75, RI2af433cd7728_76, RI2af433cd77a0_77,
    RI2af433cd7818_78, RI2af433cd7890_79, RI2af433cd7908_80,
    RI2af433cd7980_81, RI2af433cd79f8_82, RI2af433cd7a70_83,
    RI2af433cd7ae8_84, RI2af433cd7b60_85, RI2af433cd7bd8_86,
    RI2af433cd7c50_87, RI2af433cd7cc8_88, RI2af433cd7d40_89,
    RI2af433cd7db8_90, RI2af433cd7e30_91, RI2af433cd7ea8_92,
    RI2af433cd7f20_93, RI2af433cd7f98_94, RI2af433cd8010_95,
    RI2af433cd8088_96, RI2af433cd8100_97, RI2af433cd8178_98,
    RI2af433cd81f0_99, RI2af433cd8268_100, RI2af433cd82e0_101,
    RI2af433cd8358_102, RI2af433cd83d0_103, RI2af433cd8448_104,
    RI2af433cd84c0_105, RI2af433cd8538_106, RI2af433cd85b0_107,
    RI2af433cd8628_108, RI2af433cd86a0_109, RI2af433cd8718_110,
    RI2af433cd8790_111, RI2af433cd8808_112, RI2af433cd8880_113,
    RI2af433cd88f8_114, RI2af433cd8970_115, RI2af433cd89e8_116,
    RI2af433cd8a60_117, RI2af433cd8ad8_118, RI2af433cd8b50_119,
    RI2af433cd8bc8_120, RI2af433cd8c40_121, RI2af433cd8cb8_122,
    RI2af433cd8d30_123, RI2af433cd8da8_124, RI2af433cd8e20_125,
    RI2af433cd8e98_126, RI2af433cd8f10_127, RI2af433cd8f88_128,
    RI2af433cd9000_129, RI2af433cd9078_130, RI2af433cd90f0_131,
    RI2af433cd9168_132, RI2af433cd91e0_133, RI2af433cd9258_134,
    RI2af433cd92d0_135, RI2af433cd9348_136, RI2af433cd93c0_137,
    RI2af433cd9438_138, RI2af433cd94b0_139, RI2af433cd9528_140,
    RI2af433cd95a0_141, RI2af433cd9618_142, RI2af433cd9690_143,
    RI2af433cd9708_144, RI2af433cd9780_145, RI2af433cd97f8_146,
    RI2af433cd9870_147, RI2af433cd98e8_148, RI2af433cd9960_149,
    RI2af433cd99d8_150, RI2af433cd9a50_151, RI2af433cd9ac8_152,
    RI2af433cd9b40_153, RI2af433cd9bb8_154, RI2af433cd9c30_155,
    RI2af433cd9ca8_156, RI2af433cd9d20_157, RI2af433cd9d98_158,
    RI2af433cd9e10_159, RI2af433cd9e88_160, RI2af433cd9f00_161,
    RI2af433cd9f78_162, RI2af433cd9ff0_163, RI2af433cda068_164,
    RI2af433cda0e0_165, RI2af433cda158_166, RI2af433cda1d0_167,
    RI2af433cda248_168, RI2af433cda2c0_169, RI2af433cda338_170,
    RI2af433cda3b0_171, RI2af433cda428_172, RI2af433cda4a0_173,
    RI2af433cda518_174, RI2af433cda590_175, RI2af433cda608_176,
    RI2af433cda680_177, RI2af433cda6f8_178, RI2af433cda770_179,
    RI2af433cda7e8_180, RI2af433cda860_181, RI2af433cda8d8_182,
    RI2af433cda950_183, RI2af433cda9c8_184, RI2af433cdaa40_185,
    RI2af433cdaab8_186, RI2af433cdab30_187, RI2af433cdaba8_188,
    RI2af433cdac20_189, RI2af433cdac98_190, RI2af433cdad10_191,
    RI2af433cdad88_192, RI2af433cdae00_193, RI2af433cdae78_194,
    RI2af433cdaef0_195, RI2af433cdaf68_196, RI2af433cdafe0_197,
    RI2af433cdb058_198, RI2af433cdb0d0_199, RI2af433cdb148_200,
    RI2af433cdb1c0_201, RI2af433cdb238_202, RI2af433cdb2b0_203,
    RI2af433cdb328_204, RI2af433cdb3a0_205, RI2af433cdb418_206,
    RI2af433cdb490_207, RI2af433cdb508_208, RI2af433cdb580_209,
    RI2af433cdb5f8_210, RI2af433cdb670_211, RI2af433cdb6e8_212,
    RI2af433cdb760_213, RI2af433cdb7d8_214, RI2af433cdb850_215,
    RI2af433cdb8c8_216, RI2af433cdb940_217;
  output eq;
  wire new_n219_, new_n220_, new_n221_, new_n222_, new_n223_, new_n224_,
    new_n225_, new_n226_, new_n227_, new_n228_, new_n229_, new_n230_,
    new_n231_, new_n232_, new_n233_, new_n234_, new_n235_, new_n236_,
    new_n237_, new_n238_, new_n239_, new_n240_, new_n241_, new_n242_,
    new_n243_, new_n244_, new_n245_, new_n246_, new_n247_, new_n248_,
    new_n249_, new_n250_, new_n251_, new_n252_, new_n253_, new_n254_,
    new_n255_, new_n256_, new_n257_, new_n258_, new_n259_, new_n260_,
    new_n261_, new_n262_, new_n263_, new_n264_, new_n265_, new_n266_,
    new_n267_, new_n268_, new_n269_, new_n270_, new_n271_, new_n272_,
    new_n273_, new_n274_, new_n275_, new_n276_, new_n277_, new_n278_,
    new_n279_, new_n280_, new_n281_, new_n282_, new_n283_, new_n284_,
    new_n285_, new_n286_, new_n287_, new_n288_, new_n289_, new_n290_,
    new_n291_, new_n292_, new_n293_, new_n294_, new_n295_, new_n296_,
    new_n297_, new_n298_, new_n299_, new_n300_, new_n301_, new_n302_,
    new_n303_, new_n304_, new_n305_, new_n306_, new_n307_, new_n308_,
    new_n309_, new_n310_, new_n311_, new_n312_, new_n313_, new_n314_,
    new_n315_, new_n316_, new_n317_, new_n318_, new_n319_, new_n320_,
    new_n321_, new_n322_, new_n323_, new_n324_, new_n325_, new_n326_,
    new_n327_, new_n328_, new_n329_, new_n330_, new_n331_, new_n332_,
    new_n333_, new_n334_, new_n335_, new_n336_, new_n337_, new_n338_,
    new_n339_, new_n340_, new_n341_, new_n342_, new_n343_, new_n344_,
    new_n345_, new_n346_, new_n347_, new_n348_, new_n349_, new_n350_,
    new_n351_, new_n352_, new_n353_, new_n354_, new_n355_, new_n356_,
    new_n357_, new_n358_, new_n359_, new_n360_, new_n361_, new_n362_,
    new_n363_, new_n364_, new_n365_, new_n366_, new_n367_, new_n368_,
    new_n369_, new_n370_, new_n371_, new_n372_, new_n373_, new_n374_,
    new_n375_, new_n376_, new_n377_, new_n378_, new_n379_, new_n380_,
    new_n381_, new_n382_, new_n383_, new_n384_, new_n385_, new_n386_,
    new_n387_, new_n388_, new_n389_, new_n390_, new_n391_, new_n392_,
    new_n393_, new_n394_, new_n395_, new_n396_, new_n397_, new_n398_,
    new_n399_, new_n400_, new_n401_, new_n402_, new_n403_, new_n404_,
    new_n405_, new_n406_, new_n407_, new_n408_, new_n409_, new_n410_,
    new_n411_, new_n412_, new_n413_, new_n414_, new_n415_, new_n416_,
    new_n417_, new_n418_, new_n419_, new_n420_, new_n421_, new_n422_,
    new_n423_, new_n424_, new_n425_, new_n426_, new_n427_, new_n428_,
    new_n429_, new_n430_, new_n431_, new_n432_, new_n433_, new_n434_,
    new_n435_, new_n436_, new_n437_, new_n438_, new_n439_, new_n440_,
    new_n441_, new_n442_, new_n443_, new_n444_, new_n445_, new_n446_,
    new_n447_, new_n448_, new_n449_, new_n450_, new_n451_, new_n452_,
    new_n453_, new_n454_, new_n455_, new_n456_, new_n457_, new_n458_,
    new_n459_, new_n460_, new_n461_, new_n462_, new_n463_, new_n464_,
    new_n465_, new_n466_, new_n467_, new_n468_, new_n469_, new_n470_,
    new_n471_, new_n472_, new_n473_, new_n474_, new_n475_, new_n476_,
    new_n477_, new_n478_, new_n479_, new_n480_, new_n481_, new_n482_,
    new_n483_, new_n484_, new_n485_, new_n486_, new_n487_, new_n488_,
    new_n489_, new_n490_, new_n491_, new_n492_, new_n493_, new_n494_,
    new_n495_, new_n496_, new_n497_, new_n498_, new_n499_, new_n500_,
    new_n501_, new_n502_, new_n503_, new_n504_, new_n505_, new_n506_,
    new_n507_, new_n508_, new_n509_, new_n510_, new_n511_, new_n512_,
    new_n513_, new_n514_, new_n515_, new_n516_, new_n517_, new_n518_,
    new_n519_, new_n520_, new_n521_, new_n522_, new_n523_, new_n524_,
    new_n525_, new_n526_, new_n527_, new_n528_, new_n529_, new_n530_,
    new_n531_, new_n532_, new_n533_, new_n534_, new_n535_, new_n536_,
    new_n537_, new_n538_, new_n539_, new_n540_, new_n541_, new_n542_,
    new_n543_, new_n544_, new_n545_, new_n546_, new_n547_, new_n548_,
    new_n549_, new_n550_, new_n551_, new_n552_, new_n553_, new_n554_,
    new_n555_, new_n556_, new_n557_, new_n558_, new_n559_, new_n560_,
    new_n561_, new_n562_, new_n563_, new_n564_, new_n565_, new_n566_,
    new_n567_, new_n568_, new_n569_, new_n570_, new_n571_, new_n572_,
    new_n573_, new_n574_, new_n575_, new_n576_, new_n577_, new_n578_,
    new_n579_, new_n580_, new_n581_, new_n582_, new_n583_, new_n584_,
    new_n585_, new_n586_, new_n587_, new_n588_, new_n589_, new_n590_,
    new_n591_, new_n592_, new_n593_, new_n594_, new_n595_, new_n596_,
    new_n597_, new_n598_, new_n599_, new_n600_, new_n601_, new_n602_,
    new_n603_, new_n604_, new_n605_, new_n606_, new_n607_, new_n608_,
    new_n609_, new_n610_, new_n611_, new_n612_, new_n613_, new_n614_,
    new_n615_, new_n616_, new_n617_, new_n618_, new_n619_, new_n620_,
    new_n621_, new_n622_, new_n623_, new_n624_, new_n625_, new_n626_,
    new_n627_, new_n628_, new_n629_, new_n630_, new_n631_, new_n632_,
    new_n633_, new_n634_, new_n635_, new_n636_, new_n637_, new_n638_,
    new_n639_, new_n640_, new_n641_, new_n642_, new_n643_, new_n644_,
    new_n645_, new_n646_, new_n647_, new_n648_, new_n649_, new_n650_,
    new_n651_, new_n652_, new_n653_, new_n654_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n749_, new_n750_, new_n751_, new_n752_,
    new_n753_, new_n754_, new_n755_, new_n756_, new_n757_, new_n758_,
    new_n759_, new_n760_, new_n761_, new_n762_, new_n763_, new_n764_,
    new_n765_, new_n766_, new_n767_, new_n768_, new_n769_, new_n770_,
    new_n771_, new_n772_, new_n773_, new_n774_, new_n775_, new_n776_,
    new_n777_, new_n778_, new_n779_, new_n780_, new_n781_, new_n782_,
    new_n783_, new_n784_, new_n785_, new_n786_, new_n787_, new_n788_,
    new_n789_, new_n790_, new_n791_, new_n792_, new_n793_, new_n794_,
    new_n795_, new_n796_, new_n797_, new_n798_, new_n799_, new_n800_,
    new_n801_, new_n802_, new_n803_, new_n804_, new_n805_, new_n806_,
    new_n807_, new_n808_, new_n809_, new_n810_, new_n811_, new_n812_,
    new_n813_, new_n814_, new_n815_, new_n816_, new_n817_, new_n818_,
    new_n819_, new_n820_, new_n821_, new_n822_, new_n823_, new_n824_,
    new_n825_, new_n826_, new_n827_, new_n828_, new_n829_, new_n830_,
    new_n831_, new_n832_, new_n833_, new_n834_, new_n835_, new_n836_,
    new_n837_, new_n838_, new_n839_, new_n840_, new_n841_, new_n842_,
    new_n843_, new_n844_, new_n845_, new_n846_, new_n847_, new_n848_,
    new_n849_, new_n850_, new_n851_, new_n852_, new_n853_, new_n854_,
    new_n855_, new_n856_, new_n857_, new_n858_, new_n859_, new_n860_,
    new_n861_, new_n862_, new_n863_, new_n864_, new_n865_, new_n866_,
    new_n867_, new_n868_, new_n869_, new_n870_, new_n871_, new_n872_,
    new_n873_, new_n874_, new_n875_, new_n876_, new_n877_, new_n878_,
    new_n879_, new_n880_, new_n881_, new_n882_, new_n883_, new_n884_,
    new_n885_, new_n886_, new_n887_, new_n888_, new_n889_, new_n890_,
    new_n891_, new_n892_, new_n893_, new_n894_, new_n895_, new_n896_,
    new_n897_, new_n898_, new_n899_, new_n900_, new_n901_, new_n902_,
    new_n903_, new_n904_, new_n905_, new_n906_, new_n907_, new_n908_,
    new_n909_, new_n910_, new_n911_, new_n912_, new_n913_, new_n914_,
    new_n915_, new_n916_, new_n917_, new_n918_, new_n919_, new_n920_,
    new_n921_, new_n922_, new_n923_, new_n924_, new_n925_, new_n926_,
    new_n927_, new_n928_, new_n929_, new_n930_, new_n931_, new_n932_,
    new_n933_, new_n934_, new_n935_, new_n936_, new_n937_, new_n938_,
    new_n939_, new_n940_, new_n941_, new_n942_, new_n943_, new_n944_,
    new_n945_, new_n946_, new_n947_, new_n948_, new_n949_, new_n950_,
    new_n951_, new_n952_, new_n953_, new_n954_, new_n955_, new_n956_,
    new_n957_, new_n958_, new_n959_, new_n960_, new_n961_, new_n962_,
    new_n963_, new_n964_, new_n965_, new_n966_, new_n967_, new_n968_,
    new_n969_, new_n970_, new_n971_, new_n972_, new_n973_, new_n974_,
    new_n975_, new_n976_, new_n977_, new_n978_, new_n979_, new_n980_,
    new_n981_, new_n982_, new_n983_, new_n984_, new_n985_, new_n986_,
    new_n987_, new_n988_, new_n989_, new_n990_, new_n991_, new_n992_,
    new_n993_, new_n994_, new_n995_, new_n996_, new_n997_, new_n998_,
    new_n999_, new_n1000_, new_n1001_, new_n1002_, new_n1003_, new_n1004_,
    new_n1005_, new_n1006_;
not  ( new_n219_, RI2af433cd5928_12 );
and  ( new_n220_, RI2af433cd58b0_11, new_n219_ );
not  ( new_n221_, RI2af433cd59a0_13 );
not  ( new_n222_, RI2af433cd5a90_15 );
and  ( new_n223_, new_n222_, RI2af433cd5b08_16 );
and  ( new_n224_, new_n223_, RI2af433cd5a18_14 );
and  ( new_n225_, new_n224_, new_n221_ );
and  ( new_n226_, new_n225_, new_n220_ );
and  ( new_n227_, new_n226_, RI2af433cd6be8_52 );
not  ( new_n228_, RI2af433cd5b08_16 );
and  ( new_n229_, RI2af433cd5a90_15, new_n228_ );
and  ( new_n230_, new_n229_, RI2af433cd5a18_14 );
and  ( new_n231_, new_n230_, RI2af433cd59a0_13 );
and  ( new_n232_, new_n231_, new_n220_ );
and  ( new_n233_, new_n232_, RI2af433cd67b0_43 );
nor  ( new_n234_, new_n233_, new_n227_ );
not  ( new_n235_, RI2af433cd5a18_14 );
and  ( new_n236_, new_n229_, new_n235_ );
and  ( new_n237_, new_n236_, RI2af433cd59a0_13 );
and  ( new_n238_, new_n237_, new_n220_ );
and  ( new_n239_, new_n238_, RI2af433cd6990_47 );
and  ( new_n240_, new_n222_, new_n228_ );
and  ( new_n241_, new_n240_, RI2af433cd5a18_14 );
and  ( new_n242_, new_n241_, new_n221_ );
and  ( new_n243_, new_n242_, new_n220_ );
and  ( new_n244_, new_n243_, RI2af433cd6c60_53 );
nor  ( new_n245_, new_n244_, new_n239_ );
and  ( new_n246_, new_n245_, new_n234_ );
and  ( new_n247_, RI2af433cd5a90_15, RI2af433cd5b08_16 );
and  ( new_n248_, new_n247_, RI2af433cd5a18_14 );
and  ( new_n249_, new_n248_, new_n221_ );
and  ( new_n250_, new_n249_, new_n220_ );
and  ( new_n251_, new_n250_, RI2af433cd6af8_50 );
nor  ( new_n252_, new_n251_, RI2af433cd5838_10 );
and  ( new_n253_, new_n236_, new_n221_ );
and  ( new_n254_, new_n253_, new_n220_ );
and  ( new_n255_, new_n254_, RI2af433cd6d50_55 );
and  ( new_n256_, new_n230_, new_n221_ );
and  ( new_n257_, new_n256_, new_n220_ );
and  ( new_n258_, new_n257_, RI2af433cd6b70_51 );
nor  ( new_n259_, new_n258_, new_n255_ );
and  ( new_n260_, new_n259_, new_n252_ );
and  ( new_n261_, new_n260_, new_n246_ );
and  ( new_n262_, new_n224_, RI2af433cd59a0_13 );
and  ( new_n263_, new_n262_, new_n220_ );
and  ( new_n264_, new_n263_, RI2af433cd6828_44 );
not  ( new_n265_, new_n264_ );
and  ( new_n266_, new_n248_, RI2af433cd59a0_13 );
and  ( new_n267_, new_n266_, new_n220_ );
and  ( new_n268_, new_n267_, RI2af433cd6738_42 );
and  ( new_n269_, new_n223_, new_n235_ );
and  ( new_n270_, new_n269_, RI2af433cd59a0_13 );
and  ( new_n271_, new_n270_, new_n220_ );
and  ( new_n272_, new_n271_, RI2af433cd6a08_48 );
nor  ( new_n273_, new_n272_, new_n268_ );
and  ( new_n274_, new_n273_, new_n265_ );
and  ( new_n275_, new_n247_, new_n235_ );
and  ( new_n276_, new_n275_, new_n221_ );
and  ( new_n277_, new_n276_, new_n220_ );
and  ( new_n278_, new_n277_, RI2af433cd6cd8_54 );
and  ( new_n279_, new_n241_, RI2af433cd59a0_13 );
and  ( new_n280_, new_n279_, new_n220_ );
and  ( new_n281_, new_n280_, RI2af433cd68a0_45 );
nor  ( new_n282_, new_n281_, new_n278_ );
and  ( new_n283_, new_n240_, new_n235_ );
and  ( new_n284_, new_n283_, RI2af433cd59a0_13 );
and  ( new_n285_, new_n284_, new_n220_ );
and  ( new_n286_, new_n285_, RI2af433cd6a80_49 );
and  ( new_n287_, new_n275_, RI2af433cd59a0_13 );
and  ( new_n288_, new_n287_, new_n220_ );
and  ( new_n289_, new_n288_, RI2af433cd6918_46 );
nor  ( new_n290_, new_n289_, new_n286_ );
and  ( new_n291_, new_n290_, new_n282_ );
and  ( new_n292_, new_n291_, new_n274_ );
and  ( new_n293_, new_n292_, new_n261_ );
and  ( new_n294_, new_n262_, RI2af433cd5928_12 );
and  ( new_n295_, new_n294_, RI2af433cd58b0_11 );
and  ( new_n296_, new_n295_, RI2af433cd60a8_28 );
and  ( new_n297_, new_n283_, new_n221_ );
and  ( new_n298_, new_n297_, RI2af433cd5928_12 );
and  ( new_n299_, new_n298_, RI2af433cd58b0_11 );
and  ( new_n300_, new_n299_, RI2af433cd66c0_41 );
nor  ( new_n301_, new_n300_, new_n296_ );
and  ( new_n302_, new_n279_, RI2af433cd5928_12 );
and  ( new_n303_, new_n302_, RI2af433cd58b0_11 );
and  ( new_n304_, new_n303_, RI2af433cd6120_29 );
and  ( new_n305_, new_n287_, RI2af433cd5928_12 );
and  ( new_n306_, new_n305_, RI2af433cd58b0_11 );
and  ( new_n307_, new_n306_, RI2af433cd6198_30 );
nor  ( new_n308_, new_n307_, new_n304_ );
and  ( new_n309_, new_n308_, new_n301_ );
and  ( new_n310_, new_n276_, RI2af433cd5928_12 );
and  ( new_n311_, new_n310_, RI2af433cd58b0_11 );
and  ( new_n312_, new_n311_, RI2af433cd6558_38 );
and  ( new_n313_, new_n266_, RI2af433cd5928_12 );
and  ( new_n314_, new_n313_, RI2af433cd58b0_11 );
and  ( new_n315_, new_n314_, RI2af433cd5fb8_26 );
nor  ( new_n316_, new_n315_, new_n312_ );
and  ( new_n317_, new_n231_, RI2af433cd5928_12 );
and  ( new_n318_, new_n317_, RI2af433cd58b0_11 );
and  ( new_n319_, new_n318_, RI2af433cd6030_27 );
and  ( new_n320_, new_n253_, RI2af433cd5928_12 );
and  ( new_n321_, new_n320_, RI2af433cd58b0_11 );
and  ( new_n322_, new_n321_, RI2af433cd65d0_39 );
nor  ( new_n323_, new_n322_, new_n319_ );
and  ( new_n324_, new_n323_, new_n316_ );
and  ( new_n325_, new_n324_, new_n309_ );
and  ( new_n326_, new_n284_, RI2af433cd5928_12 );
and  ( new_n327_, new_n326_, RI2af433cd58b0_11 );
and  ( new_n328_, new_n327_, RI2af433cd6300_33 );
and  ( new_n329_, new_n249_, RI2af433cd5928_12 );
and  ( new_n330_, new_n329_, RI2af433cd58b0_11 );
and  ( new_n331_, new_n330_, RI2af433cd6378_34 );
nor  ( new_n332_, new_n331_, new_n328_ );
and  ( new_n333_, new_n225_, RI2af433cd5928_12 );
and  ( new_n334_, new_n333_, RI2af433cd58b0_11 );
and  ( new_n335_, new_n334_, RI2af433cd6468_36 );
and  ( new_n336_, new_n270_, RI2af433cd5928_12 );
and  ( new_n337_, new_n336_, RI2af433cd58b0_11 );
and  ( new_n338_, new_n337_, RI2af433cd6288_32 );
nor  ( new_n339_, new_n338_, new_n335_ );
and  ( new_n340_, new_n339_, new_n332_ );
and  ( new_n341_, new_n237_, RI2af433cd5928_12 );
and  ( new_n342_, new_n341_, RI2af433cd58b0_11 );
and  ( new_n343_, new_n342_, RI2af433cd6210_31 );
and  ( new_n344_, new_n242_, RI2af433cd5928_12 );
and  ( new_n345_, new_n344_, RI2af433cd58b0_11 );
and  ( new_n346_, new_n345_, RI2af433cd64e0_37 );
nor  ( new_n347_, new_n346_, new_n343_ );
and  ( new_n348_, new_n269_, new_n221_ );
and  ( new_n349_, new_n348_, RI2af433cd5928_12 );
and  ( new_n350_, new_n349_, RI2af433cd58b0_11 );
and  ( new_n351_, new_n350_, RI2af433cd6648_40 );
and  ( new_n352_, new_n256_, RI2af433cd5928_12 );
and  ( new_n353_, new_n352_, RI2af433cd58b0_11 );
and  ( new_n354_, new_n353_, RI2af433cd63f0_35 );
nor  ( new_n355_, new_n354_, new_n351_ );
and  ( new_n356_, new_n355_, new_n347_ );
and  ( new_n357_, new_n356_, new_n340_ );
and  ( new_n358_, new_n357_, new_n325_ );
and  ( new_n359_, new_n358_, new_n293_ );
not  ( new_n360_, new_n359_ );
not  ( new_n361_, RI2af433cd5658_6 );
nor  ( new_n362_, RI2af433cd56d0_7, RI2af433cd5748_8 );
and  ( new_n363_, new_n362_, new_n361_ );
and  ( new_n364_, new_n363_, RI2af433cd57c0_9 );
not  ( new_n365_, new_n364_ );
not  ( new_n366_, RI2af433cd58b0_11 );
and  ( new_n367_, new_n366_, new_n219_ );
and  ( new_n368_, new_n367_, new_n297_ );
and  ( new_n369_, new_n368_, RI2af433cd5f40_25 );
not  ( new_n370_, new_n369_ );
not  ( new_n371_, RI2af433cd5838_10 );
and  ( new_n372_, new_n367_, new_n348_ );
and  ( new_n373_, new_n372_, RI2af433cd5ec8_24 );
nor  ( new_n374_, new_n373_, new_n371_ );
and  ( new_n375_, new_n374_, new_n370_ );
nor  ( new_n376_, new_n375_, new_n365_ );
and  ( new_n377_, new_n376_, new_n360_ );
and  ( new_n378_, new_n367_, new_n284_ );
and  ( new_n379_, new_n378_, RI2af433cd7980_81 );
and  ( new_n380_, new_n367_, new_n256_ );
and  ( new_n381_, new_n380_, RI2af433cd7a70_83 );
nor  ( new_n382_, new_n381_, new_n379_ );
and  ( new_n383_, new_n368_, RI2af433cd7d40_89 );
and  ( new_n384_, new_n367_, new_n253_ );
and  ( new_n385_, new_n384_, RI2af433cd7c50_87 );
nor  ( new_n386_, new_n385_, new_n383_ );
and  ( new_n387_, new_n386_, new_n382_ );
and  ( new_n388_, new_n367_, new_n242_ );
and  ( new_n389_, new_n388_, RI2af433cd7b60_85 );
nor  ( new_n390_, new_n389_, RI2af433cd5838_10 );
and  ( new_n391_, new_n372_, RI2af433cd7cc8_88 );
and  ( new_n392_, new_n367_, new_n276_ );
and  ( new_n393_, new_n392_, RI2af433cd7bd8_86 );
nor  ( new_n394_, new_n393_, new_n391_ );
and  ( new_n395_, new_n367_, new_n225_ );
and  ( new_n396_, new_n395_, RI2af433cd7ae8_84 );
and  ( new_n397_, new_n367_, new_n249_ );
and  ( new_n398_, new_n397_, RI2af433cd79f8_82 );
nor  ( new_n399_, new_n398_, new_n396_ );
and  ( new_n400_, new_n399_, new_n394_ );
and  ( new_n401_, new_n400_, new_n390_ );
and  ( new_n402_, new_n401_, new_n387_ );
not  ( new_n403_, new_n402_ );
and  ( new_n404_, new_n397_, RI2af433cd5bf8_18 );
and  ( new_n405_, new_n378_, RI2af433cd5b80_17 );
nor  ( new_n406_, new_n405_, new_n404_ );
and  ( new_n407_, new_n380_, RI2af433cd5c70_19 );
and  ( new_n408_, new_n392_, RI2af433cd5dd8_22 );
nor  ( new_n409_, new_n408_, new_n407_ );
and  ( new_n410_, new_n409_, new_n406_ );
and  ( new_n411_, new_n384_, RI2af433cd5e50_23 );
nor  ( new_n412_, new_n411_, new_n371_ );
and  ( new_n413_, new_n395_, RI2af433cd5ce8_20 );
and  ( new_n414_, new_n388_, RI2af433cd5d60_21 );
nor  ( new_n415_, new_n414_, new_n413_ );
and  ( new_n416_, new_n415_, new_n412_ );
and  ( new_n417_, new_n416_, new_n410_ );
nor  ( new_n418_, new_n417_, new_n365_ );
and  ( new_n419_, new_n418_, new_n403_ );
nor  ( new_n420_, new_n419_, new_n377_ );
nor  ( new_n421_, RI2af433cd5568_4, RI2af433cd55e0_5 );
not  ( new_n422_, RI2af433cc8a70_1 );
nor  ( new_n423_, RI2af433cd5478_2, RI2af433cd54f0_3 );
and  ( new_n424_, new_n423_, new_n422_ );
and  ( new_n425_, new_n424_, new_n421_ );
not  ( new_n426_, new_n425_ );
or   ( new_n427_, new_n426_, new_n420_ );
not  ( new_n428_, RI2af433cd57c0_9 );
and  ( new_n429_, new_n363_, new_n428_ );
and  ( new_n430_, new_n429_, RI2af433cd5838_10 );
not  ( new_n431_, new_n430_ );
and  ( new_n432_, new_n318_, RI2af433cd7e30_91 );
not  ( new_n433_, new_n432_ );
and  ( new_n434_, new_n314_, RI2af433cd7db8_90 );
and  ( new_n435_, new_n295_, RI2af433cd7ea8_92 );
nor  ( new_n436_, new_n435_, new_n434_ );
and  ( new_n437_, new_n436_, new_n433_ );
nor  ( new_n438_, new_n437_, new_n431_ );
not  ( new_n439_, new_n438_ );
and  ( new_n440_, new_n280_, RI2af433cd86a0_109 );
and  ( new_n441_, new_n226_, RI2af433cd89e8_116 );
nor  ( new_n442_, new_n441_, new_n440_ );
and  ( new_n443_, new_n257_, RI2af433cd8970_115 );
and  ( new_n444_, new_n250_, RI2af433cd88f8_114 );
nor  ( new_n445_, new_n444_, new_n443_ );
and  ( new_n446_, new_n445_, new_n442_ );
nor  ( new_n447_, new_n446_, new_n431_ );
not  ( new_n448_, new_n447_ );
and  ( new_n449_, new_n297_, new_n220_ );
and  ( new_n450_, new_n429_, new_n371_ );
and  ( new_n451_, new_n450_, RI2af433cdaa40_185 );
and  ( new_n452_, new_n451_, new_n449_ );
and  ( new_n453_, new_n302_, new_n366_ );
and  ( new_n454_, new_n450_, RI2af433cdac20_189 );
and  ( new_n455_, new_n454_, new_n453_ );
nor  ( new_n456_, new_n455_, new_n452_ );
and  ( new_n457_, new_n367_, new_n266_ );
and  ( new_n458_, new_n450_, RI2af433cdb238_202 );
and  ( new_n459_, new_n458_, new_n457_ );
and  ( new_n460_, new_n367_, new_n231_ );
and  ( new_n461_, new_n450_, RI2af433cdb2b0_203 );
and  ( new_n462_, new_n461_, new_n460_ );
nor  ( new_n463_, new_n462_, new_n459_ );
and  ( new_n464_, new_n463_, new_n456_ );
and  ( new_n465_, new_n464_, new_n448_ );
and  ( new_n466_, new_n465_, new_n439_ );
not  ( new_n467_, new_n450_ );
and  ( new_n468_, new_n341_, new_n366_ );
and  ( new_n469_, new_n468_, RI2af433cdad10_191 );
not  ( new_n470_, new_n469_ );
and  ( new_n471_, new_n294_, new_n366_ );
and  ( new_n472_, new_n471_, RI2af433cdaba8_188 );
not  ( new_n473_, new_n472_ );
and  ( new_n474_, new_n367_, new_n270_ );
and  ( new_n475_, new_n474_, RI2af433cdb508_208 );
and  ( new_n476_, new_n348_, new_n220_ );
and  ( new_n477_, new_n476_, RI2af433cda9c8_184 );
nor  ( new_n478_, new_n477_, new_n475_ );
and  ( new_n479_, new_n478_, new_n473_ );
and  ( new_n480_, new_n479_, new_n470_ );
nor  ( new_n481_, new_n480_, new_n467_ );
and  ( new_n482_, new_n367_, new_n279_ );
and  ( new_n483_, new_n482_, RI2af433cdb3a0_205 );
and  ( new_n484_, new_n367_, new_n237_ );
and  ( new_n485_, new_n484_, RI2af433cdb490_207 );
nor  ( new_n486_, new_n485_, new_n483_ );
and  ( new_n487_, new_n367_, new_n287_ );
and  ( new_n488_, new_n487_, RI2af433cdb418_206 );
and  ( new_n489_, new_n367_, new_n262_ );
and  ( new_n490_, new_n489_, RI2af433cdb328_204 );
nor  ( new_n491_, new_n490_, new_n488_ );
and  ( new_n492_, new_n491_, new_n486_ );
and  ( new_n493_, new_n298_, new_n366_ );
and  ( new_n494_, new_n493_, RI2af433cdb1c0_201 );
and  ( new_n495_, new_n349_, new_n366_ );
and  ( new_n496_, new_n495_, RI2af433cdb148_200 );
nor  ( new_n497_, new_n496_, new_n494_ );
and  ( new_n498_, new_n497_, new_n492_ );
nor  ( new_n499_, new_n498_, new_n467_ );
nor  ( new_n500_, new_n499_, new_n481_ );
and  ( new_n501_, new_n500_, new_n466_ );
and  ( new_n502_, new_n395_, RI2af433cdb6e8_212 );
not  ( new_n503_, new_n502_ );
and  ( new_n504_, new_n378_, RI2af433cdb580_209 );
and  ( new_n505_, new_n388_, RI2af433cdb760_213 );
nor  ( new_n506_, new_n505_, new_n504_ );
and  ( new_n507_, new_n506_, new_n503_ );
and  ( new_n508_, new_n397_, RI2af433cdb5f8_210 );
and  ( new_n509_, new_n384_, RI2af433cdb850_215 );
nor  ( new_n510_, new_n509_, new_n508_ );
and  ( new_n511_, new_n392_, RI2af433cdb7d8_214 );
and  ( new_n512_, new_n380_, RI2af433cdb670_211 );
nor  ( new_n513_, new_n512_, new_n511_ );
and  ( new_n514_, new_n513_, new_n510_ );
and  ( new_n515_, new_n514_, new_n507_ );
nor  ( new_n516_, new_n515_, new_n467_ );
not  ( new_n517_, new_n516_ );
and  ( new_n518_, new_n482_, RI2af433cd95a0_141 );
not  ( new_n519_, new_n518_ );
and  ( new_n520_, new_n487_, RI2af433cd9618_142 );
and  ( new_n521_, new_n484_, RI2af433cd9690_143 );
nor  ( new_n522_, new_n521_, new_n520_ );
and  ( new_n523_, new_n522_, new_n519_ );
nor  ( new_n524_, new_n523_, new_n431_ );
not  ( new_n525_, new_n524_ );
and  ( new_n526_, new_n430_, RI2af433cd84c0_105 );
and  ( new_n527_, new_n526_, new_n299_ );
and  ( new_n528_, new_n368_, RI2af433cdb940_217 );
and  ( new_n529_, new_n528_, new_n450_ );
nor  ( new_n530_, new_n529_, new_n527_ );
and  ( new_n531_, new_n530_, new_n525_ );
and  ( new_n532_, new_n531_, new_n517_ );
and  ( new_n533_, new_n254_, RI2af433cda950_183 );
and  ( new_n534_, new_n277_, RI2af433cda8d8_182 );
nor  ( new_n535_, new_n534_, new_n533_ );
and  ( new_n536_, new_n243_, RI2af433cda860_181 );
and  ( new_n537_, new_n226_, RI2af433cda7e8_180 );
nor  ( new_n538_, new_n537_, new_n536_ );
and  ( new_n539_, new_n538_, new_n535_ );
nor  ( new_n540_, new_n539_, new_n467_ );
not  ( new_n541_, new_n540_ );
and  ( new_n542_, new_n257_, RI2af433cda770_179 );
and  ( new_n543_, new_n250_, RI2af433cda6f8_178 );
nor  ( new_n544_, new_n543_, new_n542_ );
and  ( new_n545_, new_n285_, RI2af433cda680_177 );
and  ( new_n546_, new_n271_, RI2af433cda608_176 );
nor  ( new_n547_, new_n546_, new_n545_ );
and  ( new_n548_, new_n547_, new_n544_ );
nor  ( new_n549_, new_n548_, new_n467_ );
not  ( new_n550_, new_n549_ );
and  ( new_n551_, new_n313_, new_n366_ );
and  ( new_n552_, new_n551_, RI2af433cdaab8_186 );
and  ( new_n553_, new_n305_, new_n366_ );
and  ( new_n554_, new_n553_, RI2af433cdac98_190 );
nor  ( new_n555_, new_n554_, new_n552_ );
nor  ( new_n556_, new_n555_, new_n467_ );
not  ( new_n557_, new_n556_ );
and  ( new_n558_, new_n557_, new_n550_ );
and  ( new_n559_, new_n558_, new_n541_ );
and  ( new_n560_, new_n559_, new_n532_ );
and  ( new_n561_, new_n560_, new_n501_ );
nor  ( new_n562_, new_n561_, new_n426_ );
not  ( new_n563_, new_n562_ );
and  ( new_n564_, new_n263_, RI2af433cd8628_108 );
and  ( new_n565_, new_n564_, new_n430_ );
and  ( new_n566_, new_n565_, new_n425_ );
and  ( new_n567_, new_n430_, new_n425_ );
and  ( new_n568_, new_n345_, RI2af433cd82e0_101 );
and  ( new_n569_, new_n568_, new_n567_ );
nor  ( new_n570_, new_n569_, new_n566_ );
and  ( new_n571_, new_n271_, RI2af433cd8808_112 );
and  ( new_n572_, new_n571_, new_n430_ );
and  ( new_n573_, new_n572_, new_n425_ );
and  ( new_n574_, new_n327_, RI2af433cd8100_97 );
and  ( new_n575_, new_n574_, new_n567_ );
nor  ( new_n576_, new_n575_, new_n573_ );
and  ( new_n577_, new_n576_, new_n570_ );
and  ( new_n578_, new_n243_, RI2af433cd8a60_117 );
and  ( new_n579_, new_n578_, new_n430_ );
and  ( new_n580_, new_n579_, new_n425_ );
and  ( new_n581_, new_n567_, RI2af433cd8da8_124 );
and  ( new_n582_, new_n581_, new_n471_ );
nor  ( new_n583_, new_n582_, new_n580_ );
and  ( new_n584_, new_n395_, RI2af433cd98e8_148 );
and  ( new_n585_, new_n584_, new_n430_ );
and  ( new_n586_, new_n585_, new_n425_ );
and  ( new_n587_, new_n336_, new_n366_ );
and  ( new_n588_, new_n567_, RI2af433cd8f88_128 );
and  ( new_n589_, new_n588_, new_n587_ );
nor  ( new_n590_, new_n589_, new_n586_ );
and  ( new_n591_, new_n590_, new_n583_ );
and  ( new_n592_, new_n591_, new_n577_ );
not  ( new_n593_, new_n342_ );
and  ( new_n594_, new_n450_, RI2af433cd9e10_159 );
and  ( new_n595_, new_n430_, RI2af433cd8010_95 );
nor  ( new_n596_, new_n595_, new_n594_ );
nor  ( new_n597_, new_n596_, new_n593_ );
not  ( new_n598_, new_n306_ );
and  ( new_n599_, new_n450_, RI2af433cd9d98_158 );
and  ( new_n600_, new_n430_, RI2af433cd7f98_94 );
nor  ( new_n601_, new_n600_, new_n599_ );
nor  ( new_n602_, new_n601_, new_n598_ );
nor  ( new_n603_, new_n602_, new_n597_ );
nor  ( new_n604_, new_n603_, new_n426_ );
not  ( new_n605_, new_n567_ );
and  ( new_n606_, new_n317_, new_n366_ );
and  ( new_n607_, new_n606_, RI2af433cd8d30_123 );
and  ( new_n608_, new_n551_, RI2af433cd8cb8_122 );
nor  ( new_n609_, new_n608_, new_n607_ );
and  ( new_n610_, new_n468_, RI2af433cd8f10_127 );
and  ( new_n611_, new_n553_, RI2af433cd8e98_126 );
nor  ( new_n612_, new_n611_, new_n610_ );
and  ( new_n613_, new_n612_, new_n609_ );
nor  ( new_n614_, new_n613_, new_n605_ );
nor  ( new_n615_, new_n614_, new_n604_ );
and  ( new_n616_, new_n615_, new_n592_ );
and  ( new_n617_, new_n450_, new_n303_ );
and  ( new_n618_, new_n425_, RI2af433cd9d20_157 );
and  ( new_n619_, new_n618_, new_n617_ );
and  ( new_n620_, new_n450_, new_n295_ );
and  ( new_n621_, new_n425_, RI2af433cd9ca8_156 );
and  ( new_n622_, new_n621_, new_n620_ );
nor  ( new_n623_, new_n622_, new_n619_ );
and  ( new_n624_, new_n450_, new_n299_ );
and  ( new_n625_, new_n425_, RI2af433cda2c0_169 );
and  ( new_n626_, new_n625_, new_n624_ );
and  ( new_n627_, new_n450_, new_n350_ );
and  ( new_n628_, new_n425_, RI2af433cda248_168 );
and  ( new_n629_, new_n628_, new_n627_ );
nor  ( new_n630_, new_n629_, new_n626_ );
and  ( new_n631_, new_n630_, new_n623_ );
and  ( new_n632_, new_n321_, RI2af433cd83d0_103 );
and  ( new_n633_, new_n311_, RI2af433cd8358_102 );
nor  ( new_n634_, new_n633_, new_n632_ );
nor  ( new_n635_, new_n634_, new_n605_ );
and  ( new_n636_, new_n352_, new_n366_ );
and  ( new_n637_, new_n636_, RI2af433cd90f0_131 );
and  ( new_n638_, new_n329_, new_n366_ );
and  ( new_n639_, new_n638_, RI2af433cd9078_130 );
nor  ( new_n640_, new_n639_, new_n637_ );
not  ( new_n641_, new_n640_ );
and  ( new_n642_, new_n641_, new_n567_ );
nor  ( new_n643_, new_n642_, new_n635_ );
and  ( new_n644_, new_n643_, new_n631_ );
and  ( new_n645_, new_n285_, RI2af433cd8880_113 );
and  ( new_n646_, new_n645_, new_n430_ );
and  ( new_n647_, new_n646_, new_n425_ );
and  ( new_n648_, new_n350_, RI2af433cd8448_104 );
and  ( new_n649_, new_n648_, new_n567_ );
nor  ( new_n650_, new_n649_, new_n647_ );
and  ( new_n651_, new_n430_, RI2af433cd8bc8_120 );
and  ( new_n652_, new_n651_, new_n476_ );
and  ( new_n653_, new_n652_, new_n425_ );
and  ( new_n654_, new_n326_, new_n366_ );
and  ( new_n655_, new_n567_, RI2af433cd9000_129 );
and  ( new_n656_, new_n655_, new_n654_ );
nor  ( new_n657_, new_n656_, new_n653_ );
and  ( new_n658_, new_n657_, new_n650_ );
and  ( new_n659_, new_n430_, RI2af433cd9528_140 );
and  ( new_n660_, new_n659_, new_n489_ );
and  ( new_n661_, new_n660_, new_n425_ );
and  ( new_n662_, new_n344_, new_n366_ );
and  ( new_n663_, new_n662_, RI2af433cd91e0_133 );
and  ( new_n664_, new_n663_, new_n567_ );
nor  ( new_n665_, new_n664_, new_n661_ );
and  ( new_n666_, new_n372_, RI2af433cdb8c8_216 );
and  ( new_n667_, new_n666_, new_n450_ );
and  ( new_n668_, new_n667_, new_n425_ );
and  ( new_n669_, new_n567_, RI2af433cd9348_136 );
and  ( new_n670_, new_n669_, new_n495_ );
nor  ( new_n671_, new_n670_, new_n668_ );
and  ( new_n672_, new_n671_, new_n665_ );
and  ( new_n673_, new_n672_, new_n658_ );
and  ( new_n674_, new_n673_, new_n644_ );
and  ( new_n675_, new_n674_, new_n616_ );
and  ( new_n676_, new_n450_, RI2af433cdae78_194 );
and  ( new_n677_, new_n676_, new_n638_ );
and  ( new_n678_, new_n450_, RI2af433cdae00_193 );
and  ( new_n679_, new_n678_, new_n654_ );
nor  ( new_n680_, new_n679_, new_n677_ );
and  ( new_n681_, new_n450_, RI2af433cdaef0_195 );
and  ( new_n682_, new_n681_, new_n636_ );
and  ( new_n683_, new_n364_, new_n371_ );
and  ( new_n684_, new_n489_, RI2af433cd7728_76 );
and  ( new_n685_, new_n684_, new_n683_ );
nor  ( new_n686_, new_n685_, new_n682_ );
and  ( new_n687_, new_n686_, new_n680_ );
and  ( new_n688_, new_n320_, new_n366_ );
and  ( new_n689_, new_n683_, RI2af433cd74d0_71 );
and  ( new_n690_, new_n689_, new_n688_ );
and  ( new_n691_, new_n310_, new_n366_ );
and  ( new_n692_, new_n683_, RI2af433cd7458_70 );
and  ( new_n693_, new_n692_, new_n691_ );
nor  ( new_n694_, new_n693_, new_n690_ );
and  ( new_n695_, new_n683_, RI2af433cd7188_64 );
and  ( new_n696_, new_n695_, new_n587_ );
and  ( new_n697_, new_n683_, RI2af433cd7200_65 );
and  ( new_n698_, new_n697_, new_n654_ );
nor  ( new_n699_, new_n698_, new_n696_ );
and  ( new_n700_, new_n699_, new_n694_ );
and  ( new_n701_, new_n700_, new_n687_ );
and  ( new_n702_, new_n333_, new_n366_ );
and  ( new_n703_, new_n450_, RI2af433cdaf68_196 );
and  ( new_n704_, new_n703_, new_n702_ );
and  ( new_n705_, new_n450_, RI2af433cdab30_187 );
and  ( new_n706_, new_n705_, new_n606_ );
nor  ( new_n707_, new_n706_, new_n704_ );
and  ( new_n708_, new_n450_, RI2af433cdafe0_197 );
and  ( new_n709_, new_n708_, new_n662_ );
and  ( new_n710_, new_n450_, RI2af433cdb058_198 );
and  ( new_n711_, new_n710_, new_n691_ );
nor  ( new_n712_, new_n711_, new_n709_ );
and  ( new_n713_, new_n712_, new_n707_ );
and  ( new_n714_, new_n450_, RI2af433cdad88_192 );
and  ( new_n715_, new_n714_, new_n587_ );
and  ( new_n716_, new_n450_, RI2af433cdb0d0_199 );
and  ( new_n717_, new_n716_, new_n688_ );
nor  ( new_n718_, new_n717_, new_n715_ );
and  ( new_n719_, new_n482_, RI2af433cd77a0_77 );
and  ( new_n720_, new_n719_, new_n683_ );
and  ( new_n721_, new_n683_, RI2af433cd7818_78 );
and  ( new_n722_, new_n721_, new_n487_ );
nor  ( new_n723_, new_n722_, new_n720_ );
and  ( new_n724_, new_n723_, new_n718_ );
and  ( new_n725_, new_n724_, new_n713_ );
and  ( new_n726_, new_n725_, new_n701_ );
nor  ( new_n727_, new_n726_, new_n426_ );
and  ( new_n728_, new_n254_, RI2af433cd8b50_119 );
and  ( new_n729_, new_n277_, RI2af433cd8ad8_118 );
nor  ( new_n730_, new_n729_, new_n728_ );
and  ( new_n731_, new_n392_, RI2af433cd99d8_150 );
and  ( new_n732_, new_n388_, RI2af433cd9960_149 );
nor  ( new_n733_, new_n732_, new_n731_ );
and  ( new_n734_, new_n449_, RI2af433cd8c40_121 );
and  ( new_n735_, new_n474_, RI2af433cd9708_144 );
nor  ( new_n736_, new_n735_, new_n734_ );
and  ( new_n737_, new_n736_, new_n733_ );
and  ( new_n738_, new_n737_, new_n730_ );
nor  ( new_n739_, new_n738_, new_n431_ );
not  ( new_n740_, new_n739_ );
not  ( new_n741_, new_n683_ );
and  ( new_n742_, new_n495_, RI2af433cd7548_72 );
and  ( new_n743_, new_n484_, RI2af433cd7890_79 );
nor  ( new_n744_, new_n743_, new_n742_ );
nor  ( new_n745_, new_n744_, new_n741_ );
not  ( new_n746_, new_n745_ );
and  ( new_n747_, new_n683_, RI2af433cd75c0_73 );
and  ( new_n748_, new_n747_, new_n493_ );
and  ( new_n749_, new_n683_, RI2af433cd7638_74 );
and  ( new_n750_, new_n749_, new_n457_ );
nor  ( new_n751_, new_n750_, new_n748_ );
and  ( new_n752_, new_n751_, new_n746_ );
and  ( new_n753_, new_n752_, new_n740_ );
nor  ( new_n754_, new_n753_, new_n426_ );
nor  ( new_n755_, new_n754_, new_n727_ );
and  ( new_n756_, new_n755_, new_n675_ );
and  ( new_n757_, new_n662_, RI2af433cd73e0_69 );
and  ( new_n758_, new_n702_, RI2af433cd7368_68 );
nor  ( new_n759_, new_n758_, new_n757_ );
nor  ( new_n760_, new_n759_, new_n741_ );
not  ( new_n761_, new_n760_ );
and  ( new_n762_, new_n449_, RI2af433cd6e40_57 );
and  ( new_n763_, new_n476_, RI2af433cd6dc8_56 );
nor  ( new_n764_, new_n763_, new_n762_ );
nor  ( new_n765_, new_n764_, new_n741_ );
not  ( new_n766_, new_n765_ );
and  ( new_n767_, new_n766_, new_n761_ );
and  ( new_n768_, new_n468_, RI2af433cd7110_63 );
and  ( new_n769_, new_n553_, RI2af433cd7098_62 );
nor  ( new_n770_, new_n769_, new_n768_ );
nor  ( new_n771_, new_n770_, new_n741_ );
and  ( new_n772_, new_n606_, RI2af433cd6f30_59 );
and  ( new_n773_, new_n551_, RI2af433cd6eb8_58 );
nor  ( new_n774_, new_n773_, new_n772_ );
nor  ( new_n775_, new_n774_, new_n741_ );
nor  ( new_n776_, new_n775_, new_n771_ );
and  ( new_n777_, new_n776_, new_n767_ );
and  ( new_n778_, new_n474_, RI2af433cd7908_80 );
and  ( new_n779_, new_n460_, RI2af433cd76b0_75 );
nor  ( new_n780_, new_n779_, new_n778_ );
nor  ( new_n781_, new_n780_, new_n741_ );
and  ( new_n782_, new_n471_, RI2af433cd6fa8_60 );
and  ( new_n783_, new_n453_, RI2af433cd7020_61 );
nor  ( new_n784_, new_n783_, new_n782_ );
nor  ( new_n785_, new_n784_, new_n741_ );
nor  ( new_n786_, new_n785_, new_n781_ );
and  ( new_n787_, new_n238_, RI2af433cda590_175 );
and  ( new_n788_, new_n288_, RI2af433cda518_174 );
nor  ( new_n789_, new_n788_, new_n787_ );
and  ( new_n790_, new_n280_, RI2af433cda4a0_173 );
and  ( new_n791_, new_n263_, RI2af433cda428_172 );
nor  ( new_n792_, new_n791_, new_n790_ );
and  ( new_n793_, new_n792_, new_n789_ );
nor  ( new_n794_, new_n793_, new_n467_ );
and  ( new_n795_, new_n380_, RI2af433cd9870_147 );
and  ( new_n796_, new_n378_, RI2af433cd9780_145 );
nor  ( new_n797_, new_n796_, new_n795_ );
and  ( new_n798_, new_n397_, RI2af433cd97f8_146 );
and  ( new_n799_, new_n384_, RI2af433cd9a50_151 );
nor  ( new_n800_, new_n799_, new_n798_ );
and  ( new_n801_, new_n800_, new_n797_ );
nor  ( new_n802_, new_n801_, new_n431_ );
nor  ( new_n803_, new_n802_, new_n794_ );
and  ( new_n804_, new_n803_, new_n786_ );
and  ( new_n805_, new_n804_, new_n777_ );
nor  ( new_n806_, new_n805_, new_n426_ );
not  ( new_n807_, new_n806_ );
and  ( new_n808_, new_n450_, new_n425_ );
not  ( new_n809_, new_n808_ );
and  ( new_n810_, new_n318_, RI2af433cd9c30_155 );
and  ( new_n811_, new_n314_, RI2af433cd9bb8_154 );
nor  ( new_n812_, new_n811_, new_n810_ );
and  ( new_n813_, new_n321_, RI2af433cda1d0_167 );
and  ( new_n814_, new_n311_, RI2af433cda158_166 );
nor  ( new_n815_, new_n814_, new_n813_ );
and  ( new_n816_, new_n815_, new_n812_ );
and  ( new_n817_, new_n353_, RI2af433cd9ff0_163 );
and  ( new_n818_, new_n330_, RI2af433cd9f78_162 );
nor  ( new_n819_, new_n818_, new_n817_ );
and  ( new_n820_, new_n327_, RI2af433cd9f00_161 );
and  ( new_n821_, new_n337_, RI2af433cd9e88_160 );
nor  ( new_n822_, new_n821_, new_n820_ );
and  ( new_n823_, new_n822_, new_n819_ );
and  ( new_n824_, new_n823_, new_n816_ );
nor  ( new_n825_, new_n824_, new_n809_ );
not  ( new_n826_, new_n825_ );
and  ( new_n827_, new_n238_, RI2af433cd8790_111 );
and  ( new_n828_, new_n288_, RI2af433cd8718_110 );
nor  ( new_n829_, new_n828_, new_n827_ );
and  ( new_n830_, new_n232_, RI2af433cd85b0_107 );
and  ( new_n831_, new_n267_, RI2af433cd8538_106 );
nor  ( new_n832_, new_n831_, new_n830_ );
and  ( new_n833_, new_n832_, new_n829_ );
nor  ( new_n834_, new_n833_, new_n605_ );
not  ( new_n835_, new_n834_ );
and  ( new_n836_, new_n345_, RI2af433cda0e0_165 );
and  ( new_n837_, new_n334_, RI2af433cda068_164 );
nor  ( new_n838_, new_n837_, new_n836_ );
nor  ( new_n839_, new_n838_, new_n809_ );
and  ( new_n840_, new_n453_, RI2af433cd8e20_125 );
not  ( new_n841_, new_n840_ );
and  ( new_n842_, new_n702_, RI2af433cd9168_132 );
not  ( new_n843_, new_n842_ );
and  ( new_n844_, new_n843_, new_n841_ );
nor  ( new_n845_, new_n844_, new_n605_ );
nor  ( new_n846_, new_n845_, new_n839_ );
and  ( new_n847_, new_n846_, new_n835_ );
and  ( new_n848_, new_n847_, new_n826_ );
and  ( new_n849_, new_n353_, RI2af433cd81f0_99 );
and  ( new_n850_, new_n330_, RI2af433cd8178_98 );
nor  ( new_n851_, new_n850_, new_n849_ );
and  ( new_n852_, new_n303_, RI2af433cd7f20_93 );
not  ( new_n853_, new_n852_ );
and  ( new_n854_, new_n334_, RI2af433cd8268_100 );
not  ( new_n855_, new_n854_ );
and  ( new_n856_, new_n855_, new_n853_ );
and  ( new_n857_, new_n856_, new_n851_ );
and  ( new_n858_, new_n493_, RI2af433cd93c0_137 );
and  ( new_n859_, new_n337_, RI2af433cd8088_96 );
nor  ( new_n860_, new_n859_, new_n858_ );
and  ( new_n861_, new_n688_, RI2af433cd92d0_135 );
and  ( new_n862_, new_n691_, RI2af433cd9258_134 );
nor  ( new_n863_, new_n862_, new_n861_ );
and  ( new_n864_, new_n863_, new_n860_ );
and  ( new_n865_, new_n864_, new_n857_ );
nor  ( new_n866_, new_n865_, new_n605_ );
and  ( new_n867_, new_n460_, RI2af433cd94b0_139 );
and  ( new_n868_, new_n457_, RI2af433cd9438_138 );
nor  ( new_n869_, new_n868_, new_n867_ );
nor  ( new_n870_, new_n869_, new_n431_ );
and  ( new_n871_, new_n232_, RI2af433cda3b0_171 );
and  ( new_n872_, new_n267_, RI2af433cda338_170 );
nor  ( new_n873_, new_n872_, new_n871_ );
nor  ( new_n874_, new_n873_, new_n467_ );
nor  ( new_n875_, new_n874_, new_n870_ );
and  ( new_n876_, new_n683_, RI2af433cd72f0_67 );
and  ( new_n877_, new_n876_, new_n636_ );
and  ( new_n878_, new_n683_, RI2af433cd7278_66 );
and  ( new_n879_, new_n878_, new_n638_ );
nor  ( new_n880_, new_n879_, new_n877_ );
not  ( new_n881_, new_n880_ );
and  ( new_n882_, new_n368_, RI2af433cd9b40_153 );
and  ( new_n883_, new_n372_, RI2af433cd9ac8_152 );
nor  ( new_n884_, new_n883_, new_n882_ );
nor  ( new_n885_, new_n884_, new_n431_ );
nor  ( new_n886_, new_n885_, new_n881_ );
and  ( new_n887_, new_n886_, new_n875_ );
nor  ( new_n888_, new_n887_, new_n426_ );
nor  ( new_n889_, new_n888_, new_n866_ );
and  ( new_n890_, new_n889_, new_n848_ );
and  ( new_n891_, new_n890_, new_n807_ );
and  ( new_n892_, new_n891_, new_n756_ );
and  ( new_n893_, new_n892_, new_n563_ );
and  ( new_n894_, new_n893_, new_n427_ );
and  ( new_n895_, new_n803_, new_n439_ );
and  ( new_n896_, new_n895_, new_n500_ );
and  ( new_n897_, new_n880_, new_n766_ );
nor  ( new_n898_, new_n829_, new_n431_ );
and  ( new_n899_, new_n620_, RI2af433cd9ca8_156 );
nor  ( new_n900_, new_n899_, new_n898_ );
and  ( new_n901_, new_n900_, new_n897_ );
and  ( new_n902_, new_n694_, new_n686_ );
not  ( new_n903_, new_n874_ );
and  ( new_n904_, new_n903_, new_n699_ );
and  ( new_n905_, new_n904_, new_n902_ );
and  ( new_n906_, new_n905_, new_n901_ );
and  ( new_n907_, new_n624_, RI2af433cda2c0_169 );
not  ( new_n908_, new_n907_ );
and  ( new_n909_, new_n617_, RI2af433cd9d20_157 );
and  ( new_n910_, new_n627_, RI2af433cda248_168 );
nor  ( new_n911_, new_n910_, new_n909_ );
and  ( new_n912_, new_n911_, new_n908_ );
and  ( new_n913_, new_n912_, new_n786_ );
and  ( new_n914_, new_n913_, new_n906_ );
and  ( new_n915_, new_n914_, new_n896_ );
nor  ( new_n916_, new_n648_, new_n632_ );
and  ( new_n917_, new_n495_, RI2af433cd9348_136 );
nor  ( new_n918_, new_n917_, new_n633_ );
and  ( new_n919_, new_n918_, new_n916_ );
nor  ( new_n920_, new_n919_, new_n431_ );
not  ( new_n921_, new_n920_ );
nor  ( new_n922_, new_n840_, new_n610_ );
and  ( new_n923_, new_n654_, RI2af433cd9000_129 );
nor  ( new_n924_, new_n923_, new_n611_ );
and  ( new_n925_, new_n924_, new_n922_ );
nor  ( new_n926_, new_n925_, new_n431_ );
and  ( new_n927_, new_n838_, new_n819_ );
nor  ( new_n928_, new_n927_, new_n467_ );
nor  ( new_n929_, new_n928_, new_n926_ );
and  ( new_n930_, new_n929_, new_n921_ );
and  ( new_n931_, new_n884_, new_n730_ );
and  ( new_n932_, new_n931_, new_n737_ );
nor  ( new_n933_, new_n932_, new_n431_ );
and  ( new_n934_, new_n306_, RI2af433cd9d98_158 );
and  ( new_n935_, new_n342_, RI2af433cd9e10_159 );
nor  ( new_n936_, new_n935_, new_n934_ );
and  ( new_n937_, new_n936_, new_n812_ );
nor  ( new_n938_, new_n937_, new_n467_ );
nor  ( new_n939_, new_n938_, new_n933_ );
and  ( new_n940_, new_n587_, RI2af433cd8f88_128 );
not  ( new_n941_, new_n940_ );
and  ( new_n942_, new_n853_, new_n843_ );
and  ( new_n943_, new_n942_, new_n941_ );
nor  ( new_n944_, new_n943_, new_n431_ );
nor  ( new_n945_, new_n663_, new_n568_ );
and  ( new_n946_, new_n306_, RI2af433cd7f98_94 );
and  ( new_n947_, new_n342_, RI2af433cd8010_95 );
nor  ( new_n948_, new_n947_, new_n946_ );
and  ( new_n949_, new_n948_, new_n945_ );
nor  ( new_n950_, new_n949_, new_n431_ );
nor  ( new_n951_, new_n950_, new_n944_ );
and  ( new_n952_, new_n951_, new_n939_ );
and  ( new_n953_, new_n952_, new_n930_ );
and  ( new_n954_, new_n953_, new_n915_ );
and  ( new_n955_, new_n471_, RI2af433cd8da8_124 );
not  ( new_n956_, new_n955_ );
and  ( new_n957_, new_n956_, new_n860_ );
and  ( new_n958_, new_n863_, new_n609_ );
and  ( new_n959_, new_n958_, new_n957_ );
nor  ( new_n960_, new_n959_, new_n431_ );
not  ( new_n961_, new_n960_ );
and  ( new_n962_, new_n641_, new_n430_ );
nor  ( new_n963_, new_n815_, new_n467_ );
nor  ( new_n964_, new_n963_, new_n962_ );
nor  ( new_n965_, new_n850_, new_n574_ );
nor  ( new_n966_, new_n965_, new_n431_ );
nor  ( new_n967_, new_n854_, new_n849_ );
nor  ( new_n968_, new_n967_, new_n431_ );
nor  ( new_n969_, new_n968_, new_n966_ );
and  ( new_n970_, new_n969_, new_n964_ );
and  ( new_n971_, new_n970_, new_n532_ );
and  ( new_n972_, new_n971_, new_n961_ );
and  ( new_n973_, new_n761_, new_n746_ );
and  ( new_n974_, new_n973_, new_n465_ );
nor  ( new_n975_, new_n667_, new_n660_ );
nor  ( new_n976_, new_n652_, new_n646_ );
and  ( new_n977_, new_n976_, new_n975_ );
nor  ( new_n978_, new_n585_, new_n579_ );
and  ( new_n979_, new_n978_, new_n680_ );
and  ( new_n980_, new_n979_, new_n977_ );
and  ( new_n981_, new_n980_, new_n725_ );
and  ( new_n982_, new_n981_, new_n974_ );
and  ( new_n983_, new_n557_, new_n541_ );
and  ( new_n984_, new_n869_, new_n832_ );
nor  ( new_n985_, new_n984_, new_n431_ );
nor  ( new_n986_, new_n822_, new_n467_ );
nor  ( new_n987_, new_n986_, new_n985_ );
and  ( new_n988_, new_n987_, new_n983_ );
nor  ( new_n989_, new_n572_, new_n565_ );
and  ( new_n990_, new_n989_, new_n751_ );
and  ( new_n991_, new_n990_, new_n550_ );
and  ( new_n992_, new_n991_, new_n776_ );
and  ( new_n993_, new_n992_, new_n988_ );
and  ( new_n994_, new_n993_, new_n982_ );
and  ( new_n995_, new_n994_, new_n972_ );
and  ( new_n996_, new_n995_, new_n954_ );
and  ( new_n997_, new_n996_, new_n420_ );
or   ( new_n998_, new_n997_, new_n894_ );
nand ( new_n999_, new_n997_, new_n893_ );
or   ( new_n1000_, new_n283_, new_n221_ );
and  ( new_n1001_, new_n1000_, new_n367_ );
or   ( new_n1002_, new_n428_, new_n371_ );
or   ( new_n1003_, new_n1002_, new_n1001_ );
and  ( new_n1004_, new_n425_, new_n363_ );
and  ( new_n1005_, new_n1004_, new_n1003_ );
and  ( new_n1006_, new_n1005_, new_n999_ );
and  ( eq, new_n1006_, new_n998_ );
endmodule


