module miter ( 
    \a[15] , \a[14] , \a[13] , \a[12] , \a[11] , \a[10] , \a[9] , \a[8] ,
    \a[7] , \a[6] , \a[5] , \a[4] , \a[3] , \a[2] , \a[1] , \a[0] ,
    \b[15] , \b[14] , \b[13] , \b[12] , \b[11] , \b[10] , \b[9] , \b[8] ,
    \b[7] , \b[6] , \b[5] , \b[4] , \b[3] , \b[2] , \b[1] , \b[0] ,
    \c[15] , \c[14] , \c[13] , \c[12] , \c[11] , \c[10] , \c[9] , \c[8] ,
    \c[7] , \c[6] , \c[5] , \c[4] , \c[3] , \c[2] , \c[1] , \c[0] ,
    \d[15] , \d[14] , \d[13] , \d[12] , \d[11] , \d[10] , \d[9] , \d[8] ,
    \d[7] , \d[6] , \d[5] , \d[4] , \d[3] , \d[2] , \d[1] , \d[0] ,
    eq  );
  input  \a[15] , \a[14] , \a[13] , \a[12] , \a[11] , \a[10] , \a[9] ,
    \a[8] , \a[7] , \a[6] , \a[5] , \a[4] , \a[3] , \a[2] , \a[1] , \a[0] ,
    \b[15] , \b[14] , \b[13] , \b[12] , \b[11] , \b[10] , \b[9] , \b[8] ,
    \b[7] , \b[6] , \b[5] , \b[4] , \b[3] , \b[2] , \b[1] , \b[0] ,
    \c[15] , \c[14] , \c[13] , \c[12] , \c[11] , \c[10] , \c[9] , \c[8] ,
    \c[7] , \c[6] , \c[5] , \c[4] , \c[3] , \c[2] , \c[1] , \c[0] ,
    \d[15] , \d[14] , \d[13] , \d[12] , \d[11] , \d[10] , \d[9] , \d[8] ,
    \d[7] , \d[6] , \d[5] , \d[4] , \d[3] , \d[2] , \d[1] , \d[0] ;
  output eq;
  wire new_n66_, new_n67_, new_n68_, new_n69_, new_n70_, new_n71_, new_n72_,
    new_n73_, new_n74_, new_n75_, new_n76_, new_n77_, new_n78_, new_n79_,
    new_n80_, new_n81_, new_n82_, new_n83_, new_n84_, new_n85_, new_n86_,
    new_n87_, new_n88_, new_n89_, new_n90_, new_n91_, new_n92_, new_n93_,
    new_n94_, new_n95_, new_n96_, new_n97_, new_n98_, new_n99_, new_n100_,
    new_n101_, new_n102_, new_n103_, new_n104_, new_n105_, new_n106_,
    new_n107_, new_n108_, new_n109_, new_n110_, new_n111_, new_n112_,
    new_n113_, new_n114_, new_n115_, new_n116_, new_n117_, new_n118_,
    new_n119_, new_n120_, new_n121_, new_n122_, new_n123_, new_n124_,
    new_n125_, new_n126_, new_n127_, new_n128_, new_n129_, new_n130_,
    new_n131_, new_n132_, new_n133_, new_n134_, new_n135_, new_n136_,
    new_n137_, new_n138_, new_n139_, new_n140_, new_n141_, new_n142_,
    new_n143_, new_n144_, new_n145_, new_n146_, new_n147_, new_n148_,
    new_n149_, new_n150_, new_n151_, new_n152_, new_n153_, new_n154_,
    new_n155_, new_n156_, new_n157_, new_n158_, new_n159_, new_n160_,
    new_n161_, new_n162_, new_n163_, new_n164_, new_n165_, new_n166_,
    new_n167_, new_n168_, new_n169_, new_n170_, new_n171_, new_n172_,
    new_n173_, new_n174_, new_n175_, new_n176_, new_n177_, new_n178_,
    new_n179_, new_n180_, new_n181_, new_n182_, new_n183_, new_n184_,
    new_n185_, new_n186_, new_n187_, new_n188_, new_n189_, new_n190_,
    new_n191_, new_n192_, new_n193_, new_n194_, new_n195_, new_n196_,
    new_n197_, new_n198_, new_n199_, new_n200_, new_n201_, new_n202_,
    new_n203_, new_n204_, new_n205_, new_n206_, new_n207_, new_n208_,
    new_n209_, new_n210_, new_n211_, new_n212_, new_n213_, new_n214_,
    new_n215_, new_n216_, new_n217_, new_n218_, new_n219_, new_n220_,
    new_n221_, new_n222_, new_n223_, new_n224_, new_n225_, new_n226_,
    new_n227_, new_n228_, new_n229_, new_n230_, new_n231_, new_n232_,
    new_n233_, new_n234_, new_n235_, new_n236_, new_n237_, new_n238_,
    new_n239_, new_n240_, new_n241_, new_n242_, new_n243_, new_n244_,
    new_n245_, new_n246_, new_n247_, new_n248_, new_n249_, new_n250_,
    new_n251_, new_n252_, new_n253_, new_n254_, new_n255_, new_n256_,
    new_n257_, new_n258_, new_n259_, new_n260_, new_n261_, new_n262_,
    new_n263_, new_n264_, new_n265_, new_n266_, new_n267_, new_n268_,
    new_n269_, new_n270_, new_n271_, new_n272_, new_n273_, new_n274_,
    new_n275_, new_n276_, new_n277_, new_n278_, new_n279_, new_n280_,
    new_n281_, new_n282_, new_n283_, new_n284_, new_n285_, new_n286_,
    new_n287_, new_n288_, new_n289_, new_n290_, new_n291_, new_n292_,
    new_n293_, new_n294_, new_n295_, new_n296_, new_n297_, new_n298_,
    new_n299_, new_n300_, new_n301_, new_n302_, new_n303_, new_n304_,
    new_n305_, new_n306_, new_n307_, new_n308_, new_n309_, new_n310_,
    new_n311_, new_n312_, new_n313_, new_n314_, new_n315_, new_n316_,
    new_n317_, new_n318_, new_n319_, new_n320_, new_n321_, new_n322_,
    new_n323_, new_n324_, new_n325_, new_n326_, new_n327_, new_n328_,
    new_n329_, new_n330_, new_n331_, new_n332_, new_n333_, new_n334_,
    new_n335_, new_n336_, new_n337_, new_n338_, new_n339_, new_n340_,
    new_n341_, new_n342_, new_n343_, new_n344_, new_n345_, new_n346_,
    new_n347_, new_n348_, new_n349_, new_n350_, new_n351_, new_n352_,
    new_n353_, new_n354_, new_n355_, new_n356_, new_n357_, new_n358_,
    new_n359_, new_n360_, new_n361_, new_n362_, new_n363_, new_n364_,
    new_n365_, new_n366_, new_n367_, new_n368_, new_n369_, new_n370_,
    new_n371_, new_n372_, new_n373_, new_n374_, new_n375_, new_n376_,
    new_n377_, new_n378_, new_n379_, new_n380_, new_n381_, new_n382_,
    new_n383_, new_n384_, new_n385_, new_n386_, new_n387_, new_n388_,
    new_n389_, new_n390_, new_n391_, new_n392_, new_n393_, new_n394_,
    new_n395_, new_n396_, new_n397_, new_n398_, new_n399_, new_n400_,
    new_n401_, new_n402_, new_n403_, new_n404_, new_n405_, new_n406_,
    new_n407_, new_n408_, new_n409_, new_n410_, new_n411_, new_n412_,
    new_n413_, new_n414_, new_n415_, new_n416_, new_n417_, new_n418_,
    new_n419_, new_n420_, new_n421_, new_n422_, new_n423_, new_n424_,
    new_n425_, new_n426_, new_n427_, new_n428_, new_n429_, new_n430_,
    new_n431_, new_n432_, new_n433_, new_n434_, new_n435_, new_n436_,
    new_n437_, new_n438_, new_n439_, new_n440_, new_n441_, new_n442_,
    new_n443_, new_n444_, new_n445_, new_n446_, new_n447_, new_n448_,
    new_n449_, new_n450_, new_n451_, new_n452_, new_n453_, new_n454_,
    new_n455_, new_n456_, new_n457_, new_n458_, new_n459_, new_n460_,
    new_n461_, new_n462_, new_n463_, new_n464_, new_n465_, new_n466_,
    new_n467_, new_n468_, new_n469_, new_n470_, new_n471_, new_n472_,
    new_n473_, new_n474_, new_n475_, new_n476_, new_n477_, new_n478_,
    new_n479_, new_n480_, new_n481_, new_n482_, new_n483_, new_n484_,
    new_n485_, new_n486_, new_n487_, new_n488_, new_n489_, new_n490_,
    new_n491_, new_n492_, new_n493_, new_n494_, new_n495_, new_n496_,
    new_n497_, new_n498_, new_n499_, new_n500_, new_n501_, new_n502_,
    new_n503_, new_n504_, new_n505_, new_n506_, new_n507_, new_n508_,
    new_n509_, new_n510_, new_n511_, new_n512_, new_n513_, new_n514_,
    new_n515_, new_n516_, new_n517_, new_n518_, new_n519_, new_n520_,
    new_n521_, new_n522_, new_n523_, new_n524_, new_n525_, new_n526_,
    new_n527_, new_n528_, new_n529_, new_n530_, new_n531_, new_n532_,
    new_n533_, new_n534_, new_n535_, new_n536_, new_n537_, new_n538_,
    new_n539_, new_n540_, new_n541_, new_n542_, new_n543_, new_n544_,
    new_n545_, new_n546_, new_n547_, new_n548_, new_n549_, new_n550_,
    new_n551_, new_n552_, new_n553_, new_n554_, new_n555_, new_n556_,
    new_n557_, new_n558_, new_n559_, new_n560_, new_n561_, new_n562_,
    new_n563_, new_n564_, new_n565_, new_n566_, new_n567_, new_n568_,
    new_n569_, new_n570_, new_n571_, new_n572_, new_n573_, new_n574_,
    new_n575_, new_n576_, new_n577_, new_n578_, new_n579_, new_n580_,
    new_n581_, new_n582_, new_n583_, new_n584_, new_n585_, new_n586_,
    new_n587_, new_n588_, new_n589_, new_n590_, new_n591_, new_n592_,
    new_n593_, new_n594_, new_n595_, new_n596_, new_n597_, new_n598_,
    new_n599_, new_n600_, new_n601_, new_n602_, new_n603_, new_n604_,
    new_n605_, new_n606_, new_n607_, new_n608_, new_n609_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n691_, new_n692_, new_n693_, new_n694_,
    new_n695_, new_n696_, new_n697_, new_n698_, new_n699_, new_n700_,
    new_n701_, new_n702_, new_n703_, new_n704_, new_n705_, new_n706_,
    new_n707_, new_n708_, new_n709_, new_n710_, new_n711_, new_n712_,
    new_n713_, new_n714_, new_n715_, new_n716_, new_n717_, new_n718_,
    new_n719_, new_n720_, new_n721_, new_n722_, new_n723_, new_n724_,
    new_n725_, new_n726_, new_n727_, new_n728_, new_n729_, new_n730_,
    new_n731_, new_n732_, new_n733_, new_n734_, new_n735_, new_n736_,
    new_n737_, new_n738_, new_n739_, new_n740_, new_n741_, new_n742_,
    new_n743_, new_n744_, new_n745_, new_n746_, new_n747_, new_n748_,
    new_n749_, new_n750_, new_n751_, new_n752_, new_n753_, new_n754_,
    new_n755_, new_n756_, new_n757_, new_n758_, new_n759_, new_n760_,
    new_n761_, new_n762_, new_n763_, new_n764_, new_n765_, new_n766_,
    new_n767_, new_n768_, new_n769_, new_n770_, new_n771_, new_n772_,
    new_n773_, new_n774_, new_n775_, new_n776_, new_n777_, new_n778_,
    new_n779_, new_n780_, new_n781_, new_n782_, new_n783_, new_n784_,
    new_n785_, new_n786_, new_n787_, new_n788_, new_n789_, new_n790_,
    new_n791_, new_n792_, new_n793_, new_n794_, new_n795_, new_n796_,
    new_n797_, new_n798_, new_n799_, new_n800_, new_n801_, new_n802_,
    new_n803_, new_n804_, new_n805_, new_n806_, new_n807_, new_n808_,
    new_n809_, new_n810_, new_n811_, new_n812_, new_n813_, new_n814_,
    new_n815_, new_n816_, new_n817_, new_n818_, new_n819_, new_n820_,
    new_n821_, new_n822_, new_n823_, new_n824_, new_n825_, new_n826_,
    new_n827_, new_n828_, new_n829_, new_n830_, new_n831_, new_n832_,
    new_n833_, new_n834_, new_n835_, new_n836_, new_n837_, new_n838_,
    new_n839_, new_n840_, new_n841_, new_n842_, new_n843_, new_n844_,
    new_n845_, new_n846_, new_n847_, new_n848_, new_n849_, new_n850_,
    new_n851_, new_n852_, new_n853_, new_n854_, new_n855_, new_n856_,
    new_n857_, new_n858_, new_n859_, new_n860_, new_n861_, new_n862_,
    new_n863_, new_n864_, new_n865_, new_n866_, new_n867_, new_n868_,
    new_n869_, new_n870_, new_n871_, new_n872_, new_n873_, new_n874_,
    new_n875_, new_n876_, new_n877_, new_n878_, new_n879_, new_n880_,
    new_n881_, new_n882_, new_n883_, new_n884_, new_n885_, new_n886_,
    new_n887_, new_n888_, new_n889_, new_n890_, new_n891_, new_n892_,
    new_n893_, new_n894_, new_n895_, new_n896_, new_n897_, new_n898_,
    new_n899_, new_n900_, new_n901_, new_n902_, new_n903_, new_n904_,
    new_n905_, new_n906_, new_n907_, new_n908_, new_n909_, new_n910_,
    new_n911_, new_n912_, new_n913_, new_n914_, new_n915_, new_n916_,
    new_n917_, new_n918_, new_n919_, new_n920_, new_n921_, new_n922_,
    new_n923_, new_n924_, new_n925_, new_n926_, new_n927_, new_n928_,
    new_n929_, new_n930_, new_n931_, new_n932_, new_n933_, new_n934_,
    new_n935_, new_n936_, new_n937_, new_n938_, new_n939_, new_n940_,
    new_n941_, new_n942_, new_n943_, new_n944_, new_n945_, new_n946_,
    new_n947_, new_n948_, new_n949_, new_n950_, new_n951_, new_n952_,
    new_n953_, new_n954_, new_n955_, new_n956_, new_n957_, new_n958_,
    new_n959_, new_n960_, new_n961_, new_n962_, new_n963_, new_n964_,
    new_n965_, new_n966_, new_n967_, new_n968_, new_n969_, new_n970_,
    new_n971_, new_n972_, new_n973_, new_n974_, new_n975_, new_n976_,
    new_n977_, new_n978_, new_n979_, new_n980_, new_n981_, new_n982_,
    new_n983_, new_n984_, new_n985_, new_n986_, new_n987_, new_n988_,
    new_n989_, new_n990_, new_n991_, new_n992_, new_n993_, new_n994_,
    new_n995_, new_n996_, new_n997_, new_n998_, new_n999_, new_n1000_,
    new_n1001_, new_n1002_, new_n1003_, new_n1004_, new_n1005_, new_n1006_,
    new_n1007_, new_n1008_, new_n1009_, new_n1010_, new_n1011_, new_n1012_,
    new_n1013_, new_n1014_, new_n1015_, new_n1016_, new_n1017_, new_n1018_,
    new_n1019_, new_n1020_, new_n1021_, new_n1022_, new_n1023_, new_n1024_,
    new_n1025_, new_n1026_, new_n1027_, new_n1028_, new_n1029_, new_n1030_,
    new_n1031_, new_n1032_, new_n1033_, new_n1034_, new_n1035_, new_n1036_,
    new_n1037_, new_n1038_, new_n1039_, new_n1040_, new_n1041_, new_n1042_,
    new_n1043_, new_n1044_, new_n1045_, new_n1046_, new_n1047_, new_n1048_,
    new_n1049_, new_n1050_, new_n1051_, new_n1052_, new_n1053_, new_n1054_,
    new_n1055_, new_n1056_, new_n1057_, new_n1058_, new_n1059_, new_n1060_,
    new_n1061_, new_n1062_, new_n1063_, new_n1064_, new_n1065_, new_n1066_,
    new_n1067_, new_n1068_, new_n1069_, new_n1070_, new_n1071_, new_n1072_,
    new_n1073_, new_n1074_, new_n1075_, new_n1076_, new_n1077_, new_n1078_,
    new_n1079_, new_n1080_, new_n1081_, new_n1082_, new_n1083_, new_n1084_,
    new_n1085_, new_n1086_, new_n1087_, new_n1088_, new_n1089_, new_n1090_,
    new_n1091_, new_n1092_, new_n1093_, new_n1094_, new_n1095_, new_n1096_,
    new_n1097_, new_n1098_, new_n1099_, new_n1100_, new_n1101_, new_n1102_,
    new_n1103_, new_n1104_, new_n1105_, new_n1106_, new_n1107_, new_n1108_,
    new_n1109_, new_n1110_, new_n1111_, new_n1112_, new_n1113_, new_n1114_,
    new_n1115_, new_n1116_, new_n1117_, new_n1118_, new_n1119_, new_n1120_,
    new_n1121_, new_n1122_, new_n1123_, new_n1124_, new_n1125_, new_n1126_,
    new_n1127_, new_n1128_, new_n1129_, new_n1130_, new_n1131_, new_n1132_,
    new_n1133_, new_n1134_, new_n1135_, new_n1136_, new_n1137_, new_n1138_,
    new_n1139_, new_n1140_, new_n1141_, new_n1142_, new_n1143_, new_n1144_,
    new_n1145_, new_n1146_, new_n1147_, new_n1148_, new_n1149_, new_n1150_,
    new_n1151_, new_n1152_, new_n1153_, new_n1154_, new_n1155_, new_n1156_,
    new_n1157_, new_n1158_, new_n1159_, new_n1160_, new_n1161_, new_n1162_,
    new_n1163_, new_n1164_, new_n1165_, new_n1166_, new_n1167_, new_n1168_,
    new_n1169_, new_n1170_, new_n1171_, new_n1172_, new_n1173_, new_n1174_,
    new_n1175_, new_n1176_, new_n1177_, new_n1178_, new_n1179_, new_n1180_,
    new_n1181_, new_n1182_, new_n1183_, new_n1184_, new_n1185_, new_n1186_,
    new_n1187_, new_n1188_, new_n1189_, new_n1190_, new_n1191_, new_n1192_,
    new_n1193_, new_n1194_, new_n1195_, new_n1196_, new_n1197_, new_n1198_,
    new_n1199_, new_n1200_, new_n1201_, new_n1202_, new_n1203_, new_n1204_,
    new_n1205_, new_n1206_, new_n1207_, new_n1208_, new_n1209_, new_n1210_,
    new_n1211_, new_n1212_, new_n1213_, new_n1214_, new_n1215_, new_n1216_,
    new_n1217_, new_n1218_, new_n1219_, new_n1220_, new_n1221_, new_n1222_,
    new_n1223_, new_n1224_, new_n1225_, new_n1226_, new_n1227_, new_n1228_,
    new_n1229_, new_n1230_, new_n1231_, new_n1232_, new_n1233_, new_n1234_,
    new_n1235_, new_n1236_, new_n1237_, new_n1238_, new_n1239_, new_n1240_,
    new_n1241_, new_n1242_, new_n1243_, new_n1244_, new_n1245_, new_n1246_,
    new_n1247_, new_n1248_, new_n1249_, new_n1250_, new_n1251_, new_n1252_,
    new_n1253_, new_n1254_, new_n1255_, new_n1256_, new_n1257_, new_n1258_,
    new_n1259_, new_n1260_, new_n1261_, new_n1262_, new_n1263_, new_n1264_,
    new_n1265_, new_n1266_, new_n1267_, new_n1268_, new_n1269_, new_n1270_,
    new_n1271_, new_n1272_, new_n1273_, new_n1274_, new_n1275_, new_n1276_,
    new_n1277_, new_n1278_, new_n1279_, new_n1280_, new_n1281_, new_n1282_,
    new_n1283_, new_n1284_, new_n1285_, new_n1286_, new_n1287_, new_n1288_,
    new_n1289_, new_n1290_, new_n1291_, new_n1292_, new_n1293_, new_n1294_,
    new_n1295_, new_n1296_, new_n1297_, new_n1298_, new_n1299_, new_n1300_,
    new_n1301_, new_n1302_, new_n1303_, new_n1304_, new_n1305_, new_n1306_,
    new_n1307_, new_n1308_, new_n1309_, new_n1310_, new_n1311_, new_n1312_,
    new_n1313_, new_n1314_, new_n1315_, new_n1316_, new_n1317_, new_n1318_,
    new_n1319_, new_n1320_, new_n1321_, new_n1322_, new_n1323_, new_n1324_,
    new_n1325_, new_n1326_, new_n1327_, new_n1328_, new_n1329_, new_n1330_,
    new_n1331_, new_n1332_, new_n1333_, new_n1334_, new_n1335_, new_n1336_,
    new_n1337_, new_n1338_, new_n1339_, new_n1340_, new_n1341_, new_n1342_,
    new_n1343_, new_n1344_, new_n1345_, new_n1346_, new_n1347_, new_n1348_,
    new_n1349_, new_n1350_, new_n1351_, new_n1352_, new_n1353_, new_n1354_,
    new_n1355_, new_n1356_, new_n1357_, new_n1358_, new_n1359_, new_n1360_,
    new_n1361_, new_n1362_, new_n1363_, new_n1364_, new_n1365_, new_n1366_,
    new_n1367_, new_n1368_, new_n1369_, new_n1370_, new_n1371_, new_n1372_,
    new_n1373_, new_n1374_, new_n1375_, new_n1376_, new_n1377_, new_n1378_,
    new_n1379_, new_n1380_, new_n1381_, new_n1382_, new_n1383_, new_n1384_,
    new_n1385_, new_n1386_, new_n1387_, new_n1388_, new_n1389_, new_n1390_,
    new_n1391_, new_n1392_, new_n1393_, new_n1394_, new_n1395_, new_n1396_,
    new_n1397_, new_n1398_, new_n1399_, new_n1400_, new_n1401_, new_n1402_,
    new_n1403_, new_n1404_, new_n1405_, new_n1406_, new_n1407_, new_n1408_,
    new_n1409_, new_n1410_, new_n1411_, new_n1412_, new_n1413_, new_n1414_,
    new_n1415_, new_n1416_, new_n1417_, new_n1418_, new_n1419_, new_n1420_,
    new_n1421_, new_n1422_, new_n1423_, new_n1424_, new_n1425_, new_n1426_,
    new_n1427_, new_n1428_, new_n1429_, new_n1430_, new_n1431_, new_n1432_,
    new_n1433_, new_n1434_, new_n1435_, new_n1436_, new_n1437_, new_n1438_,
    new_n1439_, new_n1440_, new_n1441_, new_n1442_, new_n1443_, new_n1444_,
    new_n1445_, new_n1446_, new_n1447_, new_n1448_, new_n1449_, new_n1450_,
    new_n1451_, new_n1452_, new_n1453_, new_n1454_, new_n1455_, new_n1456_,
    new_n1457_, new_n1458_, new_n1459_, new_n1460_, new_n1461_, new_n1462_,
    new_n1463_, new_n1464_, new_n1465_, new_n1466_, new_n1467_, new_n1468_,
    new_n1469_, new_n1470_, new_n1471_, new_n1472_, new_n1473_, new_n1474_,
    new_n1475_, new_n1476_, new_n1477_, new_n1478_, new_n1479_, new_n1480_,
    new_n1481_, new_n1482_, new_n1483_, new_n1484_, new_n1485_, new_n1486_,
    new_n1487_, new_n1488_, new_n1489_, new_n1490_, new_n1491_, new_n1492_,
    new_n1493_, new_n1494_, new_n1495_, new_n1496_, new_n1497_, new_n1498_,
    new_n1499_, new_n1500_, new_n1501_, new_n1502_, new_n1503_, new_n1504_,
    new_n1505_, new_n1506_, new_n1507_, new_n1508_, new_n1509_, new_n1510_,
    new_n1511_, new_n1512_, new_n1513_, new_n1514_, new_n1515_, new_n1516_,
    new_n1517_, new_n1518_, new_n1519_, new_n1520_, new_n1521_, new_n1522_,
    new_n1523_, new_n1524_, new_n1525_, new_n1526_, new_n1527_, new_n1528_,
    new_n1529_, new_n1530_, new_n1531_, new_n1532_, new_n1533_, new_n1534_,
    new_n1535_, new_n1536_, new_n1537_, new_n1538_, new_n1539_, new_n1540_,
    new_n1541_, new_n1542_, new_n1543_, new_n1544_, new_n1545_, new_n1546_,
    new_n1547_, new_n1548_, new_n1549_, new_n1550_, new_n1551_, new_n1552_,
    new_n1553_, new_n1554_, new_n1555_, new_n1556_, new_n1557_, new_n1558_,
    new_n1559_, new_n1560_, new_n1561_, new_n1562_, new_n1563_, new_n1564_,
    new_n1565_, new_n1566_, new_n1567_, new_n1568_, new_n1569_, new_n1570_,
    new_n1571_, new_n1572_, new_n1573_, new_n1574_, new_n1575_, new_n1576_,
    new_n1577_, new_n1578_, new_n1579_, new_n1580_, new_n1581_, new_n1582_,
    new_n1583_, new_n1584_, new_n1585_, new_n1586_, new_n1587_, new_n1588_,
    new_n1589_, new_n1590_, new_n1591_, new_n1592_, new_n1593_, new_n1594_,
    new_n1595_, new_n1596_, new_n1597_, new_n1598_, new_n1599_, new_n1600_,
    new_n1601_, new_n1602_, new_n1603_, new_n1604_, new_n1605_, new_n1606_,
    new_n1607_, new_n1608_, new_n1609_, new_n1610_, new_n1611_, new_n1612_,
    new_n1613_, new_n1614_, new_n1615_, new_n1616_, new_n1617_, new_n1618_,
    new_n1619_, new_n1620_, new_n1621_, new_n1622_, new_n1623_, new_n1624_,
    new_n1625_, new_n1626_, new_n1627_, new_n1628_, new_n1629_, new_n1630_,
    new_n1631_, new_n1632_, new_n1633_, new_n1634_, new_n1635_, new_n1636_,
    new_n1637_, new_n1638_, new_n1639_, new_n1640_, new_n1641_, new_n1642_,
    new_n1643_, new_n1644_, new_n1645_, new_n1646_, new_n1647_, new_n1648_,
    new_n1649_, new_n1650_, new_n1651_, new_n1652_, new_n1653_, new_n1654_,
    new_n1655_, new_n1656_, new_n1657_, new_n1658_, new_n1659_, new_n1660_,
    new_n1661_, new_n1662_, new_n1663_, new_n1664_, new_n1665_, new_n1666_,
    new_n1667_, new_n1668_, new_n1669_, new_n1670_, new_n1671_, new_n1672_,
    new_n1673_, new_n1674_, new_n1675_, new_n1676_, new_n1677_, new_n1678_,
    new_n1679_, new_n1680_, new_n1681_, new_n1682_, new_n1683_, new_n1684_,
    new_n1685_, new_n1686_, new_n1687_, new_n1688_, new_n1689_, new_n1690_,
    new_n1691_, new_n1692_, new_n1693_, new_n1694_, new_n1695_, new_n1696_,
    new_n1697_, new_n1698_, new_n1699_, new_n1700_, new_n1701_, new_n1702_,
    new_n1703_, new_n1704_, new_n1705_, new_n1706_, new_n1707_, new_n1708_,
    new_n1709_, new_n1710_, new_n1711_, new_n1712_, new_n1713_, new_n1714_,
    new_n1715_, new_n1716_, new_n1717_, new_n1718_, new_n1719_, new_n1720_,
    new_n1721_, new_n1722_, new_n1723_, new_n1724_, new_n1725_, new_n1726_,
    new_n1727_, new_n1728_, new_n1729_, new_n1730_, new_n1731_, new_n1732_,
    new_n1733_, new_n1734_, new_n1735_, new_n1736_, new_n1737_, new_n1738_,
    new_n1739_, new_n1740_, new_n1741_, new_n1742_, new_n1743_, new_n1744_,
    new_n1745_, new_n1746_, new_n1747_, new_n1748_, new_n1749_, new_n1750_,
    new_n1751_, new_n1752_, new_n1753_, new_n1754_, new_n1755_, new_n1756_,
    new_n1757_, new_n1758_, new_n1759_, new_n1760_, new_n1761_, new_n1762_,
    new_n1763_, new_n1764_, new_n1765_, new_n1766_, new_n1767_, new_n1768_,
    new_n1769_, new_n1770_, new_n1771_, new_n1772_, new_n1773_, new_n1774_,
    new_n1775_, new_n1776_, new_n1777_, new_n1778_, new_n1779_, new_n1780_,
    new_n1781_, new_n1782_, new_n1783_, new_n1784_, new_n1785_, new_n1786_,
    new_n1787_, new_n1788_, new_n1789_, new_n1790_, new_n1791_, new_n1792_,
    new_n1793_, new_n1794_, new_n1795_, new_n1796_, new_n1797_, new_n1798_,
    new_n1799_, new_n1800_, new_n1801_, new_n1802_, new_n1803_, new_n1804_,
    new_n1805_, new_n1806_, new_n1807_, new_n1808_, new_n1809_, new_n1810_,
    new_n1811_, new_n1812_, new_n1813_, new_n1814_, new_n1815_, new_n1816_,
    new_n1817_, new_n1818_, new_n1819_, new_n1820_, new_n1821_, new_n1822_,
    new_n1823_, new_n1824_, new_n1825_, new_n1826_, new_n1827_, new_n1828_,
    new_n1829_, new_n1830_, new_n1831_, new_n1832_, new_n1833_, new_n1834_,
    new_n1835_, new_n1836_, new_n1837_, new_n1838_, new_n1839_, new_n1840_,
    new_n1841_, new_n1842_, new_n1843_, new_n1844_, new_n1845_, new_n1846_,
    new_n1847_, new_n1848_, new_n1849_, new_n1850_, new_n1851_, new_n1852_,
    new_n1853_, new_n1854_, new_n1855_, new_n1856_, new_n1857_, new_n1858_,
    new_n1859_, new_n1860_, new_n1861_, new_n1862_, new_n1863_, new_n1864_,
    new_n1865_, new_n1866_, new_n1867_, new_n1868_, new_n1869_, new_n1870_,
    new_n1871_, new_n1872_, new_n1873_, new_n1874_, new_n1875_, new_n1876_,
    new_n1877_, new_n1878_, new_n1879_, new_n1880_, new_n1881_, new_n1882_,
    new_n1883_, new_n1884_, new_n1885_, new_n1886_, new_n1887_, new_n1888_,
    new_n1889_, new_n1890_, new_n1891_, new_n1892_, new_n1893_, new_n1894_,
    new_n1895_, new_n1896_, new_n1897_, new_n1898_, new_n1899_, new_n1900_,
    new_n1901_, new_n1902_, new_n1903_, new_n1904_, new_n1905_, new_n1906_,
    new_n1907_, new_n1908_, new_n1909_, new_n1910_, new_n1911_, new_n1912_,
    new_n1913_, new_n1914_, new_n1915_, new_n1916_, new_n1917_, new_n1918_,
    new_n1919_, new_n1920_, new_n1921_, new_n1922_, new_n1923_, new_n1924_,
    new_n1925_, new_n1926_, new_n1927_, new_n1928_, new_n1929_, new_n1930_,
    new_n1931_, new_n1932_, new_n1933_, new_n1934_, new_n1935_, new_n1936_,
    new_n1937_, new_n1938_, new_n1939_, new_n1940_, new_n1941_, new_n1942_,
    new_n1943_, new_n1944_, new_n1945_, new_n1946_, new_n1947_, new_n1948_,
    new_n1949_, new_n1950_, new_n1951_, new_n1952_, new_n1953_, new_n1954_,
    new_n1955_, new_n1956_, new_n1957_, new_n1958_, new_n1959_, new_n1960_,
    new_n1961_, new_n1962_, new_n1963_, new_n1964_, new_n1965_, new_n1966_,
    new_n1967_, new_n1968_, new_n1969_, new_n1970_, new_n1971_, new_n1972_,
    new_n1973_, new_n1974_, new_n1975_, new_n1976_, new_n1977_, new_n1978_,
    new_n1979_, new_n1980_, new_n1981_, new_n1982_, new_n1983_, new_n1984_,
    new_n1985_, new_n1986_, new_n1987_, new_n1988_, new_n1989_, new_n1990_,
    new_n1991_, new_n1992_, new_n1993_, new_n1994_, new_n1995_, new_n1996_,
    new_n1997_, new_n1998_, new_n1999_, new_n2000_, new_n2001_, new_n2002_,
    new_n2003_, new_n2004_, new_n2005_, new_n2006_, new_n2007_, new_n2008_,
    new_n2009_, new_n2010_, new_n2011_, new_n2012_, new_n2013_, new_n2014_,
    new_n2015_, new_n2016_, new_n2017_, new_n2018_, new_n2019_, new_n2020_,
    new_n2021_, new_n2022_, new_n2023_, new_n2024_, new_n2025_, new_n2026_,
    new_n2027_, new_n2028_, new_n2029_, new_n2030_, new_n2031_, new_n2032_,
    new_n2033_, new_n2034_, new_n2035_, new_n2036_, new_n2037_, new_n2038_,
    new_n2039_, new_n2040_, new_n2041_, new_n2042_, new_n2043_, new_n2044_,
    new_n2045_, new_n2046_, new_n2047_, new_n2048_, new_n2049_, new_n2050_,
    new_n2051_, new_n2052_, new_n2053_, new_n2054_, new_n2055_, new_n2056_,
    new_n2057_, new_n2058_, new_n2059_, new_n2060_, new_n2061_, new_n2062_,
    new_n2063_, new_n2064_, new_n2065_, new_n2066_, new_n2067_, new_n2068_,
    new_n2069_, new_n2070_, new_n2071_, new_n2072_, new_n2073_, new_n2074_,
    new_n2075_, new_n2076_, new_n2077_, new_n2078_, new_n2079_, new_n2080_,
    new_n2081_, new_n2082_, new_n2083_, new_n2084_, new_n2085_, new_n2086_,
    new_n2087_, new_n2088_, new_n2089_, new_n2090_, new_n2091_, new_n2092_,
    new_n2093_, new_n2094_, new_n2095_, new_n2096_, new_n2097_, new_n2098_,
    new_n2099_, new_n2100_, new_n2101_, new_n2102_, new_n2103_, new_n2104_,
    new_n2105_, new_n2106_, new_n2107_, new_n2108_, new_n2109_, new_n2110_,
    new_n2111_, new_n2112_, new_n2113_, new_n2114_, new_n2115_, new_n2116_,
    new_n2117_, new_n2118_, new_n2119_, new_n2120_, new_n2121_, new_n2122_,
    new_n2123_, new_n2124_, new_n2125_, new_n2126_, new_n2127_, new_n2128_,
    new_n2129_, new_n2130_, new_n2131_, new_n2132_, new_n2133_, new_n2134_,
    new_n2135_, new_n2136_, new_n2137_, new_n2138_, new_n2139_, new_n2140_,
    new_n2141_, new_n2142_, new_n2143_, new_n2144_, new_n2145_, new_n2146_,
    new_n2147_, new_n2148_, new_n2149_, new_n2150_, new_n2151_, new_n2152_,
    new_n2153_, new_n2154_, new_n2155_, new_n2156_, new_n2157_, new_n2158_,
    new_n2159_, new_n2160_, new_n2161_, new_n2162_, new_n2163_, new_n2164_,
    new_n2165_, new_n2166_, new_n2167_, new_n2168_, new_n2169_, new_n2170_,
    new_n2171_, new_n2172_, new_n2173_, new_n2174_, new_n2175_, new_n2176_,
    new_n2177_, new_n2178_, new_n2179_, new_n2180_, new_n2181_, new_n2182_,
    new_n2183_, new_n2184_, new_n2185_, new_n2186_, new_n2187_, new_n2188_,
    new_n2189_, new_n2190_, new_n2191_, new_n2192_, new_n2193_, new_n2194_,
    new_n2195_, new_n2196_, new_n2197_, new_n2198_, new_n2199_, new_n2200_,
    new_n2201_, new_n2202_, new_n2203_, new_n2204_, new_n2205_, new_n2206_,
    new_n2207_, new_n2208_, new_n2209_, new_n2210_, new_n2211_, new_n2212_,
    new_n2213_, new_n2214_, new_n2215_, new_n2216_, new_n2217_, new_n2218_,
    new_n2219_, new_n2220_, new_n2221_, new_n2222_, new_n2223_, new_n2224_,
    new_n2225_, new_n2226_, new_n2227_, new_n2228_, new_n2229_, new_n2230_,
    new_n2231_, new_n2232_, new_n2233_, new_n2234_, new_n2235_, new_n2236_,
    new_n2237_, new_n2238_, new_n2239_, new_n2240_, new_n2241_, new_n2242_,
    new_n2243_, new_n2244_, new_n2245_, new_n2246_, new_n2247_, new_n2248_,
    new_n2249_, new_n2250_, new_n2251_, new_n2252_, new_n2253_, new_n2254_,
    new_n2255_, new_n2256_, new_n2257_, new_n2258_, new_n2259_, new_n2260_,
    new_n2261_, new_n2262_, new_n2263_, new_n2264_, new_n2265_, new_n2266_,
    new_n2267_, new_n2268_, new_n2269_, new_n2270_, new_n2271_, new_n2272_,
    new_n2273_, new_n2274_, new_n2275_, new_n2276_, new_n2277_, new_n2278_,
    new_n2279_, new_n2280_, new_n2281_, new_n2282_, new_n2283_, new_n2284_,
    new_n2285_, new_n2286_, new_n2287_, new_n2288_, new_n2289_, new_n2290_,
    new_n2291_, new_n2292_, new_n2293_, new_n2294_, new_n2295_, new_n2296_,
    new_n2297_, new_n2298_, new_n2299_, new_n2300_, new_n2301_, new_n2302_,
    new_n2303_, new_n2304_, new_n2305_, new_n2306_, new_n2307_, new_n2308_,
    new_n2309_, new_n2310_, new_n2311_, new_n2312_, new_n2313_, new_n2314_,
    new_n2315_, new_n2316_, new_n2317_, new_n2318_, new_n2319_, new_n2320_,
    new_n2321_, new_n2322_, new_n2323_, new_n2324_, new_n2325_, new_n2326_,
    new_n2327_, new_n2328_, new_n2329_, new_n2330_, new_n2331_, new_n2332_,
    new_n2333_, new_n2334_, new_n2335_, new_n2336_, new_n2337_, new_n2338_,
    new_n2339_, new_n2340_, new_n2341_, new_n2342_, new_n2343_, new_n2344_,
    new_n2345_, new_n2346_, new_n2347_, new_n2348_, new_n2349_, new_n2350_,
    new_n2351_, new_n2352_, new_n2353_, new_n2354_, new_n2355_, new_n2356_,
    new_n2357_, new_n2358_, new_n2359_, new_n2360_, new_n2361_, new_n2362_,
    new_n2363_, new_n2364_, new_n2365_, new_n2366_, new_n2367_, new_n2368_,
    new_n2369_, new_n2370_, new_n2371_, new_n2372_, new_n2373_, new_n2374_,
    new_n2375_, new_n2376_, new_n2377_, new_n2378_, new_n2379_, new_n2380_,
    new_n2381_, new_n2382_, new_n2383_, new_n2384_, new_n2385_, new_n2386_,
    new_n2387_, new_n2388_, new_n2389_, new_n2390_, new_n2391_, new_n2392_,
    new_n2393_, new_n2394_, new_n2395_, new_n2396_, new_n2397_, new_n2398_,
    new_n2399_, new_n2400_, new_n2401_, new_n2402_, new_n2403_, new_n2404_,
    new_n2405_, new_n2406_, new_n2407_, new_n2408_, new_n2409_, new_n2410_,
    new_n2411_, new_n2412_, new_n2413_, new_n2414_, new_n2415_, new_n2416_,
    new_n2417_, new_n2418_, new_n2419_, new_n2420_, new_n2421_, new_n2422_,
    new_n2423_, new_n2424_, new_n2425_, new_n2426_, new_n2427_, new_n2428_,
    new_n2429_, new_n2430_, new_n2431_, new_n2432_, new_n2433_, new_n2434_,
    new_n2435_, new_n2436_, new_n2437_, new_n2438_, new_n2439_, new_n2440_,
    new_n2441_, new_n2442_, new_n2443_, new_n2444_, new_n2445_, new_n2446_,
    new_n2447_, new_n2448_, new_n2449_, new_n2450_, new_n2451_, new_n2452_,
    new_n2453_, new_n2454_, new_n2455_, new_n2456_, new_n2457_, new_n2458_,
    new_n2459_, new_n2460_, new_n2461_, new_n2462_, new_n2463_, new_n2464_,
    new_n2465_, new_n2466_, new_n2467_, new_n2468_, new_n2469_, new_n2470_,
    new_n2471_, new_n2472_, new_n2473_, new_n2474_, new_n2475_, new_n2476_,
    new_n2477_, new_n2478_, new_n2479_, new_n2480_, new_n2481_, new_n2482_,
    new_n2483_, new_n2484_, new_n2485_, new_n2486_, new_n2487_, new_n2488_,
    new_n2489_, new_n2490_, new_n2491_, new_n2492_, new_n2493_, new_n2494_,
    new_n2495_, new_n2496_, new_n2497_, new_n2498_, new_n2499_, new_n2500_,
    new_n2501_, new_n2502_, new_n2503_, new_n2504_, new_n2505_, new_n2506_,
    new_n2507_, new_n2508_, new_n2509_, new_n2510_, new_n2511_, new_n2512_,
    new_n2513_, new_n2514_, new_n2515_, new_n2516_, new_n2517_, new_n2518_,
    new_n2519_, new_n2520_, new_n2521_, new_n2522_, new_n2523_, new_n2524_,
    new_n2525_, new_n2526_, new_n2527_, new_n2528_, new_n2529_, new_n2530_,
    new_n2531_, new_n2532_, new_n2533_, new_n2534_, new_n2535_, new_n2536_,
    new_n2537_, new_n2538_, new_n2539_, new_n2540_, new_n2541_, new_n2542_,
    new_n2543_, new_n2544_, new_n2545_, new_n2546_, new_n2547_, new_n2548_,
    new_n2549_, new_n2550_, new_n2551_, new_n2552_, new_n2553_, new_n2554_,
    new_n2555_, new_n2556_, new_n2557_, new_n2558_, new_n2559_, new_n2560_,
    new_n2561_, new_n2562_, new_n2563_, new_n2564_, new_n2565_, new_n2566_,
    new_n2567_, new_n2568_, new_n2569_, new_n2570_, new_n2571_, new_n2572_,
    new_n2573_, new_n2574_, new_n2575_, new_n2576_, new_n2577_, new_n2578_,
    new_n2579_, new_n2580_, new_n2581_, new_n2582_, new_n2583_, new_n2584_,
    new_n2585_, new_n2586_, new_n2587_, new_n2588_, new_n2589_, new_n2590_,
    new_n2591_, new_n2592_, new_n2593_, new_n2594_, new_n2595_, new_n2596_,
    new_n2597_, new_n2598_, new_n2599_, new_n2600_, new_n2601_, new_n2602_,
    new_n2603_, new_n2604_, new_n2605_, new_n2606_, new_n2607_, new_n2608_,
    new_n2609_, new_n2610_, new_n2611_, new_n2612_, new_n2613_, new_n2614_,
    new_n2615_, new_n2616_, new_n2617_, new_n2618_, new_n2619_, new_n2620_,
    new_n2621_, new_n2622_, new_n2623_, new_n2624_, new_n2625_, new_n2626_,
    new_n2627_, new_n2628_, new_n2629_, new_n2630_, new_n2631_, new_n2632_,
    new_n2633_, new_n2634_, new_n2635_, new_n2636_, new_n2637_, new_n2638_,
    new_n2639_, new_n2640_, new_n2641_, new_n2642_, new_n2643_, new_n2644_,
    new_n2645_, new_n2646_, new_n2647_, new_n2648_, new_n2649_, new_n2650_,
    new_n2651_, new_n2652_, new_n2653_, new_n2654_, new_n2655_, new_n2656_,
    new_n2657_, new_n2658_, new_n2659_, new_n2660_, new_n2661_, new_n2662_,
    new_n2663_, new_n2664_, new_n2665_, new_n2666_, new_n2667_, new_n2668_,
    new_n2669_, new_n2670_, new_n2671_, new_n2672_, new_n2673_, new_n2674_,
    new_n2675_, new_n2676_, new_n2677_, new_n2678_, new_n2679_, new_n2680_,
    new_n2681_, new_n2682_, new_n2683_, new_n2684_, new_n2685_, new_n2686_,
    new_n2687_, new_n2688_, new_n2689_, new_n2690_, new_n2691_, new_n2692_,
    new_n2693_, new_n2694_, new_n2695_, new_n2696_, new_n2697_, new_n2698_,
    new_n2699_, new_n2700_, new_n2701_, new_n2702_, new_n2703_, new_n2704_,
    new_n2705_, new_n2706_, new_n2707_, new_n2708_, new_n2709_, new_n2710_,
    new_n2711_, new_n2712_, new_n2713_, new_n2714_, new_n2715_, new_n2716_,
    new_n2717_, new_n2718_, new_n2719_, new_n2720_, new_n2721_, new_n2722_,
    new_n2723_, new_n2724_, new_n2725_, new_n2726_, new_n2727_, new_n2728_,
    new_n2729_, new_n2730_, new_n2731_, new_n2732_, new_n2733_, new_n2734_,
    new_n2735_, new_n2736_, new_n2737_, new_n2738_, new_n2739_, new_n2740_,
    new_n2741_, new_n2742_, new_n2743_, new_n2744_, new_n2745_, new_n2746_,
    new_n2747_, new_n2748_, new_n2749_, new_n2750_, new_n2751_, new_n2752_,
    new_n2753_, new_n2754_, new_n2755_, new_n2756_, new_n2757_, new_n2758_,
    new_n2759_, new_n2760_, new_n2761_, new_n2762_, new_n2763_, new_n2764_,
    new_n2765_, new_n2766_, new_n2767_, new_n2768_, new_n2769_, new_n2770_,
    new_n2771_, new_n2772_, new_n2773_, new_n2774_, new_n2775_, new_n2776_,
    new_n2777_, new_n2778_, new_n2779_, new_n2780_, new_n2781_, new_n2782_,
    new_n2783_, new_n2784_, new_n2785_, new_n2786_, new_n2787_, new_n2788_,
    new_n2789_, new_n2790_, new_n2791_, new_n2792_, new_n2793_, new_n2794_,
    new_n2795_, new_n2796_, new_n2797_, new_n2798_, new_n2799_, new_n2800_,
    new_n2801_, new_n2802_, new_n2803_, new_n2804_, new_n2805_, new_n2806_,
    new_n2807_, new_n2808_, new_n2809_, new_n2810_, new_n2811_, new_n2812_,
    new_n2813_, new_n2814_, new_n2815_, new_n2816_, new_n2817_, new_n2818_,
    new_n2819_, new_n2820_, new_n2821_, new_n2822_, new_n2823_, new_n2824_,
    new_n2825_, new_n2826_, new_n2827_, new_n2828_, new_n2829_, new_n2830_,
    new_n2831_, new_n2832_, new_n2833_, new_n2834_, new_n2835_, new_n2836_,
    new_n2837_, new_n2838_, new_n2839_, new_n2840_, new_n2841_, new_n2842_,
    new_n2843_, new_n2844_, new_n2845_, new_n2846_, new_n2847_, new_n2848_,
    new_n2849_, new_n2850_, new_n2851_, new_n2852_, new_n2853_, new_n2854_,
    new_n2855_, new_n2856_, new_n2857_, new_n2858_, new_n2859_, new_n2860_,
    new_n2861_, new_n2862_, new_n2863_, new_n2864_, new_n2865_, new_n2866_,
    new_n2867_, new_n2868_, new_n2869_, new_n2870_, new_n2871_, new_n2872_,
    new_n2873_, new_n2874_, new_n2875_, new_n2876_, new_n2877_, new_n2878_,
    new_n2879_, new_n2880_, new_n2881_, new_n2882_, new_n2883_, new_n2884_,
    new_n2885_, new_n2886_, new_n2887_, new_n2888_, new_n2889_, new_n2890_,
    new_n2891_, new_n2892_, new_n2893_, new_n2894_, new_n2895_, new_n2896_,
    new_n2897_, new_n2898_, new_n2899_, new_n2900_, new_n2901_, new_n2902_,
    new_n2903_, new_n2904_, new_n2905_, new_n2906_, new_n2907_, new_n2908_,
    new_n2909_, new_n2910_, new_n2911_, new_n2912_, new_n2913_, new_n2914_,
    new_n2915_, new_n2916_, new_n2917_, new_n2918_, new_n2919_, new_n2920_,
    new_n2921_, new_n2922_, new_n2923_, new_n2924_, new_n2925_, new_n2926_,
    new_n2927_, new_n2928_, new_n2929_, new_n2930_, new_n2931_, new_n2932_,
    new_n2933_, new_n2934_, new_n2935_, new_n2936_, new_n2937_, new_n2938_,
    new_n2939_, new_n2940_, new_n2941_, new_n2942_, new_n2943_, new_n2944_,
    new_n2945_, new_n2946_, new_n2947_, new_n2948_, new_n2949_, new_n2950_,
    new_n2951_, new_n2952_, new_n2953_, new_n2954_, new_n2955_, new_n2956_,
    new_n2957_, new_n2958_, new_n2959_, new_n2960_, new_n2961_, new_n2962_,
    new_n2963_, new_n2964_, new_n2965_, new_n2966_, new_n2967_, new_n2968_,
    new_n2969_, new_n2970_, new_n2971_, new_n2972_, new_n2973_, new_n2974_,
    new_n2975_, new_n2976_, new_n2977_, new_n2978_, new_n2979_, new_n2980_,
    new_n2981_, new_n2982_, new_n2983_, new_n2984_, new_n2985_, new_n2986_,
    new_n2987_, new_n2988_, new_n2989_, new_n2990_, new_n2991_, new_n2992_,
    new_n2993_, new_n2994_, new_n2995_, new_n2996_, new_n2997_, new_n2998_,
    new_n2999_, new_n3000_, new_n3001_, new_n3002_, new_n3003_, new_n3004_,
    new_n3005_, new_n3006_, new_n3007_, new_n3008_, new_n3009_, new_n3010_,
    new_n3011_, new_n3012_, new_n3013_, new_n3014_, new_n3015_, new_n3016_,
    new_n3017_, new_n3018_, new_n3019_, new_n3020_, new_n3021_, new_n3022_,
    new_n3023_, new_n3024_, new_n3025_, new_n3026_, new_n3027_, new_n3028_,
    new_n3029_, new_n3030_, new_n3031_, new_n3032_, new_n3033_, new_n3034_,
    new_n3035_, new_n3036_, new_n3037_, new_n3038_, new_n3039_, new_n3040_,
    new_n3041_, new_n3042_, new_n3043_, new_n3044_, new_n3045_, new_n3046_,
    new_n3047_, new_n3048_, new_n3049_, new_n3050_, new_n3051_, new_n3052_,
    new_n3053_, new_n3054_, new_n3055_, new_n3056_, new_n3057_, new_n3058_,
    new_n3059_, new_n3060_, new_n3061_, new_n3062_, new_n3063_, new_n3064_,
    new_n3065_, new_n3066_, new_n3067_, new_n3068_, new_n3069_, new_n3070_,
    new_n3071_, new_n3072_, new_n3073_, new_n3074_, new_n3075_, new_n3076_,
    new_n3077_, new_n3078_, new_n3079_, new_n3080_, new_n3081_, new_n3082_,
    new_n3083_, new_n3084_, new_n3085_, new_n3086_, new_n3087_, new_n3088_,
    new_n3089_, new_n3090_, new_n3091_, new_n3092_, new_n3093_, new_n3094_,
    new_n3095_, new_n3096_, new_n3097_, new_n3098_, new_n3099_, new_n3100_,
    new_n3101_, new_n3102_, new_n3103_, new_n3104_, new_n3105_, new_n3106_,
    new_n3107_, new_n3108_, new_n3109_, new_n3110_, new_n3111_, new_n3112_,
    new_n3113_, new_n3114_, new_n3115_, new_n3116_, new_n3117_, new_n3118_,
    new_n3119_, new_n3120_, new_n3121_, new_n3122_, new_n3123_, new_n3124_,
    new_n3125_, new_n3126_, new_n3127_, new_n3128_, new_n3129_, new_n3130_,
    new_n3131_, new_n3132_, new_n3133_, new_n3134_, new_n3135_, new_n3136_,
    new_n3137_, new_n3138_, new_n3139_, new_n3140_, new_n3141_, new_n3142_,
    new_n3143_, new_n3144_, new_n3145_, new_n3146_, new_n3147_, new_n3148_,
    new_n3149_, new_n3150_, new_n3151_, new_n3152_, new_n3153_, new_n3154_,
    new_n3155_, new_n3156_, new_n3157_, new_n3158_, new_n3159_, new_n3160_,
    new_n3161_, new_n3162_, new_n3163_, new_n3164_, new_n3165_, new_n3166_,
    new_n3167_, new_n3168_, new_n3169_, new_n3170_, new_n3171_, new_n3172_,
    new_n3173_, new_n3174_, new_n3175_, new_n3176_, new_n3177_, new_n3178_,
    new_n3179_, new_n3180_, new_n3181_, new_n3182_, new_n3183_, new_n3184_,
    new_n3185_, new_n3186_, new_n3187_, new_n3188_, new_n3189_, new_n3190_,
    new_n3191_, new_n3192_, new_n3193_, new_n3194_, new_n3195_, new_n3196_,
    new_n3197_, new_n3198_, new_n3199_, new_n3200_, new_n3201_, new_n3202_,
    new_n3203_, new_n3204_, new_n3205_, new_n3206_, new_n3207_, new_n3208_,
    new_n3209_, new_n3210_, new_n3211_, new_n3212_, new_n3213_, new_n3214_,
    new_n3215_, new_n3216_, new_n3217_, new_n3218_, new_n3219_, new_n3220_,
    new_n3221_, new_n3222_, new_n3223_, new_n3224_, new_n3225_, new_n3226_,
    new_n3227_, new_n3228_, new_n3229_, new_n3230_, new_n3231_, new_n3232_,
    new_n3233_, new_n3234_, new_n3235_, new_n3236_, new_n3237_, new_n3238_,
    new_n3239_, new_n3240_, new_n3241_, new_n3242_, new_n3243_, new_n3244_,
    new_n3245_, new_n3246_, new_n3247_, new_n3248_, new_n3249_, new_n3250_,
    new_n3251_, new_n3252_, new_n3253_, new_n3254_, new_n3255_, new_n3256_,
    new_n3257_, new_n3258_, new_n3259_, new_n3260_, new_n3261_, new_n3262_,
    new_n3263_, new_n3264_, new_n3265_, new_n3266_, new_n3267_, new_n3268_,
    new_n3269_, new_n3270_, new_n3271_, new_n3272_, new_n3273_, new_n3274_,
    new_n3275_, new_n3276_, new_n3277_, new_n3278_, new_n3279_, new_n3280_,
    new_n3281_, new_n3282_, new_n3283_, new_n3284_, new_n3285_, new_n3286_,
    new_n3287_, new_n3288_, new_n3289_, new_n3290_, new_n3291_, new_n3292_,
    new_n3293_, new_n3294_, new_n3295_, new_n3296_, new_n3297_, new_n3298_,
    new_n3299_, new_n3300_, new_n3301_, new_n3302_, new_n3303_, new_n3304_,
    new_n3305_, new_n3306_, new_n3307_, new_n3308_, new_n3309_, new_n3310_,
    new_n3311_, new_n3312_, new_n3313_, new_n3314_, new_n3315_, new_n3316_,
    new_n3317_, new_n3318_, new_n3319_, new_n3320_, new_n3321_, new_n3322_,
    new_n3323_, new_n3324_, new_n3325_, new_n3326_, new_n3327_, new_n3328_,
    new_n3329_, new_n3330_, new_n3331_, new_n3332_, new_n3333_, new_n3334_,
    new_n3335_, new_n3336_, new_n3337_, new_n3338_, new_n3339_, new_n3340_,
    new_n3341_, new_n3342_, new_n3343_, new_n3344_, new_n3345_, new_n3346_,
    new_n3347_, new_n3348_, new_n3349_, new_n3350_, new_n3351_, new_n3352_,
    new_n3353_, new_n3354_, new_n3355_, new_n3356_, new_n3357_, new_n3358_,
    new_n3359_, new_n3360_, new_n3361_, new_n3362_, new_n3363_, new_n3364_,
    new_n3365_, new_n3366_, new_n3367_, new_n3368_, new_n3369_, new_n3370_,
    new_n3371_, new_n3372_, new_n3373_, new_n3374_, new_n3375_, new_n3376_,
    new_n3377_, new_n3378_, new_n3379_, new_n3380_, new_n3381_, new_n3382_,
    new_n3383_, new_n3384_, new_n3385_, new_n3386_, new_n3387_, new_n3388_,
    new_n3389_, new_n3390_, new_n3391_, new_n3392_, new_n3393_, new_n3394_,
    new_n3395_, new_n3396_, new_n3397_, new_n3398_, new_n3399_, new_n3400_,
    new_n3401_, new_n3402_, new_n3403_, new_n3404_, new_n3405_, new_n3406_,
    new_n3407_, new_n3408_, new_n3409_, new_n3410_, new_n3411_, new_n3412_,
    new_n3413_, new_n3414_, new_n3415_, new_n3416_, new_n3417_, new_n3418_,
    new_n3419_, new_n3420_, new_n3421_, new_n3422_, new_n3423_, new_n3424_,
    new_n3425_, new_n3426_, new_n3427_, new_n3428_, new_n3429_, new_n3430_,
    new_n3431_, new_n3432_, new_n3433_, new_n3434_, new_n3435_, new_n3436_,
    new_n3437_, new_n3438_, new_n3439_, new_n3440_, new_n3441_, new_n3442_,
    new_n3443_, new_n3444_, new_n3445_, new_n3446_, new_n3447_, new_n3448_,
    new_n3449_, new_n3450_, new_n3451_, new_n3452_, new_n3453_, new_n3454_,
    new_n3455_, new_n3456_, new_n3457_, new_n3458_, new_n3459_, new_n3460_,
    new_n3461_, new_n3462_, new_n3463_, new_n3464_, new_n3465_, new_n3466_,
    new_n3467_, new_n3468_, new_n3469_, new_n3470_, new_n3471_, new_n3472_,
    new_n3473_, new_n3474_, new_n3475_, new_n3476_, new_n3477_, new_n3478_,
    new_n3479_, new_n3480_, new_n3481_, new_n3482_, new_n3483_, new_n3484_,
    new_n3485_, new_n3486_, new_n3487_, new_n3488_, new_n3489_, new_n3490_,
    new_n3491_, new_n3492_, new_n3493_, new_n3494_, new_n3495_, new_n3496_,
    new_n3497_, new_n3498_, new_n3499_, new_n3500_, new_n3501_, new_n3502_,
    new_n3503_, new_n3504_, new_n3505_, new_n3506_, new_n3507_, new_n3508_,
    new_n3509_, new_n3510_, new_n3511_, new_n3512_, new_n3513_, new_n3514_,
    new_n3515_, new_n3516_, new_n3517_, new_n3518_, new_n3519_, new_n3520_,
    new_n3521_, new_n3522_, new_n3523_, new_n3524_, new_n3525_, new_n3526_,
    new_n3527_, new_n3528_, new_n3529_, new_n3530_, new_n3531_, new_n3532_,
    new_n3533_, new_n3534_, new_n3535_, new_n3536_, new_n3537_, new_n3538_,
    new_n3539_, new_n3540_, new_n3541_, new_n3542_, new_n3543_, new_n3544_,
    new_n3545_, new_n3546_, new_n3547_, new_n3548_, new_n3549_, new_n3550_,
    new_n3551_, new_n3552_, new_n3553_, new_n3554_, new_n3555_, new_n3556_,
    new_n3557_, new_n3558_, new_n3559_, new_n3560_, new_n3561_, new_n3562_,
    new_n3563_, new_n3564_, new_n3565_, new_n3566_, new_n3567_, new_n3568_,
    new_n3569_, new_n3570_, new_n3571_, new_n3572_, new_n3573_, new_n3574_,
    new_n3575_, new_n3576_, new_n3577_, new_n3578_, new_n3579_, new_n3580_,
    new_n3581_, new_n3582_, new_n3583_, new_n3584_, new_n3585_, new_n3586_,
    new_n3587_, new_n3588_, new_n3589_, new_n3590_, new_n3591_, new_n3592_,
    new_n3593_, new_n3594_, new_n3595_, new_n3596_, new_n3597_, new_n3598_,
    new_n3599_, new_n3600_, new_n3601_, new_n3602_, new_n3603_, new_n3604_,
    new_n3605_, new_n3606_, new_n3607_, new_n3608_, new_n3609_, new_n3610_,
    new_n3611_, new_n3612_, new_n3613_, new_n3614_, new_n3615_, new_n3616_,
    new_n3617_, new_n3618_, new_n3619_, new_n3620_, new_n3621_, new_n3622_,
    new_n3623_, new_n3624_, new_n3625_, new_n3626_, new_n3627_, new_n3628_,
    new_n3629_, new_n3630_, new_n3631_, new_n3632_, new_n3633_, new_n3634_,
    new_n3635_, new_n3636_, new_n3637_, new_n3638_, new_n3639_, new_n3640_,
    new_n3641_, new_n3642_, new_n3643_, new_n3644_, new_n3645_, new_n3646_,
    new_n3647_, new_n3648_, new_n3649_, new_n3650_, new_n3651_, new_n3652_,
    new_n3653_, new_n3654_, new_n3655_, new_n3656_, new_n3657_, new_n3658_,
    new_n3659_, new_n3660_, new_n3661_, new_n3662_, new_n3663_, new_n3664_,
    new_n3665_, new_n3666_, new_n3667_, new_n3668_, new_n3669_, new_n3670_,
    new_n3671_, new_n3672_, new_n3673_, new_n3674_, new_n3675_, new_n3676_,
    new_n3677_, new_n3678_, new_n3679_, new_n3680_, new_n3681_, new_n3682_,
    new_n3683_, new_n3684_, new_n3685_, new_n3686_, new_n3687_, new_n3688_,
    new_n3689_, new_n3690_, new_n3691_, new_n3692_, new_n3693_, new_n3694_,
    new_n3695_, new_n3696_, new_n3697_, new_n3698_, new_n3699_, new_n3700_,
    new_n3701_, new_n3702_, new_n3703_, new_n3704_, new_n3705_, new_n3706_,
    new_n3707_, new_n3708_, new_n3709_, new_n3710_, new_n3711_, new_n3712_,
    new_n3713_, new_n3714_, new_n3715_, new_n3716_, new_n3717_, new_n3718_,
    new_n3719_, new_n3720_, new_n3721_, new_n3722_, new_n3723_, new_n3724_,
    new_n3725_, new_n3726_, new_n3727_, new_n3728_, new_n3729_, new_n3730_,
    new_n3731_, new_n3732_, new_n3733_, new_n3734_, new_n3735_, new_n3736_,
    new_n3737_, new_n3738_, new_n3739_, new_n3740_, new_n3741_, new_n3742_,
    new_n3743_, new_n3744_, new_n3745_, new_n3746_, new_n3747_, new_n3748_,
    new_n3749_, new_n3750_, new_n3751_, new_n3752_, new_n3753_, new_n3754_,
    new_n3755_, new_n3756_, new_n3757_, new_n3758_, new_n3759_, new_n3760_,
    new_n3761_, new_n3762_, new_n3763_, new_n3764_, new_n3765_, new_n3766_,
    new_n3767_, new_n3768_, new_n3769_, new_n3770_, new_n3771_, new_n3772_,
    new_n3773_, new_n3774_, new_n3775_, new_n3776_, new_n3777_, new_n3778_,
    new_n3779_, new_n3780_, new_n3781_, new_n3782_, new_n3783_, new_n3784_,
    new_n3785_, new_n3786_, new_n3787_, new_n3788_, new_n3789_, new_n3790_,
    new_n3791_, new_n3792_, new_n3793_, new_n3794_, new_n3795_, new_n3796_,
    new_n3797_, new_n3798_, new_n3799_, new_n3800_, new_n3801_, new_n3802_,
    new_n3803_, new_n3804_, new_n3805_, new_n3806_, new_n3807_, new_n3808_,
    new_n3809_, new_n3810_, new_n3811_, new_n3812_, new_n3813_, new_n3814_,
    new_n3815_, new_n3816_, new_n3817_, new_n3818_, new_n3819_, new_n3820_,
    new_n3821_, new_n3822_, new_n3823_, new_n3824_, new_n3825_, new_n3826_,
    new_n3827_, new_n3828_, new_n3829_, new_n3830_, new_n3831_, new_n3832_,
    new_n3833_, new_n3834_, new_n3835_, new_n3836_, new_n3837_, new_n3838_,
    new_n3839_, new_n3840_, new_n3841_, new_n3842_, new_n3843_, new_n3844_,
    new_n3845_, new_n3846_, new_n3847_, new_n3848_, new_n3849_, new_n3850_,
    new_n3851_, new_n3852_, new_n3853_, new_n3854_, new_n3855_, new_n3856_,
    new_n3857_, new_n3858_, new_n3859_, new_n3860_, new_n3861_, new_n3862_,
    new_n3863_, new_n3864_, new_n3865_, new_n3866_, new_n3867_, new_n3868_,
    new_n3869_, new_n3870_, new_n3871_, new_n3872_, new_n3873_, new_n3874_,
    new_n3875_, new_n3876_, new_n3877_, new_n3878_, new_n3879_, new_n3880_,
    new_n3881_, new_n3882_, new_n3883_, new_n3884_, new_n3885_, new_n3886_,
    new_n3887_, new_n3888_, new_n3889_, new_n3890_, new_n3891_, new_n3892_,
    new_n3893_, new_n3894_, new_n3895_, new_n3896_, new_n3897_, new_n3898_,
    new_n3899_, new_n3900_, new_n3901_, new_n3902_, new_n3903_, new_n3904_,
    new_n3905_, new_n3906_, new_n3907_, new_n3908_, new_n3909_, new_n3910_,
    new_n3911_, new_n3912_, new_n3913_, new_n3914_, new_n3915_, new_n3916_,
    new_n3917_, new_n3918_, new_n3919_, new_n3920_, new_n3921_, new_n3922_,
    new_n3923_, new_n3924_, new_n3925_, new_n3926_, new_n3927_, new_n3928_,
    new_n3929_, new_n3930_, new_n3931_, new_n3932_, new_n3933_, new_n3934_,
    new_n3935_, new_n3936_, new_n3937_, new_n3938_, new_n3939_, new_n3940_,
    new_n3941_, new_n3942_, new_n3943_, new_n3944_, new_n3945_, new_n3946_,
    new_n3947_, new_n3948_, new_n3949_, new_n3950_, new_n3951_, new_n3952_,
    new_n3953_, new_n3954_, new_n3955_, new_n3956_, new_n3957_, new_n3958_,
    new_n3959_, new_n3960_, new_n3961_, new_n3962_, new_n3963_, new_n3964_,
    new_n3965_, new_n3966_, new_n3967_, new_n3968_, new_n3969_, new_n3970_,
    new_n3971_, new_n3972_, new_n3973_, new_n3974_, new_n3975_, new_n3976_,
    new_n3977_, new_n3978_, new_n3979_, new_n3980_, new_n3981_, new_n3982_,
    new_n3983_, new_n3984_, new_n3985_, new_n3986_, new_n3987_, new_n3988_,
    new_n3989_, new_n3990_, new_n3991_, new_n3992_, new_n3993_, new_n3994_,
    new_n3995_, new_n3996_, new_n3997_, new_n3998_, new_n3999_, new_n4000_,
    new_n4001_, new_n4002_, new_n4003_, new_n4004_, new_n4005_, new_n4006_,
    new_n4007_, new_n4008_, new_n4009_, new_n4010_, new_n4011_, new_n4012_,
    new_n4013_, new_n4014_, new_n4015_, new_n4016_, new_n4017_, new_n4018_,
    new_n4019_, new_n4020_, new_n4021_, new_n4022_, new_n4023_, new_n4024_,
    new_n4025_, new_n4026_, new_n4027_, new_n4028_, new_n4029_, new_n4030_,
    new_n4031_, new_n4032_, new_n4033_, new_n4034_, new_n4035_, new_n4036_,
    new_n4037_, new_n4038_, new_n4039_, new_n4040_, new_n4041_, new_n4042_,
    new_n4043_, new_n4044_, new_n4045_, new_n4046_, new_n4047_, new_n4048_,
    new_n4049_, new_n4050_, new_n4051_, new_n4052_, new_n4053_, new_n4054_,
    new_n4055_, new_n4056_, new_n4057_, new_n4058_, new_n4059_, new_n4060_,
    new_n4061_, new_n4062_, new_n4063_, new_n4064_, new_n4065_, new_n4066_,
    new_n4067_, new_n4068_, new_n4069_, new_n4070_, new_n4071_, new_n4072_,
    new_n4073_, new_n4074_, new_n4075_, new_n4076_, new_n4077_, new_n4078_,
    new_n4079_, new_n4080_, new_n4081_, new_n4082_, new_n4083_, new_n4084_,
    new_n4085_, new_n4086_, new_n4087_, new_n4088_, new_n4089_, new_n4090_,
    new_n4091_, new_n4092_, new_n4093_, new_n4094_, new_n4095_, new_n4096_,
    new_n4097_, new_n4098_, new_n4099_, new_n4100_, new_n4101_, new_n4102_,
    new_n4103_, new_n4104_, new_n4105_, new_n4106_, new_n4107_, new_n4108_,
    new_n4109_, new_n4110_, new_n4111_, new_n4112_, new_n4113_, new_n4114_,
    new_n4115_, new_n4116_, new_n4117_, new_n4118_, new_n4119_, new_n4120_,
    new_n4121_, new_n4122_, new_n4123_, new_n4124_, new_n4125_, new_n4126_,
    new_n4127_, new_n4128_, new_n4129_, new_n4130_, new_n4131_, new_n4132_,
    new_n4133_, new_n4134_, new_n4135_, new_n4136_, new_n4137_, new_n4138_,
    new_n4139_, new_n4140_, new_n4141_, new_n4142_, new_n4143_, new_n4144_,
    new_n4145_, new_n4146_, new_n4147_, new_n4148_, new_n4149_, new_n4150_,
    new_n4151_, new_n4152_, new_n4153_, new_n4154_, new_n4155_, new_n4156_,
    new_n4157_, new_n4158_, new_n4159_, new_n4160_, new_n4161_, new_n4162_,
    new_n4163_, new_n4164_, new_n4165_, new_n4166_, new_n4167_, new_n4168_,
    new_n4169_, new_n4170_, new_n4171_, new_n4172_, new_n4173_, new_n4174_,
    new_n4175_, new_n4176_, new_n4177_, new_n4178_, new_n4179_, new_n4180_,
    new_n4181_, new_n4182_, new_n4183_, new_n4184_, new_n4185_, new_n4186_,
    new_n4187_, new_n4188_, new_n4189_, new_n4190_, new_n4191_, new_n4192_,
    new_n4193_, new_n4194_, new_n4195_, new_n4196_, new_n4197_, new_n4198_,
    new_n4199_, new_n4200_, new_n4201_, new_n4202_, new_n4203_, new_n4204_,
    new_n4205_, new_n4206_, new_n4207_, new_n4208_, new_n4209_, new_n4210_,
    new_n4211_, new_n4212_, new_n4213_, new_n4214_, new_n4215_, new_n4216_,
    new_n4217_, new_n4218_, new_n4219_, new_n4220_, new_n4221_, new_n4222_,
    new_n4223_, new_n4224_, new_n4225_, new_n4226_, new_n4227_, new_n4228_,
    new_n4229_, new_n4230_, new_n4231_, new_n4232_, new_n4233_, new_n4234_,
    new_n4235_, new_n4236_, new_n4237_, new_n4238_, new_n4239_, new_n4240_,
    new_n4241_, new_n4242_, new_n4243_, new_n4244_, new_n4245_, new_n4246_,
    new_n4247_, new_n4248_, new_n4249_, new_n4250_, new_n4251_, new_n4252_,
    new_n4253_, new_n4254_, new_n4255_, new_n4256_, new_n4257_, new_n4258_,
    new_n4259_, new_n4260_, new_n4261_, new_n4262_, new_n4263_, new_n4264_,
    new_n4265_, new_n4266_, new_n4267_, new_n4268_, new_n4269_, new_n4270_,
    new_n4271_, new_n4272_, new_n4273_, new_n4274_, new_n4275_, new_n4276_,
    new_n4277_, new_n4278_, new_n4279_, new_n4280_, new_n4281_, new_n4282_,
    new_n4283_, new_n4284_, new_n4285_, new_n4286_, new_n4287_, new_n4288_,
    new_n4289_, new_n4290_, new_n4291_, new_n4292_, new_n4293_, new_n4294_,
    new_n4295_, new_n4296_, new_n4297_, new_n4298_, new_n4299_, new_n4300_,
    new_n4301_, new_n4302_, new_n4303_, new_n4304_, new_n4305_, new_n4306_,
    new_n4307_, new_n4308_, new_n4309_, new_n4310_, new_n4311_, new_n4312_,
    new_n4313_, new_n4314_, new_n4315_, new_n4316_, new_n4317_, new_n4318_,
    new_n4319_, new_n4320_, new_n4321_, new_n4322_, new_n4323_, new_n4324_,
    new_n4325_, new_n4326_, new_n4327_, new_n4328_, new_n4329_, new_n4330_,
    new_n4331_, new_n4332_, new_n4333_, new_n4334_, new_n4335_, new_n4336_,
    new_n4337_, new_n4338_, new_n4339_, new_n4340_, new_n4341_, new_n4342_,
    new_n4343_, new_n4344_, new_n4345_, new_n4346_, new_n4347_, new_n4348_,
    new_n4349_, new_n4350_, new_n4351_, new_n4352_, new_n4353_, new_n4354_,
    new_n4355_, new_n4356_, new_n4357_, new_n4358_, new_n4359_, new_n4360_,
    new_n4361_, new_n4362_, new_n4363_, new_n4364_, new_n4365_, new_n4366_,
    new_n4367_, new_n4368_, new_n4369_, new_n4370_, new_n4371_, new_n4372_,
    new_n4373_, new_n4374_, new_n4375_, new_n4376_, new_n4377_, new_n4378_,
    new_n4379_, new_n4380_, new_n4381_, new_n4382_, new_n4383_, new_n4384_,
    new_n4385_, new_n4386_, new_n4387_, new_n4388_, new_n4389_, new_n4390_,
    new_n4391_, new_n4392_, new_n4393_, new_n4394_, new_n4395_, new_n4396_,
    new_n4397_, new_n4398_, new_n4399_, new_n4400_, new_n4401_, new_n4402_,
    new_n4403_, new_n4404_, new_n4405_, new_n4406_, new_n4407_, new_n4408_,
    new_n4409_, new_n4410_, new_n4411_, new_n4412_, new_n4413_, new_n4414_,
    new_n4415_, new_n4416_, new_n4417_, new_n4418_, new_n4419_, new_n4420_,
    new_n4421_, new_n4422_, new_n4423_, new_n4424_, new_n4425_, new_n4426_,
    new_n4427_, new_n4428_, new_n4429_, new_n4430_, new_n4431_, new_n4432_,
    new_n4433_, new_n4434_, new_n4435_, new_n4436_, new_n4437_, new_n4438_,
    new_n4439_, new_n4440_, new_n4441_, new_n4442_, new_n4443_, new_n4444_,
    new_n4445_, new_n4446_, new_n4447_, new_n4448_, new_n4449_, new_n4450_,
    new_n4451_, new_n4452_, new_n4453_, new_n4454_, new_n4455_, new_n4456_,
    new_n4457_, new_n4458_, new_n4459_, new_n4460_, new_n4461_, new_n4462_,
    new_n4463_, new_n4464_, new_n4465_, new_n4466_, new_n4467_, new_n4468_,
    new_n4469_, new_n4470_, new_n4471_, new_n4472_, new_n4473_, new_n4474_,
    new_n4475_, new_n4476_, new_n4477_, new_n4478_, new_n4479_, new_n4480_,
    new_n4481_, new_n4482_, new_n4483_, new_n4484_, new_n4485_, new_n4486_,
    new_n4487_, new_n4488_, new_n4489_, new_n4490_, new_n4491_, new_n4492_,
    new_n4493_, new_n4494_, new_n4495_, new_n4496_, new_n4497_, new_n4498_,
    new_n4499_, new_n4500_, new_n4501_, new_n4502_, new_n4503_, new_n4504_,
    new_n4505_, new_n4506_, new_n4507_, new_n4508_, new_n4509_, new_n4510_,
    new_n4511_, new_n4512_, new_n4513_, new_n4514_, new_n4515_, new_n4516_,
    new_n4517_, new_n4518_, new_n4519_, new_n4520_, new_n4521_, new_n4522_,
    new_n4523_, new_n4524_, new_n4525_, new_n4526_, new_n4527_, new_n4528_,
    new_n4529_, new_n4530_, new_n4531_, new_n4532_, new_n4533_, new_n4534_,
    new_n4535_, new_n4536_, new_n4537_, new_n4538_, new_n4539_, new_n4540_,
    new_n4541_, new_n4542_, new_n4543_, new_n4544_, new_n4545_, new_n4546_,
    new_n4547_, new_n4548_, new_n4549_, new_n4550_, new_n4551_, new_n4552_,
    new_n4553_, new_n4554_, new_n4555_, new_n4556_, new_n4557_, new_n4558_,
    new_n4559_, new_n4560_, new_n4561_, new_n4562_, new_n4563_, new_n4564_,
    new_n4565_, new_n4566_, new_n4567_, new_n4568_, new_n4569_, new_n4570_,
    new_n4571_, new_n4572_, new_n4573_, new_n4574_, new_n4575_, new_n4576_,
    new_n4577_, new_n4578_, new_n4579_, new_n4580_, new_n4581_, new_n4582_,
    new_n4583_, new_n4584_, new_n4585_, new_n4586_, new_n4587_, new_n4588_,
    new_n4589_, new_n4590_, new_n4591_, new_n4592_, new_n4593_, new_n4594_,
    new_n4595_, new_n4596_, new_n4597_, new_n4598_, new_n4599_, new_n4600_,
    new_n4601_, new_n4602_, new_n4603_, new_n4604_, new_n4605_, new_n4606_,
    new_n4607_, new_n4608_, new_n4609_, new_n4610_, new_n4611_, new_n4612_,
    new_n4613_, new_n4614_, new_n4615_, new_n4616_, new_n4617_, new_n4618_,
    new_n4619_, new_n4620_, new_n4621_, new_n4622_, new_n4623_, new_n4624_,
    new_n4625_, new_n4626_, new_n4627_, new_n4628_, new_n4629_, new_n4630_,
    new_n4631_, new_n4632_, new_n4633_, new_n4634_, new_n4635_, new_n4636_,
    new_n4637_, new_n4638_, new_n4639_, new_n4640_, new_n4641_, new_n4642_,
    new_n4643_, new_n4644_, new_n4645_, new_n4646_, new_n4647_, new_n4648_,
    new_n4649_, new_n4650_, new_n4651_, new_n4652_, new_n4653_, new_n4654_,
    new_n4655_, new_n4656_, new_n4657_, new_n4658_, new_n4659_, new_n4660_,
    new_n4661_, new_n4662_, new_n4663_, new_n4664_, new_n4665_, new_n4666_,
    new_n4667_, new_n4668_, new_n4669_, new_n4670_, new_n4671_, new_n4672_,
    new_n4673_, new_n4674_, new_n4675_, new_n4676_, new_n4677_, new_n4678_,
    new_n4679_, new_n4680_, new_n4681_, new_n4682_, new_n4683_, new_n4684_,
    new_n4685_, new_n4686_, new_n4687_, new_n4688_, new_n4689_, new_n4690_,
    new_n4691_, new_n4692_, new_n4693_, new_n4694_, new_n4695_, new_n4696_,
    new_n4697_, new_n4698_, new_n4699_, new_n4700_, new_n4701_, new_n4702_,
    new_n4703_, new_n4704_, new_n4705_, new_n4706_, new_n4707_, new_n4708_,
    new_n4709_, new_n4710_, new_n4711_, new_n4712_, new_n4713_, new_n4714_,
    new_n4715_, new_n4716_, new_n4717_, new_n4718_, new_n4719_, new_n4720_,
    new_n4721_, new_n4722_, new_n4723_, new_n4724_, new_n4725_, new_n4726_,
    new_n4727_, new_n4728_, new_n4729_, new_n4730_, new_n4731_, new_n4732_,
    new_n4733_, new_n4734_, new_n4735_, new_n4736_, new_n4737_, new_n4738_,
    new_n4739_, new_n4740_, new_n4741_, new_n4742_, new_n4743_, new_n4744_,
    new_n4745_, new_n4746_, new_n4747_, new_n4748_, new_n4749_, new_n4750_,
    new_n4751_, new_n4752_, new_n4753_, new_n4754_, new_n4755_, new_n4756_,
    new_n4757_, new_n4758_, new_n4759_, new_n4760_, new_n4761_, new_n4762_,
    new_n4763_, new_n4764_, new_n4765_, new_n4766_, new_n4767_, new_n4768_,
    new_n4769_, new_n4770_, new_n4771_, new_n4772_, new_n4773_, new_n4774_,
    new_n4775_, new_n4776_, new_n4777_, new_n4778_, new_n4779_, new_n4780_,
    new_n4781_, new_n4782_, new_n4783_, new_n4784_, new_n4785_, new_n4786_,
    new_n4787_, new_n4788_, new_n4789_, new_n4790_, new_n4791_, new_n4792_,
    new_n4793_, new_n4794_, new_n4795_, new_n4796_, new_n4797_, new_n4798_,
    new_n4799_, new_n4800_, new_n4801_, new_n4802_, new_n4803_, new_n4804_,
    new_n4805_, new_n4806_, new_n4807_, new_n4808_, new_n4809_, new_n4810_,
    new_n4811_, new_n4812_, new_n4813_, new_n4814_, new_n4815_, new_n4816_,
    new_n4817_, new_n4818_, new_n4819_, new_n4820_, new_n4821_, new_n4822_,
    new_n4823_, new_n4824_, new_n4825_, new_n4826_, new_n4827_, new_n4828_,
    new_n4829_, new_n4830_, new_n4831_, new_n4832_, new_n4833_, new_n4834_,
    new_n4835_, new_n4836_, new_n4837_, new_n4838_, new_n4839_, new_n4840_,
    new_n4841_, new_n4842_, new_n4843_, new_n4844_, new_n4845_, new_n4846_,
    new_n4847_, new_n4848_, new_n4849_, new_n4850_, new_n4851_, new_n4852_,
    new_n4853_, new_n4854_, new_n4855_, new_n4856_, new_n4857_, new_n4858_,
    new_n4859_, new_n4860_, new_n4861_, new_n4862_, new_n4863_, new_n4864_,
    new_n4865_, new_n4866_, new_n4867_, new_n4868_, new_n4869_, new_n4870_,
    new_n4871_, new_n4872_, new_n4873_, new_n4874_, new_n4875_, new_n4876_,
    new_n4877_, new_n4878_, new_n4879_, new_n4880_, new_n4881_, new_n4882_,
    new_n4883_, new_n4884_, new_n4885_, new_n4886_, new_n4887_, new_n4888_,
    new_n4889_, new_n4890_, new_n4891_, new_n4892_, new_n4893_, new_n4894_,
    new_n4895_, new_n4896_, new_n4897_, new_n4898_, new_n4899_, new_n4900_,
    new_n4901_, new_n4902_, new_n4903_, new_n4904_, new_n4905_, new_n4906_,
    new_n4907_, new_n4908_, new_n4909_, new_n4910_, new_n4911_, new_n4912_,
    new_n4913_, new_n4914_, new_n4915_, new_n4916_, new_n4917_, new_n4918_,
    new_n4919_, new_n4920_, new_n4921_, new_n4922_, new_n4923_, new_n4924_,
    new_n4925_, new_n4926_, new_n4927_, new_n4928_, new_n4929_, new_n4930_,
    new_n4931_, new_n4932_, new_n4933_, new_n4934_, new_n4935_, new_n4936_,
    new_n4937_, new_n4938_, new_n4939_, new_n4940_, new_n4941_, new_n4942_,
    new_n4943_, new_n4944_, new_n4945_, new_n4946_, new_n4947_, new_n4948_,
    new_n4949_, new_n4950_, new_n4951_, new_n4952_, new_n4953_, new_n4954_,
    new_n4955_, new_n4956_, new_n4957_, new_n4958_, new_n4959_, new_n4960_,
    new_n4961_, new_n4962_, new_n4963_, new_n4964_, new_n4965_, new_n4966_,
    new_n4967_, new_n4968_, new_n4969_, new_n4970_, new_n4971_, new_n4972_,
    new_n4973_, new_n4974_, new_n4975_, new_n4976_, new_n4977_, new_n4978_,
    new_n4979_, new_n4980_, new_n4981_, new_n4982_, new_n4983_, new_n4984_,
    new_n4985_, new_n4986_, new_n4987_, new_n4988_, new_n4989_, new_n4990_,
    new_n4991_, new_n4992_, new_n4993_, new_n4994_, new_n4995_, new_n4996_,
    new_n4997_, new_n4998_, new_n4999_, new_n5000_, new_n5001_, new_n5002_,
    new_n5003_, new_n5004_, new_n5005_, new_n5006_, new_n5007_, new_n5008_,
    new_n5009_, new_n5010_, new_n5011_, new_n5012_, new_n5013_, new_n5014_,
    new_n5015_, new_n5016_, new_n5017_, new_n5018_, new_n5019_, new_n5020_,
    new_n5021_, new_n5022_, new_n5023_, new_n5024_, new_n5025_, new_n5026_,
    new_n5027_, new_n5028_, new_n5029_, new_n5030_, new_n5031_, new_n5032_,
    new_n5033_, new_n5034_, new_n5035_, new_n5036_, new_n5037_, new_n5038_,
    new_n5039_, new_n5040_, new_n5041_, new_n5042_, new_n5043_, new_n5044_,
    new_n5045_, new_n5046_, new_n5047_, new_n5048_, new_n5049_, new_n5050_,
    new_n5051_, new_n5052_, new_n5053_, new_n5054_, new_n5055_, new_n5056_,
    new_n5057_, new_n5058_, new_n5059_, new_n5060_, new_n5061_, new_n5062_,
    new_n5063_, new_n5064_, new_n5065_, new_n5066_, new_n5067_, new_n5068_,
    new_n5069_, new_n5070_, new_n5071_, new_n5072_, new_n5073_, new_n5074_,
    new_n5075_, new_n5076_, new_n5077_, new_n5078_, new_n5079_, new_n5080_,
    new_n5081_, new_n5082_, new_n5083_, new_n5084_, new_n5085_, new_n5086_,
    new_n5087_, new_n5088_, new_n5089_, new_n5090_, new_n5091_, new_n5092_,
    new_n5093_, new_n5094_, new_n5095_, new_n5096_, new_n5097_, new_n5098_,
    new_n5099_, new_n5100_, new_n5101_, new_n5102_, new_n5103_, new_n5104_,
    new_n5105_, new_n5106_, new_n5107_, new_n5108_, new_n5109_, new_n5110_,
    new_n5111_, new_n5112_, new_n5113_, new_n5114_, new_n5115_, new_n5116_,
    new_n5117_, new_n5118_, new_n5119_, new_n5120_, new_n5121_, new_n5122_,
    new_n5123_, new_n5124_, new_n5125_, new_n5126_, new_n5127_, new_n5128_,
    new_n5129_, new_n5130_, new_n5131_, new_n5132_, new_n5133_, new_n5134_,
    new_n5135_, new_n5136_, new_n5137_, new_n5138_, new_n5139_, new_n5140_,
    new_n5141_, new_n5142_, new_n5143_, new_n5144_, new_n5145_, new_n5146_,
    new_n5147_, new_n5148_, new_n5149_, new_n5150_, new_n5151_, new_n5152_,
    new_n5153_, new_n5154_, new_n5155_, new_n5156_, new_n5157_, new_n5158_,
    new_n5159_, new_n5160_, new_n5161_, new_n5162_, new_n5163_, new_n5164_,
    new_n5165_, new_n5166_, new_n5167_, new_n5168_, new_n5169_, new_n5170_,
    new_n5171_, new_n5172_, new_n5173_, new_n5174_, new_n5175_, new_n5176_,
    new_n5177_, new_n5178_, new_n5179_, new_n5180_, new_n5181_, new_n5182_,
    new_n5183_, new_n5184_, new_n5185_, new_n5186_, new_n5187_, new_n5188_,
    new_n5189_, new_n5190_, new_n5191_, new_n5192_, new_n5193_, new_n5194_,
    new_n5195_, new_n5196_, new_n5197_, new_n5198_, new_n5199_, new_n5200_,
    new_n5201_, new_n5202_, new_n5203_, new_n5204_, new_n5205_, new_n5206_,
    new_n5207_, new_n5208_, new_n5209_, new_n5210_, new_n5211_, new_n5212_,
    new_n5213_, new_n5214_, new_n5215_, new_n5216_, new_n5217_, new_n5218_,
    new_n5219_, new_n5220_, new_n5221_, new_n5222_, new_n5223_, new_n5224_,
    new_n5225_, new_n5226_, new_n5227_, new_n5228_, new_n5229_, new_n5230_,
    new_n5231_, new_n5232_, new_n5233_, new_n5234_, new_n5235_, new_n5236_,
    new_n5237_, new_n5238_, new_n5239_, new_n5240_, new_n5241_, new_n5242_,
    new_n5243_, new_n5244_, new_n5245_, new_n5246_, new_n5247_, new_n5248_,
    new_n5249_, new_n5250_, new_n5251_, new_n5252_, new_n5253_, new_n5254_,
    new_n5255_, new_n5256_, new_n5257_, new_n5258_, new_n5259_, new_n5260_,
    new_n5261_, new_n5262_, new_n5263_, new_n5264_, new_n5265_, new_n5266_,
    new_n5267_, new_n5268_, new_n5269_, new_n5270_, new_n5271_, new_n5272_,
    new_n5273_, new_n5274_, new_n5275_, new_n5276_, new_n5277_, new_n5278_,
    new_n5279_, new_n5280_, new_n5281_, new_n5282_, new_n5283_, new_n5284_,
    new_n5285_, new_n5286_, new_n5287_, new_n5288_, new_n5289_, new_n5290_,
    new_n5291_, new_n5292_, new_n5293_, new_n5294_, new_n5295_, new_n5296_,
    new_n5297_, new_n5298_, new_n5299_, new_n5300_, new_n5301_, new_n5302_,
    new_n5303_, new_n5304_, new_n5305_, new_n5306_, new_n5307_, new_n5308_,
    new_n5309_, new_n5310_, new_n5311_, new_n5312_, new_n5313_, new_n5314_,
    new_n5315_, new_n5316_, new_n5317_, new_n5318_, new_n5319_, new_n5320_,
    new_n5321_, new_n5322_, new_n5323_, new_n5324_, new_n5325_, new_n5326_,
    new_n5327_, new_n5328_, new_n5329_, new_n5330_, new_n5331_, new_n5332_,
    new_n5333_, new_n5334_, new_n5335_, new_n5336_, new_n5337_, new_n5338_,
    new_n5339_, new_n5340_, new_n5341_, new_n5342_, new_n5343_, new_n5344_,
    new_n5345_, new_n5346_, new_n5347_, new_n5348_, new_n5349_, new_n5350_,
    new_n5351_, new_n5352_, new_n5353_, new_n5354_, new_n5355_, new_n5356_,
    new_n5357_, new_n5358_, new_n5359_, new_n5360_, new_n5361_, new_n5362_,
    new_n5363_, new_n5364_, new_n5365_, new_n5366_, new_n5367_, new_n5368_,
    new_n5369_, new_n5370_, new_n5371_, new_n5372_, new_n5373_, new_n5374_,
    new_n5375_, new_n5376_, new_n5377_, new_n5378_, new_n5379_, new_n5380_,
    new_n5381_, new_n5382_, new_n5383_, new_n5384_, new_n5385_, new_n5386_,
    new_n5387_, new_n5388_, new_n5389_, new_n5390_, new_n5391_, new_n5392_,
    new_n5393_, new_n5394_, new_n5395_, new_n5396_, new_n5397_, new_n5398_,
    new_n5399_, new_n5400_, new_n5401_, new_n5402_, new_n5403_, new_n5404_,
    new_n5405_, new_n5406_, new_n5407_, new_n5408_, new_n5409_, new_n5410_,
    new_n5411_, new_n5412_, new_n5413_, new_n5414_, new_n5415_, new_n5416_,
    new_n5417_, new_n5418_, new_n5419_, new_n5420_, new_n5421_, new_n5422_,
    new_n5423_, new_n5424_, new_n5425_, new_n5426_, new_n5427_, new_n5428_,
    new_n5429_, new_n5430_, new_n5431_, new_n5432_, new_n5433_, new_n5434_,
    new_n5435_, new_n5436_, new_n5437_, new_n5438_, new_n5439_, new_n5440_,
    new_n5441_, new_n5442_, new_n5443_, new_n5444_, new_n5445_, new_n5446_,
    new_n5447_, new_n5448_, new_n5449_, new_n5450_, new_n5451_, new_n5452_,
    new_n5453_, new_n5454_, new_n5455_, new_n5456_, new_n5457_, new_n5458_,
    new_n5459_, new_n5460_, new_n5461_, new_n5462_, new_n5463_, new_n5464_,
    new_n5465_, new_n5466_, new_n5467_, new_n5468_, new_n5469_, new_n5470_,
    new_n5471_, new_n5472_, new_n5473_, new_n5474_, new_n5475_, new_n5476_,
    new_n5477_, new_n5478_, new_n5479_, new_n5480_, new_n5481_, new_n5482_,
    new_n5483_, new_n5484_, new_n5485_, new_n5486_, new_n5487_, new_n5488_,
    new_n5489_, new_n5490_, new_n5491_, new_n5492_, new_n5493_, new_n5494_,
    new_n5495_, new_n5496_, new_n5497_, new_n5498_, new_n5499_, new_n5500_,
    new_n5501_, new_n5502_, new_n5503_, new_n5504_, new_n5505_, new_n5506_,
    new_n5507_, new_n5508_, new_n5509_, new_n5510_, new_n5511_, new_n5512_,
    new_n5513_, new_n5514_, new_n5515_, new_n5516_, new_n5517_, new_n5518_,
    new_n5519_, new_n5520_, new_n5521_, new_n5522_, new_n5523_, new_n5524_,
    new_n5525_, new_n5526_, new_n5527_, new_n5528_, new_n5529_, new_n5530_,
    new_n5531_, new_n5532_, new_n5533_, new_n5534_, new_n5535_, new_n5536_,
    new_n5537_, new_n5538_, new_n5539_, new_n5540_, new_n5541_, new_n5542_,
    new_n5543_, new_n5544_, new_n5545_, new_n5546_, new_n5547_, new_n5548_,
    new_n5549_, new_n5550_, new_n5551_, new_n5552_, new_n5553_, new_n5554_,
    new_n5555_, new_n5556_, new_n5557_, new_n5558_, new_n5559_, new_n5560_,
    new_n5561_, new_n5562_, new_n5563_, new_n5564_, new_n5565_, new_n5566_,
    new_n5567_, new_n5568_, new_n5569_, new_n5570_, new_n5571_, new_n5572_,
    new_n5573_, new_n5574_, new_n5575_, new_n5576_, new_n5577_, new_n5578_,
    new_n5579_, new_n5580_, new_n5581_, new_n5582_, new_n5583_, new_n5584_,
    new_n5585_, new_n5586_, new_n5587_, new_n5588_, new_n5589_, new_n5590_,
    new_n5591_, new_n5592_, new_n5593_, new_n5594_, new_n5595_, new_n5596_,
    new_n5597_, new_n5598_, new_n5599_, new_n5600_, new_n5601_, new_n5602_,
    new_n5603_, new_n5604_, new_n5605_, new_n5606_, new_n5607_, new_n5608_,
    new_n5609_, new_n5610_, new_n5611_, new_n5612_, new_n5613_, new_n5614_,
    new_n5615_, new_n5616_, new_n5617_, new_n5618_, new_n5619_, new_n5620_,
    new_n5621_, new_n5622_, new_n5623_, new_n5624_, new_n5625_, new_n5626_,
    new_n5627_, new_n5628_, new_n5629_, new_n5630_, new_n5631_, new_n5632_,
    new_n5633_, new_n5634_, new_n5635_, new_n5636_, new_n5637_, new_n5638_,
    new_n5639_, new_n5640_, new_n5641_, new_n5642_, new_n5643_, new_n5644_,
    new_n5645_, new_n5646_, new_n5647_, new_n5648_, new_n5649_, new_n5650_,
    new_n5651_, new_n5652_, new_n5653_, new_n5654_, new_n5655_, new_n5656_,
    new_n5657_, new_n5658_, new_n5659_, new_n5660_, new_n5661_, new_n5662_,
    new_n5663_, new_n5664_, new_n5665_, new_n5666_, new_n5667_, new_n5668_,
    new_n5669_, new_n5670_, new_n5671_, new_n5672_, new_n5673_, new_n5674_,
    new_n5675_, new_n5676_, new_n5677_, new_n5678_, new_n5679_, new_n5680_,
    new_n5681_, new_n5682_, new_n5683_, new_n5684_, new_n5685_, new_n5686_,
    new_n5687_, new_n5688_, new_n5689_, new_n5690_, new_n5691_, new_n5692_,
    new_n5693_, new_n5694_, new_n5695_, new_n5696_, new_n5697_, new_n5698_,
    new_n5699_, new_n5700_, new_n5701_, new_n5702_, new_n5703_, new_n5704_,
    new_n5705_, new_n5706_, new_n5707_, new_n5708_, new_n5709_, new_n5710_,
    new_n5711_, new_n5712_, new_n5713_, new_n5714_, new_n5715_, new_n5716_,
    new_n5717_, new_n5718_, new_n5719_, new_n5720_, new_n5721_, new_n5722_,
    new_n5723_, new_n5724_, new_n5725_, new_n5726_, new_n5727_, new_n5728_,
    new_n5729_, new_n5730_, new_n5731_, new_n5732_, new_n5733_, new_n5734_,
    new_n5735_, new_n5736_, new_n5737_, new_n5738_, new_n5739_, new_n5740_,
    new_n5741_, new_n5742_, new_n5743_, new_n5744_, new_n5745_, new_n5746_,
    new_n5747_, new_n5748_, new_n5749_, new_n5750_, new_n5751_, new_n5752_,
    new_n5753_, new_n5754_, new_n5755_, new_n5756_, new_n5757_, new_n5758_,
    new_n5759_, new_n5760_, new_n5761_, new_n5762_, new_n5763_, new_n5764_,
    new_n5765_, new_n5766_, new_n5767_, new_n5768_, new_n5769_, new_n5770_,
    new_n5771_, new_n5772_, new_n5773_, new_n5774_, new_n5775_, new_n5776_,
    new_n5777_, new_n5778_, new_n5779_, new_n5780_, new_n5781_, new_n5782_,
    new_n5783_, new_n5784_, new_n5785_, new_n5786_, new_n5787_, new_n5788_,
    new_n5789_, new_n5790_, new_n5791_, new_n5792_, new_n5793_, new_n5794_,
    new_n5795_, new_n5796_, new_n5797_, new_n5798_, new_n5799_, new_n5800_,
    new_n5801_, new_n5802_, new_n5803_, new_n5804_, new_n5805_, new_n5806_,
    new_n5807_, new_n5808_, new_n5809_, new_n5810_, new_n5811_, new_n5812_,
    new_n5813_, new_n5814_, new_n5815_, new_n5816_, new_n5817_, new_n5818_,
    new_n5819_, new_n5820_, new_n5821_, new_n5822_, new_n5823_, new_n5824_,
    new_n5825_, new_n5826_, new_n5827_, new_n5828_, new_n5829_, new_n5830_,
    new_n5831_, new_n5832_, new_n5833_, new_n5834_, new_n5835_, new_n5836_,
    new_n5837_, new_n5838_, new_n5839_, new_n5840_, new_n5841_, new_n5842_,
    new_n5843_, new_n5844_, new_n5845_, new_n5846_, new_n5847_, new_n5848_,
    new_n5849_, new_n5850_, new_n5851_, new_n5852_, new_n5853_, new_n5854_,
    new_n5855_, new_n5856_, new_n5857_, new_n5858_, new_n5859_, new_n5860_,
    new_n5861_, new_n5862_, new_n5863_, new_n5864_, new_n5865_, new_n5866_,
    new_n5867_, new_n5868_, new_n5869_, new_n5870_, new_n5871_, new_n5872_,
    new_n5873_, new_n5874_, new_n5875_, new_n5876_, new_n5877_, new_n5878_,
    new_n5879_, new_n5880_, new_n5881_, new_n5882_, new_n5883_, new_n5884_,
    new_n5885_, new_n5886_, new_n5887_, new_n5888_, new_n5889_, new_n5890_,
    new_n5891_, new_n5892_, new_n5893_, new_n5894_, new_n5895_, new_n5896_,
    new_n5897_, new_n5898_, new_n5899_, new_n5900_, new_n5901_, new_n5902_,
    new_n5903_, new_n5904_, new_n5905_, new_n5906_, new_n5907_, new_n5908_,
    new_n5909_, new_n5910_, new_n5911_, new_n5912_, new_n5913_, new_n5914_,
    new_n5915_, new_n5916_, new_n5917_, new_n5918_, new_n5919_, new_n5920_,
    new_n5921_, new_n5922_, new_n5923_, new_n5924_, new_n5925_, new_n5926_,
    new_n5927_, new_n5928_, new_n5929_, new_n5930_, new_n5931_, new_n5932_,
    new_n5933_, new_n5934_, new_n5935_, new_n5936_, new_n5937_, new_n5938_,
    new_n5939_, new_n5940_, new_n5941_, new_n5942_, new_n5943_, new_n5944_,
    new_n5945_, new_n5946_, new_n5947_, new_n5948_, new_n5949_, new_n5950_,
    new_n5951_, new_n5952_, new_n5953_, new_n5954_, new_n5955_, new_n5956_,
    new_n5957_, new_n5958_, new_n5959_, new_n5960_, new_n5961_, new_n5962_,
    new_n5963_, new_n5964_, new_n5965_, new_n5966_, new_n5967_, new_n5968_,
    new_n5969_, new_n5970_, new_n5971_, new_n5972_, new_n5973_, new_n5974_,
    new_n5975_, new_n5976_, new_n5977_, new_n5978_, new_n5979_, new_n5980_,
    new_n5981_, new_n5982_, new_n5983_, new_n5984_, new_n5985_, new_n5986_,
    new_n5987_, new_n5988_, new_n5989_, new_n5990_, new_n5991_, new_n5992_,
    new_n5993_, new_n5994_, new_n5995_, new_n5996_, new_n5997_, new_n5998_,
    new_n5999_, new_n6000_, new_n6001_, new_n6002_, new_n6003_, new_n6004_,
    new_n6005_, new_n6006_, new_n6007_, new_n6008_, new_n6009_, new_n6010_,
    new_n6011_, new_n6012_, new_n6013_, new_n6014_, new_n6015_, new_n6016_,
    new_n6017_, new_n6018_, new_n6019_, new_n6020_, new_n6021_, new_n6022_,
    new_n6023_, new_n6024_, new_n6025_, new_n6026_, new_n6027_, new_n6028_,
    new_n6029_, new_n6030_, new_n6031_, new_n6032_, new_n6033_, new_n6034_,
    new_n6035_, new_n6036_, new_n6037_, new_n6038_, new_n6039_, new_n6040_,
    new_n6041_, new_n6042_, new_n6043_, new_n6044_, new_n6045_, new_n6046_,
    new_n6047_, new_n6048_, new_n6049_, new_n6050_, new_n6051_, new_n6052_,
    new_n6053_, new_n6054_, new_n6055_, new_n6056_, new_n6057_, new_n6058_,
    new_n6059_, new_n6060_, new_n6061_, new_n6062_, new_n6063_, new_n6064_,
    new_n6065_, new_n6066_, new_n6067_, new_n6068_, new_n6069_, new_n6070_,
    new_n6071_, new_n6072_, new_n6073_, new_n6074_, new_n6075_, new_n6076_,
    new_n6077_, new_n6078_, new_n6079_, new_n6080_, new_n6081_, new_n6082_,
    new_n6083_, new_n6084_, new_n6085_, new_n6086_, new_n6087_, new_n6088_,
    new_n6089_, new_n6090_, new_n6091_, new_n6092_, new_n6093_, new_n6094_,
    new_n6095_, new_n6096_, new_n6097_, new_n6098_, new_n6099_, new_n6100_,
    new_n6101_, new_n6102_, new_n6103_, new_n6104_, new_n6105_, new_n6106_,
    new_n6107_, new_n6108_, new_n6109_, new_n6110_, new_n6111_, new_n6112_,
    new_n6113_, new_n6114_, new_n6115_, new_n6116_, new_n6117_, new_n6118_,
    new_n6119_, new_n6120_, new_n6121_, new_n6122_, new_n6123_, new_n6124_,
    new_n6125_, new_n6126_, new_n6127_, new_n6128_, new_n6129_, new_n6130_,
    new_n6131_, new_n6132_, new_n6133_, new_n6134_, new_n6135_, new_n6136_,
    new_n6137_, new_n6138_, new_n6139_, new_n6140_, new_n6141_, new_n6142_,
    new_n6143_, new_n6144_, new_n6145_, new_n6146_, new_n6147_, new_n6148_,
    new_n6149_, new_n6150_, new_n6151_, new_n6152_, new_n6153_, new_n6154_,
    new_n6155_, new_n6156_, new_n6157_, new_n6158_, new_n6159_, new_n6160_,
    new_n6161_, new_n6162_, new_n6163_, new_n6164_, new_n6165_, new_n6166_,
    new_n6167_, new_n6168_, new_n6169_, new_n6170_, new_n6171_, new_n6172_,
    new_n6173_, new_n6174_, new_n6175_, new_n6176_, new_n6177_, new_n6178_,
    new_n6179_, new_n6180_, new_n6181_, new_n6182_, new_n6183_, new_n6184_,
    new_n6185_, new_n6186_, new_n6187_, new_n6188_, new_n6189_, new_n6190_,
    new_n6191_, new_n6192_, new_n6193_, new_n6194_, new_n6195_, new_n6196_,
    new_n6197_, new_n6198_, new_n6199_, new_n6200_, new_n6201_, new_n6202_,
    new_n6203_, new_n6204_, new_n6205_, new_n6206_, new_n6207_, new_n6208_,
    new_n6209_, new_n6210_, new_n6211_, new_n6212_, new_n6213_, new_n6214_,
    new_n6215_, new_n6216_, new_n6217_, new_n6218_, new_n6219_, new_n6220_,
    new_n6221_, new_n6222_, new_n6223_, new_n6224_, new_n6225_, new_n6226_,
    new_n6227_, new_n6228_, new_n6229_, new_n6230_, new_n6231_, new_n6232_,
    new_n6233_, new_n6234_, new_n6235_, new_n6236_, new_n6237_, new_n6238_,
    new_n6239_, new_n6240_, new_n6241_, new_n6242_, new_n6243_, new_n6244_,
    new_n6245_, new_n6246_, new_n6247_, new_n6248_, new_n6249_, new_n6250_,
    new_n6251_, new_n6252_, new_n6253_, new_n6254_, new_n6255_, new_n6256_,
    new_n6257_, new_n6258_, new_n6259_, new_n6260_, new_n6261_, new_n6262_,
    new_n6263_, new_n6264_, new_n6265_, new_n6266_, new_n6267_, new_n6268_,
    new_n6269_, new_n6270_, new_n6271_, new_n6272_, new_n6273_, new_n6274_,
    new_n6275_, new_n6276_, new_n6277_, new_n6278_, new_n6279_, new_n6280_,
    new_n6281_, new_n6282_, new_n6283_, new_n6284_, new_n6285_, new_n6286_,
    new_n6287_, new_n6288_, new_n6289_, new_n6290_, new_n6291_, new_n6292_,
    new_n6293_, new_n6294_, new_n6295_, new_n6296_, new_n6297_, new_n6298_,
    new_n6299_, new_n6300_, new_n6301_, new_n6302_, new_n6303_, new_n6304_,
    new_n6305_, new_n6306_, new_n6307_, new_n6308_, new_n6309_, new_n6310_,
    new_n6311_, new_n6312_, new_n6313_, new_n6314_, new_n6315_, new_n6316_,
    new_n6317_, new_n6318_, new_n6319_, new_n6320_, new_n6321_, new_n6322_,
    new_n6323_, new_n6324_, new_n6325_, new_n6326_, new_n6327_, new_n6328_,
    new_n6329_, new_n6330_, new_n6331_, new_n6332_, new_n6333_, new_n6334_,
    new_n6335_, new_n6336_, new_n6337_, new_n6338_, new_n6339_, new_n6340_,
    new_n6341_, new_n6342_, new_n6343_, new_n6344_, new_n6345_, new_n6346_,
    new_n6347_, new_n6348_, new_n6349_, new_n6350_, new_n6351_, new_n6352_,
    new_n6353_, new_n6354_, new_n6355_, new_n6356_, new_n6357_, new_n6358_,
    new_n6359_, new_n6360_, new_n6361_, new_n6362_, new_n6363_, new_n6364_,
    new_n6365_, new_n6366_, new_n6367_, new_n6368_, new_n6369_, new_n6370_,
    new_n6371_, new_n6372_, new_n6373_, new_n6374_, new_n6375_, new_n6376_,
    new_n6377_, new_n6378_, new_n6379_, new_n6380_, new_n6381_, new_n6382_,
    new_n6383_, new_n6384_, new_n6385_, new_n6386_, new_n6387_, new_n6388_,
    new_n6389_, new_n6390_, new_n6391_, new_n6392_, new_n6393_, new_n6394_,
    new_n6395_, new_n6396_, new_n6397_, new_n6398_, new_n6399_, new_n6400_,
    new_n6401_, new_n6402_, new_n6403_, new_n6404_, new_n6405_, new_n6406_,
    new_n6407_, new_n6408_, new_n6409_, new_n6410_, new_n6411_, new_n6412_,
    new_n6413_, new_n6414_, new_n6415_, new_n6416_, new_n6417_, new_n6418_,
    new_n6419_, new_n6420_, new_n6421_, new_n6422_, new_n6423_, new_n6424_,
    new_n6425_, new_n6426_, new_n6427_, new_n6428_, new_n6429_, new_n6430_,
    new_n6431_, new_n6432_, new_n6433_, new_n6434_, new_n6435_, new_n6436_,
    new_n6437_, new_n6438_, new_n6439_, new_n6440_, new_n6441_, new_n6442_,
    new_n6443_, new_n6444_, new_n6445_, new_n6446_, new_n6447_, new_n6448_,
    new_n6449_, new_n6450_, new_n6451_, new_n6452_, new_n6453_, new_n6454_,
    new_n6455_, new_n6456_, new_n6457_, new_n6458_, new_n6459_, new_n6460_,
    new_n6461_, new_n6462_, new_n6463_, new_n6464_, new_n6465_, new_n6466_,
    new_n6467_, new_n6468_, new_n6469_, new_n6470_, new_n6471_, new_n6472_,
    new_n6473_, new_n6474_, new_n6475_, new_n6476_, new_n6477_, new_n6478_,
    new_n6479_, new_n6480_, new_n6481_, new_n6482_, new_n6483_, new_n6484_,
    new_n6485_, new_n6486_, new_n6487_, new_n6488_, new_n6489_, new_n6490_,
    new_n6491_, new_n6492_, new_n6493_, new_n6494_, new_n6495_, new_n6496_,
    new_n6497_, new_n6498_, new_n6499_, new_n6500_, new_n6501_, new_n6502_,
    new_n6503_, new_n6504_, new_n6505_, new_n6506_, new_n6507_, new_n6508_,
    new_n6509_, new_n6510_, new_n6511_, new_n6512_, new_n6513_, new_n6514_,
    new_n6515_, new_n6516_, new_n6517_, new_n6518_, new_n6519_, new_n6520_,
    new_n6521_, new_n6522_, new_n6523_, new_n6524_, new_n6525_, new_n6526_,
    new_n6527_, new_n6528_, new_n6529_, new_n6530_, new_n6531_, new_n6532_,
    new_n6533_, new_n6534_, new_n6535_, new_n6536_, new_n6537_, new_n6538_,
    new_n6539_, new_n6540_, new_n6541_, new_n6542_, new_n6543_, new_n6544_,
    new_n6545_, new_n6546_, new_n6547_, new_n6548_, new_n6549_, new_n6550_,
    new_n6551_, new_n6552_, new_n6553_, new_n6554_, new_n6555_, new_n6556_,
    new_n6557_, new_n6558_, new_n6559_, new_n6560_, new_n6561_, new_n6562_,
    new_n6563_, new_n6564_, new_n6565_, new_n6566_, new_n6567_, new_n6568_,
    new_n6569_, new_n6570_, new_n6571_, new_n6572_, new_n6573_, new_n6574_,
    new_n6575_, new_n6576_, new_n6577_, new_n6578_, new_n6579_, new_n6580_,
    new_n6581_, new_n6582_, new_n6583_, new_n6584_, new_n6585_, new_n6586_,
    new_n6587_, new_n6588_, new_n6589_, new_n6590_, new_n6591_, new_n6592_,
    new_n6593_, new_n6594_, new_n6595_, new_n6596_, new_n6597_, new_n6598_,
    new_n6599_, new_n6600_, new_n6601_, new_n6602_, new_n6603_, new_n6604_,
    new_n6605_, new_n6606_, new_n6607_, new_n6608_, new_n6609_, new_n6610_,
    new_n6611_, new_n6612_, new_n6613_, new_n6614_, new_n6615_, new_n6616_,
    new_n6617_, new_n6618_, new_n6619_, new_n6620_, new_n6621_, new_n6622_,
    new_n6623_, new_n6624_, new_n6625_, new_n6626_, new_n6627_, new_n6628_,
    new_n6629_, new_n6630_, new_n6631_, new_n6632_, new_n6633_, new_n6634_,
    new_n6635_, new_n6636_, new_n6637_, new_n6638_, new_n6639_, new_n6640_,
    new_n6641_, new_n6642_, new_n6643_, new_n6644_, new_n6645_, new_n6646_,
    new_n6647_, new_n6648_, new_n6649_, new_n6650_, new_n6651_, new_n6652_,
    new_n6653_, new_n6654_, new_n6655_, new_n6656_, new_n6657_, new_n6658_,
    new_n6659_, new_n6660_, new_n6661_, new_n6662_, new_n6663_, new_n6664_,
    new_n6665_, new_n6666_, new_n6667_, new_n6668_, new_n6669_, new_n6670_,
    new_n6671_, new_n6672_, new_n6673_, new_n6674_, new_n6675_, new_n6676_,
    new_n6677_, new_n6678_, new_n6679_, new_n6680_, new_n6681_, new_n6682_,
    new_n6683_, new_n6684_, new_n6685_, new_n6686_, new_n6687_, new_n6688_,
    new_n6689_, new_n6690_, new_n6691_, new_n6692_, new_n6693_, new_n6694_,
    new_n6695_, new_n6696_, new_n6697_, new_n6698_, new_n6699_, new_n6700_,
    new_n6701_, new_n6702_, new_n6703_, new_n6704_, new_n6705_, new_n6706_,
    new_n6707_, new_n6708_, new_n6709_, new_n6710_, new_n6711_, new_n6712_,
    new_n6713_, new_n6714_, new_n6715_, new_n6716_, new_n6717_, new_n6718_,
    new_n6719_, new_n6720_, new_n6721_, new_n6722_, new_n6723_, new_n6724_,
    new_n6725_, new_n6726_, new_n6727_, new_n6728_, new_n6729_, new_n6730_,
    new_n6731_, new_n6732_, new_n6733_, new_n6734_, new_n6735_, new_n6736_,
    new_n6737_, new_n6738_, new_n6739_, new_n6740_, new_n6741_, new_n6742_,
    new_n6743_, new_n6744_, new_n6745_, new_n6746_, new_n6747_, new_n6748_,
    new_n6749_, new_n6750_, new_n6751_, new_n6752_, new_n6753_, new_n6754_,
    new_n6755_, new_n6756_, new_n6757_, new_n6758_, new_n6759_, new_n6760_,
    new_n6761_, new_n6762_, new_n6763_, new_n6764_, new_n6765_, new_n6766_,
    new_n6767_, new_n6768_, new_n6769_, new_n6770_, new_n6771_, new_n6772_,
    new_n6773_, new_n6774_, new_n6775_, new_n6776_, new_n6777_, new_n6778_,
    new_n6779_, new_n6780_, new_n6781_, new_n6782_, new_n6783_, new_n6784_,
    new_n6785_, new_n6786_, new_n6787_, new_n6788_, new_n6789_, new_n6790_,
    new_n6791_, new_n6792_, new_n6793_, new_n6794_, new_n6795_, new_n6796_,
    new_n6797_, new_n6798_, new_n6799_, new_n6800_, new_n6801_, new_n6802_,
    new_n6803_, new_n6804_, new_n6805_, new_n6806_, new_n6807_, new_n6808_,
    new_n6809_, new_n6810_, new_n6811_, new_n6812_, new_n6813_, new_n6814_,
    new_n6815_, new_n6816_, new_n6817_, new_n6818_, new_n6819_, new_n6820_,
    new_n6821_, new_n6822_, new_n6823_, new_n6824_, new_n6825_, new_n6826_,
    new_n6827_, new_n6828_, new_n6829_, new_n6830_, new_n6831_, new_n6832_,
    new_n6833_, new_n6834_, new_n6835_, new_n6836_, new_n6837_, new_n6838_,
    new_n6839_, new_n6840_, new_n6841_, new_n6842_, new_n6843_, new_n6844_,
    new_n6845_, new_n6846_, new_n6847_, new_n6848_, new_n6849_, new_n6850_,
    new_n6851_, new_n6852_, new_n6853_, new_n6854_, new_n6855_, new_n6856_,
    new_n6857_, new_n6858_, new_n6859_, new_n6860_, new_n6861_, new_n6862_,
    new_n6863_, new_n6864_, new_n6865_, new_n6866_, new_n6867_, new_n6868_,
    new_n6869_, new_n6870_, new_n6871_, new_n6872_, new_n6873_, new_n6874_,
    new_n6875_, new_n6876_, new_n6877_, new_n6878_, new_n6879_, new_n6880_,
    new_n6881_, new_n6882_, new_n6883_, new_n6884_, new_n6885_, new_n6886_,
    new_n6887_, new_n6888_, new_n6889_, new_n6890_, new_n6891_, new_n6892_,
    new_n6893_, new_n6894_, new_n6895_, new_n6896_, new_n6897_, new_n6898_,
    new_n6899_, new_n6900_, new_n6901_, new_n6902_, new_n6903_, new_n6904_,
    new_n6905_, new_n6906_, new_n6907_, new_n6908_, new_n6909_, new_n6910_,
    new_n6911_, new_n6912_, new_n6913_, new_n6914_, new_n6915_, new_n6916_,
    new_n6917_, new_n6918_, new_n6919_, new_n6920_, new_n6921_, new_n6922_,
    new_n6923_, new_n6924_, new_n6925_, new_n6926_, new_n6927_, new_n6928_,
    new_n6929_, new_n6930_, new_n6931_, new_n6932_, new_n6933_, new_n6934_,
    new_n6935_, new_n6936_, new_n6937_, new_n6938_, new_n6939_, new_n6940_,
    new_n6941_, new_n6942_, new_n6943_, new_n6944_, new_n6945_, new_n6946_,
    new_n6947_, new_n6948_, new_n6949_, new_n6950_, new_n6951_, new_n6952_,
    new_n6953_, new_n6954_, new_n6955_, new_n6956_, new_n6957_, new_n6958_,
    new_n6959_, new_n6960_, new_n6961_, new_n6962_, new_n6963_, new_n6964_,
    new_n6965_, new_n6966_, new_n6967_, new_n6968_, new_n6969_, new_n6970_,
    new_n6971_, new_n6972_, new_n6973_, new_n6974_, new_n6975_, new_n6976_,
    new_n6977_, new_n6978_, new_n6979_, new_n6980_, new_n6981_, new_n6982_,
    new_n6983_, new_n6984_, new_n6985_, new_n6986_, new_n6987_, new_n6988_,
    new_n6989_, new_n6990_, new_n6991_, new_n6992_, new_n6993_, new_n6994_,
    new_n6995_, new_n6996_, new_n6997_, new_n6998_, new_n6999_, new_n7000_,
    new_n7001_, new_n7002_, new_n7003_, new_n7004_, new_n7005_, new_n7006_,
    new_n7007_, new_n7008_, new_n7009_, new_n7010_, new_n7011_, new_n7012_,
    new_n7013_, new_n7014_, new_n7015_, new_n7016_, new_n7017_, new_n7018_,
    new_n7019_, new_n7020_, new_n7021_, new_n7022_, new_n7023_, new_n7024_,
    new_n7025_, new_n7026_, new_n7027_, new_n7028_, new_n7029_, new_n7030_,
    new_n7031_, new_n7032_, new_n7033_, new_n7034_, new_n7035_, new_n7036_,
    new_n7037_, new_n7038_, new_n7039_, new_n7040_, new_n7041_, new_n7042_,
    new_n7043_, new_n7044_, new_n7045_, new_n7046_, new_n7047_, new_n7048_,
    new_n7049_, new_n7050_, new_n7051_, new_n7052_, new_n7053_, new_n7054_,
    new_n7055_, new_n7056_, new_n7057_, new_n7058_, new_n7059_, new_n7060_,
    new_n7061_, new_n7062_, new_n7063_, new_n7064_, new_n7065_, new_n7066_,
    new_n7067_, new_n7068_, new_n7069_, new_n7070_, new_n7071_, new_n7072_,
    new_n7073_, new_n7074_, new_n7075_, new_n7076_, new_n7077_, new_n7078_,
    new_n7079_, new_n7080_, new_n7081_, new_n7082_, new_n7083_, new_n7084_,
    new_n7085_, new_n7086_, new_n7087_, new_n7088_, new_n7089_, new_n7090_,
    new_n7091_, new_n7092_, new_n7093_, new_n7094_, new_n7095_, new_n7096_,
    new_n7097_, new_n7098_, new_n7099_, new_n7100_, new_n7101_, new_n7102_,
    new_n7103_, new_n7104_, new_n7105_, new_n7106_, new_n7107_, new_n7108_,
    new_n7109_, new_n7110_, new_n7111_, new_n7112_, new_n7113_, new_n7114_,
    new_n7115_, new_n7116_, new_n7117_, new_n7118_, new_n7119_, new_n7120_,
    new_n7121_, new_n7122_, new_n7123_, new_n7124_, new_n7125_, new_n7126_,
    new_n7127_, new_n7128_, new_n7129_, new_n7130_, new_n7131_, new_n7132_,
    new_n7133_, new_n7134_, new_n7135_, new_n7136_, new_n7137_, new_n7138_,
    new_n7139_, new_n7140_, new_n7141_, new_n7142_, new_n7143_, new_n7144_,
    new_n7145_, new_n7146_, new_n7147_, new_n7148_, new_n7149_, new_n7150_,
    new_n7151_, new_n7152_, new_n7153_, new_n7154_, new_n7155_, new_n7156_,
    new_n7157_, new_n7158_, new_n7159_, new_n7160_, new_n7161_, new_n7162_,
    new_n7163_, new_n7164_, new_n7165_, new_n7166_, new_n7167_, new_n7168_,
    new_n7169_, new_n7170_, new_n7171_, new_n7172_, new_n7173_, new_n7174_,
    new_n7175_, new_n7176_, new_n7177_, new_n7178_, new_n7179_, new_n7180_,
    new_n7181_, new_n7182_, new_n7183_, new_n7184_, new_n7185_, new_n7186_,
    new_n7187_, new_n7188_, new_n7189_, new_n7190_, new_n7191_, new_n7192_,
    new_n7193_, new_n7194_, new_n7195_, new_n7196_, new_n7197_, new_n7198_,
    new_n7199_, new_n7200_, new_n7201_, new_n7202_, new_n7203_, new_n7204_,
    new_n7205_, new_n7206_, new_n7207_, new_n7208_, new_n7209_, new_n7210_,
    new_n7211_, new_n7212_, new_n7213_, new_n7214_, new_n7215_, new_n7216_,
    new_n7217_, new_n7218_, new_n7219_, new_n7220_, new_n7221_, new_n7222_,
    new_n7223_, new_n7224_, new_n7225_, new_n7226_, new_n7227_, new_n7228_,
    new_n7229_, new_n7230_, new_n7231_, new_n7232_, new_n7233_, new_n7234_,
    new_n7235_, new_n7236_, new_n7237_, new_n7238_, new_n7239_, new_n7240_,
    new_n7241_, new_n7242_, new_n7243_, new_n7244_, new_n7245_, new_n7246_,
    new_n7247_, new_n7248_, new_n7249_, new_n7250_, new_n7251_, new_n7252_,
    new_n7253_, new_n7254_, new_n7255_, new_n7256_, new_n7257_, new_n7258_,
    new_n7259_, new_n7260_, new_n7261_, new_n7262_, new_n7263_, new_n7264_,
    new_n7265_, new_n7266_, new_n7267_, new_n7268_, new_n7269_, new_n7270_,
    new_n7271_, new_n7272_, new_n7273_, new_n7274_, new_n7275_, new_n7276_,
    new_n7277_, new_n7278_, new_n7279_, new_n7280_, new_n7281_, new_n7282_,
    new_n7283_, new_n7284_, new_n7285_, new_n7286_, new_n7287_, new_n7288_,
    new_n7289_, new_n7290_, new_n7291_, new_n7292_, new_n7293_, new_n7294_,
    new_n7295_, new_n7296_, new_n7297_, new_n7298_, new_n7299_, new_n7300_,
    new_n7301_, new_n7302_, new_n7303_, new_n7304_, new_n7305_, new_n7306_,
    new_n7307_, new_n7308_, new_n7309_, new_n7310_, new_n7311_, new_n7312_,
    new_n7313_, new_n7314_, new_n7315_, new_n7316_, new_n7317_, new_n7318_,
    new_n7319_, new_n7320_, new_n7321_, new_n7322_, new_n7323_, new_n7324_,
    new_n7325_, new_n7326_, new_n7327_, new_n7328_, new_n7329_, new_n7330_,
    new_n7331_, new_n7332_, new_n7333_, new_n7334_, new_n7335_, new_n7336_,
    new_n7337_, new_n7338_, new_n7339_, new_n7340_, new_n7341_, new_n7342_,
    new_n7343_, new_n7344_, new_n7345_, new_n7346_, new_n7347_, new_n7348_,
    new_n7349_, new_n7350_, new_n7351_, new_n7352_, new_n7353_, new_n7354_,
    new_n7355_, new_n7356_, new_n7357_, new_n7358_, new_n7359_, new_n7360_,
    new_n7361_, new_n7362_, new_n7363_, new_n7364_, new_n7365_, new_n7366_,
    new_n7367_, new_n7368_, new_n7369_, new_n7370_, new_n7371_, new_n7372_,
    new_n7373_, new_n7374_, new_n7375_, new_n7376_, new_n7377_, new_n7378_,
    new_n7379_, new_n7380_, new_n7381_, new_n7382_, new_n7383_, new_n7384_,
    new_n7385_, new_n7386_, new_n7387_, new_n7388_, new_n7389_, new_n7390_,
    new_n7391_, new_n7392_, new_n7393_, new_n7394_, new_n7395_, new_n7396_,
    new_n7397_, new_n7398_, new_n7399_, new_n7400_, new_n7401_, new_n7402_,
    new_n7403_, new_n7404_, new_n7405_, new_n7406_, new_n7407_, new_n7408_,
    new_n7409_, new_n7410_, new_n7411_, new_n7412_, new_n7413_, new_n7414_,
    new_n7415_, new_n7416_, new_n7417_, new_n7418_, new_n7419_, new_n7420_,
    new_n7421_, new_n7422_, new_n7423_, new_n7424_, new_n7425_, new_n7426_,
    new_n7427_, new_n7428_, new_n7429_, new_n7430_, new_n7431_, new_n7432_,
    new_n7433_, new_n7434_, new_n7435_, new_n7436_, new_n7437_, new_n7438_,
    new_n7439_, new_n7440_, new_n7441_, new_n7442_, new_n7443_, new_n7444_,
    new_n7445_, new_n7446_, new_n7447_, new_n7448_, new_n7449_, new_n7450_,
    new_n7451_, new_n7452_, new_n7453_, new_n7454_, new_n7455_, new_n7456_,
    new_n7457_, new_n7458_, new_n7459_, new_n7460_, new_n7461_, new_n7462_,
    new_n7463_, new_n7464_, new_n7465_, new_n7466_, new_n7467_, new_n7468_,
    new_n7469_, new_n7470_, new_n7471_, new_n7472_, new_n7473_, new_n7474_,
    new_n7475_, new_n7476_, new_n7477_, new_n7478_, new_n7479_, new_n7480_,
    new_n7481_, new_n7482_, new_n7483_, new_n7484_, new_n7485_, new_n7486_,
    new_n7487_, new_n7488_, new_n7489_, new_n7490_, new_n7491_, new_n7492_,
    new_n7493_, new_n7494_, new_n7495_, new_n7496_, new_n7497_, new_n7498_,
    new_n7499_, new_n7500_, new_n7501_, new_n7502_, new_n7503_, new_n7504_,
    new_n7505_, new_n7506_, new_n7507_, new_n7508_, new_n7509_, new_n7510_,
    new_n7511_, new_n7512_, new_n7513_, new_n7514_, new_n7515_, new_n7516_,
    new_n7517_, new_n7518_, new_n7519_, new_n7520_, new_n7521_, new_n7522_,
    new_n7523_, new_n7524_, new_n7525_, new_n7526_, new_n7527_, new_n7528_,
    new_n7529_, new_n7530_, new_n7531_, new_n7532_, new_n7533_, new_n7534_,
    new_n7535_, new_n7536_, new_n7537_, new_n7538_, new_n7539_, new_n7540_,
    new_n7541_, new_n7542_, new_n7543_, new_n7544_, new_n7545_, new_n7546_,
    new_n7547_, new_n7548_, new_n7549_, new_n7550_, new_n7551_, new_n7552_,
    new_n7553_, new_n7554_, new_n7555_, new_n7556_, new_n7557_, new_n7558_,
    new_n7559_, new_n7560_, new_n7561_, new_n7562_, new_n7563_, new_n7564_,
    new_n7565_, new_n7566_, new_n7567_, new_n7568_, new_n7569_, new_n7570_,
    new_n7571_, new_n7572_, new_n7573_, new_n7574_, new_n7575_, new_n7576_,
    new_n7577_, new_n7578_, new_n7579_, new_n7580_, new_n7581_, new_n7582_,
    new_n7583_, new_n7584_, new_n7585_, new_n7586_, new_n7587_, new_n7588_,
    new_n7589_, new_n7590_, new_n7591_, new_n7592_, new_n7593_, new_n7594_,
    new_n7595_, new_n7596_, new_n7597_, new_n7598_, new_n7599_, new_n7600_,
    new_n7601_, new_n7602_, new_n7603_, new_n7604_, new_n7605_, new_n7606_,
    new_n7607_, new_n7608_, new_n7609_, new_n7610_, new_n7611_, new_n7612_,
    new_n7613_, new_n7614_, new_n7615_, new_n7616_, new_n7617_, new_n7618_,
    new_n7619_, new_n7620_, new_n7621_, new_n7622_, new_n7623_, new_n7624_,
    new_n7625_, new_n7626_, new_n7627_, new_n7628_, new_n7629_, new_n7630_,
    new_n7631_, new_n7632_, new_n7633_, new_n7634_, new_n7635_, new_n7636_,
    new_n7637_, new_n7638_, new_n7639_, new_n7640_, new_n7641_, new_n7642_,
    new_n7643_, new_n7644_, new_n7645_, new_n7646_, new_n7647_, new_n7648_,
    new_n7649_, new_n7650_, new_n7651_, new_n7652_, new_n7653_, new_n7654_,
    new_n7655_, new_n7656_, new_n7657_, new_n7658_, new_n7659_, new_n7660_,
    new_n7661_, new_n7662_, new_n7663_, new_n7664_, new_n7665_, new_n7666_,
    new_n7667_, new_n7668_, new_n7669_, new_n7670_, new_n7671_, new_n7672_,
    new_n7673_, new_n7674_, new_n7675_, new_n7676_, new_n7677_, new_n7678_,
    new_n7679_, new_n7680_, new_n7681_, new_n7682_, new_n7683_, new_n7684_,
    new_n7685_, new_n7686_, new_n7687_, new_n7688_, new_n7689_, new_n7690_,
    new_n7691_, new_n7692_, new_n7693_, new_n7694_, new_n7695_, new_n7696_,
    new_n7697_, new_n7698_, new_n7699_, new_n7700_, new_n7701_, new_n7702_,
    new_n7703_, new_n7704_, new_n7705_, new_n7706_, new_n7707_, new_n7708_,
    new_n7709_, new_n7710_, new_n7711_, new_n7712_, new_n7713_, new_n7714_,
    new_n7715_, new_n7716_, new_n7717_, new_n7718_, new_n7719_, new_n7720_,
    new_n7721_, new_n7722_, new_n7723_, new_n7724_, new_n7725_, new_n7726_,
    new_n7727_, new_n7728_, new_n7729_, new_n7730_, new_n7731_, new_n7732_,
    new_n7733_, new_n7734_, new_n7735_, new_n7736_, new_n7737_, new_n7738_,
    new_n7739_, new_n7740_, new_n7741_, new_n7742_, new_n7743_, new_n7744_,
    new_n7745_, new_n7746_, new_n7747_, new_n7748_, new_n7749_, new_n7750_,
    new_n7751_, new_n7752_, new_n7753_, new_n7754_, new_n7755_, new_n7756_,
    new_n7757_, new_n7758_, new_n7759_, new_n7760_, new_n7761_, new_n7762_,
    new_n7763_, new_n7764_, new_n7765_, new_n7766_, new_n7767_, new_n7768_,
    new_n7769_, new_n7770_, new_n7771_, new_n7772_, new_n7773_, new_n7774_,
    new_n7775_, new_n7776_, new_n7777_, new_n7778_, new_n7779_, new_n7780_,
    new_n7781_, new_n7782_, new_n7783_, new_n7784_, new_n7785_, new_n7786_,
    new_n7787_, new_n7788_, new_n7789_, new_n7790_, new_n7791_, new_n7792_,
    new_n7793_, new_n7794_, new_n7795_, new_n7796_, new_n7797_, new_n7798_,
    new_n7799_, new_n7800_, new_n7801_, new_n7802_, new_n7803_, new_n7804_,
    new_n7805_, new_n7806_, new_n7807_, new_n7808_, new_n7809_, new_n7810_,
    new_n7811_, new_n7812_, new_n7813_, new_n7814_, new_n7815_, new_n7816_,
    new_n7817_, new_n7818_, new_n7819_, new_n7820_, new_n7821_, new_n7822_,
    new_n7823_, new_n7824_, new_n7825_, new_n7826_, new_n7827_, new_n7828_,
    new_n7829_, new_n7830_, new_n7831_, new_n7832_, new_n7833_, new_n7834_,
    new_n7835_, new_n7836_, new_n7837_, new_n7838_, new_n7839_, new_n7840_,
    new_n7841_, new_n7842_, new_n7843_, new_n7844_, new_n7845_, new_n7846_,
    new_n7847_, new_n7848_, new_n7849_, new_n7850_, new_n7851_, new_n7852_,
    new_n7853_, new_n7854_, new_n7855_, new_n7856_, new_n7857_, new_n7858_,
    new_n7859_, new_n7860_, new_n7861_, new_n7862_, new_n7863_, new_n7864_,
    new_n7865_, new_n7866_, new_n7867_, new_n7868_, new_n7869_, new_n7870_,
    new_n7871_, new_n7872_, new_n7873_, new_n7874_, new_n7875_, new_n7876_,
    new_n7877_, new_n7878_, new_n7879_, new_n7880_, new_n7881_, new_n7882_,
    new_n7883_, new_n7884_, new_n7885_, new_n7886_, new_n7887_, new_n7888_,
    new_n7889_, new_n7890_, new_n7891_, new_n7892_, new_n7893_, new_n7894_,
    new_n7895_, new_n7896_, new_n7897_, new_n7898_, new_n7899_, new_n7900_,
    new_n7901_, new_n7902_, new_n7903_, new_n7904_, new_n7905_, new_n7906_,
    new_n7907_, new_n7908_, new_n7909_, new_n7910_, new_n7911_, new_n7912_,
    new_n7913_, new_n7914_, new_n7915_, new_n7916_, new_n7917_, new_n7918_,
    new_n7919_, new_n7920_, new_n7921_, new_n7922_, new_n7923_, new_n7924_,
    new_n7925_, new_n7926_, new_n7927_, new_n7928_, new_n7929_, new_n7930_,
    new_n7931_, new_n7932_, new_n7933_, new_n7934_, new_n7935_, new_n7936_,
    new_n7937_, new_n7938_, new_n7939_, new_n7940_, new_n7941_, new_n7942_,
    new_n7943_, new_n7944_, new_n7945_, new_n7946_, new_n7947_, new_n7948_,
    new_n7949_, new_n7950_, new_n7951_, new_n7952_, new_n7953_, new_n7954_,
    new_n7955_, new_n7956_, new_n7957_, new_n7958_, new_n7959_, new_n7960_,
    new_n7961_, new_n7962_, new_n7963_, new_n7964_, new_n7965_, new_n7966_,
    new_n7967_, new_n7968_, new_n7969_, new_n7970_, new_n7971_, new_n7972_,
    new_n7973_, new_n7974_, new_n7975_, new_n7976_, new_n7977_, new_n7978_,
    new_n7979_, new_n7980_, new_n7981_, new_n7982_, new_n7983_, new_n7984_,
    new_n7985_, new_n7986_, new_n7987_, new_n7988_, new_n7989_, new_n7990_,
    new_n7991_, new_n7992_, new_n7993_, new_n7994_, new_n7995_, new_n7996_,
    new_n7997_, new_n7998_, new_n7999_, new_n8000_, new_n8001_, new_n8002_,
    new_n8003_, new_n8004_, new_n8005_, new_n8006_, new_n8007_, new_n8008_,
    new_n8009_, new_n8010_, new_n8011_, new_n8012_, new_n8013_, new_n8014_,
    new_n8015_, new_n8016_, new_n8017_, new_n8018_, new_n8019_, new_n8020_,
    new_n8021_, new_n8022_, new_n8023_, new_n8024_, new_n8025_, new_n8026_,
    new_n8027_, new_n8028_, new_n8029_, new_n8030_, new_n8031_, new_n8032_,
    new_n8033_, new_n8034_, new_n8035_, new_n8036_, new_n8037_, new_n8038_,
    new_n8039_, new_n8040_, new_n8041_, new_n8042_, new_n8043_, new_n8044_,
    new_n8045_, new_n8046_, new_n8047_, new_n8048_, new_n8049_, new_n8050_,
    new_n8051_, new_n8052_, new_n8053_, new_n8054_, new_n8055_, new_n8056_,
    new_n8057_, new_n8058_, new_n8059_, new_n8060_, new_n8061_, new_n8062_,
    new_n8063_, new_n8064_, new_n8065_, new_n8066_, new_n8067_, new_n8068_,
    new_n8069_, new_n8070_, new_n8071_, new_n8072_, new_n8073_, new_n8074_,
    new_n8075_, new_n8076_, new_n8077_, new_n8078_, new_n8079_, new_n8080_,
    new_n8081_, new_n8082_, new_n8083_, new_n8084_, new_n8085_, new_n8086_,
    new_n8087_, new_n8088_, new_n8089_, new_n8090_, new_n8091_, new_n8092_,
    new_n8093_, new_n8094_, new_n8095_, new_n8096_, new_n8097_, new_n8098_,
    new_n8099_, new_n8100_, new_n8101_, new_n8102_, new_n8103_, new_n8104_,
    new_n8105_, new_n8106_, new_n8107_, new_n8108_, new_n8109_, new_n8110_,
    new_n8111_, new_n8112_, new_n8113_, new_n8114_, new_n8115_, new_n8116_,
    new_n8117_, new_n8118_, new_n8119_, new_n8120_, new_n8121_, new_n8122_,
    new_n8123_, new_n8124_, new_n8125_, new_n8126_, new_n8127_, new_n8128_,
    new_n8129_, new_n8130_, new_n8131_, new_n8132_, new_n8133_, new_n8134_,
    new_n8135_, new_n8136_, new_n8137_, new_n8138_, new_n8139_, new_n8140_,
    new_n8141_, new_n8142_, new_n8143_, new_n8144_, new_n8145_, new_n8146_,
    new_n8147_, new_n8148_, new_n8149_, new_n8150_, new_n8151_, new_n8152_,
    new_n8153_, new_n8154_, new_n8155_, new_n8156_, new_n8157_, new_n8158_,
    new_n8159_, new_n8160_, new_n8161_, new_n8162_, new_n8163_, new_n8164_,
    new_n8165_, new_n8166_, new_n8167_, new_n8168_, new_n8169_, new_n8170_,
    new_n8171_, new_n8172_, new_n8173_, new_n8174_, new_n8175_, new_n8176_,
    new_n8177_, new_n8178_, new_n8179_, new_n8180_, new_n8181_, new_n8182_,
    new_n8183_, new_n8184_, new_n8185_, new_n8186_, new_n8187_, new_n8188_,
    new_n8189_, new_n8190_, new_n8191_, new_n8192_, new_n8193_, new_n8194_,
    new_n8195_, new_n8196_, new_n8197_, new_n8198_, new_n8199_, new_n8200_,
    new_n8201_, new_n8202_, new_n8203_, new_n8204_, new_n8205_, new_n8206_,
    new_n8207_, new_n8208_, new_n8209_, new_n8210_, new_n8211_, new_n8212_,
    new_n8213_, new_n8214_, new_n8215_, new_n8216_, new_n8217_, new_n8218_,
    new_n8219_, new_n8220_, new_n8221_, new_n8222_, new_n8223_, new_n8224_,
    new_n8225_, new_n8226_, new_n8227_, new_n8228_, new_n8229_, new_n8230_,
    new_n8231_, new_n8232_, new_n8233_, new_n8234_, new_n8235_, new_n8236_,
    new_n8237_, new_n8238_, new_n8239_, new_n8240_, new_n8241_, new_n8242_,
    new_n8243_, new_n8244_, new_n8245_, new_n8246_, new_n8247_, new_n8248_,
    new_n8249_, new_n8250_, new_n8251_, new_n8252_, new_n8253_, new_n8254_,
    new_n8255_, new_n8256_, new_n8257_, new_n8258_, new_n8259_, new_n8260_,
    new_n8261_, new_n8262_, new_n8263_, new_n8264_, new_n8265_, new_n8266_,
    new_n8267_, new_n8268_, new_n8269_, new_n8270_, new_n8271_, new_n8272_,
    new_n8273_, new_n8274_, new_n8275_, new_n8276_, new_n8277_, new_n8278_,
    new_n8279_, new_n8280_, new_n8281_, new_n8282_, new_n8283_, new_n8284_,
    new_n8285_, new_n8286_, new_n8287_, new_n8288_, new_n8289_, new_n8290_,
    new_n8291_, new_n8292_, new_n8293_, new_n8294_, new_n8295_, new_n8296_,
    new_n8297_, new_n8298_, new_n8299_, new_n8300_, new_n8301_, new_n8302_,
    new_n8303_, new_n8304_, new_n8305_, new_n8306_, new_n8307_, new_n8308_,
    new_n8309_, new_n8310_, new_n8311_, new_n8312_, new_n8313_, new_n8314_,
    new_n8315_, new_n8316_, new_n8317_, new_n8318_, new_n8319_, new_n8320_,
    new_n8321_, new_n8322_, new_n8323_, new_n8324_, new_n8325_, new_n8326_,
    new_n8327_, new_n8328_, new_n8329_, new_n8330_, new_n8331_, new_n8332_,
    new_n8333_, new_n8334_, new_n8335_, new_n8336_, new_n8337_, new_n8338_,
    new_n8339_, new_n8340_, new_n8341_, new_n8342_, new_n8343_, new_n8344_,
    new_n8345_, new_n8346_, new_n8347_, new_n8348_, new_n8349_, new_n8350_,
    new_n8351_, new_n8352_, new_n8353_, new_n8354_, new_n8355_, new_n8356_,
    new_n8357_, new_n8358_, new_n8359_, new_n8360_, new_n8361_, new_n8362_,
    new_n8363_, new_n8364_, new_n8365_, new_n8366_, new_n8367_, new_n8368_,
    new_n8369_, new_n8370_, new_n8371_, new_n8372_, new_n8373_, new_n8374_,
    new_n8375_, new_n8376_, new_n8377_, new_n8378_, new_n8379_, new_n8380_,
    new_n8381_, new_n8382_, new_n8383_, new_n8384_, new_n8385_, new_n8386_,
    new_n8387_, new_n8388_, new_n8389_, new_n8390_, new_n8391_, new_n8392_,
    new_n8393_, new_n8394_, new_n8395_, new_n8396_, new_n8397_, new_n8398_,
    new_n8399_, new_n8400_, new_n8401_, new_n8402_, new_n8403_, new_n8404_,
    new_n8405_, new_n8406_, new_n8407_, new_n8408_, new_n8409_, new_n8410_,
    new_n8411_, new_n8412_, new_n8413_, new_n8414_, new_n8415_, new_n8416_,
    new_n8417_, new_n8418_, new_n8419_, new_n8420_, new_n8421_, new_n8422_,
    new_n8423_, new_n8424_, new_n8425_, new_n8426_, new_n8427_, new_n8428_,
    new_n8429_, new_n8430_, new_n8431_, new_n8432_, new_n8433_, new_n8434_,
    new_n8435_, new_n8436_, new_n8437_, new_n8438_, new_n8439_, new_n8440_,
    new_n8441_, new_n8442_, new_n8443_, new_n8444_, new_n8445_, new_n8446_,
    new_n8447_, new_n8448_, new_n8449_, new_n8450_, new_n8451_, new_n8452_,
    new_n8453_, new_n8454_, new_n8455_, new_n8456_, new_n8457_, new_n8458_,
    new_n8459_, new_n8460_, new_n8461_, new_n8462_, new_n8463_, new_n8464_,
    new_n8465_, new_n8466_, new_n8467_, new_n8468_, new_n8469_, new_n8470_,
    new_n8471_, new_n8472_, new_n8473_, new_n8474_, new_n8475_, new_n8476_,
    new_n8477_, new_n8478_, new_n8479_, new_n8480_, new_n8481_, new_n8482_,
    new_n8483_, new_n8484_, new_n8485_, new_n8486_, new_n8487_, new_n8488_,
    new_n8489_, new_n8490_, new_n8491_, new_n8492_, new_n8493_, new_n8494_,
    new_n8495_, new_n8496_, new_n8497_, new_n8498_, new_n8499_, new_n8500_,
    new_n8501_, new_n8502_, new_n8503_, new_n8504_, new_n8505_, new_n8506_,
    new_n8507_, new_n8508_, new_n8509_, new_n8510_, new_n8511_, new_n8512_,
    new_n8513_, new_n8514_, new_n8515_, new_n8516_, new_n8517_, new_n8518_,
    new_n8519_, new_n8520_, new_n8521_, new_n8522_, new_n8523_, new_n8524_,
    new_n8525_, new_n8526_, new_n8527_, new_n8528_, new_n8529_, new_n8530_,
    new_n8531_, new_n8532_, new_n8533_, new_n8534_, new_n8535_, new_n8536_,
    new_n8537_, new_n8538_, new_n8539_, new_n8540_, new_n8541_, new_n8542_,
    new_n8543_, new_n8544_, new_n8545_, new_n8546_, new_n8547_, new_n8548_,
    new_n8549_, new_n8550_, new_n8551_, new_n8552_, new_n8553_, new_n8554_,
    new_n8555_, new_n8556_, new_n8557_, new_n8558_, new_n8559_, new_n8560_,
    new_n8561_, new_n8562_, new_n8563_, new_n8564_, new_n8565_, new_n8566_,
    new_n8567_, new_n8568_, new_n8569_, new_n8570_, new_n8571_, new_n8572_,
    new_n8573_, new_n8574_, new_n8575_, new_n8576_, new_n8577_, new_n8578_,
    new_n8579_, new_n8580_, new_n8581_, new_n8582_, new_n8583_, new_n8584_,
    new_n8585_, new_n8586_, new_n8587_, new_n8588_, new_n8589_, new_n8590_,
    new_n8591_, new_n8592_, new_n8593_, new_n8594_, new_n8595_, new_n8596_,
    new_n8597_, new_n8598_, new_n8599_, new_n8600_, new_n8601_, new_n8602_,
    new_n8603_, new_n8604_, new_n8605_, new_n8606_, new_n8607_, new_n8608_,
    new_n8609_, new_n8610_, new_n8611_, new_n8612_, new_n8613_, new_n8614_,
    new_n8615_, new_n8616_, new_n8617_, new_n8618_, new_n8619_, new_n8620_,
    new_n8621_, new_n8622_, new_n8623_, new_n8624_, new_n8625_, new_n8626_,
    new_n8627_, new_n8628_, new_n8629_, new_n8630_, new_n8631_, new_n8632_,
    new_n8633_, new_n8634_, new_n8635_, new_n8636_, new_n8637_, new_n8638_,
    new_n8639_, new_n8640_, new_n8641_, new_n8642_, new_n8643_, new_n8644_,
    new_n8645_, new_n8646_, new_n8647_, new_n8648_, new_n8649_, new_n8650_,
    new_n8651_, new_n8652_, new_n8653_, new_n8654_, new_n8655_, new_n8656_,
    new_n8657_, new_n8658_, new_n8659_, new_n8660_, new_n8661_, new_n8662_,
    new_n8663_, new_n8664_, new_n8665_, new_n8666_, new_n8667_, new_n8668_,
    new_n8669_, new_n8670_, new_n8671_, new_n8672_, new_n8673_, new_n8674_,
    new_n8675_, new_n8676_, new_n8677_, new_n8678_, new_n8679_, new_n8680_,
    new_n8681_, new_n8682_, new_n8683_, new_n8684_, new_n8685_, new_n8686_,
    new_n8687_, new_n8688_, new_n8689_, new_n8690_, new_n8691_, new_n8692_,
    new_n8693_, new_n8694_, new_n8695_, new_n8696_, new_n8697_, new_n8698_,
    new_n8699_, new_n8700_, new_n8701_, new_n8702_, new_n8703_, new_n8704_,
    new_n8705_, new_n8706_, new_n8707_, new_n8708_, new_n8709_, new_n8710_,
    new_n8711_, new_n8712_, new_n8713_, new_n8714_, new_n8715_, new_n8716_,
    new_n8717_, new_n8718_, new_n8719_, new_n8720_, new_n8721_, new_n8722_,
    new_n8723_, new_n8724_, new_n8725_, new_n8726_, new_n8727_, new_n8728_,
    new_n8729_, new_n8730_, new_n8731_, new_n8732_, new_n8733_, new_n8734_,
    new_n8735_, new_n8736_, new_n8737_, new_n8738_, new_n8739_, new_n8740_,
    new_n8741_, new_n8742_, new_n8743_, new_n8744_, new_n8745_, new_n8746_,
    new_n8747_, new_n8748_, new_n8749_, new_n8750_, new_n8751_, new_n8752_,
    new_n8753_, new_n8754_, new_n8755_, new_n8756_, new_n8757_, new_n8758_,
    new_n8759_, new_n8760_, new_n8761_, new_n8762_, new_n8763_, new_n8764_,
    new_n8765_, new_n8766_, new_n8767_, new_n8768_, new_n8769_, new_n8770_,
    new_n8771_, new_n8772_, new_n8773_, new_n8774_, new_n8775_, new_n8776_,
    new_n8777_, new_n8778_, new_n8779_, new_n8780_, new_n8781_, new_n8782_,
    new_n8783_, new_n8784_, new_n8785_, new_n8786_, new_n8787_, new_n8788_,
    new_n8789_, new_n8790_, new_n8791_, new_n8792_, new_n8793_, new_n8794_,
    new_n8795_, new_n8796_, new_n8797_, new_n8798_, new_n8799_, new_n8800_,
    new_n8801_, new_n8802_, new_n8803_, new_n8804_, new_n8805_, new_n8806_,
    new_n8807_, new_n8808_, new_n8809_, new_n8810_, new_n8811_, new_n8812_,
    new_n8813_, new_n8814_, new_n8815_, new_n8816_, new_n8817_, new_n8818_,
    new_n8819_, new_n8820_, new_n8821_, new_n8822_, new_n8823_, new_n8824_,
    new_n8825_, new_n8826_, new_n8827_, new_n8828_, new_n8829_, new_n8830_,
    new_n8831_, new_n8832_, new_n8833_, new_n8834_, new_n8835_, new_n8836_,
    new_n8837_, new_n8838_, new_n8839_, new_n8840_, new_n8841_, new_n8842_,
    new_n8843_, new_n8844_, new_n8845_, new_n8846_, new_n8847_, new_n8848_,
    new_n8849_, new_n8850_, new_n8851_, new_n8852_, new_n8853_, new_n8854_,
    new_n8855_, new_n8856_, new_n8857_, new_n8858_, new_n8859_, new_n8860_,
    new_n8861_, new_n8862_, new_n8863_, new_n8864_, new_n8865_, new_n8866_,
    new_n8867_, new_n8868_, new_n8869_, new_n8870_, new_n8871_, new_n8872_,
    new_n8873_, new_n8874_, new_n8875_, new_n8876_, new_n8877_, new_n8878_,
    new_n8879_, new_n8880_, new_n8881_, new_n8882_, new_n8883_, new_n8884_,
    new_n8885_, new_n8886_, new_n8887_, new_n8888_, new_n8889_, new_n8890_,
    new_n8891_, new_n8892_, new_n8893_, new_n8894_, new_n8895_, new_n8896_,
    new_n8897_, new_n8898_, new_n8899_, new_n8900_, new_n8901_, new_n8902_,
    new_n8903_, new_n8904_, new_n8905_, new_n8906_, new_n8907_, new_n8908_,
    new_n8909_, new_n8910_, new_n8911_, new_n8912_, new_n8913_, new_n8914_,
    new_n8915_, new_n8916_, new_n8917_, new_n8918_, new_n8919_, new_n8920_,
    new_n8921_, new_n8922_, new_n8923_, new_n8924_, new_n8925_, new_n8926_,
    new_n8927_, new_n8928_, new_n8929_, new_n8930_, new_n8931_, new_n8932_,
    new_n8933_, new_n8934_, new_n8935_, new_n8936_, new_n8937_, new_n8938_,
    new_n8939_, new_n8940_, new_n8941_, new_n8942_, new_n8943_, new_n8944_,
    new_n8945_, new_n8946_, new_n8947_, new_n8948_, new_n8949_, new_n8950_,
    new_n8951_, new_n8952_, new_n8953_, new_n8954_, new_n8955_, new_n8956_,
    new_n8957_, new_n8958_, new_n8959_, new_n8960_, new_n8961_, new_n8962_,
    new_n8963_, new_n8964_, new_n8965_, new_n8966_, new_n8967_, new_n8968_,
    new_n8969_, new_n8970_, new_n8971_, new_n8972_, new_n8973_, new_n8974_,
    new_n8975_, new_n8976_, new_n8977_, new_n8978_, new_n8979_, new_n8980_,
    new_n8981_, new_n8982_, new_n8983_, new_n8984_, new_n8985_, new_n8986_,
    new_n8987_, new_n8988_, new_n8989_, new_n8990_, new_n8991_, new_n8992_,
    new_n8993_, new_n8994_, new_n8995_, new_n8996_, new_n8997_, new_n8998_,
    new_n8999_, new_n9000_, new_n9001_, new_n9002_, new_n9003_, new_n9004_,
    new_n9005_, new_n9006_, new_n9007_, new_n9008_, new_n9009_, new_n9010_,
    new_n9011_, new_n9012_, new_n9013_, new_n9014_, new_n9015_, new_n9016_,
    new_n9017_, new_n9018_, new_n9019_, new_n9020_, new_n9021_, new_n9022_,
    new_n9023_, new_n9024_, new_n9025_, new_n9026_, new_n9027_, new_n9028_,
    new_n9029_, new_n9030_, new_n9031_, new_n9032_, new_n9033_, new_n9034_,
    new_n9035_, new_n9036_, new_n9037_, new_n9038_, new_n9039_, new_n9040_,
    new_n9041_, new_n9042_, new_n9043_, new_n9044_, new_n9045_, new_n9046_,
    new_n9047_, new_n9048_, new_n9049_, new_n9050_, new_n9051_, new_n9052_,
    new_n9053_, new_n9054_, new_n9055_, new_n9056_, new_n9057_, new_n9058_,
    new_n9059_, new_n9060_, new_n9061_, new_n9062_, new_n9063_, new_n9064_,
    new_n9065_, new_n9066_, new_n9067_, new_n9068_, new_n9069_, new_n9070_,
    new_n9071_, new_n9072_, new_n9073_, new_n9074_, new_n9075_, new_n9076_,
    new_n9077_, new_n9078_, new_n9079_, new_n9080_, new_n9081_, new_n9082_,
    new_n9083_, new_n9084_, new_n9085_, new_n9086_, new_n9087_, new_n9088_,
    new_n9089_, new_n9090_, new_n9091_, new_n9092_, new_n9093_, new_n9094_,
    new_n9095_, new_n9096_, new_n9097_, new_n9098_, new_n9099_, new_n9100_,
    new_n9101_, new_n9102_, new_n9103_, new_n9104_, new_n9105_, new_n9106_,
    new_n9107_, new_n9108_, new_n9109_, new_n9110_, new_n9111_, new_n9112_,
    new_n9113_, new_n9114_, new_n9115_, new_n9116_, new_n9117_, new_n9118_,
    new_n9119_, new_n9120_, new_n9121_, new_n9122_, new_n9123_, new_n9124_,
    new_n9125_, new_n9126_, new_n9127_, new_n9128_, new_n9129_, new_n9130_,
    new_n9131_, new_n9132_, new_n9133_, new_n9134_, new_n9135_, new_n9136_,
    new_n9137_, new_n9138_, new_n9139_, new_n9140_, new_n9141_, new_n9142_,
    new_n9143_, new_n9144_, new_n9145_, new_n9146_, new_n9147_, new_n9148_,
    new_n9149_, new_n9150_, new_n9151_, new_n9152_, new_n9153_, new_n9154_,
    new_n9155_, new_n9156_, new_n9157_, new_n9158_, new_n9159_, new_n9160_,
    new_n9161_, new_n9162_, new_n9163_, new_n9164_, new_n9165_, new_n9166_,
    new_n9167_, new_n9168_, new_n9169_, new_n9170_, new_n9171_, new_n9172_,
    new_n9173_, new_n9174_, new_n9175_, new_n9176_, new_n9177_, new_n9178_,
    new_n9179_, new_n9180_, new_n9181_, new_n9182_, new_n9183_, new_n9184_,
    new_n9185_, new_n9186_, new_n9187_, new_n9188_, new_n9189_, new_n9190_,
    new_n9191_, new_n9192_, new_n9193_, new_n9194_, new_n9195_, new_n9196_,
    new_n9197_, new_n9198_, new_n9199_, new_n9200_, new_n9201_, new_n9202_,
    new_n9203_, new_n9204_, new_n9205_, new_n9206_, new_n9207_, new_n9208_,
    new_n9209_, new_n9210_, new_n9211_, new_n9212_, new_n9213_, new_n9214_,
    new_n9215_, new_n9216_, new_n9217_, new_n9218_, new_n9219_, new_n9220_,
    new_n9221_, new_n9222_, new_n9223_, new_n9224_, new_n9225_, new_n9226_,
    new_n9227_, new_n9228_, new_n9229_, new_n9230_, new_n9231_, new_n9232_,
    new_n9233_, new_n9234_, new_n9235_, new_n9236_, new_n9237_, new_n9238_,
    new_n9239_, new_n9240_, new_n9241_, new_n9242_, new_n9243_, new_n9244_,
    new_n9245_, new_n9246_, new_n9247_, new_n9248_, new_n9249_, new_n9250_,
    new_n9251_, new_n9252_, new_n9253_, new_n9254_, new_n9255_, new_n9256_,
    new_n9257_, new_n9258_, new_n9259_, new_n9260_, new_n9261_, new_n9262_,
    new_n9263_, new_n9264_, new_n9265_, new_n9266_, new_n9267_, new_n9268_,
    new_n9269_, new_n9270_, new_n9271_, new_n9272_, new_n9273_, new_n9274_,
    new_n9275_, new_n9276_, new_n9277_, new_n9278_, new_n9279_, new_n9280_,
    new_n9281_, new_n9282_, new_n9283_, new_n9284_, new_n9285_, new_n9286_,
    new_n9287_, new_n9288_, new_n9289_, new_n9290_, new_n9291_, new_n9292_,
    new_n9293_, new_n9294_, new_n9295_, new_n9296_, new_n9297_, new_n9298_,
    new_n9299_, new_n9300_, new_n9301_, new_n9302_, new_n9303_, new_n9304_,
    new_n9305_, new_n9306_, new_n9307_, new_n9308_, new_n9309_, new_n9310_,
    new_n9311_, new_n9312_, new_n9313_, new_n9314_, new_n9315_, new_n9316_,
    new_n9317_, new_n9318_, new_n9319_, new_n9320_, new_n9321_, new_n9322_,
    new_n9323_, new_n9324_, new_n9325_, new_n9326_, new_n9327_, new_n9328_,
    new_n9329_, new_n9330_, new_n9331_, new_n9332_, new_n9333_, new_n9334_,
    new_n9335_, new_n9336_, new_n9337_, new_n9338_, new_n9339_, new_n9340_,
    new_n9341_, new_n9342_, new_n9343_, new_n9344_, new_n9345_, new_n9346_,
    new_n9347_, new_n9348_, new_n9349_, new_n9350_, new_n9351_, new_n9352_,
    new_n9353_, new_n9354_, new_n9355_, new_n9356_, new_n9357_, new_n9358_,
    new_n9359_, new_n9360_, new_n9361_, new_n9362_, new_n9363_, new_n9364_,
    new_n9365_, new_n9366_, new_n9367_, new_n9368_, new_n9369_, new_n9370_,
    new_n9371_, new_n9372_, new_n9373_, new_n9374_, new_n9375_, new_n9376_,
    new_n9377_, new_n9378_, new_n9379_, new_n9380_, new_n9381_, new_n9382_,
    new_n9383_, new_n9384_, new_n9385_, new_n9386_, new_n9387_, new_n9388_,
    new_n9389_, new_n9390_, new_n9391_, new_n9392_, new_n9393_, new_n9394_,
    new_n9395_, new_n9396_, new_n9397_, new_n9398_, new_n9399_, new_n9400_,
    new_n9401_, new_n9402_, new_n9403_, new_n9404_, new_n9405_, new_n9406_,
    new_n9407_, new_n9408_, new_n9409_, new_n9410_, new_n9411_, new_n9412_,
    new_n9413_, new_n9414_, new_n9415_, new_n9416_, new_n9417_, new_n9418_,
    new_n9419_, new_n9420_, new_n9421_, new_n9422_, new_n9423_, new_n9424_,
    new_n9425_, new_n9426_, new_n9427_, new_n9428_, new_n9429_, new_n9430_,
    new_n9431_, new_n9432_, new_n9433_, new_n9434_, new_n9435_, new_n9436_,
    new_n9437_, new_n9438_, new_n9439_, new_n9440_, new_n9441_, new_n9442_,
    new_n9443_, new_n9444_, new_n9445_, new_n9446_, new_n9447_, new_n9448_,
    new_n9449_, new_n9450_, new_n9451_, new_n9452_, new_n9453_, new_n9454_,
    new_n9455_, new_n9456_, new_n9457_, new_n9458_, new_n9459_, new_n9460_,
    new_n9461_, new_n9462_, new_n9463_, new_n9464_, new_n9465_, new_n9466_,
    new_n9467_, new_n9468_, new_n9469_, new_n9470_, new_n9471_, new_n9472_,
    new_n9473_, new_n9474_, new_n9475_, new_n9476_, new_n9477_, new_n9478_,
    new_n9479_, new_n9480_, new_n9481_, new_n9482_, new_n9483_, new_n9484_,
    new_n9485_, new_n9486_, new_n9487_, new_n9488_, new_n9489_, new_n9490_,
    new_n9491_, new_n9492_, new_n9493_, new_n9494_, new_n9495_, new_n9496_,
    new_n9497_, new_n9498_, new_n9499_, new_n9500_, new_n9501_, new_n9502_,
    new_n9503_, new_n9504_, new_n9505_, new_n9506_, new_n9507_, new_n9508_,
    new_n9509_, new_n9510_, new_n9511_, new_n9512_, new_n9513_, new_n9514_,
    new_n9515_, new_n9516_, new_n9517_, new_n9518_, new_n9519_, new_n9520_,
    new_n9521_, new_n9522_, new_n9523_, new_n9524_, new_n9525_, new_n9526_,
    new_n9527_, new_n9528_, new_n9529_, new_n9530_, new_n9531_, new_n9532_,
    new_n9533_, new_n9534_, new_n9535_, new_n9536_, new_n9537_, new_n9538_,
    new_n9539_, new_n9540_, new_n9541_, new_n9542_, new_n9543_, new_n9544_,
    new_n9545_, new_n9546_, new_n9547_, new_n9548_, new_n9549_, new_n9550_,
    new_n9551_, new_n9552_, new_n9553_, new_n9554_, new_n9555_, new_n9556_,
    new_n9557_, new_n9558_, new_n9559_, new_n9560_, new_n9561_, new_n9562_,
    new_n9563_, new_n9564_, new_n9565_, new_n9566_, new_n9567_, new_n9568_,
    new_n9569_, new_n9570_, new_n9571_, new_n9572_, new_n9573_, new_n9574_,
    new_n9575_, new_n9576_, new_n9577_, new_n9578_, new_n9579_, new_n9580_,
    new_n9581_, new_n9582_, new_n9583_, new_n9584_, new_n9585_, new_n9586_,
    new_n9587_, new_n9588_, new_n9589_, new_n9590_, new_n9591_, new_n9592_,
    new_n9593_, new_n9594_, new_n9595_, new_n9596_, new_n9597_, new_n9598_,
    new_n9599_, new_n9600_, new_n9601_, new_n9602_, new_n9603_, new_n9604_,
    new_n9605_, new_n9606_, new_n9607_, new_n9608_, new_n9609_, new_n9610_,
    new_n9611_, new_n9612_, new_n9613_, new_n9614_, new_n9615_, new_n9616_,
    new_n9617_, new_n9618_, new_n9619_, new_n9620_, new_n9621_, new_n9622_,
    new_n9623_, new_n9624_, new_n9625_, new_n9626_, new_n9627_, new_n9628_,
    new_n9629_, new_n9630_, new_n9631_, new_n9632_, new_n9633_, new_n9634_,
    new_n9635_, new_n9636_, new_n9637_, new_n9638_, new_n9639_, new_n9640_,
    new_n9641_, new_n9642_, new_n9643_, new_n9644_, new_n9645_, new_n9646_,
    new_n9647_, new_n9648_, new_n9649_, new_n9650_, new_n9651_, new_n9652_,
    new_n9653_, new_n9654_, new_n9655_, new_n9656_, new_n9657_, new_n9658_,
    new_n9659_, new_n9660_, new_n9661_, new_n9662_, new_n9663_, new_n9664_,
    new_n9665_, new_n9666_, new_n9667_, new_n9668_, new_n9669_, new_n9670_,
    new_n9671_, new_n9672_, new_n9673_, new_n9674_, new_n9675_, new_n9676_,
    new_n9677_, new_n9678_, new_n9679_, new_n9680_, new_n9681_, new_n9682_,
    new_n9683_, new_n9684_, new_n9685_, new_n9686_, new_n9687_, new_n9688_,
    new_n9689_, new_n9690_, new_n9691_, new_n9692_, new_n9693_, new_n9694_,
    new_n9695_, new_n9696_, new_n9697_, new_n9698_, new_n9699_, new_n9700_,
    new_n9701_, new_n9702_, new_n9703_, new_n9704_, new_n9705_, new_n9706_,
    new_n9707_, new_n9708_, new_n9709_, new_n9710_, new_n9711_, new_n9712_,
    new_n9713_, new_n9714_, new_n9715_, new_n9716_, new_n9717_, new_n9718_,
    new_n9719_, new_n9720_, new_n9721_, new_n9722_, new_n9723_, new_n9724_,
    new_n9725_, new_n9726_, new_n9727_, new_n9728_, new_n9729_, new_n9730_,
    new_n9731_, new_n9732_, new_n9733_, new_n9734_, new_n9735_, new_n9736_,
    new_n9737_, new_n9738_, new_n9739_, new_n9740_, new_n9741_, new_n9742_,
    new_n9743_, new_n9744_, new_n9745_, new_n9746_, new_n9747_, new_n9748_,
    new_n9749_, new_n9750_, new_n9751_, new_n9752_, new_n9753_, new_n9754_,
    new_n9755_, new_n9756_, new_n9757_, new_n9758_, new_n9759_, new_n9760_,
    new_n9761_, new_n9762_, new_n9763_, new_n9764_, new_n9765_, new_n9766_,
    new_n9767_, new_n9768_, new_n9769_, new_n9770_, new_n9771_, new_n9772_,
    new_n9773_, new_n9774_, new_n9775_, new_n9776_, new_n9777_, new_n9778_,
    new_n9779_, new_n9780_, new_n9781_, new_n9782_, new_n9783_, new_n9784_,
    new_n9785_, new_n9786_, new_n9787_, new_n9788_, new_n9789_, new_n9790_,
    new_n9791_, new_n9792_, new_n9793_, new_n9794_, new_n9795_, new_n9796_,
    new_n9797_, new_n9798_, new_n9799_, new_n9800_, new_n9801_, new_n9802_,
    new_n9803_, new_n9804_, new_n9805_, new_n9806_, new_n9807_, new_n9808_,
    new_n9809_, new_n9810_, new_n9811_, new_n9812_, new_n9813_, new_n9814_,
    new_n9815_, new_n9816_, new_n9817_, new_n9818_, new_n9819_, new_n9820_,
    new_n9821_, new_n9822_, new_n9823_, new_n9824_, new_n9825_, new_n9826_,
    new_n9827_, new_n9828_, new_n9829_, new_n9830_, new_n9831_, new_n9832_,
    new_n9833_, new_n9834_, new_n9835_, new_n9836_, new_n9837_, new_n9838_,
    new_n9839_, new_n9840_, new_n9841_, new_n9842_, new_n9843_, new_n9844_,
    new_n9845_, new_n9846_, new_n9847_, new_n9848_, new_n9849_, new_n9850_,
    new_n9851_, new_n9852_, new_n9853_, new_n9854_, new_n9855_, new_n9856_,
    new_n9857_, new_n9858_, new_n9859_, new_n9860_, new_n9861_, new_n9862_,
    new_n9863_, new_n9864_, new_n9865_, new_n9866_, new_n9867_, new_n9868_,
    new_n9869_, new_n9870_, new_n9871_, new_n9872_, new_n9873_, new_n9874_,
    new_n9875_, new_n9876_, new_n9877_, new_n9878_, new_n9879_, new_n9880_,
    new_n9881_, new_n9882_, new_n9883_, new_n9884_, new_n9885_, new_n9886_,
    new_n9887_, new_n9888_, new_n9889_, new_n9890_, new_n9891_, new_n9892_,
    new_n9893_, new_n9894_, new_n9895_, new_n9896_, new_n9897_, new_n9898_,
    new_n9899_, new_n9900_, new_n9901_, new_n9902_, new_n9903_, new_n9904_,
    new_n9905_, new_n9906_, new_n9907_, new_n9908_, new_n9909_, new_n9910_,
    new_n9911_, new_n9912_, new_n9913_, new_n9914_, new_n9915_, new_n9916_,
    new_n9917_, new_n9918_, new_n9919_, new_n9920_, new_n9921_, new_n9922_,
    new_n9923_, new_n9924_, new_n9925_, new_n9926_, new_n9927_, new_n9928_,
    new_n9929_, new_n9930_, new_n9931_, new_n9932_, new_n9933_, new_n9934_,
    new_n9935_, new_n9936_, new_n9937_, new_n9938_, new_n9939_, new_n9940_,
    new_n9941_, new_n9942_, new_n9943_, new_n9944_, new_n9945_, new_n9946_,
    new_n9947_, new_n9948_, new_n9949_, new_n9950_, new_n9951_, new_n9952_,
    new_n9953_, new_n9954_, new_n9955_, new_n9956_, new_n9957_, new_n9958_,
    new_n9959_, new_n9960_, new_n9961_, new_n9962_, new_n9963_, new_n9964_,
    new_n9965_, new_n9966_, new_n9967_, new_n9968_, new_n9969_, new_n9970_,
    new_n9971_, new_n9972_, new_n9973_, new_n9974_, new_n9975_, new_n9976_,
    new_n9977_, new_n9978_, new_n9979_, new_n9980_, new_n9981_, new_n9982_,
    new_n9983_, new_n9984_, new_n9985_, new_n9986_, new_n9987_, new_n9988_,
    new_n9989_, new_n9990_, new_n9991_, new_n9992_, new_n9993_, new_n9994_,
    new_n9995_, new_n9996_, new_n9997_, new_n9998_, new_n9999_,
    new_n10000_, new_n10001_, new_n10002_, new_n10003_, new_n10004_,
    new_n10005_, new_n10006_, new_n10007_, new_n10008_, new_n10009_,
    new_n10010_, new_n10011_, new_n10012_, new_n10013_, new_n10014_,
    new_n10015_, new_n10016_, new_n10017_, new_n10018_, new_n10019_,
    new_n10020_, new_n10021_, new_n10022_, new_n10023_, new_n10024_,
    new_n10025_, new_n10026_, new_n10027_, new_n10028_, new_n10029_,
    new_n10030_, new_n10031_, new_n10032_, new_n10033_, new_n10034_,
    new_n10035_, new_n10036_, new_n10037_, new_n10038_, new_n10039_,
    new_n10040_, new_n10041_, new_n10042_, new_n10043_, new_n10044_,
    new_n10045_, new_n10046_, new_n10047_, new_n10048_, new_n10049_,
    new_n10050_, new_n10051_, new_n10052_, new_n10053_, new_n10054_,
    new_n10055_, new_n10056_, new_n10057_, new_n10058_, new_n10059_,
    new_n10060_, new_n10061_, new_n10062_, new_n10063_, new_n10064_,
    new_n10065_, new_n10066_, new_n10067_, new_n10068_, new_n10069_,
    new_n10070_, new_n10071_, new_n10072_, new_n10073_, new_n10074_,
    new_n10075_, new_n10076_, new_n10077_, new_n10078_, new_n10079_,
    new_n10080_, new_n10081_, new_n10082_, new_n10083_, new_n10084_,
    new_n10085_, new_n10086_, new_n10087_, new_n10088_, new_n10089_,
    new_n10090_, new_n10091_, new_n10092_, new_n10093_, new_n10094_,
    new_n10095_, new_n10096_, new_n10097_, new_n10098_, new_n10099_,
    new_n10100_, new_n10101_, new_n10102_, new_n10103_, new_n10104_,
    new_n10105_, new_n10106_, new_n10107_, new_n10108_, new_n10109_,
    new_n10110_, new_n10111_, new_n10112_, new_n10113_, new_n10114_,
    new_n10115_, new_n10116_, new_n10117_, new_n10118_, new_n10119_,
    new_n10120_, new_n10121_, new_n10122_, new_n10123_, new_n10124_,
    new_n10125_, new_n10126_, new_n10127_, new_n10128_, new_n10129_,
    new_n10130_, new_n10131_, new_n10132_, new_n10133_, new_n10134_,
    new_n10135_, new_n10136_, new_n10137_, new_n10138_, new_n10139_,
    new_n10140_, new_n10141_, new_n10142_, new_n10143_, new_n10144_,
    new_n10145_, new_n10146_, new_n10147_, new_n10148_, new_n10149_,
    new_n10150_, new_n10151_, new_n10152_, new_n10153_, new_n10154_,
    new_n10155_, new_n10156_, new_n10157_, new_n10158_, new_n10159_,
    new_n10160_, new_n10161_, new_n10162_, new_n10163_, new_n10164_,
    new_n10165_, new_n10166_, new_n10167_, new_n10168_, new_n10169_,
    new_n10170_, new_n10171_, new_n10172_, new_n10173_, new_n10174_,
    new_n10175_, new_n10176_, new_n10177_, new_n10178_, new_n10179_,
    new_n10180_, new_n10181_, new_n10182_, new_n10183_, new_n10184_,
    new_n10185_, new_n10186_, new_n10187_, new_n10188_, new_n10189_,
    new_n10190_, new_n10191_, new_n10192_, new_n10193_, new_n10194_,
    new_n10195_, new_n10196_, new_n10197_, new_n10198_, new_n10199_,
    new_n10200_, new_n10201_, new_n10202_, new_n10203_, new_n10204_,
    new_n10205_, new_n10206_, new_n10207_, new_n10208_, new_n10209_,
    new_n10210_, new_n10211_, new_n10212_, new_n10213_, new_n10214_,
    new_n10215_, new_n10216_, new_n10217_, new_n10218_, new_n10219_,
    new_n10220_, new_n10221_, new_n10222_, new_n10223_, new_n10224_,
    new_n10225_, new_n10226_, new_n10227_, new_n10228_, new_n10229_,
    new_n10230_, new_n10231_, new_n10232_, new_n10233_, new_n10234_,
    new_n10235_, new_n10236_, new_n10237_, new_n10238_, new_n10239_,
    new_n10240_, new_n10241_, new_n10242_, new_n10243_, new_n10244_,
    new_n10245_, new_n10246_, new_n10247_, new_n10248_, new_n10249_,
    new_n10250_, new_n10251_, new_n10252_, new_n10253_, new_n10254_,
    new_n10255_, new_n10256_, new_n10257_, new_n10258_, new_n10259_,
    new_n10260_, new_n10261_, new_n10262_, new_n10263_, new_n10264_,
    new_n10265_, new_n10266_, new_n10267_, new_n10268_, new_n10269_,
    new_n10270_, new_n10271_, new_n10272_, new_n10273_, new_n10274_,
    new_n10275_, new_n10276_, new_n10277_, new_n10278_, new_n10279_,
    new_n10280_, new_n10281_, new_n10282_, new_n10283_, new_n10284_,
    new_n10285_, new_n10286_, new_n10287_, new_n10288_, new_n10289_,
    new_n10290_, new_n10291_, new_n10292_, new_n10293_, new_n10294_,
    new_n10295_, new_n10296_, new_n10297_, new_n10298_, new_n10299_,
    new_n10300_, new_n10301_, new_n10302_, new_n10303_, new_n10304_,
    new_n10305_, new_n10306_, new_n10307_, new_n10308_, new_n10309_,
    new_n10310_, new_n10311_, new_n10312_, new_n10313_, new_n10314_,
    new_n10315_, new_n10316_, new_n10317_, new_n10318_, new_n10319_,
    new_n10320_, new_n10321_, new_n10322_, new_n10323_, new_n10324_,
    new_n10325_, new_n10326_, new_n10327_, new_n10328_, new_n10329_,
    new_n10330_, new_n10331_, new_n10332_, new_n10333_, new_n10334_,
    new_n10335_, new_n10336_, new_n10337_, new_n10338_, new_n10339_,
    new_n10340_, new_n10341_, new_n10342_, new_n10343_, new_n10344_,
    new_n10345_, new_n10346_, new_n10347_, new_n10348_, new_n10349_,
    new_n10350_, new_n10351_, new_n10352_, new_n10353_, new_n10354_,
    new_n10355_, new_n10356_, new_n10357_, new_n10358_, new_n10359_,
    new_n10360_, new_n10361_, new_n10362_, new_n10363_, new_n10364_,
    new_n10365_, new_n10366_, new_n10367_, new_n10368_, new_n10369_,
    new_n10370_, new_n10371_, new_n10372_, new_n10373_, new_n10374_,
    new_n10375_, new_n10376_, new_n10377_, new_n10378_, new_n10379_,
    new_n10380_, new_n10381_, new_n10382_, new_n10383_, new_n10384_,
    new_n10385_, new_n10386_, new_n10387_, new_n10388_, new_n10389_,
    new_n10390_, new_n10391_, new_n10392_, new_n10393_, new_n10394_,
    new_n10395_, new_n10396_, new_n10397_, new_n10398_, new_n10399_,
    new_n10400_, new_n10401_, new_n10402_, new_n10403_, new_n10404_,
    new_n10405_, new_n10406_, new_n10407_, new_n10408_, new_n10409_,
    new_n10410_, new_n10411_, new_n10412_, new_n10413_, new_n10414_,
    new_n10415_, new_n10416_, new_n10417_, new_n10418_, new_n10419_,
    new_n10420_, new_n10421_, new_n10422_, new_n10423_, new_n10424_,
    new_n10425_, new_n10426_, new_n10427_, new_n10428_, new_n10429_,
    new_n10430_, new_n10431_, new_n10432_, new_n10433_, new_n10434_,
    new_n10435_, new_n10436_, new_n10437_, new_n10438_, new_n10439_,
    new_n10440_, new_n10441_, new_n10442_, new_n10443_, new_n10444_,
    new_n10445_, new_n10446_, new_n10447_, new_n10448_, new_n10449_,
    new_n10450_, new_n10451_, new_n10452_, new_n10453_, new_n10454_,
    new_n10455_, new_n10456_, new_n10457_, new_n10458_, new_n10459_,
    new_n10460_, new_n10461_, new_n10462_, new_n10463_, new_n10464_,
    new_n10465_, new_n10466_, new_n10467_, new_n10468_, new_n10469_,
    new_n10470_, new_n10471_, new_n10472_, new_n10473_, new_n10474_,
    new_n10475_, new_n10476_, new_n10477_, new_n10478_, new_n10479_,
    new_n10480_, new_n10481_, new_n10482_, new_n10483_, new_n10484_,
    new_n10485_, new_n10486_, new_n10487_, new_n10488_, new_n10489_,
    new_n10490_, new_n10491_, new_n10492_, new_n10493_, new_n10494_,
    new_n10495_, new_n10496_, new_n10497_, new_n10498_, new_n10499_,
    new_n10500_, new_n10501_, new_n10502_, new_n10503_, new_n10504_,
    new_n10505_, new_n10506_, new_n10507_, new_n10508_, new_n10509_,
    new_n10510_, new_n10511_, new_n10512_, new_n10513_, new_n10514_,
    new_n10515_, new_n10516_, new_n10517_, new_n10518_, new_n10519_,
    new_n10520_, new_n10521_, new_n10522_, new_n10523_, new_n10524_,
    new_n10525_, new_n10526_, new_n10527_, new_n10528_, new_n10529_,
    new_n10530_, new_n10531_, new_n10532_, new_n10533_, new_n10534_,
    new_n10535_, new_n10536_, new_n10537_, new_n10538_, new_n10539_,
    new_n10540_, new_n10541_, new_n10542_, new_n10543_, new_n10544_,
    new_n10545_, new_n10546_, new_n10547_, new_n10548_, new_n10549_,
    new_n10550_, new_n10551_, new_n10552_, new_n10553_, new_n10554_,
    new_n10555_, new_n10556_, new_n10557_, new_n10558_, new_n10559_,
    new_n10560_, new_n10561_, new_n10562_, new_n10563_, new_n10564_,
    new_n10565_, new_n10566_, new_n10567_, new_n10568_, new_n10569_,
    new_n10570_, new_n10571_, new_n10572_, new_n10573_, new_n10574_,
    new_n10575_, new_n10576_, new_n10577_, new_n10578_, new_n10579_,
    new_n10580_, new_n10581_, new_n10582_, new_n10583_, new_n10584_,
    new_n10585_, new_n10586_, new_n10587_, new_n10588_, new_n10589_,
    new_n10590_, new_n10591_, new_n10592_, new_n10593_, new_n10594_,
    new_n10595_, new_n10596_, new_n10597_, new_n10598_, new_n10599_,
    new_n10600_, new_n10601_, new_n10602_, new_n10603_, new_n10604_,
    new_n10605_, new_n10606_, new_n10607_, new_n10608_, new_n10609_,
    new_n10610_, new_n10611_, new_n10612_, new_n10613_, new_n10614_,
    new_n10615_, new_n10616_, new_n10617_, new_n10618_, new_n10619_,
    new_n10620_, new_n10621_, new_n10622_, new_n10623_, new_n10624_,
    new_n10625_, new_n10626_, new_n10627_, new_n10628_, new_n10629_,
    new_n10630_, new_n10631_, new_n10632_, new_n10633_, new_n10634_,
    new_n10635_, new_n10636_, new_n10637_, new_n10638_, new_n10639_,
    new_n10640_, new_n10641_, new_n10642_, new_n10643_, new_n10644_,
    new_n10645_, new_n10646_, new_n10647_, new_n10648_, new_n10649_,
    new_n10650_, new_n10651_, new_n10652_, new_n10653_, new_n10654_,
    new_n10655_, new_n10656_, new_n10657_, new_n10658_, new_n10659_,
    new_n10660_, new_n10661_, new_n10662_, new_n10663_, new_n10664_,
    new_n10665_, new_n10666_, new_n10667_, new_n10668_, new_n10669_,
    new_n10670_, new_n10671_, new_n10672_, new_n10673_, new_n10674_,
    new_n10675_, new_n10676_, new_n10677_, new_n10678_, new_n10679_,
    new_n10680_, new_n10681_, new_n10682_, new_n10683_, new_n10684_,
    new_n10685_, new_n10686_, new_n10687_, new_n10688_, new_n10689_,
    new_n10690_, new_n10691_, new_n10692_, new_n10693_, new_n10694_,
    new_n10695_, new_n10696_, new_n10697_, new_n10698_, new_n10699_,
    new_n10700_, new_n10701_, new_n10702_, new_n10703_, new_n10704_,
    new_n10705_, new_n10706_, new_n10707_, new_n10708_, new_n10709_,
    new_n10710_, new_n10711_, new_n10712_, new_n10713_, new_n10714_,
    new_n10715_, new_n10716_, new_n10717_, new_n10718_, new_n10719_,
    new_n10720_, new_n10721_, new_n10722_, new_n10723_, new_n10724_,
    new_n10725_, new_n10726_, new_n10727_, new_n10728_, new_n10729_,
    new_n10730_, new_n10731_, new_n10732_, new_n10733_, new_n10734_,
    new_n10735_, new_n10736_, new_n10737_, new_n10738_, new_n10739_,
    new_n10740_, new_n10741_, new_n10742_, new_n10743_, new_n10744_,
    new_n10745_, new_n10746_, new_n10747_, new_n10748_, new_n10749_,
    new_n10750_, new_n10751_, new_n10752_, new_n10753_, new_n10754_,
    new_n10755_, new_n10756_, new_n10757_, new_n10758_, new_n10759_,
    new_n10760_, new_n10761_, new_n10762_, new_n10763_, new_n10764_,
    new_n10765_, new_n10766_, new_n10767_, new_n10768_, new_n10769_,
    new_n10770_, new_n10771_, new_n10772_, new_n10773_, new_n10774_,
    new_n10775_, new_n10776_, new_n10777_, new_n10778_, new_n10779_,
    new_n10780_, new_n10781_, new_n10782_, new_n10783_, new_n10784_,
    new_n10785_, new_n10786_, new_n10787_, new_n10788_, new_n10789_,
    new_n10790_, new_n10791_, new_n10792_, new_n10793_, new_n10794_,
    new_n10795_, new_n10796_, new_n10797_, new_n10798_, new_n10799_,
    new_n10800_, new_n10801_, new_n10802_, new_n10803_, new_n10804_,
    new_n10805_, new_n10806_, new_n10807_, new_n10808_, new_n10809_,
    new_n10810_, new_n10811_, new_n10812_, new_n10813_, new_n10814_,
    new_n10815_, new_n10816_, new_n10817_, new_n10818_, new_n10819_,
    new_n10820_, new_n10821_, new_n10822_, new_n10823_, new_n10824_,
    new_n10825_, new_n10826_, new_n10827_, new_n10828_, new_n10829_,
    new_n10830_, new_n10831_, new_n10832_, new_n10833_, new_n10834_,
    new_n10835_, new_n10836_, new_n10837_, new_n10838_, new_n10839_,
    new_n10840_, new_n10841_, new_n10842_, new_n10843_, new_n10844_,
    new_n10845_, new_n10846_, new_n10847_, new_n10848_, new_n10849_,
    new_n10850_, new_n10851_, new_n10852_, new_n10853_, new_n10854_,
    new_n10855_, new_n10856_, new_n10857_, new_n10858_, new_n10859_,
    new_n10860_, new_n10861_, new_n10862_, new_n10863_, new_n10864_,
    new_n10865_, new_n10866_, new_n10867_, new_n10868_, new_n10869_,
    new_n10870_, new_n10871_, new_n10872_, new_n10873_, new_n10874_,
    new_n10875_, new_n10876_, new_n10877_, new_n10878_, new_n10879_,
    new_n10880_, new_n10881_, new_n10882_, new_n10883_, new_n10884_,
    new_n10885_, new_n10886_, new_n10887_, new_n10888_, new_n10889_,
    new_n10890_, new_n10891_, new_n10892_, new_n10893_, new_n10894_,
    new_n10895_, new_n10896_, new_n10897_, new_n10898_, new_n10899_,
    new_n10900_, new_n10901_, new_n10902_, new_n10903_, new_n10904_,
    new_n10905_, new_n10906_, new_n10907_, new_n10908_, new_n10909_,
    new_n10910_, new_n10911_, new_n10912_, new_n10913_, new_n10914_,
    new_n10915_, new_n10916_, new_n10917_, new_n10918_, new_n10919_,
    new_n10920_, new_n10921_, new_n10922_, new_n10923_, new_n10924_,
    new_n10925_, new_n10926_, new_n10927_, new_n10928_, new_n10929_,
    new_n10930_, new_n10931_, new_n10932_, new_n10933_, new_n10934_,
    new_n10935_, new_n10936_, new_n10937_, new_n10938_, new_n10939_,
    new_n10940_, new_n10941_, new_n10942_, new_n10943_, new_n10944_,
    new_n10945_, new_n10946_, new_n10947_, new_n10948_, new_n10949_,
    new_n10950_, new_n10951_, new_n10952_, new_n10953_, new_n10954_,
    new_n10955_, new_n10956_, new_n10957_, new_n10958_, new_n10959_,
    new_n10960_, new_n10961_, new_n10962_, new_n10963_, new_n10964_,
    new_n10965_, new_n10966_, new_n10967_, new_n10968_, new_n10969_,
    new_n10970_, new_n10971_, new_n10972_, new_n10973_, new_n10974_,
    new_n10975_, new_n10976_, new_n10977_, new_n10978_, new_n10979_,
    new_n10980_, new_n10981_, new_n10982_, new_n10983_, new_n10984_,
    new_n10985_, new_n10986_, new_n10987_, new_n10988_, new_n10989_,
    new_n10990_, new_n10991_, new_n10992_, new_n10993_, new_n10994_,
    new_n10995_, new_n10996_, new_n10997_, new_n10998_, new_n10999_,
    new_n11000_, new_n11001_, new_n11002_, new_n11003_, new_n11004_,
    new_n11005_, new_n11006_, new_n11007_, new_n11008_, new_n11009_,
    new_n11010_, new_n11011_, new_n11012_, new_n11013_, new_n11014_,
    new_n11015_, new_n11016_, new_n11017_, new_n11018_, new_n11019_,
    new_n11020_, new_n11021_, new_n11022_, new_n11023_, new_n11024_,
    new_n11025_, new_n11026_, new_n11027_, new_n11028_, new_n11029_,
    new_n11030_, new_n11031_, new_n11032_, new_n11033_, new_n11034_,
    new_n11035_, new_n11036_, new_n11037_, new_n11038_, new_n11039_,
    new_n11040_, new_n11041_, new_n11042_, new_n11043_, new_n11044_,
    new_n11045_, new_n11046_, new_n11047_, new_n11048_, new_n11049_,
    new_n11050_, new_n11051_, new_n11052_, new_n11053_, new_n11054_,
    new_n11055_, new_n11056_, new_n11057_, new_n11058_, new_n11059_,
    new_n11060_, new_n11061_, new_n11062_, new_n11063_, new_n11064_,
    new_n11065_, new_n11066_, new_n11067_, new_n11068_, new_n11069_,
    new_n11070_, new_n11071_, new_n11072_, new_n11073_, new_n11074_,
    new_n11075_, new_n11076_, new_n11077_, new_n11078_, new_n11079_,
    new_n11080_, new_n11081_, new_n11082_, new_n11083_, new_n11084_,
    new_n11085_, new_n11086_, new_n11087_, new_n11088_, new_n11089_,
    new_n11090_, new_n11091_, new_n11092_, new_n11093_, new_n11094_,
    new_n11095_, new_n11096_, new_n11097_, new_n11098_, new_n11099_,
    new_n11100_, new_n11101_, new_n11102_, new_n11103_, new_n11104_,
    new_n11105_, new_n11106_, new_n11107_, new_n11108_, new_n11109_,
    new_n11110_, new_n11111_, new_n11112_, new_n11113_, new_n11114_,
    new_n11115_, new_n11116_, new_n11117_, new_n11118_, new_n11119_,
    new_n11120_, new_n11121_, new_n11122_, new_n11123_, new_n11124_,
    new_n11125_, new_n11126_, new_n11127_, new_n11128_, new_n11129_,
    new_n11130_, new_n11131_, new_n11132_, new_n11133_, new_n11134_,
    new_n11135_, new_n11136_, new_n11137_, new_n11138_, new_n11139_,
    new_n11140_, new_n11141_, new_n11142_, new_n11143_, new_n11144_,
    new_n11145_, new_n11146_, new_n11147_, new_n11148_, new_n11149_,
    new_n11150_, new_n11151_, new_n11152_, new_n11153_, new_n11154_,
    new_n11155_, new_n11156_, new_n11157_, new_n11158_, new_n11159_,
    new_n11160_, new_n11161_, new_n11162_, new_n11163_, new_n11164_,
    new_n11165_, new_n11166_, new_n11167_, new_n11168_, new_n11169_,
    new_n11170_, new_n11171_, new_n11172_, new_n11173_, new_n11174_,
    new_n11175_, new_n11176_, new_n11177_, new_n11178_, new_n11179_,
    new_n11180_, new_n11181_, new_n11182_, new_n11183_, new_n11184_,
    new_n11185_, new_n11186_, new_n11187_, new_n11188_, new_n11189_,
    new_n11190_, new_n11191_, new_n11192_, new_n11193_, new_n11194_,
    new_n11195_, new_n11196_, new_n11197_, new_n11198_, new_n11199_,
    new_n11200_, new_n11201_, new_n11202_, new_n11203_, new_n11204_,
    new_n11205_, new_n11206_, new_n11207_, new_n11208_, new_n11209_,
    new_n11210_, new_n11211_, new_n11212_, new_n11213_, new_n11214_,
    new_n11215_, new_n11216_, new_n11217_, new_n11218_, new_n11219_,
    new_n11220_, new_n11221_, new_n11222_, new_n11223_, new_n11224_,
    new_n11225_, new_n11226_, new_n11227_, new_n11228_, new_n11229_,
    new_n11230_, new_n11231_, new_n11232_, new_n11233_, new_n11234_,
    new_n11235_, new_n11236_, new_n11237_, new_n11238_, new_n11239_,
    new_n11240_, new_n11241_, new_n11242_, new_n11243_, new_n11244_,
    new_n11245_, new_n11246_, new_n11247_, new_n11248_, new_n11249_,
    new_n11250_, new_n11251_, new_n11252_, new_n11253_, new_n11254_,
    new_n11255_, new_n11256_, new_n11257_, new_n11258_, new_n11259_,
    new_n11260_, new_n11261_, new_n11262_, new_n11263_, new_n11264_,
    new_n11265_, new_n11266_, new_n11267_, new_n11268_, new_n11269_,
    new_n11270_, new_n11271_, new_n11272_, new_n11273_, new_n11274_,
    new_n11275_, new_n11276_, new_n11277_, new_n11278_, new_n11279_,
    new_n11280_, new_n11281_, new_n11282_, new_n11283_, new_n11284_,
    new_n11285_, new_n11286_, new_n11287_, new_n11288_, new_n11289_,
    new_n11290_, new_n11291_, new_n11292_, new_n11293_, new_n11294_,
    new_n11295_, new_n11296_, new_n11297_, new_n11298_, new_n11299_,
    new_n11300_, new_n11301_, new_n11302_, new_n11303_, new_n11304_,
    new_n11305_, new_n11306_, new_n11307_, new_n11308_, new_n11309_,
    new_n11310_, new_n11311_, new_n11312_, new_n11313_, new_n11314_,
    new_n11315_, new_n11316_, new_n11317_, new_n11318_, new_n11319_,
    new_n11320_, new_n11321_, new_n11322_, new_n11323_, new_n11324_,
    new_n11325_, new_n11326_, new_n11327_, new_n11328_, new_n11329_,
    new_n11330_, new_n11331_, new_n11332_, new_n11333_, new_n11334_,
    new_n11335_, new_n11336_, new_n11337_, new_n11338_, new_n11339_,
    new_n11340_, new_n11341_, new_n11342_, new_n11343_, new_n11344_,
    new_n11345_, new_n11346_, new_n11347_, new_n11348_, new_n11349_,
    new_n11350_, new_n11351_, new_n11352_, new_n11353_, new_n11354_,
    new_n11355_, new_n11356_, new_n11357_, new_n11358_, new_n11359_,
    new_n11360_, new_n11361_, new_n11362_, new_n11363_, new_n11364_,
    new_n11365_, new_n11366_, new_n11367_, new_n11368_, new_n11369_,
    new_n11370_, new_n11371_, new_n11372_, new_n11373_, new_n11374_,
    new_n11375_, new_n11376_, new_n11377_, new_n11378_, new_n11379_,
    new_n11380_, new_n11381_, new_n11382_, new_n11383_, new_n11384_,
    new_n11385_, new_n11386_, new_n11387_, new_n11388_, new_n11389_,
    new_n11390_, new_n11391_, new_n11392_, new_n11393_, new_n11394_,
    new_n11395_, new_n11396_, new_n11397_, new_n11398_, new_n11399_,
    new_n11400_, new_n11401_, new_n11402_, new_n11403_, new_n11404_,
    new_n11405_, new_n11406_, new_n11407_, new_n11408_, new_n11409_,
    new_n11410_, new_n11411_, new_n11412_, new_n11413_, new_n11414_,
    new_n11415_, new_n11416_, new_n11417_, new_n11418_, new_n11419_,
    new_n11420_, new_n11421_, new_n11422_, new_n11423_, new_n11424_,
    new_n11425_, new_n11426_, new_n11427_, new_n11428_, new_n11429_,
    new_n11430_, new_n11431_, new_n11432_, new_n11433_, new_n11434_,
    new_n11435_, new_n11436_, new_n11437_, new_n11438_, new_n11439_,
    new_n11440_, new_n11441_, new_n11442_, new_n11443_, new_n11444_,
    new_n11445_, new_n11446_, new_n11447_, new_n11448_, new_n11449_,
    new_n11450_, new_n11451_, new_n11452_, new_n11453_, new_n11454_,
    new_n11455_, new_n11456_, new_n11457_, new_n11458_, new_n11459_,
    new_n11460_, new_n11461_, new_n11462_, new_n11463_, new_n11464_,
    new_n11465_, new_n11466_, new_n11467_, new_n11468_, new_n11469_,
    new_n11470_, new_n11471_, new_n11472_, new_n11473_, new_n11474_,
    new_n11475_, new_n11476_, new_n11477_, new_n11478_, new_n11479_,
    new_n11480_, new_n11481_, new_n11482_, new_n11483_, new_n11484_,
    new_n11485_, new_n11486_, new_n11487_, new_n11488_, new_n11489_,
    new_n11490_, new_n11491_, new_n11492_, new_n11493_, new_n11494_,
    new_n11495_, new_n11496_, new_n11497_, new_n11498_, new_n11499_,
    new_n11500_, new_n11501_, new_n11502_, new_n11503_, new_n11504_,
    new_n11505_, new_n11506_, new_n11507_, new_n11508_, new_n11509_,
    new_n11510_, new_n11511_, new_n11512_, new_n11513_, new_n11514_;
not  ( new_n66_, \d[5]  );
xor  ( new_n67_, \d[4] , new_n66_ );
xor  ( new_n68_, \d[3] , \d[4]  );
nor  ( new_n69_, new_n68_, new_n67_ );
xor  ( new_n70_, \d[5] , \a[10]  );
and  ( new_n71_, new_n70_, new_n69_ );
xor  ( new_n72_, \d[5] , \a[11]  );
and  ( new_n73_, new_n72_, new_n68_ );
nor  ( new_n74_, new_n73_, new_n71_ );
not  ( new_n75_, \d[11]  );
xor  ( new_n76_, \d[10] , new_n75_ );
xor  ( new_n77_, \d[9] , \d[10]  );
nor  ( new_n78_, new_n77_, new_n76_ );
xor  ( new_n79_, \d[11] , \a[4]  );
nand ( new_n80_, new_n79_, new_n78_ );
xor  ( new_n81_, \d[11] , \a[5]  );
nand ( new_n82_, new_n81_, new_n77_ );
and  ( new_n83_, new_n82_, new_n80_ );
xor  ( new_n84_, new_n83_, new_n74_ );
not  ( new_n85_, \a[12]  );
not  ( new_n86_, \d[0]  );
and  ( new_n87_, new_n86_, \d[1]  );
and  ( new_n88_, new_n87_, new_n85_ );
not  ( new_n89_, \a[13]  );
not  ( new_n90_, \d[1]  );
and  ( new_n91_, new_n90_, new_n89_ );
not  ( new_n92_, new_n91_ );
and  ( new_n93_, \d[1] , \a[13]  );
nor  ( new_n94_, new_n93_, new_n86_ );
and  ( new_n95_, new_n94_, new_n92_ );
nor  ( new_n96_, new_n95_, new_n88_ );
not  ( new_n97_, new_n96_ );
not  ( new_n98_, \a[0]  );
not  ( new_n99_, \d[12]  );
and  ( new_n100_, new_n75_, new_n99_ );
nor  ( new_n101_, new_n100_, new_n98_ );
not  ( new_n102_, new_n101_ );
not  ( new_n103_, \d[13]  );
and  ( new_n104_, \d[11] , \d[12]  );
nor  ( new_n105_, new_n104_, new_n103_ );
and  ( new_n106_, new_n105_, new_n102_ );
nand ( new_n107_, new_n106_, new_n97_ );
not  ( new_n108_, \a[1]  );
xor  ( new_n109_, \d[13] , new_n108_ );
xor  ( new_n110_, \d[11] , \d[12]  );
xor  ( new_n111_, \d[12] , new_n103_ );
or   ( new_n112_, new_n111_, new_n110_ );
or   ( new_n113_, new_n112_, new_n109_ );
not  ( new_n114_, new_n110_ );
not  ( new_n115_, \a[2]  );
xor  ( new_n116_, \d[13] , new_n115_ );
or   ( new_n117_, new_n116_, new_n114_ );
and  ( new_n118_, new_n117_, new_n113_ );
or   ( new_n119_, new_n118_, new_n107_ );
and  ( new_n120_, new_n118_, new_n107_ );
xor  ( new_n121_, \d[11] , \a[3]  );
and  ( new_n122_, new_n121_, new_n78_ );
and  ( new_n123_, new_n79_, new_n77_ );
nor  ( new_n124_, new_n123_, new_n122_ );
or   ( new_n125_, new_n124_, new_n120_ );
and  ( new_n126_, new_n125_, new_n119_ );
xnor ( new_n127_, new_n126_, new_n84_ );
not  ( new_n128_, \d[7]  );
xor  ( new_n129_, \d[6] , new_n128_ );
xor  ( new_n130_, \d[5] , \d[6]  );
nor  ( new_n131_, new_n130_, new_n129_ );
not  ( new_n132_, new_n131_ );
not  ( new_n133_, \a[8]  );
xor  ( new_n134_, \d[7] , new_n133_ );
or   ( new_n135_, new_n134_, new_n132_ );
not  ( new_n136_, new_n130_ );
not  ( new_n137_, \a[9]  );
xor  ( new_n138_, \d[7] , new_n137_ );
or   ( new_n139_, new_n138_, new_n136_ );
and  ( new_n140_, new_n139_, new_n135_ );
xor  ( new_n141_, new_n140_, new_n127_ );
xor  ( new_n142_, \d[13] , \d[14]  );
and  ( new_n143_, new_n142_, \a[0]  );
not  ( new_n144_, new_n143_ );
xor  ( new_n145_, \d[1] , \a[14]  );
and  ( new_n146_, new_n145_, \d[0]  );
and  ( new_n147_, new_n87_, new_n89_ );
nor  ( new_n148_, new_n147_, new_n146_ );
nor  ( new_n149_, new_n148_, new_n144_ );
not  ( new_n150_, \d[3]  );
xor  ( new_n151_, \d[2] , new_n150_ );
xor  ( new_n152_, \d[1] , \d[2]  );
nor  ( new_n153_, new_n152_, new_n151_ );
xor  ( new_n154_, \d[3] , \a[11]  );
and  ( new_n155_, new_n154_, new_n153_ );
xor  ( new_n156_, \d[3] , \a[12]  );
and  ( new_n157_, new_n156_, new_n152_ );
or   ( new_n158_, new_n157_, new_n155_ );
xor  ( new_n159_, new_n148_, new_n144_ );
and  ( new_n160_, new_n159_, new_n158_ );
or   ( new_n161_, new_n160_, new_n149_ );
or   ( new_n162_, new_n116_, new_n112_ );
not  ( new_n163_, \a[3]  );
xor  ( new_n164_, \d[13] , new_n163_ );
or   ( new_n165_, new_n164_, new_n114_ );
and  ( new_n166_, new_n165_, new_n162_ );
xor  ( new_n167_, new_n166_, new_n161_ );
xnor ( new_n168_, new_n167_, new_n141_ );
and  ( new_n169_, new_n128_, \d[8]  );
and  ( new_n170_, new_n128_, \d[9]  );
not  ( new_n171_, \d[9]  );
and  ( new_n172_, \d[8] , new_n171_ );
nor  ( new_n173_, new_n172_, new_n170_ );
nor  ( new_n174_, new_n173_, new_n169_ );
not  ( new_n175_, new_n174_ );
not  ( new_n176_, \a[5]  );
xor  ( new_n177_, \d[9] , new_n176_ );
or   ( new_n178_, new_n177_, new_n175_ );
not  ( new_n179_, \d[8]  );
xor  ( new_n180_, \d[7] , new_n179_ );
not  ( new_n181_, new_n180_ );
xor  ( new_n182_, \d[9] , \a[6]  );
nand ( new_n183_, new_n182_, new_n181_ );
and  ( new_n184_, new_n183_, new_n178_ );
not  ( new_n185_, \a[7]  );
xor  ( new_n186_, \d[7] , new_n185_ );
or   ( new_n187_, new_n186_, new_n132_ );
or   ( new_n188_, new_n134_, new_n136_ );
and  ( new_n189_, new_n188_, new_n187_ );
or   ( new_n190_, new_n189_, new_n184_ );
xor  ( new_n191_, \d[5] , \a[9]  );
and  ( new_n192_, new_n191_, new_n69_ );
and  ( new_n193_, new_n70_, new_n68_ );
nor  ( new_n194_, new_n193_, new_n192_ );
not  ( new_n195_, new_n194_ );
xor  ( new_n196_, new_n189_, new_n184_ );
nand ( new_n197_, new_n196_, new_n195_ );
and  ( new_n198_, new_n197_, new_n190_ );
or   ( new_n199_, new_n145_, \d[0]  );
and  ( new_n200_, \d[0] , \a[15]  );
xor  ( new_n201_, new_n200_, \d[1]  );
and  ( new_n202_, new_n201_, new_n199_ );
xor  ( new_n203_, new_n202_, new_n198_ );
xor  ( new_n204_, new_n196_, new_n195_ );
xnor ( new_n205_, new_n118_, new_n107_ );
xor  ( new_n206_, new_n205_, new_n124_ );
and  ( new_n207_, new_n206_, new_n204_ );
or   ( new_n208_, new_n206_, new_n204_ );
or   ( new_n209_, new_n114_, new_n98_ );
xor  ( new_n210_, \d[7] , new_n176_ );
or   ( new_n211_, new_n210_, new_n132_ );
not  ( new_n212_, \a[6]  );
xor  ( new_n213_, \d[7] , new_n212_ );
or   ( new_n214_, new_n213_, new_n136_ );
and  ( new_n215_, new_n214_, new_n211_ );
nor  ( new_n216_, new_n215_, new_n209_ );
xor  ( new_n217_, \d[3] , \a[9]  );
and  ( new_n218_, new_n217_, new_n153_ );
xor  ( new_n219_, \d[3] , \a[10]  );
and  ( new_n220_, new_n219_, new_n152_ );
nor  ( new_n221_, new_n220_, new_n218_ );
not  ( new_n222_, new_n221_ );
xor  ( new_n223_, new_n215_, new_n209_ );
and  ( new_n224_, new_n223_, new_n222_ );
or   ( new_n225_, new_n224_, new_n216_ );
xor  ( new_n226_, new_n106_, new_n97_ );
and  ( new_n227_, new_n226_, new_n225_ );
nor  ( new_n228_, new_n226_, new_n225_ );
xor  ( new_n229_, \d[9] , new_n163_ );
or   ( new_n230_, new_n229_, new_n175_ );
not  ( new_n231_, \a[4]  );
xor  ( new_n232_, \d[9] , new_n231_ );
or   ( new_n233_, new_n232_, new_n180_ );
and  ( new_n234_, new_n233_, new_n230_ );
not  ( new_n235_, new_n87_ );
or   ( new_n236_, new_n235_, \a[11]  );
and  ( new_n237_, new_n90_, new_n85_ );
and  ( new_n238_, \d[1] , \a[12]  );
or   ( new_n239_, new_n238_, new_n86_ );
or   ( new_n240_, new_n239_, new_n237_ );
and  ( new_n241_, new_n240_, new_n236_ );
nor  ( new_n242_, new_n241_, new_n234_ );
xor  ( new_n243_, \d[11] , \a[1]  );
and  ( new_n244_, new_n243_, new_n78_ );
xor  ( new_n245_, \d[11] , \a[2]  );
and  ( new_n246_, new_n245_, new_n77_ );
nor  ( new_n247_, new_n246_, new_n244_ );
and  ( new_n248_, new_n241_, new_n234_ );
nor  ( new_n249_, new_n248_, new_n247_ );
nor  ( new_n250_, new_n249_, new_n242_ );
nor  ( new_n251_, new_n250_, new_n228_ );
or   ( new_n252_, new_n251_, new_n227_ );
and  ( new_n253_, new_n252_, new_n208_ );
or   ( new_n254_, new_n253_, new_n207_ );
not  ( new_n255_, \d[15]  );
not  ( new_n256_, \d[14]  );
and  ( new_n257_, new_n256_, new_n98_ );
nor  ( new_n258_, new_n257_, new_n255_ );
and  ( new_n259_, \d[14] , \a[0]  );
not  ( new_n260_, new_n259_ );
and  ( new_n261_, new_n260_, new_n255_ );
or   ( new_n262_, new_n261_, new_n142_ );
or   ( new_n263_, new_n262_, new_n258_ );
xor  ( new_n264_, \d[15] , \a[1]  );
nand ( new_n265_, new_n264_, new_n142_ );
and  ( new_n266_, new_n265_, new_n263_ );
xor  ( new_n267_, new_n266_, new_n254_ );
xor  ( new_n268_, new_n267_, new_n203_ );
xor  ( new_n269_, new_n268_, new_n168_ );
nand ( new_n270_, new_n245_, new_n78_ );
nand ( new_n271_, new_n121_, new_n77_ );
and  ( new_n272_, new_n271_, new_n270_ );
or   ( new_n273_, new_n114_, new_n109_ );
and  ( new_n274_, new_n99_, \d[13]  );
and  ( new_n275_, \d[12] , \a[0]  );
nor  ( new_n276_, new_n275_, new_n274_ );
and  ( new_n277_, \d[13] , \a[0]  );
or   ( new_n278_, new_n277_, new_n110_ );
or   ( new_n279_, new_n278_, new_n276_ );
and  ( new_n280_, new_n279_, new_n273_ );
nor  ( new_n281_, new_n280_, new_n272_ );
xor  ( new_n282_, \d[5] , \a[8]  );
and  ( new_n283_, new_n282_, new_n69_ );
and  ( new_n284_, new_n191_, new_n68_ );
or   ( new_n285_, new_n284_, new_n283_ );
xor  ( new_n286_, new_n280_, new_n272_ );
and  ( new_n287_, new_n286_, new_n285_ );
or   ( new_n288_, new_n287_, new_n281_ );
xor  ( new_n289_, new_n159_, new_n158_ );
and  ( new_n290_, new_n289_, new_n288_ );
xnor ( new_n291_, new_n289_, new_n288_ );
or   ( new_n292_, new_n232_, new_n175_ );
or   ( new_n293_, new_n180_, new_n177_ );
and  ( new_n294_, new_n293_, new_n292_ );
or   ( new_n295_, new_n213_, new_n132_ );
or   ( new_n296_, new_n186_, new_n136_ );
and  ( new_n297_, new_n296_, new_n295_ );
nor  ( new_n298_, new_n297_, new_n294_ );
and  ( new_n299_, new_n219_, new_n153_ );
and  ( new_n300_, new_n154_, new_n152_ );
nor  ( new_n301_, new_n300_, new_n299_ );
and  ( new_n302_, new_n297_, new_n294_ );
nor  ( new_n303_, new_n302_, new_n301_ );
nor  ( new_n304_, new_n303_, new_n298_ );
nor  ( new_n305_, new_n304_, new_n291_ );
or   ( new_n306_, new_n305_, new_n290_ );
and  ( new_n307_, new_n182_, new_n174_ );
xor  ( new_n308_, \d[9] , \a[7]  );
and  ( new_n309_, new_n308_, new_n181_ );
or   ( new_n310_, new_n309_, new_n307_ );
nand ( new_n311_, new_n156_, new_n153_ );
not  ( new_n312_, new_n152_ );
xor  ( new_n313_, \d[3] , new_n89_ );
or   ( new_n314_, new_n313_, new_n312_ );
and  ( new_n315_, new_n314_, new_n311_ );
xor  ( new_n316_, new_n315_, new_n310_ );
xor  ( new_n317_, new_n316_, new_n306_ );
xnor ( new_n318_, new_n317_, new_n269_ );
not  ( new_n319_, new_n318_ );
xor  ( new_n320_, new_n226_, new_n225_ );
xor  ( new_n321_, new_n320_, new_n250_ );
xor  ( new_n322_, \d[3] , \a[8]  );
and  ( new_n323_, new_n322_, new_n153_ );
and  ( new_n324_, new_n217_, new_n152_ );
nor  ( new_n325_, new_n324_, new_n323_ );
not  ( new_n326_, \d[10]  );
and  ( new_n327_, new_n171_, new_n98_ );
or   ( new_n328_, new_n327_, new_n326_ );
and  ( new_n329_, \d[9] , \a[0]  );
nor  ( new_n330_, new_n329_, new_n75_ );
nand ( new_n331_, new_n330_, new_n328_ );
nor  ( new_n332_, new_n331_, new_n325_ );
not  ( new_n333_, new_n332_ );
not  ( new_n334_, new_n69_ );
xor  ( new_n335_, \d[5] , new_n185_ );
or   ( new_n336_, new_n335_, new_n334_ );
nand ( new_n337_, new_n282_, new_n68_ );
and  ( new_n338_, new_n337_, new_n336_ );
nor  ( new_n339_, new_n338_, new_n333_ );
xor  ( new_n340_, new_n338_, new_n333_ );
not  ( new_n341_, new_n340_ );
xor  ( new_n342_, \d[7] , \a[4]  );
nand ( new_n343_, new_n342_, new_n131_ );
or   ( new_n344_, new_n210_, new_n136_ );
and  ( new_n345_, new_n344_, new_n343_ );
xor  ( new_n346_, \d[9] , new_n115_ );
or   ( new_n347_, new_n346_, new_n175_ );
or   ( new_n348_, new_n229_, new_n180_ );
and  ( new_n349_, new_n348_, new_n347_ );
or   ( new_n350_, new_n349_, new_n345_ );
and  ( new_n351_, new_n349_, new_n345_ );
not  ( new_n352_, \a[10]  );
and  ( new_n353_, new_n87_, new_n352_ );
not  ( new_n354_, \a[11]  );
and  ( new_n355_, new_n90_, new_n354_ );
not  ( new_n356_, new_n355_ );
and  ( new_n357_, \d[1] , \a[11]  );
nor  ( new_n358_, new_n357_, new_n86_ );
and  ( new_n359_, new_n358_, new_n356_ );
nor  ( new_n360_, new_n359_, new_n353_ );
or   ( new_n361_, new_n360_, new_n351_ );
and  ( new_n362_, new_n361_, new_n350_ );
nor  ( new_n363_, new_n362_, new_n341_ );
nor  ( new_n364_, new_n363_, new_n339_ );
xor  ( new_n365_, new_n286_, new_n285_ );
xor  ( new_n366_, new_n365_, new_n364_ );
xnor ( new_n367_, new_n297_, new_n294_ );
xor  ( new_n368_, new_n367_, new_n301_ );
xor  ( new_n369_, new_n368_, new_n366_ );
nor  ( new_n370_, new_n369_, new_n321_ );
and  ( new_n371_, new_n369_, new_n321_ );
xor  ( new_n372_, new_n223_, new_n222_ );
xnor ( new_n373_, new_n241_, new_n234_ );
nand ( new_n374_, new_n373_, new_n247_ );
not  ( new_n375_, new_n249_ );
or   ( new_n376_, new_n375_, new_n242_ );
and  ( new_n377_, new_n376_, new_n374_ );
and  ( new_n378_, new_n377_, new_n372_ );
xnor ( new_n379_, new_n377_, new_n372_ );
xor  ( new_n380_, \d[5] , \a[6]  );
nand ( new_n381_, new_n380_, new_n69_ );
not  ( new_n382_, new_n68_ );
or   ( new_n383_, new_n335_, new_n382_ );
and  ( new_n384_, new_n383_, new_n381_ );
nand ( new_n385_, new_n243_, new_n77_ );
and  ( new_n386_, new_n326_, \d[11]  );
and  ( new_n387_, \d[10] , \a[0]  );
nor  ( new_n388_, new_n387_, new_n386_ );
and  ( new_n389_, \d[11] , \a[0]  );
or   ( new_n390_, new_n389_, new_n77_ );
or   ( new_n391_, new_n390_, new_n388_ );
and  ( new_n392_, new_n391_, new_n385_ );
or   ( new_n393_, new_n392_, new_n384_ );
and  ( new_n394_, new_n392_, new_n384_ );
xnor ( new_n395_, new_n331_, new_n325_ );
or   ( new_n396_, new_n395_, new_n394_ );
and  ( new_n397_, new_n396_, new_n393_ );
nor  ( new_n398_, new_n397_, new_n379_ );
nor  ( new_n399_, new_n398_, new_n378_ );
nor  ( new_n400_, new_n399_, new_n371_ );
nor  ( new_n401_, new_n400_, new_n370_ );
xor  ( new_n402_, new_n304_, new_n291_ );
xor  ( new_n403_, new_n206_, new_n204_ );
xor  ( new_n404_, new_n403_, new_n252_ );
xor  ( new_n405_, new_n404_, new_n402_ );
not  ( new_n406_, new_n364_ );
and  ( new_n407_, new_n365_, new_n406_ );
or   ( new_n408_, new_n365_, new_n406_ );
and  ( new_n409_, new_n368_, new_n408_ );
nor  ( new_n410_, new_n409_, new_n407_ );
xor  ( new_n411_, new_n410_, new_n405_ );
nor  ( new_n412_, new_n411_, new_n401_ );
and  ( new_n413_, new_n411_, new_n401_ );
xor  ( new_n414_, new_n362_, new_n341_ );
not  ( new_n415_, new_n414_ );
or   ( new_n416_, new_n346_, new_n180_ );
xor  ( new_n417_, \d[9] , \a[1]  );
nand ( new_n418_, new_n417_, new_n174_ );
and  ( new_n419_, new_n418_, new_n416_ );
or   ( new_n420_, new_n235_, \a[9]  );
and  ( new_n421_, new_n90_, new_n352_ );
and  ( new_n422_, \d[1] , \a[10]  );
or   ( new_n423_, new_n422_, new_n86_ );
or   ( new_n424_, new_n423_, new_n421_ );
and  ( new_n425_, new_n424_, new_n420_ );
nor  ( new_n426_, new_n425_, new_n419_ );
xor  ( new_n427_, \d[5] , \a[5]  );
and  ( new_n428_, new_n427_, new_n69_ );
and  ( new_n429_, new_n380_, new_n68_ );
nor  ( new_n430_, new_n429_, new_n428_ );
and  ( new_n431_, new_n425_, new_n419_ );
nor  ( new_n432_, new_n431_, new_n430_ );
or   ( new_n433_, new_n432_, new_n426_ );
xnor ( new_n434_, new_n349_, new_n345_ );
xor  ( new_n435_, new_n434_, new_n360_ );
nand ( new_n436_, new_n435_, new_n433_ );
nor  ( new_n437_, new_n435_, new_n433_ );
xor  ( new_n438_, \d[3] , \a[7]  );
and  ( new_n439_, new_n438_, new_n153_ );
and  ( new_n440_, new_n322_, new_n152_ );
or   ( new_n441_, new_n440_, new_n439_ );
and  ( new_n442_, new_n77_, \a[0]  );
and  ( new_n443_, new_n442_, new_n441_ );
nor  ( new_n444_, new_n442_, new_n441_ );
xor  ( new_n445_, \d[7] , \a[3]  );
and  ( new_n446_, new_n445_, new_n131_ );
and  ( new_n447_, new_n342_, new_n130_ );
nor  ( new_n448_, new_n447_, new_n446_ );
nor  ( new_n449_, new_n448_, new_n444_ );
nor  ( new_n450_, new_n449_, new_n443_ );
or   ( new_n451_, new_n450_, new_n437_ );
and  ( new_n452_, new_n451_, new_n436_ );
nor  ( new_n453_, new_n452_, new_n415_ );
xor  ( new_n454_, new_n452_, new_n415_ );
xor  ( new_n455_, new_n397_, new_n379_ );
and  ( new_n456_, new_n455_, new_n454_ );
or   ( new_n457_, new_n456_, new_n453_ );
xnor ( new_n458_, new_n369_, new_n321_ );
xor  ( new_n459_, new_n458_, new_n399_ );
nor  ( new_n460_, new_n459_, new_n457_ );
and  ( new_n461_, new_n459_, new_n457_ );
xor  ( new_n462_, new_n455_, new_n454_ );
not  ( new_n463_, new_n462_ );
xor  ( new_n464_, new_n392_, new_n384_ );
xor  ( new_n465_, new_n464_, new_n395_ );
xor  ( new_n466_, \d[3] , \a[6]  );
and  ( new_n467_, new_n466_, new_n153_ );
and  ( new_n468_, new_n438_, new_n152_ );
or   ( new_n469_, new_n468_, new_n467_ );
and  ( new_n470_, new_n128_, new_n98_ );
or   ( new_n471_, new_n470_, new_n179_ );
and  ( new_n472_, \d[7] , \a[0]  );
not  ( new_n473_, new_n472_ );
and  ( new_n474_, new_n473_, \d[9]  );
and  ( new_n475_, new_n474_, new_n471_ );
and  ( new_n476_, new_n475_, new_n469_ );
xnor ( new_n477_, new_n442_, new_n441_ );
xor  ( new_n478_, new_n477_, new_n448_ );
nand ( new_n479_, new_n478_, new_n476_ );
nor  ( new_n480_, new_n478_, new_n476_ );
xor  ( new_n481_, \d[7] , \a[2]  );
and  ( new_n482_, new_n481_, new_n131_ );
and  ( new_n483_, new_n445_, new_n130_ );
nor  ( new_n484_, new_n483_, new_n482_ );
or   ( new_n485_, new_n235_, \a[8]  );
and  ( new_n486_, new_n90_, new_n137_ );
and  ( new_n487_, \d[1] , \a[9]  );
or   ( new_n488_, new_n487_, new_n86_ );
or   ( new_n489_, new_n488_, new_n486_ );
and  ( new_n490_, new_n489_, new_n485_ );
nor  ( new_n491_, new_n490_, new_n484_ );
and  ( new_n492_, new_n490_, new_n484_ );
and  ( new_n493_, new_n417_, new_n181_ );
xor  ( new_n494_, \d[9] , \a[0]  );
and  ( new_n495_, new_n494_, new_n174_ );
nor  ( new_n496_, new_n495_, new_n493_ );
nor  ( new_n497_, new_n496_, new_n492_ );
nor  ( new_n498_, new_n497_, new_n491_ );
or   ( new_n499_, new_n498_, new_n480_ );
and  ( new_n500_, new_n499_, new_n479_ );
or   ( new_n501_, new_n500_, new_n465_ );
nand ( new_n502_, new_n500_, new_n465_ );
xor  ( new_n503_, new_n435_, new_n433_ );
xnor ( new_n504_, new_n503_, new_n450_ );
nand ( new_n505_, new_n504_, new_n502_ );
and  ( new_n506_, new_n505_, new_n501_ );
nor  ( new_n507_, new_n506_, new_n463_ );
and  ( new_n508_, new_n506_, new_n463_ );
xor  ( new_n509_, \d[5] , \a[4]  );
and  ( new_n510_, new_n509_, new_n69_ );
and  ( new_n511_, new_n427_, new_n68_ );
or   ( new_n512_, new_n511_, new_n510_ );
xor  ( new_n513_, new_n475_, new_n469_ );
nor  ( new_n514_, new_n513_, new_n512_ );
or   ( new_n515_, new_n180_, new_n98_ );
or   ( new_n516_, new_n235_, \a[7]  );
and  ( new_n517_, new_n90_, new_n133_ );
and  ( new_n518_, \d[1] , \a[8]  );
or   ( new_n519_, new_n518_, new_n86_ );
or   ( new_n520_, new_n519_, new_n517_ );
and  ( new_n521_, new_n520_, new_n516_ );
and  ( new_n522_, new_n521_, new_n515_ );
xor  ( new_n523_, \d[7] , \a[1]  );
nand ( new_n524_, new_n523_, new_n131_ );
nand ( new_n525_, new_n481_, new_n130_ );
and  ( new_n526_, new_n525_, new_n524_ );
xor  ( new_n527_, new_n521_, new_n515_ );
and  ( new_n528_, new_n527_, new_n526_ );
or   ( new_n529_, new_n528_, new_n522_ );
xor  ( new_n530_, new_n513_, new_n512_ );
and  ( new_n531_, new_n530_, new_n529_ );
nor  ( new_n532_, new_n531_, new_n514_ );
xnor ( new_n533_, new_n425_, new_n419_ );
nand ( new_n534_, new_n533_, new_n430_ );
not  ( new_n535_, new_n426_ );
nand ( new_n536_, new_n432_, new_n535_ );
and  ( new_n537_, new_n536_, new_n534_ );
nor  ( new_n538_, new_n537_, new_n532_ );
xor  ( new_n539_, new_n537_, new_n532_ );
not  ( new_n540_, new_n539_ );
xnor ( new_n541_, new_n478_, new_n476_ );
xor  ( new_n542_, new_n541_, new_n498_ );
nor  ( new_n543_, new_n542_, new_n540_ );
nor  ( new_n544_, new_n543_, new_n538_ );
xor  ( new_n545_, new_n500_, new_n465_ );
xor  ( new_n546_, new_n545_, new_n504_ );
and  ( new_n547_, new_n546_, new_n544_ );
nor  ( new_n548_, new_n546_, new_n544_ );
xor  ( new_n549_, new_n542_, new_n540_ );
xnor ( new_n550_, new_n490_, new_n484_ );
and  ( new_n551_, new_n550_, new_n496_ );
not  ( new_n552_, new_n491_ );
and  ( new_n553_, new_n497_, new_n552_ );
or   ( new_n554_, new_n553_, new_n551_ );
and  ( new_n555_, new_n87_, new_n212_ );
and  ( new_n556_, new_n90_, new_n185_ );
not  ( new_n557_, new_n556_ );
and  ( new_n558_, \d[1] , \a[7]  );
nor  ( new_n559_, new_n558_, new_n86_ );
and  ( new_n560_, new_n559_, new_n557_ );
nor  ( new_n561_, new_n560_, new_n555_ );
not  ( new_n562_, new_n561_ );
not  ( new_n563_, \d[6]  );
and  ( new_n564_, new_n66_, new_n563_ );
or   ( new_n565_, new_n564_, new_n98_ );
or   ( new_n566_, new_n66_, new_n563_ );
and  ( new_n567_, new_n566_, \d[7]  );
and  ( new_n568_, new_n567_, new_n565_ );
nand ( new_n569_, new_n568_, new_n562_ );
xor  ( new_n570_, \d[5] , new_n163_ );
or   ( new_n571_, new_n570_, new_n334_ );
nand ( new_n572_, new_n509_, new_n68_ );
and  ( new_n573_, new_n572_, new_n571_ );
or   ( new_n574_, new_n573_, new_n569_ );
and  ( new_n575_, new_n573_, new_n569_ );
xor  ( new_n576_, \d[3] , \a[5]  );
and  ( new_n577_, new_n576_, new_n153_ );
and  ( new_n578_, new_n466_, new_n152_ );
nor  ( new_n579_, new_n578_, new_n577_ );
or   ( new_n580_, new_n579_, new_n575_ );
and  ( new_n581_, new_n580_, new_n574_ );
or   ( new_n582_, new_n581_, new_n554_ );
and  ( new_n583_, new_n581_, new_n554_ );
xor  ( new_n584_, new_n530_, new_n529_ );
or   ( new_n585_, new_n584_, new_n583_ );
and  ( new_n586_, new_n585_, new_n582_ );
nor  ( new_n587_, new_n586_, new_n549_ );
and  ( new_n588_, new_n586_, new_n549_ );
xor  ( new_n589_, new_n527_, new_n526_ );
xor  ( new_n590_, \d[3] , \a[4]  );
nand ( new_n591_, new_n590_, new_n153_ );
nand ( new_n592_, new_n576_, new_n152_ );
and  ( new_n593_, new_n592_, new_n591_ );
xor  ( new_n594_, \d[5] , new_n115_ );
or   ( new_n595_, new_n594_, new_n334_ );
or   ( new_n596_, new_n570_, new_n382_ );
and  ( new_n597_, new_n596_, new_n595_ );
nor  ( new_n598_, new_n597_, new_n593_ );
and  ( new_n599_, new_n597_, new_n593_ );
and  ( new_n600_, new_n523_, new_n130_ );
and  ( new_n601_, new_n563_, \d[7]  );
and  ( new_n602_, \d[6] , \a[0]  );
nor  ( new_n603_, new_n602_, new_n601_ );
not  ( new_n604_, new_n603_ );
and  ( new_n605_, new_n473_, new_n136_ );
and  ( new_n606_, new_n605_, new_n604_ );
nor  ( new_n607_, new_n606_, new_n600_ );
nor  ( new_n608_, new_n607_, new_n599_ );
nor  ( new_n609_, new_n608_, new_n598_ );
and  ( new_n610_, new_n609_, new_n589_ );
nor  ( new_n611_, new_n609_, new_n589_ );
xor  ( new_n612_, new_n573_, new_n569_ );
xnor ( new_n613_, new_n612_, new_n579_ );
nor  ( new_n614_, new_n613_, new_n611_ );
nor  ( new_n615_, new_n614_, new_n610_ );
not  ( new_n616_, new_n615_ );
xor  ( new_n617_, new_n581_, new_n554_ );
xor  ( new_n618_, new_n617_, new_n584_ );
nor  ( new_n619_, new_n618_, new_n616_ );
and  ( new_n620_, new_n618_, new_n616_ );
xor  ( new_n621_, new_n568_, new_n562_ );
not  ( new_n622_, new_n621_ );
or   ( new_n623_, new_n136_, new_n98_ );
or   ( new_n624_, new_n235_, \a[5]  );
and  ( new_n625_, new_n90_, new_n212_ );
and  ( new_n626_, \d[1] , \a[6]  );
or   ( new_n627_, new_n626_, new_n86_ );
or   ( new_n628_, new_n627_, new_n625_ );
and  ( new_n629_, new_n628_, new_n624_ );
or   ( new_n630_, new_n629_, new_n623_ );
and  ( new_n631_, new_n629_, new_n623_ );
xor  ( new_n632_, \d[3] , \a[3]  );
and  ( new_n633_, new_n632_, new_n153_ );
and  ( new_n634_, new_n590_, new_n152_ );
nor  ( new_n635_, new_n634_, new_n633_ );
or   ( new_n636_, new_n635_, new_n631_ );
and  ( new_n637_, new_n636_, new_n630_ );
and  ( new_n638_, new_n637_, new_n622_ );
xor  ( new_n639_, new_n637_, new_n622_ );
not  ( new_n640_, new_n639_ );
xnor ( new_n641_, new_n597_, new_n593_ );
nand ( new_n642_, new_n641_, new_n607_ );
not  ( new_n643_, new_n608_ );
or   ( new_n644_, new_n643_, new_n598_ );
and  ( new_n645_, new_n644_, new_n642_ );
nor  ( new_n646_, new_n645_, new_n640_ );
nor  ( new_n647_, new_n646_, new_n638_ );
not  ( new_n648_, new_n647_ );
xnor ( new_n649_, new_n609_, new_n589_ );
xor  ( new_n650_, new_n649_, new_n613_ );
nor  ( new_n651_, new_n650_, new_n648_ );
and  ( new_n652_, new_n650_, new_n648_ );
xor  ( new_n653_, new_n645_, new_n640_ );
and  ( new_n654_, new_n87_, new_n231_ );
or   ( new_n655_, \d[1] , \a[5]  );
and  ( new_n656_, \d[1] , \a[5]  );
nor  ( new_n657_, new_n656_, new_n86_ );
and  ( new_n658_, new_n657_, new_n655_ );
or   ( new_n659_, new_n658_, new_n654_ );
not  ( new_n660_, \d[4]  );
and  ( new_n661_, new_n150_, new_n660_ );
or   ( new_n662_, new_n661_, new_n98_ );
or   ( new_n663_, new_n150_, new_n660_ );
and  ( new_n664_, new_n663_, \d[5]  );
and  ( new_n665_, new_n664_, new_n662_ );
nand ( new_n666_, new_n665_, new_n659_ );
xor  ( new_n667_, \d[5] , new_n108_ );
or   ( new_n668_, new_n667_, new_n334_ );
or   ( new_n669_, new_n594_, new_n382_ );
and  ( new_n670_, new_n669_, new_n668_ );
or   ( new_n671_, new_n670_, new_n666_ );
nand ( new_n672_, new_n670_, new_n666_ );
xor  ( new_n673_, new_n629_, new_n623_ );
xnor ( new_n674_, new_n673_, new_n635_ );
nand ( new_n675_, new_n674_, new_n672_ );
and  ( new_n676_, new_n675_, new_n671_ );
nor  ( new_n677_, new_n676_, new_n653_ );
and  ( new_n678_, new_n676_, new_n653_ );
xor  ( new_n679_, \d[3] , \a[2]  );
and  ( new_n680_, new_n679_, new_n153_ );
and  ( new_n681_, new_n632_, new_n152_ );
nor  ( new_n682_, new_n681_, new_n680_ );
or   ( new_n683_, new_n667_, new_n382_ );
and  ( new_n684_, new_n660_, \d[5]  );
and  ( new_n685_, \d[4] , \a[0]  );
nor  ( new_n686_, new_n685_, new_n684_ );
and  ( new_n687_, \d[5] , \a[0]  );
or   ( new_n688_, new_n687_, new_n68_ );
or   ( new_n689_, new_n688_, new_n686_ );
and  ( new_n690_, new_n689_, new_n683_ );
nor  ( new_n691_, new_n690_, new_n682_ );
xor  ( new_n692_, new_n690_, new_n682_ );
xor  ( new_n693_, new_n665_, new_n659_ );
and  ( new_n694_, new_n693_, new_n692_ );
nor  ( new_n695_, new_n694_, new_n691_ );
not  ( new_n696_, new_n695_ );
xor  ( new_n697_, new_n670_, new_n666_ );
xor  ( new_n698_, new_n697_, new_n674_ );
and  ( new_n699_, new_n698_, new_n696_ );
xor  ( new_n700_, new_n698_, new_n696_ );
xnor ( new_n701_, new_n693_, new_n692_ );
or   ( new_n702_, new_n382_, new_n98_ );
or   ( new_n703_, new_n235_, \a[3]  );
and  ( new_n704_, new_n90_, new_n231_ );
and  ( new_n705_, \d[1] , \a[4]  );
or   ( new_n706_, new_n705_, new_n86_ );
or   ( new_n707_, new_n706_, new_n704_ );
and  ( new_n708_, new_n707_, new_n703_ );
or   ( new_n709_, new_n708_, new_n702_ );
and  ( new_n710_, new_n708_, new_n702_ );
xor  ( new_n711_, \d[3] , \a[1]  );
and  ( new_n712_, new_n711_, new_n153_ );
and  ( new_n713_, new_n679_, new_n152_ );
nor  ( new_n714_, new_n713_, new_n712_ );
or   ( new_n715_, new_n714_, new_n710_ );
and  ( new_n716_, new_n715_, new_n709_ );
or   ( new_n717_, new_n716_, new_n701_ );
and  ( new_n718_, new_n716_, new_n701_ );
and  ( new_n719_, new_n87_, new_n115_ );
and  ( new_n720_, new_n90_, new_n163_ );
not  ( new_n721_, new_n720_ );
and  ( new_n722_, \d[1] , \a[3]  );
nor  ( new_n723_, new_n722_, new_n86_ );
and  ( new_n724_, new_n723_, new_n721_ );
nor  ( new_n725_, new_n724_, new_n719_ );
not  ( new_n726_, \d[2]  );
and  ( new_n727_, new_n90_, new_n726_ );
or   ( new_n728_, new_n727_, new_n98_ );
or   ( new_n729_, new_n90_, new_n726_ );
and  ( new_n730_, new_n729_, \d[3]  );
nand ( new_n731_, new_n730_, new_n728_ );
nor  ( new_n732_, new_n731_, new_n725_ );
xnor ( new_n733_, new_n708_, new_n702_ );
xor  ( new_n734_, new_n733_, new_n714_ );
and  ( new_n735_, new_n734_, new_n732_ );
nor  ( new_n736_, new_n734_, new_n732_ );
xnor ( new_n737_, new_n731_, new_n725_ );
nand ( new_n738_, new_n711_, new_n152_ );
and  ( new_n739_, new_n726_, \d[3]  );
and  ( new_n740_, \d[2] , \a[0]  );
nor  ( new_n741_, new_n740_, new_n739_ );
and  ( new_n742_, \d[3] , \a[0]  );
or   ( new_n743_, new_n742_, new_n152_ );
or   ( new_n744_, new_n743_, new_n741_ );
and  ( new_n745_, new_n744_, new_n738_ );
nor  ( new_n746_, new_n745_, new_n737_ );
and  ( new_n747_, new_n745_, new_n737_ );
or   ( new_n748_, new_n312_, new_n98_ );
or   ( new_n749_, new_n235_, \a[1]  );
and  ( new_n750_, new_n90_, new_n115_ );
and  ( new_n751_, \d[1] , \a[2]  );
or   ( new_n752_, new_n751_, new_n86_ );
or   ( new_n753_, new_n752_, new_n750_ );
and  ( new_n754_, new_n753_, new_n749_ );
nor  ( new_n755_, new_n754_, new_n748_ );
and  ( new_n756_, new_n754_, new_n748_ );
and  ( new_n757_, \d[0] , \a[1]  );
not  ( new_n758_, new_n757_ );
and  ( new_n759_, \d[1] , new_n98_ );
and  ( new_n760_, new_n759_, new_n758_ );
not  ( new_n761_, new_n760_ );
nor  ( new_n762_, new_n761_, new_n756_ );
nor  ( new_n763_, new_n762_, new_n755_ );
nor  ( new_n764_, new_n763_, new_n747_ );
nor  ( new_n765_, new_n764_, new_n746_ );
nor  ( new_n766_, new_n765_, new_n736_ );
nor  ( new_n767_, new_n766_, new_n735_ );
or   ( new_n768_, new_n767_, new_n718_ );
nand ( new_n769_, new_n768_, new_n717_ );
and  ( new_n770_, new_n769_, new_n700_ );
nor  ( new_n771_, new_n770_, new_n699_ );
nor  ( new_n772_, new_n771_, new_n678_ );
nor  ( new_n773_, new_n772_, new_n677_ );
nor  ( new_n774_, new_n773_, new_n652_ );
nor  ( new_n775_, new_n774_, new_n651_ );
nor  ( new_n776_, new_n775_, new_n620_ );
nor  ( new_n777_, new_n776_, new_n619_ );
nor  ( new_n778_, new_n777_, new_n588_ );
nor  ( new_n779_, new_n778_, new_n587_ );
nor  ( new_n780_, new_n779_, new_n548_ );
nor  ( new_n781_, new_n780_, new_n547_ );
nor  ( new_n782_, new_n781_, new_n508_ );
nor  ( new_n783_, new_n782_, new_n507_ );
not  ( new_n784_, new_n783_ );
nor  ( new_n785_, new_n784_, new_n461_ );
nor  ( new_n786_, new_n785_, new_n460_ );
not  ( new_n787_, new_n786_ );
nor  ( new_n788_, new_n787_, new_n413_ );
nor  ( new_n789_, new_n788_, new_n412_ );
and  ( new_n790_, new_n404_, new_n402_ );
nor  ( new_n791_, new_n404_, new_n402_ );
nor  ( new_n792_, new_n410_, new_n791_ );
or   ( new_n793_, new_n792_, new_n790_ );
or   ( new_n794_, new_n257_, new_n103_ );
and  ( new_n795_, new_n260_, \d[15]  );
and  ( new_n796_, new_n795_, new_n794_ );
xor  ( new_n797_, new_n796_, new_n793_ );
xnor ( new_n798_, new_n797_, new_n789_ );
and  ( new_n799_, new_n798_, new_n319_ );
not  ( new_n800_, new_n799_ );
xor  ( new_n801_, \b[3] , \b[4]  );
not  ( new_n802_, new_n801_ );
or   ( new_n803_, new_n802_, new_n98_ );
not  ( new_n804_, \b[0]  );
and  ( new_n805_, new_n804_, \b[1]  );
not  ( new_n806_, new_n805_ );
or   ( new_n807_, new_n806_, \a[3]  );
not  ( new_n808_, \b[1]  );
and  ( new_n809_, new_n808_, new_n231_ );
and  ( new_n810_, \b[1] , \a[4]  );
or   ( new_n811_, new_n810_, new_n804_ );
or   ( new_n812_, new_n811_, new_n809_ );
and  ( new_n813_, new_n812_, new_n807_ );
or   ( new_n814_, new_n813_, new_n803_ );
not  ( new_n815_, \b[3]  );
xor  ( new_n816_, \b[2] , new_n815_ );
xor  ( new_n817_, \b[1] , \b[2]  );
nor  ( new_n818_, new_n817_, new_n816_ );
xor  ( new_n819_, \b[3] , \a[1]  );
nand ( new_n820_, new_n819_, new_n818_ );
xor  ( new_n821_, \b[3] , \a[2]  );
nand ( new_n822_, new_n821_, new_n817_ );
and  ( new_n823_, new_n822_, new_n820_ );
and  ( new_n824_, new_n813_, new_n803_ );
or   ( new_n825_, new_n824_, new_n823_ );
and  ( new_n826_, new_n825_, new_n814_ );
and  ( new_n827_, new_n821_, new_n818_ );
xor  ( new_n828_, \b[3] , \a[3]  );
and  ( new_n829_, new_n828_, new_n817_ );
nor  ( new_n830_, new_n829_, new_n827_ );
not  ( new_n831_, new_n830_ );
not  ( new_n832_, \b[4]  );
and  ( new_n833_, new_n815_, new_n832_ );
or   ( new_n834_, new_n833_, new_n98_ );
or   ( new_n835_, new_n815_, new_n832_ );
and  ( new_n836_, new_n835_, \b[5]  );
and  ( new_n837_, new_n836_, new_n834_ );
xor  ( new_n838_, new_n837_, new_n831_ );
or   ( new_n839_, new_n806_, \a[4]  );
and  ( new_n840_, new_n808_, new_n176_ );
and  ( new_n841_, \b[1] , \a[5]  );
or   ( new_n842_, new_n841_, new_n804_ );
or   ( new_n843_, new_n842_, new_n840_ );
and  ( new_n844_, new_n843_, new_n839_ );
xor  ( new_n845_, \b[5] , new_n108_ );
or   ( new_n846_, new_n845_, new_n802_ );
not  ( new_n847_, \b[5]  );
xor  ( new_n848_, \b[4] , new_n847_ );
nor  ( new_n849_, new_n848_, new_n801_ );
not  ( new_n850_, new_n849_ );
xor  ( new_n851_, \b[5] , new_n98_ );
or   ( new_n852_, new_n851_, new_n850_ );
and  ( new_n853_, new_n852_, new_n846_ );
xnor ( new_n854_, new_n853_, new_n844_ );
xor  ( new_n855_, new_n854_, new_n838_ );
nor  ( new_n856_, new_n855_, new_n826_ );
and  ( new_n857_, new_n855_, new_n826_ );
and  ( new_n858_, new_n805_, new_n115_ );
and  ( new_n859_, new_n808_, new_n163_ );
not  ( new_n860_, new_n859_ );
and  ( new_n861_, \b[1] , \a[3]  );
nor  ( new_n862_, new_n861_, new_n804_ );
and  ( new_n863_, new_n862_, new_n860_ );
nor  ( new_n864_, new_n863_, new_n858_ );
not  ( new_n865_, \b[2]  );
and  ( new_n866_, new_n808_, new_n865_ );
or   ( new_n867_, new_n866_, new_n98_ );
or   ( new_n868_, new_n808_, new_n865_ );
and  ( new_n869_, new_n868_, \b[3]  );
nand ( new_n870_, new_n869_, new_n867_ );
or   ( new_n871_, new_n870_, new_n864_ );
xor  ( new_n872_, new_n813_, new_n803_ );
xor  ( new_n873_, new_n872_, new_n823_ );
nor  ( new_n874_, new_n873_, new_n871_ );
and  ( new_n875_, new_n873_, new_n871_ );
xnor ( new_n876_, new_n870_, new_n864_ );
nand ( new_n877_, new_n819_, new_n817_ );
or   ( new_n878_, \b[2] , new_n815_ );
and  ( new_n879_, \b[2] , \a[0]  );
not  ( new_n880_, new_n879_ );
and  ( new_n881_, new_n880_, new_n878_ );
and  ( new_n882_, \b[3] , \a[0]  );
or   ( new_n883_, new_n882_, new_n817_ );
or   ( new_n884_, new_n883_, new_n881_ );
and  ( new_n885_, new_n884_, new_n877_ );
nor  ( new_n886_, new_n885_, new_n876_ );
and  ( new_n887_, new_n885_, new_n876_ );
and  ( new_n888_, new_n805_, new_n108_ );
and  ( new_n889_, new_n808_, new_n115_ );
not  ( new_n890_, new_n889_ );
and  ( new_n891_, \b[1] , \a[2]  );
nor  ( new_n892_, new_n891_, new_n804_ );
and  ( new_n893_, new_n892_, new_n890_ );
nor  ( new_n894_, new_n893_, new_n888_ );
not  ( new_n895_, new_n817_ );
or   ( new_n896_, new_n895_, new_n98_ );
and  ( new_n897_, \b[0] , \a[1]  );
or   ( new_n898_, new_n808_, \a[0]  );
or   ( new_n899_, new_n898_, new_n897_ );
and  ( new_n900_, new_n899_, new_n896_ );
nor  ( new_n901_, new_n900_, new_n894_ );
not  ( new_n902_, new_n901_ );
nor  ( new_n903_, new_n902_, new_n887_ );
nor  ( new_n904_, new_n903_, new_n886_ );
nor  ( new_n905_, new_n904_, new_n875_ );
nor  ( new_n906_, new_n905_, new_n874_ );
nor  ( new_n907_, new_n906_, new_n857_ );
nor  ( new_n908_, new_n907_, new_n856_ );
nor  ( new_n909_, new_n853_, new_n844_ );
nand ( new_n910_, new_n853_, new_n844_ );
and  ( new_n911_, new_n910_, new_n838_ );
or   ( new_n912_, new_n911_, new_n909_ );
and  ( new_n913_, new_n828_, new_n818_ );
xor  ( new_n914_, \b[3] , \a[4]  );
and  ( new_n915_, new_n914_, new_n817_ );
nor  ( new_n916_, new_n915_, new_n913_ );
not  ( new_n917_, new_n916_ );
xor  ( new_n918_, \b[5] , \b[6]  );
not  ( new_n919_, new_n918_ );
or   ( new_n920_, new_n919_, new_n98_ );
or   ( new_n921_, new_n850_, new_n845_ );
xor  ( new_n922_, \b[5] , \a[2]  );
nand ( new_n923_, new_n922_, new_n801_ );
and  ( new_n924_, new_n923_, new_n921_ );
xor  ( new_n925_, new_n924_, new_n920_ );
xor  ( new_n926_, new_n925_, new_n917_ );
nand ( new_n927_, new_n837_, new_n831_ );
or   ( new_n928_, new_n806_, \a[5]  );
and  ( new_n929_, new_n808_, new_n212_ );
and  ( new_n930_, \b[1] , \a[6]  );
or   ( new_n931_, new_n930_, new_n804_ );
or   ( new_n932_, new_n931_, new_n929_ );
and  ( new_n933_, new_n932_, new_n928_ );
xor  ( new_n934_, new_n933_, new_n927_ );
xor  ( new_n935_, new_n934_, new_n926_ );
xor  ( new_n936_, new_n935_, new_n912_ );
xnor ( new_n937_, new_n936_, new_n908_ );
not  ( new_n938_, new_n937_ );
nor  ( new_n939_, new_n798_, new_n319_ );
nor  ( new_n940_, new_n939_, new_n938_ );
and  ( new_n941_, new_n940_, new_n800_ );
not  ( new_n942_, new_n941_ );
not  ( new_n943_, \c[5]  );
xor  ( new_n944_, \c[4] , new_n943_ );
xor  ( new_n945_, \c[3] , \c[4]  );
nor  ( new_n946_, new_n945_, new_n944_ );
xor  ( new_n947_, \c[5] , \b[8]  );
and  ( new_n948_, new_n947_, new_n946_ );
xor  ( new_n949_, \c[5] , \b[9]  );
and  ( new_n950_, new_n949_, new_n945_ );
nor  ( new_n951_, new_n950_, new_n948_ );
not  ( new_n952_, \c[11]  );
xor  ( new_n953_, \c[10] , new_n952_ );
xor  ( new_n954_, \c[9] , \c[10]  );
nor  ( new_n955_, new_n954_, new_n953_ );
xor  ( new_n956_, \c[11] , \b[2]  );
nand ( new_n957_, new_n956_, new_n955_ );
not  ( new_n958_, new_n954_ );
xor  ( new_n959_, \c[11] , new_n815_ );
or   ( new_n960_, new_n959_, new_n958_ );
and  ( new_n961_, new_n960_, new_n957_ );
or   ( new_n962_, new_n961_, new_n951_ );
xnor ( new_n963_, new_n961_, new_n951_ );
xor  ( new_n964_, \c[11] , \c[12]  );
not  ( new_n965_, new_n964_ );
xor  ( new_n966_, \c[13] , new_n808_ );
or   ( new_n967_, new_n966_, new_n965_ );
and  ( new_n968_, \c[12] , \b[0]  );
not  ( new_n969_, \c[12]  );
and  ( new_n970_, new_n969_, \c[13]  );
nor  ( new_n971_, new_n970_, new_n968_ );
and  ( new_n972_, \c[13] , \b[0]  );
or   ( new_n973_, new_n972_, new_n964_ );
or   ( new_n974_, new_n973_, new_n971_ );
and  ( new_n975_, new_n974_, new_n967_ );
or   ( new_n976_, new_n975_, new_n963_ );
nand ( new_n977_, new_n976_, new_n962_ );
not  ( new_n978_, \c[3]  );
xor  ( new_n979_, \c[2] , new_n978_ );
xor  ( new_n980_, \c[1] , \c[2]  );
nor  ( new_n981_, new_n980_, new_n979_ );
xor  ( new_n982_, \c[3] , \b[11]  );
and  ( new_n983_, new_n982_, new_n981_ );
xor  ( new_n984_, \c[3] , \b[12]  );
and  ( new_n985_, new_n984_, new_n980_ );
or   ( new_n986_, new_n985_, new_n983_ );
xor  ( new_n987_, \c[13] , \c[14]  );
and  ( new_n988_, new_n987_, \b[0]  );
not  ( new_n989_, new_n988_ );
xor  ( new_n990_, \c[1] , \b[14]  );
and  ( new_n991_, new_n990_, \c[0]  );
not  ( new_n992_, \b[13]  );
not  ( new_n993_, \c[0]  );
and  ( new_n994_, new_n993_, \c[1]  );
and  ( new_n995_, new_n994_, new_n992_ );
nor  ( new_n996_, new_n995_, new_n991_ );
xor  ( new_n997_, new_n996_, new_n989_ );
xor  ( new_n998_, new_n997_, new_n986_ );
xnor ( new_n999_, new_n998_, new_n977_ );
not  ( new_n1000_, \c[7]  );
and  ( new_n1001_, new_n1000_, \c[8]  );
and  ( new_n1002_, new_n1000_, \c[9]  );
not  ( new_n1003_, \c[9]  );
and  ( new_n1004_, \c[8] , new_n1003_ );
nor  ( new_n1005_, new_n1004_, new_n1002_ );
nor  ( new_n1006_, new_n1005_, new_n1001_ );
not  ( new_n1007_, new_n1006_ );
xor  ( new_n1008_, \c[9] , new_n832_ );
or   ( new_n1009_, new_n1008_, new_n1007_ );
not  ( new_n1010_, \c[8]  );
xor  ( new_n1011_, \c[7] , new_n1010_ );
xor  ( new_n1012_, \c[9] , new_n847_ );
or   ( new_n1013_, new_n1012_, new_n1011_ );
and  ( new_n1014_, new_n1013_, new_n1009_ );
xor  ( new_n1015_, \c[6] , new_n1000_ );
xor  ( new_n1016_, \c[5] , \c[6]  );
nor  ( new_n1017_, new_n1016_, new_n1015_ );
not  ( new_n1018_, new_n1017_ );
not  ( new_n1019_, \b[6]  );
xor  ( new_n1020_, \c[7] , new_n1019_ );
or   ( new_n1021_, new_n1020_, new_n1018_ );
not  ( new_n1022_, new_n1016_ );
not  ( new_n1023_, \b[7]  );
xor  ( new_n1024_, \c[7] , new_n1023_ );
or   ( new_n1025_, new_n1024_, new_n1022_ );
and  ( new_n1026_, new_n1025_, new_n1021_ );
or   ( new_n1027_, new_n1026_, new_n1014_ );
xor  ( new_n1028_, \c[3] , \b[10]  );
nand ( new_n1029_, new_n1028_, new_n981_ );
nand ( new_n1030_, new_n982_, new_n980_ );
and  ( new_n1031_, new_n1030_, new_n1029_ );
and  ( new_n1032_, new_n1026_, new_n1014_ );
or   ( new_n1033_, new_n1032_, new_n1031_ );
and  ( new_n1034_, new_n1033_, new_n1027_ );
xnor ( new_n1035_, new_n1034_, new_n999_ );
nand ( new_n1036_, new_n949_, new_n946_ );
not  ( new_n1037_, new_n945_ );
not  ( new_n1038_, \b[10]  );
xor  ( new_n1039_, \c[5] , new_n1038_ );
or   ( new_n1040_, new_n1039_, new_n1037_ );
nand ( new_n1041_, new_n1040_, new_n1036_ );
not  ( new_n1042_, new_n1011_ );
xor  ( new_n1043_, \c[9] , \b[6]  );
nand ( new_n1044_, new_n1043_, new_n1042_ );
or   ( new_n1045_, new_n1012_, new_n1007_ );
and  ( new_n1046_, new_n1045_, new_n1044_ );
or   ( new_n1047_, new_n1024_, new_n1018_ );
xor  ( new_n1048_, \c[7] , \b[8]  );
nand ( new_n1049_, new_n1048_, new_n1016_ );
and  ( new_n1050_, new_n1049_, new_n1047_ );
xor  ( new_n1051_, new_n1050_, new_n1046_ );
xor  ( new_n1052_, new_n1051_, new_n1041_ );
not  ( new_n1053_, \b[12]  );
and  ( new_n1054_, new_n994_, new_n1053_ );
or   ( new_n1055_, \c[1] , \b[13]  );
and  ( new_n1056_, \c[1] , \b[13]  );
nor  ( new_n1057_, new_n1056_, new_n993_ );
and  ( new_n1058_, new_n1057_, new_n1055_ );
or   ( new_n1059_, new_n1058_, new_n1054_ );
and  ( new_n1060_, new_n952_, new_n969_ );
or   ( new_n1061_, new_n1060_, new_n804_ );
or   ( new_n1062_, new_n952_, new_n969_ );
and  ( new_n1063_, new_n1062_, \c[13]  );
and  ( new_n1064_, new_n1063_, new_n1061_ );
nand ( new_n1065_, new_n1064_, new_n1059_ );
not  ( new_n1066_, \c[13]  );
xor  ( new_n1067_, \c[12] , new_n1066_ );
or   ( new_n1068_, new_n1067_, new_n964_ );
or   ( new_n1069_, new_n1068_, new_n966_ );
xor  ( new_n1070_, \c[13] , new_n865_ );
or   ( new_n1071_, new_n1070_, new_n965_ );
and  ( new_n1072_, new_n1071_, new_n1069_ );
xnor ( new_n1073_, new_n1072_, new_n1065_ );
not  ( new_n1074_, new_n955_ );
or   ( new_n1075_, new_n959_, new_n1074_ );
xor  ( new_n1076_, \c[11] , new_n832_ );
or   ( new_n1077_, new_n1076_, new_n958_ );
and  ( new_n1078_, new_n1077_, new_n1075_ );
xor  ( new_n1079_, new_n1078_, new_n1073_ );
xor  ( new_n1080_, new_n1079_, new_n1052_ );
or   ( new_n1081_, new_n965_, new_n804_ );
xor  ( new_n1082_, \c[7] , new_n847_ );
or   ( new_n1083_, new_n1082_, new_n1018_ );
or   ( new_n1084_, new_n1020_, new_n1022_ );
and  ( new_n1085_, new_n1084_, new_n1083_ );
nor  ( new_n1086_, new_n1085_, new_n1081_ );
xor  ( new_n1087_, \c[3] , \b[9]  );
and  ( new_n1088_, new_n1087_, new_n981_ );
and  ( new_n1089_, new_n1028_, new_n980_ );
nor  ( new_n1090_, new_n1089_, new_n1088_ );
not  ( new_n1091_, new_n1090_ );
xor  ( new_n1092_, new_n1085_, new_n1081_ );
and  ( new_n1093_, new_n1092_, new_n1091_ );
or   ( new_n1094_, new_n1093_, new_n1086_ );
xor  ( new_n1095_, new_n1064_, new_n1059_ );
and  ( new_n1096_, new_n1095_, new_n1094_ );
nor  ( new_n1097_, new_n1095_, new_n1094_ );
xor  ( new_n1098_, \c[9] , new_n815_ );
or   ( new_n1099_, new_n1098_, new_n1007_ );
or   ( new_n1100_, new_n1011_, new_n1008_ );
and  ( new_n1101_, new_n1100_, new_n1099_ );
not  ( new_n1102_, new_n994_ );
or   ( new_n1103_, new_n1102_, \b[11]  );
not  ( new_n1104_, \c[1]  );
and  ( new_n1105_, new_n1104_, new_n1053_ );
and  ( new_n1106_, \c[1] , \b[12]  );
or   ( new_n1107_, new_n1106_, new_n993_ );
or   ( new_n1108_, new_n1107_, new_n1105_ );
and  ( new_n1109_, new_n1108_, new_n1103_ );
nor  ( new_n1110_, new_n1109_, new_n1101_ );
xor  ( new_n1111_, \c[11] , \b[1]  );
and  ( new_n1112_, new_n1111_, new_n955_ );
and  ( new_n1113_, new_n956_, new_n954_ );
nor  ( new_n1114_, new_n1113_, new_n1112_ );
and  ( new_n1115_, new_n1109_, new_n1101_ );
nor  ( new_n1116_, new_n1115_, new_n1114_ );
nor  ( new_n1117_, new_n1116_, new_n1110_ );
nor  ( new_n1118_, new_n1117_, new_n1097_ );
nor  ( new_n1119_, new_n1118_, new_n1096_ );
xor  ( new_n1120_, new_n1119_, new_n1080_ );
nor  ( new_n1121_, new_n1120_, new_n1035_ );
and  ( new_n1122_, new_n1120_, new_n1035_ );
xor  ( new_n1123_, \c[3] , \b[8]  );
and  ( new_n1124_, new_n1123_, new_n981_ );
and  ( new_n1125_, new_n1087_, new_n980_ );
nor  ( new_n1126_, new_n1125_, new_n1124_ );
not  ( new_n1127_, \c[10]  );
and  ( new_n1128_, new_n1003_, new_n804_ );
or   ( new_n1129_, new_n1128_, new_n1127_ );
and  ( new_n1130_, \c[9] , \b[0]  );
nor  ( new_n1131_, new_n1130_, new_n952_ );
nand ( new_n1132_, new_n1131_, new_n1129_ );
nor  ( new_n1133_, new_n1132_, new_n1126_ );
not  ( new_n1134_, new_n1133_ );
not  ( new_n1135_, new_n946_ );
xor  ( new_n1136_, \c[5] , new_n1023_ );
or   ( new_n1137_, new_n1136_, new_n1135_ );
nand ( new_n1138_, new_n947_, new_n945_ );
and  ( new_n1139_, new_n1138_, new_n1137_ );
nor  ( new_n1140_, new_n1139_, new_n1134_ );
xor  ( new_n1141_, new_n1139_, new_n1134_ );
not  ( new_n1142_, new_n1141_ );
xor  ( new_n1143_, \c[7] , \b[4]  );
nand ( new_n1144_, new_n1143_, new_n1017_ );
or   ( new_n1145_, new_n1082_, new_n1022_ );
and  ( new_n1146_, new_n1145_, new_n1144_ );
xor  ( new_n1147_, \c[9] , new_n865_ );
or   ( new_n1148_, new_n1147_, new_n1007_ );
or   ( new_n1149_, new_n1098_, new_n1011_ );
and  ( new_n1150_, new_n1149_, new_n1148_ );
or   ( new_n1151_, new_n1150_, new_n1146_ );
and  ( new_n1152_, new_n1150_, new_n1146_ );
and  ( new_n1153_, new_n994_, new_n1038_ );
not  ( new_n1154_, \b[11]  );
and  ( new_n1155_, new_n1104_, new_n1154_ );
not  ( new_n1156_, new_n1155_ );
and  ( new_n1157_, \c[1] , \b[11]  );
nor  ( new_n1158_, new_n1157_, new_n993_ );
and  ( new_n1159_, new_n1158_, new_n1156_ );
nor  ( new_n1160_, new_n1159_, new_n1153_ );
or   ( new_n1161_, new_n1160_, new_n1152_ );
and  ( new_n1162_, new_n1161_, new_n1151_ );
nor  ( new_n1163_, new_n1162_, new_n1142_ );
or   ( new_n1164_, new_n1163_, new_n1140_ );
xor  ( new_n1165_, new_n975_, new_n963_ );
and  ( new_n1166_, new_n1165_, new_n1164_ );
nor  ( new_n1167_, new_n1165_, new_n1164_ );
xor  ( new_n1168_, new_n1026_, new_n1014_ );
xnor ( new_n1169_, new_n1168_, new_n1031_ );
not  ( new_n1170_, new_n1169_ );
nor  ( new_n1171_, new_n1170_, new_n1167_ );
nor  ( new_n1172_, new_n1171_, new_n1166_ );
nor  ( new_n1173_, new_n1172_, new_n1122_ );
nor  ( new_n1174_, new_n1173_, new_n1121_ );
nor  ( new_n1175_, new_n996_, new_n989_ );
and  ( new_n1176_, new_n997_, new_n986_ );
or   ( new_n1177_, new_n1176_, new_n1175_ );
or   ( new_n1178_, new_n1070_, new_n1068_ );
xor  ( new_n1179_, \c[13] , new_n815_ );
or   ( new_n1180_, new_n1179_, new_n965_ );
and  ( new_n1181_, new_n1180_, new_n1178_ );
xor  ( new_n1182_, new_n1181_, new_n1177_ );
xnor ( new_n1183_, new_n1182_, new_n1174_ );
xor  ( new_n1184_, new_n1095_, new_n1094_ );
xor  ( new_n1185_, new_n1184_, new_n1117_ );
xor  ( new_n1186_, new_n1165_, new_n1164_ );
xor  ( new_n1187_, new_n1186_, new_n1170_ );
nor  ( new_n1188_, new_n1187_, new_n1185_ );
and  ( new_n1189_, new_n1187_, new_n1185_ );
xor  ( new_n1190_, new_n1092_, new_n1091_ );
xnor ( new_n1191_, new_n1109_, new_n1101_ );
nand ( new_n1192_, new_n1191_, new_n1114_ );
not  ( new_n1193_, new_n1116_ );
or   ( new_n1194_, new_n1193_, new_n1110_ );
and  ( new_n1195_, new_n1194_, new_n1192_ );
and  ( new_n1196_, new_n1195_, new_n1190_ );
xnor ( new_n1197_, new_n1195_, new_n1190_ );
xor  ( new_n1198_, \c[5] , \b[6]  );
nand ( new_n1199_, new_n1198_, new_n946_ );
or   ( new_n1200_, new_n1136_, new_n1037_ );
and  ( new_n1201_, new_n1200_, new_n1199_ );
nand ( new_n1202_, new_n1111_, new_n954_ );
and  ( new_n1203_, new_n1127_, \c[11]  );
and  ( new_n1204_, \c[10] , \b[0]  );
nor  ( new_n1205_, new_n1204_, new_n1203_ );
and  ( new_n1206_, \c[11] , \b[0]  );
or   ( new_n1207_, new_n1206_, new_n954_ );
or   ( new_n1208_, new_n1207_, new_n1205_ );
and  ( new_n1209_, new_n1208_, new_n1202_ );
or   ( new_n1210_, new_n1209_, new_n1201_ );
and  ( new_n1211_, new_n1209_, new_n1201_ );
xnor ( new_n1212_, new_n1132_, new_n1126_ );
or   ( new_n1213_, new_n1212_, new_n1211_ );
and  ( new_n1214_, new_n1213_, new_n1210_ );
nor  ( new_n1215_, new_n1214_, new_n1197_ );
nor  ( new_n1216_, new_n1215_, new_n1196_ );
nor  ( new_n1217_, new_n1216_, new_n1189_ );
nor  ( new_n1218_, new_n1217_, new_n1188_ );
xor  ( new_n1219_, new_n1120_, new_n1035_ );
xor  ( new_n1220_, new_n1219_, new_n1172_ );
nor  ( new_n1221_, new_n1220_, new_n1218_ );
and  ( new_n1222_, new_n1220_, new_n1218_ );
xor  ( new_n1223_, new_n1162_, new_n1142_ );
not  ( new_n1224_, new_n1223_ );
xor  ( new_n1225_, \c[5] , \b[5]  );
and  ( new_n1226_, new_n1225_, new_n946_ );
and  ( new_n1227_, new_n1198_, new_n945_ );
or   ( new_n1228_, new_n1227_, new_n1226_ );
or   ( new_n1229_, new_n1147_, new_n1011_ );
xor  ( new_n1230_, \c[9] , \b[1]  );
nand ( new_n1231_, new_n1230_, new_n1006_ );
and  ( new_n1232_, new_n1231_, new_n1229_ );
or   ( new_n1233_, new_n1102_, \b[9]  );
and  ( new_n1234_, new_n1104_, new_n1038_ );
and  ( new_n1235_, \c[1] , \b[10]  );
or   ( new_n1236_, new_n1235_, new_n993_ );
or   ( new_n1237_, new_n1236_, new_n1234_ );
and  ( new_n1238_, new_n1237_, new_n1233_ );
nand ( new_n1239_, new_n1238_, new_n1232_ );
and  ( new_n1240_, new_n1239_, new_n1228_ );
nor  ( new_n1241_, new_n1238_, new_n1232_ );
or   ( new_n1242_, new_n1241_, new_n1240_ );
xnor ( new_n1243_, new_n1150_, new_n1146_ );
xor  ( new_n1244_, new_n1243_, new_n1160_ );
nand ( new_n1245_, new_n1244_, new_n1242_ );
nor  ( new_n1246_, new_n1244_, new_n1242_ );
and  ( new_n1247_, new_n1123_, new_n980_ );
xor  ( new_n1248_, \c[3] , \b[7]  );
and  ( new_n1249_, new_n1248_, new_n981_ );
or   ( new_n1250_, new_n1249_, new_n1247_ );
and  ( new_n1251_, new_n954_, \b[0]  );
and  ( new_n1252_, new_n1251_, new_n1250_ );
nor  ( new_n1253_, new_n1251_, new_n1250_ );
xor  ( new_n1254_, \c[7] , \b[3]  );
and  ( new_n1255_, new_n1254_, new_n1017_ );
and  ( new_n1256_, new_n1143_, new_n1016_ );
nor  ( new_n1257_, new_n1256_, new_n1255_ );
nor  ( new_n1258_, new_n1257_, new_n1253_ );
nor  ( new_n1259_, new_n1258_, new_n1252_ );
or   ( new_n1260_, new_n1259_, new_n1246_ );
and  ( new_n1261_, new_n1260_, new_n1245_ );
nor  ( new_n1262_, new_n1261_, new_n1224_ );
xor  ( new_n1263_, new_n1261_, new_n1224_ );
xor  ( new_n1264_, new_n1214_, new_n1197_ );
and  ( new_n1265_, new_n1264_, new_n1263_ );
nor  ( new_n1266_, new_n1265_, new_n1262_ );
not  ( new_n1267_, new_n1266_ );
xnor ( new_n1268_, new_n1187_, new_n1185_ );
xor  ( new_n1269_, new_n1268_, new_n1216_ );
nor  ( new_n1270_, new_n1269_, new_n1267_ );
and  ( new_n1271_, new_n1269_, new_n1267_ );
xor  ( new_n1272_, new_n1264_, new_n1263_ );
not  ( new_n1273_, new_n1272_ );
xor  ( new_n1274_, new_n1209_, new_n1201_ );
xor  ( new_n1275_, new_n1274_, new_n1212_ );
xor  ( new_n1276_, \c[3] , \b[6]  );
and  ( new_n1277_, new_n1276_, new_n981_ );
and  ( new_n1278_, new_n1248_, new_n980_ );
or   ( new_n1279_, new_n1278_, new_n1277_ );
and  ( new_n1280_, new_n1000_, new_n804_ );
or   ( new_n1281_, new_n1280_, new_n1010_ );
and  ( new_n1282_, \c[7] , \b[0]  );
not  ( new_n1283_, new_n1282_ );
and  ( new_n1284_, new_n1283_, \c[9]  );
and  ( new_n1285_, new_n1284_, new_n1281_ );
and  ( new_n1286_, new_n1285_, new_n1279_ );
xnor ( new_n1287_, new_n1251_, new_n1250_ );
xor  ( new_n1288_, new_n1287_, new_n1257_ );
nand ( new_n1289_, new_n1288_, new_n1286_ );
nor  ( new_n1290_, new_n1288_, new_n1286_ );
xor  ( new_n1291_, \c[7] , \b[2]  );
and  ( new_n1292_, new_n1291_, new_n1017_ );
and  ( new_n1293_, new_n1254_, new_n1016_ );
nor  ( new_n1294_, new_n1293_, new_n1292_ );
or   ( new_n1295_, new_n1102_, \b[8]  );
not  ( new_n1296_, \b[9]  );
and  ( new_n1297_, new_n1104_, new_n1296_ );
and  ( new_n1298_, \c[1] , \b[9]  );
or   ( new_n1299_, new_n1298_, new_n993_ );
or   ( new_n1300_, new_n1299_, new_n1297_ );
and  ( new_n1301_, new_n1300_, new_n1295_ );
nor  ( new_n1302_, new_n1301_, new_n1294_ );
and  ( new_n1303_, new_n1301_, new_n1294_ );
and  ( new_n1304_, new_n1230_, new_n1042_ );
xor  ( new_n1305_, \c[9] , \b[0]  );
and  ( new_n1306_, new_n1305_, new_n1006_ );
nor  ( new_n1307_, new_n1306_, new_n1304_ );
nor  ( new_n1308_, new_n1307_, new_n1303_ );
nor  ( new_n1309_, new_n1308_, new_n1302_ );
or   ( new_n1310_, new_n1309_, new_n1290_ );
and  ( new_n1311_, new_n1310_, new_n1289_ );
or   ( new_n1312_, new_n1311_, new_n1275_ );
nand ( new_n1313_, new_n1311_, new_n1275_ );
xor  ( new_n1314_, new_n1244_, new_n1242_ );
xnor ( new_n1315_, new_n1314_, new_n1259_ );
nand ( new_n1316_, new_n1315_, new_n1313_ );
and  ( new_n1317_, new_n1316_, new_n1312_ );
nor  ( new_n1318_, new_n1317_, new_n1273_ );
and  ( new_n1319_, new_n1317_, new_n1273_ );
xor  ( new_n1320_, \c[5] , \b[4]  );
and  ( new_n1321_, new_n1320_, new_n946_ );
and  ( new_n1322_, new_n1225_, new_n945_ );
or   ( new_n1323_, new_n1322_, new_n1321_ );
xor  ( new_n1324_, new_n1285_, new_n1279_ );
nor  ( new_n1325_, new_n1324_, new_n1323_ );
or   ( new_n1326_, new_n1011_, new_n804_ );
or   ( new_n1327_, new_n1102_, \b[7]  );
not  ( new_n1328_, \b[8]  );
and  ( new_n1329_, new_n1104_, new_n1328_ );
and  ( new_n1330_, \c[1] , \b[8]  );
or   ( new_n1331_, new_n1330_, new_n993_ );
or   ( new_n1332_, new_n1331_, new_n1329_ );
and  ( new_n1333_, new_n1332_, new_n1327_ );
and  ( new_n1334_, new_n1333_, new_n1326_ );
xor  ( new_n1335_, \c[7] , \b[1]  );
nand ( new_n1336_, new_n1335_, new_n1017_ );
nand ( new_n1337_, new_n1291_, new_n1016_ );
and  ( new_n1338_, new_n1337_, new_n1336_ );
xor  ( new_n1339_, new_n1333_, new_n1326_ );
and  ( new_n1340_, new_n1339_, new_n1338_ );
nor  ( new_n1341_, new_n1340_, new_n1334_ );
not  ( new_n1342_, new_n1341_ );
xor  ( new_n1343_, new_n1324_, new_n1323_ );
and  ( new_n1344_, new_n1343_, new_n1342_ );
nor  ( new_n1345_, new_n1344_, new_n1325_ );
xor  ( new_n1346_, new_n1238_, new_n1232_ );
xor  ( new_n1347_, new_n1346_, new_n1228_ );
nor  ( new_n1348_, new_n1347_, new_n1345_ );
xor  ( new_n1349_, new_n1347_, new_n1345_ );
not  ( new_n1350_, new_n1349_ );
xnor ( new_n1351_, new_n1288_, new_n1286_ );
xor  ( new_n1352_, new_n1351_, new_n1309_ );
nor  ( new_n1353_, new_n1352_, new_n1350_ );
nor  ( new_n1354_, new_n1353_, new_n1348_ );
xor  ( new_n1355_, new_n1311_, new_n1275_ );
xor  ( new_n1356_, new_n1355_, new_n1315_ );
and  ( new_n1357_, new_n1356_, new_n1354_ );
nor  ( new_n1358_, new_n1356_, new_n1354_ );
xor  ( new_n1359_, new_n1352_, new_n1350_ );
xnor ( new_n1360_, new_n1301_, new_n1294_ );
and  ( new_n1361_, new_n1360_, new_n1307_ );
not  ( new_n1362_, new_n1302_ );
and  ( new_n1363_, new_n1308_, new_n1362_ );
or   ( new_n1364_, new_n1363_, new_n1361_ );
and  ( new_n1365_, new_n994_, new_n1019_ );
and  ( new_n1366_, new_n1104_, new_n1023_ );
not  ( new_n1367_, new_n1366_ );
and  ( new_n1368_, \c[1] , \b[7]  );
nor  ( new_n1369_, new_n1368_, new_n993_ );
and  ( new_n1370_, new_n1369_, new_n1367_ );
nor  ( new_n1371_, new_n1370_, new_n1365_ );
not  ( new_n1372_, new_n1371_ );
not  ( new_n1373_, \c[6]  );
and  ( new_n1374_, new_n943_, new_n1373_ );
or   ( new_n1375_, new_n1374_, new_n804_ );
or   ( new_n1376_, new_n943_, new_n1373_ );
and  ( new_n1377_, new_n1376_, \c[7]  );
and  ( new_n1378_, new_n1377_, new_n1375_ );
nand ( new_n1379_, new_n1378_, new_n1372_ );
xor  ( new_n1380_, \c[5] , new_n815_ );
or   ( new_n1381_, new_n1380_, new_n1135_ );
nand ( new_n1382_, new_n1320_, new_n945_ );
and  ( new_n1383_, new_n1382_, new_n1381_ );
or   ( new_n1384_, new_n1383_, new_n1379_ );
and  ( new_n1385_, new_n1383_, new_n1379_ );
xor  ( new_n1386_, \c[3] , \b[5]  );
and  ( new_n1387_, new_n1386_, new_n981_ );
and  ( new_n1388_, new_n1276_, new_n980_ );
nor  ( new_n1389_, new_n1388_, new_n1387_ );
or   ( new_n1390_, new_n1389_, new_n1385_ );
and  ( new_n1391_, new_n1390_, new_n1384_ );
or   ( new_n1392_, new_n1391_, new_n1364_ );
and  ( new_n1393_, new_n1391_, new_n1364_ );
xor  ( new_n1394_, new_n1343_, new_n1342_ );
or   ( new_n1395_, new_n1394_, new_n1393_ );
and  ( new_n1396_, new_n1395_, new_n1392_ );
nor  ( new_n1397_, new_n1396_, new_n1359_ );
and  ( new_n1398_, new_n1396_, new_n1359_ );
xor  ( new_n1399_, new_n1391_, new_n1364_ );
xor  ( new_n1400_, new_n1399_, new_n1394_ );
not  ( new_n1401_, new_n1400_ );
xor  ( new_n1402_, new_n1339_, new_n1338_ );
xor  ( new_n1403_, \c[3] , \b[4]  );
nand ( new_n1404_, new_n1403_, new_n981_ );
nand ( new_n1405_, new_n1386_, new_n980_ );
and  ( new_n1406_, new_n1405_, new_n1404_ );
xor  ( new_n1407_, \c[5] , new_n865_ );
or   ( new_n1408_, new_n1407_, new_n1135_ );
or   ( new_n1409_, new_n1380_, new_n1037_ );
and  ( new_n1410_, new_n1409_, new_n1408_ );
nor  ( new_n1411_, new_n1410_, new_n1406_ );
and  ( new_n1412_, new_n1410_, new_n1406_ );
and  ( new_n1413_, new_n1335_, new_n1016_ );
and  ( new_n1414_, new_n1373_, \c[7]  );
and  ( new_n1415_, \c[6] , \b[0]  );
nor  ( new_n1416_, new_n1415_, new_n1414_ );
not  ( new_n1417_, new_n1416_ );
and  ( new_n1418_, new_n1283_, new_n1022_ );
and  ( new_n1419_, new_n1418_, new_n1417_ );
nor  ( new_n1420_, new_n1419_, new_n1413_ );
nor  ( new_n1421_, new_n1420_, new_n1412_ );
nor  ( new_n1422_, new_n1421_, new_n1411_ );
nand ( new_n1423_, new_n1422_, new_n1402_ );
nor  ( new_n1424_, new_n1422_, new_n1402_ );
xor  ( new_n1425_, new_n1383_, new_n1379_ );
xnor ( new_n1426_, new_n1425_, new_n1389_ );
or   ( new_n1427_, new_n1426_, new_n1424_ );
and  ( new_n1428_, new_n1427_, new_n1423_ );
and  ( new_n1429_, new_n1428_, new_n1401_ );
nor  ( new_n1430_, new_n1428_, new_n1401_ );
xor  ( new_n1431_, new_n1378_, new_n1372_ );
or   ( new_n1432_, new_n1022_, new_n804_ );
or   ( new_n1433_, new_n1102_, \b[5]  );
and  ( new_n1434_, new_n1104_, new_n1019_ );
and  ( new_n1435_, \c[1] , \b[6]  );
or   ( new_n1436_, new_n1435_, new_n993_ );
or   ( new_n1437_, new_n1436_, new_n1434_ );
and  ( new_n1438_, new_n1437_, new_n1433_ );
or   ( new_n1439_, new_n1438_, new_n1432_ );
and  ( new_n1440_, new_n1438_, new_n1432_ );
xor  ( new_n1441_, \c[3] , \b[3]  );
and  ( new_n1442_, new_n1441_, new_n981_ );
and  ( new_n1443_, new_n1403_, new_n980_ );
nor  ( new_n1444_, new_n1443_, new_n1442_ );
or   ( new_n1445_, new_n1444_, new_n1440_ );
nand ( new_n1446_, new_n1445_, new_n1439_ );
nor  ( new_n1447_, new_n1446_, new_n1431_ );
xnor ( new_n1448_, new_n1446_, new_n1431_ );
xnor ( new_n1449_, new_n1410_, new_n1406_ );
nand ( new_n1450_, new_n1449_, new_n1420_ );
not  ( new_n1451_, new_n1421_ );
or   ( new_n1452_, new_n1451_, new_n1411_ );
and  ( new_n1453_, new_n1452_, new_n1450_ );
nor  ( new_n1454_, new_n1453_, new_n1448_ );
nor  ( new_n1455_, new_n1454_, new_n1447_ );
not  ( new_n1456_, new_n1455_ );
xnor ( new_n1457_, new_n1422_, new_n1402_ );
xor  ( new_n1458_, new_n1457_, new_n1426_ );
nor  ( new_n1459_, new_n1458_, new_n1456_ );
and  ( new_n1460_, new_n1458_, new_n1456_ );
xor  ( new_n1461_, new_n1453_, new_n1448_ );
and  ( new_n1462_, new_n994_, new_n832_ );
or   ( new_n1463_, \c[1] , \b[5]  );
and  ( new_n1464_, \c[1] , \b[5]  );
nor  ( new_n1465_, new_n1464_, new_n993_ );
and  ( new_n1466_, new_n1465_, new_n1463_ );
or   ( new_n1467_, new_n1466_, new_n1462_ );
not  ( new_n1468_, \c[4]  );
and  ( new_n1469_, new_n978_, new_n1468_ );
or   ( new_n1470_, new_n1469_, new_n804_ );
or   ( new_n1471_, new_n978_, new_n1468_ );
and  ( new_n1472_, new_n1471_, \c[5]  );
and  ( new_n1473_, new_n1472_, new_n1470_ );
nand ( new_n1474_, new_n1473_, new_n1467_ );
xor  ( new_n1475_, \c[5] , new_n808_ );
or   ( new_n1476_, new_n1475_, new_n1135_ );
or   ( new_n1477_, new_n1407_, new_n1037_ );
and  ( new_n1478_, new_n1477_, new_n1476_ );
or   ( new_n1479_, new_n1478_, new_n1474_ );
nand ( new_n1480_, new_n1478_, new_n1474_ );
xor  ( new_n1481_, new_n1438_, new_n1432_ );
xnor ( new_n1482_, new_n1481_, new_n1444_ );
nand ( new_n1483_, new_n1482_, new_n1480_ );
and  ( new_n1484_, new_n1483_, new_n1479_ );
nor  ( new_n1485_, new_n1484_, new_n1461_ );
and  ( new_n1486_, new_n1484_, new_n1461_ );
xor  ( new_n1487_, \c[3] , \b[2]  );
and  ( new_n1488_, new_n1487_, new_n981_ );
and  ( new_n1489_, new_n1441_, new_n980_ );
nor  ( new_n1490_, new_n1489_, new_n1488_ );
or   ( new_n1491_, new_n1475_, new_n1037_ );
and  ( new_n1492_, new_n1468_, \c[5]  );
and  ( new_n1493_, \c[4] , \b[0]  );
nor  ( new_n1494_, new_n1493_, new_n1492_ );
and  ( new_n1495_, \c[5] , \b[0]  );
or   ( new_n1496_, new_n1495_, new_n945_ );
or   ( new_n1497_, new_n1496_, new_n1494_ );
and  ( new_n1498_, new_n1497_, new_n1491_ );
nor  ( new_n1499_, new_n1498_, new_n1490_ );
xor  ( new_n1500_, new_n1498_, new_n1490_ );
xor  ( new_n1501_, new_n1473_, new_n1467_ );
and  ( new_n1502_, new_n1501_, new_n1500_ );
nor  ( new_n1503_, new_n1502_, new_n1499_ );
not  ( new_n1504_, new_n1503_ );
xor  ( new_n1505_, new_n1478_, new_n1474_ );
xor  ( new_n1506_, new_n1505_, new_n1482_ );
and  ( new_n1507_, new_n1506_, new_n1504_ );
xor  ( new_n1508_, new_n1506_, new_n1504_ );
xnor ( new_n1509_, new_n1501_, new_n1500_ );
or   ( new_n1510_, new_n1037_, new_n804_ );
or   ( new_n1511_, new_n1102_, \b[3]  );
and  ( new_n1512_, new_n1104_, new_n832_ );
and  ( new_n1513_, \c[1] , \b[4]  );
or   ( new_n1514_, new_n1513_, new_n993_ );
or   ( new_n1515_, new_n1514_, new_n1512_ );
and  ( new_n1516_, new_n1515_, new_n1511_ );
or   ( new_n1517_, new_n1516_, new_n1510_ );
and  ( new_n1518_, new_n1516_, new_n1510_ );
xor  ( new_n1519_, \c[3] , \b[1]  );
and  ( new_n1520_, new_n1519_, new_n981_ );
and  ( new_n1521_, new_n1487_, new_n980_ );
nor  ( new_n1522_, new_n1521_, new_n1520_ );
or   ( new_n1523_, new_n1522_, new_n1518_ );
and  ( new_n1524_, new_n1523_, new_n1517_ );
or   ( new_n1525_, new_n1524_, new_n1509_ );
and  ( new_n1526_, new_n1524_, new_n1509_ );
and  ( new_n1527_, new_n994_, new_n865_ );
and  ( new_n1528_, new_n1104_, new_n815_ );
not  ( new_n1529_, new_n1528_ );
and  ( new_n1530_, \c[1] , \b[3]  );
nor  ( new_n1531_, new_n1530_, new_n993_ );
and  ( new_n1532_, new_n1531_, new_n1529_ );
nor  ( new_n1533_, new_n1532_, new_n1527_ );
not  ( new_n1534_, \c[2]  );
and  ( new_n1535_, new_n1104_, new_n1534_ );
or   ( new_n1536_, new_n1535_, new_n804_ );
or   ( new_n1537_, new_n1104_, new_n1534_ );
and  ( new_n1538_, new_n1537_, \c[3]  );
nand ( new_n1539_, new_n1538_, new_n1536_ );
nor  ( new_n1540_, new_n1539_, new_n1533_ );
xnor ( new_n1541_, new_n1516_, new_n1510_ );
xor  ( new_n1542_, new_n1541_, new_n1522_ );
and  ( new_n1543_, new_n1542_, new_n1540_ );
nor  ( new_n1544_, new_n1542_, new_n1540_ );
xnor ( new_n1545_, new_n1539_, new_n1533_ );
nand ( new_n1546_, new_n1519_, new_n980_ );
and  ( new_n1547_, new_n1534_, \c[3]  );
and  ( new_n1548_, \c[2] , \b[0]  );
nor  ( new_n1549_, new_n1548_, new_n1547_ );
and  ( new_n1550_, \c[3] , \b[0]  );
or   ( new_n1551_, new_n1550_, new_n980_ );
or   ( new_n1552_, new_n1551_, new_n1549_ );
and  ( new_n1553_, new_n1552_, new_n1546_ );
nor  ( new_n1554_, new_n1553_, new_n1545_ );
and  ( new_n1555_, new_n1553_, new_n1545_ );
not  ( new_n1556_, new_n980_ );
or   ( new_n1557_, new_n1556_, new_n804_ );
or   ( new_n1558_, new_n1102_, \b[1]  );
and  ( new_n1559_, new_n1104_, new_n865_ );
and  ( new_n1560_, \c[1] , \b[2]  );
or   ( new_n1561_, new_n1560_, new_n993_ );
or   ( new_n1562_, new_n1561_, new_n1559_ );
and  ( new_n1563_, new_n1562_, new_n1558_ );
nor  ( new_n1564_, new_n1563_, new_n1557_ );
and  ( new_n1565_, new_n1563_, new_n1557_ );
and  ( new_n1566_, \c[0] , \b[1]  );
not  ( new_n1567_, new_n1566_ );
and  ( new_n1568_, \c[1] , new_n804_ );
and  ( new_n1569_, new_n1568_, new_n1567_ );
not  ( new_n1570_, new_n1569_ );
nor  ( new_n1571_, new_n1570_, new_n1565_ );
nor  ( new_n1572_, new_n1571_, new_n1564_ );
nor  ( new_n1573_, new_n1572_, new_n1555_ );
nor  ( new_n1574_, new_n1573_, new_n1554_ );
nor  ( new_n1575_, new_n1574_, new_n1544_ );
nor  ( new_n1576_, new_n1575_, new_n1543_ );
or   ( new_n1577_, new_n1576_, new_n1526_ );
nand ( new_n1578_, new_n1577_, new_n1525_ );
and  ( new_n1579_, new_n1578_, new_n1508_ );
nor  ( new_n1580_, new_n1579_, new_n1507_ );
nor  ( new_n1581_, new_n1580_, new_n1486_ );
nor  ( new_n1582_, new_n1581_, new_n1485_ );
nor  ( new_n1583_, new_n1582_, new_n1460_ );
nor  ( new_n1584_, new_n1583_, new_n1459_ );
nor  ( new_n1585_, new_n1584_, new_n1430_ );
nor  ( new_n1586_, new_n1585_, new_n1429_ );
nor  ( new_n1587_, new_n1586_, new_n1398_ );
nor  ( new_n1588_, new_n1587_, new_n1397_ );
nor  ( new_n1589_, new_n1588_, new_n1358_ );
nor  ( new_n1590_, new_n1589_, new_n1357_ );
nor  ( new_n1591_, new_n1590_, new_n1319_ );
nor  ( new_n1592_, new_n1591_, new_n1318_ );
not  ( new_n1593_, new_n1592_ );
nor  ( new_n1594_, new_n1593_, new_n1271_ );
nor  ( new_n1595_, new_n1594_, new_n1270_ );
not  ( new_n1596_, new_n1595_ );
nor  ( new_n1597_, new_n1596_, new_n1222_ );
nor  ( new_n1598_, new_n1597_, new_n1221_ );
and  ( new_n1599_, new_n1048_, new_n1017_ );
xor  ( new_n1600_, \c[7] , \b[9]  );
and  ( new_n1601_, new_n1600_, new_n1016_ );
or   ( new_n1602_, new_n1601_, new_n1599_ );
nand ( new_n1603_, new_n998_, new_n977_ );
or   ( new_n1604_, new_n1034_, new_n999_ );
and  ( new_n1605_, new_n1604_, new_n1603_ );
and  ( new_n1606_, new_n1043_, new_n1006_ );
xor  ( new_n1607_, \c[9] , \b[7]  );
and  ( new_n1608_, new_n1607_, new_n1042_ );
or   ( new_n1609_, new_n1608_, new_n1606_ );
nand ( new_n1610_, new_n984_, new_n981_ );
xor  ( new_n1611_, \c[3] , new_n992_ );
or   ( new_n1612_, new_n1611_, new_n1556_ );
and  ( new_n1613_, new_n1612_, new_n1610_ );
xor  ( new_n1614_, new_n1613_, new_n1609_ );
xor  ( new_n1615_, new_n1614_, new_n1605_ );
or   ( new_n1616_, new_n1050_, new_n1046_ );
nand ( new_n1617_, new_n1051_, new_n1041_ );
and  ( new_n1618_, new_n1617_, new_n1616_ );
or   ( new_n1619_, new_n990_, \c[0]  );
and  ( new_n1620_, \c[0] , \b[15]  );
xor  ( new_n1621_, new_n1620_, \c[1]  );
and  ( new_n1622_, new_n1621_, new_n1619_ );
xor  ( new_n1623_, new_n1622_, new_n1618_ );
not  ( new_n1624_, \c[14]  );
and  ( new_n1625_, new_n1624_, new_n804_ );
or   ( new_n1626_, new_n1625_, new_n1066_ );
and  ( new_n1627_, \c[14] , \b[0]  );
not  ( new_n1628_, new_n1627_ );
and  ( new_n1629_, new_n1628_, \c[15]  );
and  ( new_n1630_, new_n1629_, new_n1626_ );
xor  ( new_n1631_, new_n1630_, new_n1623_ );
xor  ( new_n1632_, new_n1631_, new_n1615_ );
or   ( new_n1633_, new_n1039_, new_n1135_ );
xor  ( new_n1634_, \c[5] , new_n1154_ );
or   ( new_n1635_, new_n1634_, new_n1037_ );
and  ( new_n1636_, new_n1635_, new_n1633_ );
or   ( new_n1637_, new_n1076_, new_n1074_ );
xor  ( new_n1638_, \c[11] , new_n847_ );
or   ( new_n1639_, new_n1638_, new_n958_ );
and  ( new_n1640_, new_n1639_, new_n1637_ );
xor  ( new_n1641_, new_n1640_, new_n1636_ );
or   ( new_n1642_, new_n1072_, new_n1065_ );
and  ( new_n1643_, new_n1072_, new_n1065_ );
or   ( new_n1644_, new_n1078_, new_n1643_ );
and  ( new_n1645_, new_n1644_, new_n1642_ );
xor  ( new_n1646_, new_n1645_, new_n1641_ );
xor  ( new_n1647_, new_n1646_, new_n1632_ );
xor  ( new_n1648_, new_n1647_, new_n1602_ );
and  ( new_n1649_, new_n1079_, new_n1052_ );
nor  ( new_n1650_, new_n1079_, new_n1052_ );
nor  ( new_n1651_, new_n1119_, new_n1650_ );
or   ( new_n1652_, new_n1651_, new_n1649_ );
not  ( new_n1653_, \c[15]  );
nor  ( new_n1654_, new_n1625_, new_n1653_ );
and  ( new_n1655_, new_n1628_, new_n1653_ );
or   ( new_n1656_, new_n1655_, new_n987_ );
or   ( new_n1657_, new_n1656_, new_n1654_ );
xor  ( new_n1658_, \c[15] , \b[1]  );
nand ( new_n1659_, new_n1658_, new_n987_ );
and  ( new_n1660_, new_n1659_, new_n1657_ );
xor  ( new_n1661_, new_n1660_, new_n1652_ );
xor  ( new_n1662_, new_n1661_, new_n1648_ );
xnor ( new_n1663_, new_n1662_, new_n1598_ );
nor  ( new_n1664_, new_n1663_, new_n1183_ );
not  ( new_n1665_, new_n1664_ );
and  ( new_n1666_, new_n922_, new_n849_ );
xor  ( new_n1667_, \b[5] , \a[3]  );
and  ( new_n1668_, new_n1667_, new_n801_ );
nor  ( new_n1669_, new_n1668_, new_n1666_ );
not  ( new_n1670_, new_n1669_ );
xor  ( new_n1671_, \b[7] , new_n98_ );
xor  ( new_n1672_, \b[6] , new_n1023_ );
nor  ( new_n1673_, new_n1672_, new_n918_ );
not  ( new_n1674_, new_n1673_ );
or   ( new_n1675_, new_n1674_, new_n1671_ );
xor  ( new_n1676_, \b[7] , new_n108_ );
or   ( new_n1677_, new_n1676_, new_n919_ );
and  ( new_n1678_, new_n1677_, new_n1675_ );
or   ( new_n1679_, new_n806_, \a[6]  );
and  ( new_n1680_, new_n808_, new_n185_ );
and  ( new_n1681_, \b[1] , \a[7]  );
or   ( new_n1682_, new_n1681_, new_n804_ );
or   ( new_n1683_, new_n1682_, new_n1680_ );
and  ( new_n1684_, new_n1683_, new_n1679_ );
xor  ( new_n1685_, new_n1684_, new_n1678_ );
xor  ( new_n1686_, new_n1685_, new_n1670_ );
nor  ( new_n1687_, new_n924_, new_n920_ );
and  ( new_n1688_, new_n925_, new_n917_ );
or   ( new_n1689_, new_n1688_, new_n1687_ );
and  ( new_n1690_, new_n914_, new_n818_ );
xor  ( new_n1691_, \b[3] , \a[5]  );
and  ( new_n1692_, new_n1691_, new_n817_ );
or   ( new_n1693_, new_n1692_, new_n1690_ );
and  ( new_n1694_, new_n847_, new_n98_ );
or   ( new_n1695_, new_n1694_, new_n1019_ );
and  ( new_n1696_, \b[5] , \a[0]  );
nor  ( new_n1697_, new_n1696_, new_n1023_ );
and  ( new_n1698_, new_n1697_, new_n1695_ );
xor  ( new_n1699_, new_n1698_, new_n1693_ );
xor  ( new_n1700_, new_n1699_, new_n1689_ );
xor  ( new_n1701_, new_n1700_, new_n1686_ );
not  ( new_n1702_, new_n1701_ );
or   ( new_n1703_, new_n933_, new_n927_ );
nand ( new_n1704_, new_n933_, new_n927_ );
nand ( new_n1705_, new_n1704_, new_n926_ );
and  ( new_n1706_, new_n1705_, new_n1703_ );
xor  ( new_n1707_, new_n1706_, new_n1702_ );
not  ( new_n1708_, new_n1707_ );
nand ( new_n1709_, new_n935_, new_n912_ );
nor  ( new_n1710_, new_n935_, new_n912_ );
or   ( new_n1711_, new_n1710_, new_n908_ );
and  ( new_n1712_, new_n1711_, new_n1709_ );
xor  ( new_n1713_, new_n1712_, new_n1708_ );
not  ( new_n1714_, new_n1713_ );
and  ( new_n1715_, new_n1663_, new_n1183_ );
nor  ( new_n1716_, new_n1715_, new_n1714_ );
and  ( new_n1717_, new_n1716_, new_n1665_ );
not  ( new_n1718_, new_n1717_ );
not  ( new_n1719_, \a[15]  );
xor  ( new_n1720_, \c[15] , new_n1719_ );
or   ( new_n1721_, \c[14] , \a[14]  );
and  ( new_n1722_, \c[14] , \a[14]  );
and  ( new_n1723_, new_n1066_, new_n89_ );
and  ( new_n1724_, \c[13] , \a[13]  );
and  ( new_n1725_, new_n969_, new_n85_ );
and  ( new_n1726_, \c[12] , \a[12]  );
and  ( new_n1727_, new_n952_, new_n354_ );
and  ( new_n1728_, \c[11] , \a[11]  );
and  ( new_n1729_, new_n1127_, new_n352_ );
and  ( new_n1730_, \c[10] , \a[10]  );
and  ( new_n1731_, new_n1003_, new_n137_ );
and  ( new_n1732_, \c[9] , \a[9]  );
and  ( new_n1733_, new_n1010_, new_n133_ );
and  ( new_n1734_, \c[8] , \a[8]  );
and  ( new_n1735_, new_n1000_, new_n185_ );
and  ( new_n1736_, \c[7] , \a[7]  );
and  ( new_n1737_, new_n1373_, new_n212_ );
and  ( new_n1738_, \c[6] , \a[6]  );
and  ( new_n1739_, new_n943_, new_n176_ );
and  ( new_n1740_, \c[5] , \a[5]  );
and  ( new_n1741_, new_n1468_, new_n231_ );
and  ( new_n1742_, \c[4] , \a[4]  );
and  ( new_n1743_, new_n978_, new_n163_ );
and  ( new_n1744_, \c[3] , \a[3]  );
and  ( new_n1745_, new_n1534_, new_n115_ );
and  ( new_n1746_, \c[2] , \a[2]  );
and  ( new_n1747_, new_n1104_, new_n108_ );
and  ( new_n1748_, \c[1] , \a[1]  );
and  ( new_n1749_, \c[0] , \a[0]  );
nor  ( new_n1750_, new_n1749_, new_n1748_ );
nor  ( new_n1751_, new_n1750_, new_n1747_ );
nor  ( new_n1752_, new_n1751_, new_n1746_ );
nor  ( new_n1753_, new_n1752_, new_n1745_ );
nor  ( new_n1754_, new_n1753_, new_n1744_ );
nor  ( new_n1755_, new_n1754_, new_n1743_ );
nor  ( new_n1756_, new_n1755_, new_n1742_ );
nor  ( new_n1757_, new_n1756_, new_n1741_ );
nor  ( new_n1758_, new_n1757_, new_n1740_ );
nor  ( new_n1759_, new_n1758_, new_n1739_ );
nor  ( new_n1760_, new_n1759_, new_n1738_ );
nor  ( new_n1761_, new_n1760_, new_n1737_ );
nor  ( new_n1762_, new_n1761_, new_n1736_ );
nor  ( new_n1763_, new_n1762_, new_n1735_ );
nor  ( new_n1764_, new_n1763_, new_n1734_ );
nor  ( new_n1765_, new_n1764_, new_n1733_ );
nor  ( new_n1766_, new_n1765_, new_n1732_ );
nor  ( new_n1767_, new_n1766_, new_n1731_ );
nor  ( new_n1768_, new_n1767_, new_n1730_ );
nor  ( new_n1769_, new_n1768_, new_n1729_ );
nor  ( new_n1770_, new_n1769_, new_n1728_ );
nor  ( new_n1771_, new_n1770_, new_n1727_ );
nor  ( new_n1772_, new_n1771_, new_n1726_ );
nor  ( new_n1773_, new_n1772_, new_n1725_ );
nor  ( new_n1774_, new_n1773_, new_n1724_ );
nor  ( new_n1775_, new_n1774_, new_n1723_ );
or   ( new_n1776_, new_n1775_, new_n1722_ );
and  ( new_n1777_, new_n1776_, new_n1721_ );
xnor ( new_n1778_, new_n1777_, new_n1720_ );
xor  ( new_n1779_, new_n873_, new_n871_ );
xnor ( new_n1780_, new_n1779_, new_n904_ );
and  ( new_n1781_, new_n1780_, new_n1778_ );
not  ( new_n1782_, new_n1781_ );
not  ( new_n1783_, \b[15]  );
xor  ( new_n1784_, \d[15] , new_n1783_ );
or   ( new_n1785_, \d[14] , \b[14]  );
and  ( new_n1786_, \d[14] , \b[14]  );
and  ( new_n1787_, new_n103_, new_n992_ );
and  ( new_n1788_, \d[13] , \b[13]  );
and  ( new_n1789_, new_n99_, new_n1053_ );
and  ( new_n1790_, \d[12] , \b[12]  );
and  ( new_n1791_, new_n75_, new_n1154_ );
and  ( new_n1792_, \d[11] , \b[11]  );
and  ( new_n1793_, new_n326_, new_n1038_ );
and  ( new_n1794_, \d[10] , \b[10]  );
and  ( new_n1795_, new_n171_, new_n1296_ );
and  ( new_n1796_, \d[9] , \b[9]  );
and  ( new_n1797_, new_n179_, new_n1328_ );
and  ( new_n1798_, \d[8] , \b[8]  );
and  ( new_n1799_, new_n128_, new_n1023_ );
and  ( new_n1800_, \d[7] , \b[7]  );
and  ( new_n1801_, new_n563_, new_n1019_ );
and  ( new_n1802_, \d[6] , \b[6]  );
and  ( new_n1803_, new_n66_, new_n847_ );
and  ( new_n1804_, \d[5] , \b[5]  );
and  ( new_n1805_, new_n660_, new_n832_ );
and  ( new_n1806_, \d[4] , \b[4]  );
and  ( new_n1807_, new_n150_, new_n815_ );
and  ( new_n1808_, \d[3] , \b[3]  );
and  ( new_n1809_, new_n726_, new_n865_ );
and  ( new_n1810_, \d[2] , \b[2]  );
and  ( new_n1811_, new_n90_, new_n808_ );
and  ( new_n1812_, \d[1] , \b[1]  );
and  ( new_n1813_, \d[0] , \b[0]  );
nor  ( new_n1814_, new_n1813_, new_n1812_ );
nor  ( new_n1815_, new_n1814_, new_n1811_ );
nor  ( new_n1816_, new_n1815_, new_n1810_ );
nor  ( new_n1817_, new_n1816_, new_n1809_ );
nor  ( new_n1818_, new_n1817_, new_n1808_ );
nor  ( new_n1819_, new_n1818_, new_n1807_ );
nor  ( new_n1820_, new_n1819_, new_n1806_ );
nor  ( new_n1821_, new_n1820_, new_n1805_ );
nor  ( new_n1822_, new_n1821_, new_n1804_ );
nor  ( new_n1823_, new_n1822_, new_n1803_ );
nor  ( new_n1824_, new_n1823_, new_n1802_ );
nor  ( new_n1825_, new_n1824_, new_n1801_ );
nor  ( new_n1826_, new_n1825_, new_n1800_ );
nor  ( new_n1827_, new_n1826_, new_n1799_ );
nor  ( new_n1828_, new_n1827_, new_n1798_ );
nor  ( new_n1829_, new_n1828_, new_n1797_ );
nor  ( new_n1830_, new_n1829_, new_n1796_ );
nor  ( new_n1831_, new_n1830_, new_n1795_ );
nor  ( new_n1832_, new_n1831_, new_n1794_ );
nor  ( new_n1833_, new_n1832_, new_n1793_ );
nor  ( new_n1834_, new_n1833_, new_n1792_ );
nor  ( new_n1835_, new_n1834_, new_n1791_ );
nor  ( new_n1836_, new_n1835_, new_n1790_ );
nor  ( new_n1837_, new_n1836_, new_n1789_ );
nor  ( new_n1838_, new_n1837_, new_n1788_ );
nor  ( new_n1839_, new_n1838_, new_n1787_ );
or   ( new_n1840_, new_n1839_, new_n1786_ );
and  ( new_n1841_, new_n1840_, new_n1785_ );
xnor ( new_n1842_, new_n1841_, new_n1784_ );
xor  ( new_n1843_, new_n855_, new_n826_ );
xnor ( new_n1844_, new_n1843_, new_n906_ );
and  ( new_n1845_, new_n1844_, new_n1842_ );
not  ( new_n1846_, new_n1845_ );
xor  ( new_n1847_, new_n885_, new_n876_ );
xor  ( new_n1848_, new_n1847_, new_n901_ );
not  ( new_n1849_, new_n1848_ );
xor  ( new_n1850_, \b[3] , \a[6]  );
and  ( new_n1851_, new_n1850_, new_n818_ );
xor  ( new_n1852_, \b[3] , \a[7]  );
and  ( new_n1853_, new_n1852_, new_n817_ );
or   ( new_n1854_, new_n1853_, new_n1851_ );
xor  ( new_n1855_, \b[7] , new_n115_ );
or   ( new_n1856_, new_n1855_, new_n1674_ );
xor  ( new_n1857_, \b[7] , \a[3]  );
nand ( new_n1858_, new_n1857_, new_n918_ );
and  ( new_n1859_, new_n1858_, new_n1856_ );
or   ( new_n1860_, new_n806_, \a[8]  );
and  ( new_n1861_, new_n808_, new_n137_ );
and  ( new_n1862_, \b[1] , \a[9]  );
or   ( new_n1863_, new_n1862_, new_n804_ );
or   ( new_n1864_, new_n1863_, new_n1861_ );
and  ( new_n1865_, new_n1864_, new_n1860_ );
xor  ( new_n1866_, new_n1865_, new_n1859_ );
xor  ( new_n1867_, new_n1866_, new_n1854_ );
xor  ( new_n1868_, \b[7] , \b[8]  );
nand ( new_n1869_, new_n1868_, \a[0]  );
or   ( new_n1870_, new_n806_, \a[7]  );
and  ( new_n1871_, new_n808_, new_n133_ );
and  ( new_n1872_, \b[1] , \a[8]  );
or   ( new_n1873_, new_n1872_, new_n804_ );
or   ( new_n1874_, new_n1873_, new_n1871_ );
and  ( new_n1875_, new_n1874_, new_n1870_ );
nor  ( new_n1876_, new_n1875_, new_n1869_ );
and  ( new_n1877_, new_n1691_, new_n818_ );
and  ( new_n1878_, new_n1850_, new_n817_ );
or   ( new_n1879_, new_n1878_, new_n1877_ );
xor  ( new_n1880_, new_n1875_, new_n1869_ );
and  ( new_n1881_, new_n1880_, new_n1879_ );
nor  ( new_n1882_, new_n1881_, new_n1876_ );
xor  ( new_n1883_, \b[9] , \a[1]  );
and  ( new_n1884_, new_n1883_, new_n1868_ );
xor  ( new_n1885_, \b[8] , new_n1296_ );
nor  ( new_n1886_, new_n1885_, new_n1868_ );
and  ( new_n1887_, new_n1886_, new_n1671_ );
or   ( new_n1888_, new_n1887_, new_n1884_ );
xor  ( new_n1889_, \b[5] , \a[4]  );
and  ( new_n1890_, new_n1889_, new_n849_ );
xor  ( new_n1891_, \b[5] , \a[5]  );
and  ( new_n1892_, new_n1891_, new_n801_ );
or   ( new_n1893_, new_n1892_, new_n1890_ );
and  ( new_n1894_, new_n1023_, new_n98_ );
or   ( new_n1895_, new_n1894_, new_n1328_ );
and  ( new_n1896_, \b[7] , \a[0]  );
nor  ( new_n1897_, new_n1896_, new_n1296_ );
and  ( new_n1898_, new_n1897_, new_n1895_ );
xor  ( new_n1899_, new_n1898_, new_n1893_ );
xnor ( new_n1900_, new_n1899_, new_n1888_ );
xor  ( new_n1901_, new_n1900_, new_n1882_ );
and  ( new_n1902_, new_n1901_, new_n1867_ );
or   ( new_n1903_, new_n1676_, new_n1674_ );
or   ( new_n1904_, new_n1855_, new_n919_ );
and  ( new_n1905_, new_n1904_, new_n1903_ );
nand ( new_n1906_, new_n1667_, new_n849_ );
nand ( new_n1907_, new_n1889_, new_n801_ );
and  ( new_n1908_, new_n1907_, new_n1906_ );
nor  ( new_n1909_, new_n1908_, new_n1905_ );
and  ( new_n1910_, new_n1698_, new_n1693_ );
xor  ( new_n1911_, new_n1908_, new_n1905_ );
and  ( new_n1912_, new_n1911_, new_n1910_ );
or   ( new_n1913_, new_n1912_, new_n1909_ );
or   ( new_n1914_, new_n1901_, new_n1867_ );
and  ( new_n1915_, new_n1914_, new_n1913_ );
or   ( new_n1916_, new_n1915_, new_n1902_ );
and  ( new_n1917_, new_n1852_, new_n818_ );
xor  ( new_n1918_, \b[3] , \a[8]  );
and  ( new_n1919_, new_n1918_, new_n817_ );
or   ( new_n1920_, new_n1919_, new_n1917_ );
and  ( new_n1921_, new_n1857_, new_n1673_ );
xor  ( new_n1922_, \b[7] , \a[4]  );
and  ( new_n1923_, new_n1922_, new_n918_ );
nor  ( new_n1924_, new_n1923_, new_n1921_ );
and  ( new_n1925_, new_n1886_, new_n1883_ );
xor  ( new_n1926_, \b[9] , \a[2]  );
and  ( new_n1927_, new_n1926_, new_n1868_ );
nor  ( new_n1928_, new_n1927_, new_n1925_ );
xor  ( new_n1929_, new_n1928_, new_n1924_ );
xor  ( new_n1930_, new_n1929_, new_n1920_ );
and  ( new_n1931_, new_n1898_, new_n1893_ );
not  ( new_n1932_, new_n1931_ );
nor  ( new_n1933_, new_n1865_, new_n1859_ );
and  ( new_n1934_, new_n1866_, new_n1854_ );
nor  ( new_n1935_, new_n1934_, new_n1933_ );
xor  ( new_n1936_, new_n1935_, new_n1932_ );
and  ( new_n1937_, new_n1891_, new_n849_ );
xor  ( new_n1938_, \b[5] , \a[6]  );
and  ( new_n1939_, new_n1938_, new_n801_ );
nor  ( new_n1940_, new_n1939_, new_n1937_ );
not  ( new_n1941_, new_n1940_ );
xor  ( new_n1942_, \b[9] , \b[10]  );
not  ( new_n1943_, new_n1942_ );
or   ( new_n1944_, new_n1943_, new_n98_ );
or   ( new_n1945_, new_n806_, \a[9]  );
and  ( new_n1946_, new_n808_, new_n352_ );
and  ( new_n1947_, \b[1] , \a[10]  );
or   ( new_n1948_, new_n1947_, new_n804_ );
or   ( new_n1949_, new_n1948_, new_n1946_ );
and  ( new_n1950_, new_n1949_, new_n1945_ );
xor  ( new_n1951_, new_n1950_, new_n1944_ );
xor  ( new_n1952_, new_n1951_, new_n1941_ );
xor  ( new_n1953_, new_n1952_, new_n1936_ );
xnor ( new_n1954_, new_n1953_, new_n1930_ );
and  ( new_n1955_, new_n1899_, new_n1888_ );
nor  ( new_n1956_, new_n1899_, new_n1888_ );
nor  ( new_n1957_, new_n1956_, new_n1882_ );
nor  ( new_n1958_, new_n1957_, new_n1955_ );
xor  ( new_n1959_, new_n1958_, new_n1954_ );
nor  ( new_n1960_, new_n1959_, new_n1916_ );
and  ( new_n1961_, new_n1959_, new_n1916_ );
nor  ( new_n1962_, new_n1684_, new_n1678_ );
and  ( new_n1963_, new_n1685_, new_n1670_ );
or   ( new_n1964_, new_n1963_, new_n1962_ );
xor  ( new_n1965_, new_n1880_, new_n1879_ );
or   ( new_n1966_, new_n1965_, new_n1964_ );
xor  ( new_n1967_, new_n1911_, new_n1910_ );
and  ( new_n1968_, new_n1965_, new_n1964_ );
or   ( new_n1969_, new_n1968_, new_n1967_ );
and  ( new_n1970_, new_n1969_, new_n1966_ );
xor  ( new_n1971_, new_n1901_, new_n1867_ );
xor  ( new_n1972_, new_n1971_, new_n1913_ );
nor  ( new_n1973_, new_n1972_, new_n1970_ );
and  ( new_n1974_, new_n1972_, new_n1970_ );
and  ( new_n1975_, new_n1699_, new_n1689_ );
and  ( new_n1976_, new_n1700_, new_n1686_ );
or   ( new_n1977_, new_n1976_, new_n1975_ );
xor  ( new_n1978_, new_n1965_, new_n1964_ );
xor  ( new_n1979_, new_n1978_, new_n1967_ );
nor  ( new_n1980_, new_n1979_, new_n1977_ );
and  ( new_n1981_, new_n1979_, new_n1977_ );
nor  ( new_n1982_, new_n1706_, new_n1702_ );
nor  ( new_n1983_, new_n1712_, new_n1708_ );
nor  ( new_n1984_, new_n1983_, new_n1982_ );
not  ( new_n1985_, new_n1984_ );
nor  ( new_n1986_, new_n1985_, new_n1981_ );
nor  ( new_n1987_, new_n1986_, new_n1980_ );
nor  ( new_n1988_, new_n1987_, new_n1974_ );
nor  ( new_n1989_, new_n1988_, new_n1973_ );
nor  ( new_n1990_, new_n1989_, new_n1961_ );
nor  ( new_n1991_, new_n1990_, new_n1960_ );
nand ( new_n1992_, new_n1918_, new_n818_ );
xor  ( new_n1993_, \b[3] , new_n137_ );
or   ( new_n1994_, new_n1993_, new_n895_ );
and  ( new_n1995_, new_n1994_, new_n1992_ );
xnor ( new_n1996_, new_n1995_, new_n1991_ );
nor  ( new_n1997_, new_n1928_, new_n1924_ );
and  ( new_n1998_, new_n1929_, new_n1920_ );
or   ( new_n1999_, new_n1998_, new_n1997_ );
or   ( new_n2000_, new_n806_, \a[10]  );
and  ( new_n2001_, new_n808_, new_n354_ );
and  ( new_n2002_, \b[1] , \a[11]  );
or   ( new_n2003_, new_n2002_, new_n804_ );
or   ( new_n2004_, new_n2003_, new_n2001_ );
and  ( new_n2005_, new_n2004_, new_n2000_ );
xor  ( new_n2006_, new_n2005_, new_n1999_ );
or   ( new_n2007_, new_n1950_, new_n1944_ );
nand ( new_n2008_, new_n1951_, new_n1941_ );
and  ( new_n2009_, new_n2008_, new_n2007_ );
and  ( new_n2010_, new_n1038_, new_n98_ );
nor  ( new_n2011_, new_n2010_, new_n1154_ );
and  ( new_n2012_, \b[10] , \a[0]  );
not  ( new_n2013_, new_n2012_ );
and  ( new_n2014_, new_n2013_, new_n1154_ );
or   ( new_n2015_, new_n2014_, new_n1942_ );
or   ( new_n2016_, new_n2015_, new_n2011_ );
xor  ( new_n2017_, \b[11] , new_n108_ );
or   ( new_n2018_, new_n2017_, new_n1943_ );
and  ( new_n2019_, new_n2018_, new_n2016_ );
xor  ( new_n2020_, new_n2019_, new_n2009_ );
or   ( new_n2021_, new_n2010_, new_n1296_ );
and  ( new_n2022_, new_n2013_, \b[11]  );
and  ( new_n2023_, new_n2022_, new_n2021_ );
xor  ( new_n2024_, new_n2023_, new_n2020_ );
xor  ( new_n2025_, new_n2024_, new_n2006_ );
and  ( new_n2026_, new_n1953_, new_n1930_ );
nor  ( new_n2027_, new_n1953_, new_n1930_ );
nor  ( new_n2028_, new_n1958_, new_n2027_ );
or   ( new_n2029_, new_n2028_, new_n2026_ );
nand ( new_n2030_, new_n1922_, new_n1673_ );
xor  ( new_n2031_, \b[7] , new_n176_ );
or   ( new_n2032_, new_n2031_, new_n919_ );
and  ( new_n2033_, new_n2032_, new_n2030_ );
xor  ( new_n2034_, new_n2033_, new_n2029_ );
xor  ( new_n2035_, new_n2034_, new_n2025_ );
nor  ( new_n2036_, new_n1935_, new_n1932_ );
and  ( new_n2037_, new_n1952_, new_n1936_ );
or   ( new_n2038_, new_n2037_, new_n2036_ );
and  ( new_n2039_, new_n1926_, new_n1886_ );
xor  ( new_n2040_, \b[9] , \a[3]  );
and  ( new_n2041_, new_n2040_, new_n1868_ );
or   ( new_n2042_, new_n2041_, new_n2039_ );
nand ( new_n2043_, new_n1938_, new_n849_ );
xor  ( new_n2044_, \b[5] , new_n185_ );
or   ( new_n2045_, new_n2044_, new_n802_ );
and  ( new_n2046_, new_n2045_, new_n2043_ );
xor  ( new_n2047_, new_n2046_, new_n2042_ );
xor  ( new_n2048_, new_n2047_, new_n2038_ );
xor  ( new_n2049_, new_n2048_, new_n2035_ );
xor  ( new_n2050_, new_n2049_, new_n1996_ );
and  ( new_n2051_, new_n2050_, new_n1849_ );
not  ( new_n2052_, new_n2051_ );
and  ( new_n2053_, new_n2052_, \d[15]  );
not  ( new_n2054_, new_n2053_ );
xor  ( new_n2055_, new_n1972_, new_n1970_ );
xnor ( new_n2056_, new_n2055_, new_n1987_ );
xor  ( new_n2057_, new_n1959_, new_n1916_ );
xnor ( new_n2058_, new_n2057_, new_n1989_ );
xor  ( new_n2059_, new_n1979_, new_n1977_ );
xor  ( new_n2060_, new_n2059_, new_n1984_ );
not  ( new_n2061_, new_n1844_ );
not  ( new_n2062_, new_n1780_ );
and  ( new_n2063_, \b[1] , \a[0]  );
xor  ( new_n2064_, new_n2063_, new_n897_ );
not  ( new_n2065_, new_n2064_ );
xor  ( new_n2066_, new_n900_, new_n894_ );
not  ( new_n2067_, new_n2066_ );
and  ( new_n2068_, new_n2067_, new_n2065_ );
and  ( new_n2069_, new_n2068_, new_n1849_ );
and  ( new_n2070_, new_n2069_, new_n2062_ );
and  ( new_n2071_, new_n2070_, new_n2061_ );
and  ( new_n2072_, new_n2071_, new_n938_ );
and  ( new_n2073_, new_n2072_, new_n1714_ );
and  ( new_n2074_, new_n2073_, new_n2060_ );
and  ( new_n2075_, new_n2074_, new_n2058_ );
not  ( new_n2076_, new_n2075_ );
and  ( new_n2077_, new_n2076_, new_n2056_ );
and  ( new_n2078_, new_n2077_, new_n2050_ );
not  ( new_n2079_, new_n2078_ );
and  ( new_n2080_, new_n2079_, \a[15]  );
not  ( new_n2081_, new_n2080_ );
and  ( new_n2082_, new_n2065_, new_n2056_ );
not  ( new_n2083_, new_n2082_ );
not  ( new_n2084_, new_n2058_ );
and  ( new_n2085_, new_n2084_, \c[15]  );
nor  ( new_n2086_, new_n2085_, new_n2083_ );
nor  ( new_n2087_, new_n2086_, new_n1783_ );
not  ( new_n2088_, new_n2087_ );
not  ( new_n2089_, new_n2060_ );
xor  ( new_n2090_, \d[1] , \a[1]  );
xor  ( new_n2091_, \d[0] , \a[0]  );
and  ( new_n2092_, new_n150_, new_n163_ );
and  ( new_n2093_, new_n726_, new_n115_ );
and  ( new_n2094_, new_n2093_, new_n2092_ );
and  ( new_n2095_, new_n2094_, new_n2091_ );
and  ( new_n2096_, new_n2095_, new_n2090_ );
and  ( new_n2097_, new_n179_, new_n133_ );
and  ( new_n2098_, new_n171_, new_n137_ );
and  ( new_n2099_, new_n2098_, new_n2097_ );
and  ( new_n2100_, new_n326_, new_n352_ );
and  ( new_n2101_, new_n255_, new_n1719_ );
and  ( new_n2102_, new_n2101_, new_n2100_ );
and  ( new_n2103_, new_n2102_, new_n2099_ );
and  ( new_n2104_, new_n66_, new_n176_ );
and  ( new_n2105_, new_n660_, new_n231_ );
and  ( new_n2106_, new_n2105_, new_n2104_ );
and  ( new_n2107_, new_n128_, new_n185_ );
and  ( new_n2108_, new_n563_, new_n212_ );
and  ( new_n2109_, new_n2108_, new_n2107_ );
and  ( new_n2110_, new_n2109_, new_n2106_ );
and  ( new_n2111_, new_n2110_, new_n2103_ );
and  ( new_n2112_, new_n2111_, new_n2096_ );
and  ( new_n2113_, new_n2112_, new_n2089_ );
nor  ( new_n2114_, new_n2113_, new_n2066_ );
nor  ( new_n2115_, new_n2114_, new_n1653_ );
not  ( new_n2116_, \a[14]  );
and  ( new_n2117_, new_n256_, new_n2116_ );
and  ( new_n2118_, new_n75_, new_n354_ );
and  ( new_n2119_, new_n2118_, new_n2117_ );
and  ( new_n2120_, new_n99_, new_n85_ );
and  ( new_n2121_, new_n103_, new_n89_ );
and  ( new_n2122_, new_n2121_, new_n2120_ );
and  ( new_n2123_, new_n2122_, new_n2119_ );
and  ( new_n2124_, new_n2123_, new_n2112_ );
nor  ( new_n2125_, new_n2124_, \d[15]  );
and  ( new_n2126_, new_n2125_, new_n2089_ );
nor  ( new_n2127_, new_n2126_, new_n2115_ );
and  ( new_n2128_, new_n2127_, new_n2088_ );
and  ( new_n2129_, new_n2128_, new_n2081_ );
and  ( new_n2130_, new_n2129_, new_n2054_ );
and  ( new_n2131_, new_n2130_, new_n1846_ );
and  ( new_n2132_, new_n2131_, new_n1782_ );
and  ( new_n2133_, new_n2132_, new_n1718_ );
and  ( new_n2134_, new_n2133_, new_n942_ );
xor  ( new_n2135_, new_n459_, new_n457_ );
xor  ( new_n2136_, new_n2135_, new_n783_ );
nor  ( new_n2137_, new_n2136_, new_n938_ );
not  ( new_n2138_, new_n2137_ );
xor  ( new_n2139_, new_n1269_, new_n1267_ );
and  ( new_n2140_, new_n2139_, new_n1593_ );
not  ( new_n2141_, new_n2140_ );
nor  ( new_n2142_, new_n2139_, new_n1593_ );
nor  ( new_n2143_, new_n2142_, new_n1714_ );
and  ( new_n2144_, new_n2143_, new_n2141_ );
not  ( new_n2145_, new_n2144_ );
not  ( new_n2146_, new_n2050_ );
not  ( new_n2147_, new_n2121_ );
and  ( new_n2148_, new_n2147_, new_n2146_ );
not  ( new_n2149_, new_n2148_ );
not  ( new_n2150_, new_n2077_ );
and  ( new_n2151_, new_n2150_, \a[13]  );
not  ( new_n2152_, new_n2151_ );
and  ( new_n2153_, new_n2084_, \c[13]  );
nor  ( new_n2154_, new_n2153_, new_n2083_ );
nor  ( new_n2155_, new_n2154_, new_n992_ );
not  ( new_n2156_, new_n2155_ );
xor  ( new_n2157_, \d[13] , \c[13]  );
and  ( new_n2158_, new_n2157_, new_n2089_ );
not  ( new_n2159_, new_n2158_ );
and  ( new_n2160_, new_n1848_, \d[13]  );
and  ( new_n2161_, new_n2066_, \c[13]  );
nor  ( new_n2162_, new_n2161_, new_n2160_ );
and  ( new_n2163_, new_n2162_, new_n2159_ );
and  ( new_n2164_, new_n2163_, new_n2156_ );
and  ( new_n2165_, new_n2164_, new_n2152_ );
and  ( new_n2166_, new_n2165_, new_n2149_ );
xor  ( new_n2167_, \c[13] , \a[13]  );
xnor ( new_n2168_, new_n2167_, new_n1773_ );
not  ( new_n2169_, new_n2168_ );
and  ( new_n2170_, new_n2169_, new_n1780_ );
xor  ( new_n2171_, \d[13] , \b[13]  );
xnor ( new_n2172_, new_n2171_, new_n1837_ );
not  ( new_n2173_, new_n2172_ );
and  ( new_n2174_, new_n2173_, new_n1844_ );
nor  ( new_n2175_, new_n2174_, new_n2170_ );
and  ( new_n2176_, new_n2175_, new_n2166_ );
and  ( new_n2177_, new_n2176_, new_n2145_ );
and  ( new_n2178_, new_n2177_, new_n2138_ );
xor  ( new_n2179_, new_n411_, new_n401_ );
and  ( new_n2180_, new_n2179_, new_n786_ );
not  ( new_n2181_, new_n2180_ );
nor  ( new_n2182_, new_n2179_, new_n786_ );
nor  ( new_n2183_, new_n2182_, new_n938_ );
and  ( new_n2184_, new_n2183_, new_n2181_ );
not  ( new_n2185_, new_n2184_ );
xor  ( new_n2186_, new_n1220_, new_n1218_ );
and  ( new_n2187_, new_n2186_, new_n1595_ );
not  ( new_n2188_, new_n2187_ );
nor  ( new_n2189_, new_n2186_, new_n1595_ );
nor  ( new_n2190_, new_n2189_, new_n1714_ );
and  ( new_n2191_, new_n2190_, new_n2188_ );
not  ( new_n2192_, new_n2191_ );
xor  ( new_n2193_, \c[14] , \a[14]  );
xnor ( new_n2194_, new_n2193_, new_n1775_ );
not  ( new_n2195_, new_n2194_ );
and  ( new_n2196_, new_n2195_, new_n1780_ );
not  ( new_n2197_, new_n2196_ );
xor  ( new_n2198_, \d[14] , \b[14]  );
xnor ( new_n2199_, new_n2198_, new_n1839_ );
not  ( new_n2200_, new_n2199_ );
and  ( new_n2201_, new_n2200_, new_n1844_ );
not  ( new_n2202_, new_n2201_ );
not  ( new_n2203_, new_n2117_ );
and  ( new_n2204_, new_n2203_, new_n2146_ );
not  ( new_n2205_, new_n2204_ );
not  ( new_n2206_, \b[14]  );
and  ( new_n2207_, new_n2084_, \c[14]  );
nor  ( new_n2208_, new_n2207_, new_n2083_ );
nor  ( new_n2209_, new_n2208_, new_n2206_ );
not  ( new_n2210_, new_n2209_ );
and  ( new_n2211_, new_n2150_, \a[14]  );
not  ( new_n2212_, new_n2211_ );
xor  ( new_n2213_, \d[14] , \c[14]  );
and  ( new_n2214_, new_n2213_, new_n2089_ );
not  ( new_n2215_, new_n2214_ );
and  ( new_n2216_, new_n1848_, \d[14]  );
and  ( new_n2217_, new_n2066_, \c[14]  );
nor  ( new_n2218_, new_n2217_, new_n2216_ );
and  ( new_n2219_, new_n2218_, new_n2215_ );
and  ( new_n2220_, new_n2219_, new_n2212_ );
and  ( new_n2221_, new_n2220_, new_n2210_ );
and  ( new_n2222_, new_n2221_, new_n2205_ );
and  ( new_n2223_, new_n2222_, new_n2202_ );
and  ( new_n2224_, new_n2223_, new_n2197_ );
and  ( new_n2225_, new_n2224_, new_n2192_ );
and  ( new_n2226_, new_n2225_, new_n2185_ );
and  ( new_n2227_, new_n2226_, new_n2178_ );
not  ( new_n2228_, new_n2227_ );
nor  ( new_n2229_, new_n2228_, new_n2134_ );
nor  ( new_n2230_, new_n2226_, new_n2178_ );
and  ( new_n2231_, new_n2230_, new_n2134_ );
nor  ( new_n2232_, new_n2231_, new_n2229_ );
not  ( new_n2233_, new_n2134_ );
and  ( new_n2234_, new_n103_, new_n1066_ );
and  ( new_n2235_, \d[13] , \c[13]  );
and  ( new_n2236_, new_n99_, new_n969_ );
and  ( new_n2237_, \d[12] , \c[12]  );
and  ( new_n2238_, new_n75_, new_n952_ );
and  ( new_n2239_, \d[11] , \c[11]  );
and  ( new_n2240_, new_n326_, new_n1127_ );
and  ( new_n2241_, \d[10] , \c[10]  );
and  ( new_n2242_, new_n171_, new_n1003_ );
and  ( new_n2243_, \d[9] , \c[9]  );
and  ( new_n2244_, new_n179_, new_n1010_ );
and  ( new_n2245_, \d[8] , \c[8]  );
and  ( new_n2246_, new_n128_, new_n1000_ );
and  ( new_n2247_, \d[7] , \c[7]  );
and  ( new_n2248_, new_n563_, new_n1373_ );
and  ( new_n2249_, \d[6] , \c[6]  );
and  ( new_n2250_, new_n66_, new_n943_ );
and  ( new_n2251_, \d[5] , \c[5]  );
and  ( new_n2252_, new_n660_, new_n1468_ );
and  ( new_n2253_, \d[4] , \c[4]  );
and  ( new_n2254_, new_n150_, new_n978_ );
and  ( new_n2255_, \d[3] , \c[3]  );
and  ( new_n2256_, new_n726_, new_n1534_ );
and  ( new_n2257_, \d[2] , \c[2]  );
and  ( new_n2258_, new_n90_, new_n1104_ );
and  ( new_n2259_, \d[1] , \c[1]  );
and  ( new_n2260_, \d[0] , \c[0]  );
nor  ( new_n2261_, new_n2260_, new_n2259_ );
nor  ( new_n2262_, new_n2261_, new_n2258_ );
nor  ( new_n2263_, new_n2262_, new_n2257_ );
nor  ( new_n2264_, new_n2263_, new_n2256_ );
nor  ( new_n2265_, new_n2264_, new_n2255_ );
nor  ( new_n2266_, new_n2265_, new_n2254_ );
nor  ( new_n2267_, new_n2266_, new_n2253_ );
nor  ( new_n2268_, new_n2267_, new_n2252_ );
nor  ( new_n2269_, new_n2268_, new_n2251_ );
nor  ( new_n2270_, new_n2269_, new_n2250_ );
nor  ( new_n2271_, new_n2270_, new_n2249_ );
nor  ( new_n2272_, new_n2271_, new_n2248_ );
nor  ( new_n2273_, new_n2272_, new_n2247_ );
nor  ( new_n2274_, new_n2273_, new_n2246_ );
nor  ( new_n2275_, new_n2274_, new_n2245_ );
nor  ( new_n2276_, new_n2275_, new_n2244_ );
nor  ( new_n2277_, new_n2276_, new_n2243_ );
nor  ( new_n2278_, new_n2277_, new_n2242_ );
nor  ( new_n2279_, new_n2278_, new_n2241_ );
nor  ( new_n2280_, new_n2279_, new_n2240_ );
nor  ( new_n2281_, new_n2280_, new_n2239_ );
nor  ( new_n2282_, new_n2281_, new_n2238_ );
nor  ( new_n2283_, new_n2282_, new_n2237_ );
nor  ( new_n2284_, new_n2283_, new_n2236_ );
nor  ( new_n2285_, new_n2284_, new_n2235_ );
nor  ( new_n2286_, new_n2285_, new_n2234_ );
not  ( new_n2287_, new_n2286_ );
xor  ( new_n2288_, new_n2287_, new_n2213_ );
xor  ( new_n2289_, new_n2288_, new_n2233_ );
nor  ( new_n2290_, new_n2289_, new_n2232_ );
and  ( new_n2291_, new_n256_, new_n1624_ );
and  ( new_n2292_, \d[14] , \c[14]  );
nor  ( new_n2293_, new_n2286_, new_n2292_ );
nor  ( new_n2294_, new_n2293_, new_n2291_ );
not  ( new_n2295_, new_n2294_ );
xor  ( new_n2296_, \d[15] , \c[15]  );
xor  ( new_n2297_, new_n2296_, new_n2295_ );
xor  ( new_n2298_, new_n2297_, new_n2233_ );
not  ( new_n2299_, new_n2178_ );
xor  ( new_n2300_, new_n2226_, new_n2299_ );
nor  ( new_n2301_, new_n2300_, new_n2298_ );
nor  ( new_n2302_, new_n2301_, new_n2290_ );
not  ( new_n2303_, new_n2302_ );
xnor ( new_n2304_, new_n2284_, new_n2157_ );
or   ( new_n2305_, new_n2304_, new_n2134_ );
or   ( new_n2306_, new_n2077_, new_n85_ );
or   ( new_n2307_, new_n2082_, new_n1053_ );
or   ( new_n2308_, new_n2060_, \c[12]  );
and  ( new_n2309_, new_n2308_, new_n1849_ );
or   ( new_n2310_, new_n2309_, new_n99_ );
and  ( new_n2311_, new_n2310_, new_n2307_ );
and  ( new_n2312_, new_n2311_, new_n2306_ );
xor  ( new_n2313_, \c[12] , \a[12]  );
xnor ( new_n2314_, new_n2313_, new_n1771_ );
or   ( new_n2315_, new_n2314_, new_n2062_ );
or   ( new_n2316_, new_n2058_, new_n1053_ );
or   ( new_n2317_, new_n2060_, \d[12]  );
and  ( new_n2318_, new_n2317_, new_n2067_ );
and  ( new_n2319_, new_n2318_, new_n2316_ );
or   ( new_n2320_, new_n2319_, new_n969_ );
xor  ( new_n2321_, \d[12] , \b[12]  );
xnor ( new_n2322_, new_n2321_, new_n1835_ );
or   ( new_n2323_, new_n2322_, new_n2061_ );
and  ( new_n2324_, new_n2323_, new_n2320_ );
and  ( new_n2325_, new_n2324_, new_n2315_ );
and  ( new_n2326_, new_n2325_, new_n2312_ );
xor  ( new_n2327_, new_n1317_, new_n1273_ );
not  ( new_n2328_, new_n2327_ );
nor  ( new_n2329_, new_n2328_, new_n1590_ );
and  ( new_n2330_, new_n2328_, new_n1590_ );
or   ( new_n2331_, new_n2330_, new_n1714_ );
or   ( new_n2332_, new_n2331_, new_n2329_ );
or   ( new_n2333_, new_n2120_, new_n2050_ );
xor  ( new_n2334_, new_n506_, new_n463_ );
not  ( new_n2335_, new_n2334_ );
nor  ( new_n2336_, new_n2335_, new_n781_ );
and  ( new_n2337_, new_n2335_, new_n781_ );
or   ( new_n2338_, new_n2337_, new_n938_ );
or   ( new_n2339_, new_n2338_, new_n2336_ );
and  ( new_n2340_, new_n2339_, new_n2333_ );
and  ( new_n2341_, new_n2340_, new_n2332_ );
and  ( new_n2342_, new_n2341_, new_n2326_ );
not  ( new_n2343_, new_n2118_ );
and  ( new_n2344_, new_n2343_, new_n2146_ );
not  ( new_n2345_, new_n2344_ );
and  ( new_n2346_, new_n2075_, \a[11]  );
not  ( new_n2347_, new_n2346_ );
xor  ( new_n2348_, \d[11] , \b[11]  );
xnor ( new_n2349_, new_n2348_, new_n1833_ );
not  ( new_n2350_, new_n2349_ );
and  ( new_n2351_, new_n2350_, new_n1844_ );
not  ( new_n2352_, new_n2351_ );
not  ( new_n2353_, new_n2056_ );
and  ( new_n2354_, new_n1154_, new_n354_ );
not  ( new_n2355_, new_n2354_ );
and  ( new_n2356_, new_n2355_, new_n2353_ );
not  ( new_n2357_, new_n2356_ );
xor  ( new_n2358_, \d[11] , \c[11]  );
and  ( new_n2359_, new_n2358_, new_n2089_ );
not  ( new_n2360_, new_n2359_ );
and  ( new_n2361_, new_n1848_, \d[11]  );
not  ( new_n2362_, new_n2361_ );
and  ( new_n2363_, new_n2064_, \b[11]  );
and  ( new_n2364_, new_n2066_, \c[11]  );
nor  ( new_n2365_, new_n2364_, new_n2363_ );
and  ( new_n2366_, new_n2365_, new_n2362_ );
and  ( new_n2367_, new_n2366_, new_n2360_ );
and  ( new_n2368_, new_n2367_, new_n2357_ );
and  ( new_n2369_, new_n2368_, new_n2352_ );
and  ( new_n2370_, \c[11] , \b[11]  );
and  ( new_n2371_, new_n2370_, new_n2084_ );
xor  ( new_n2372_, \c[11] , \a[11]  );
xnor ( new_n2373_, new_n2372_, new_n1769_ );
not  ( new_n2374_, new_n2373_ );
and  ( new_n2375_, new_n2374_, new_n1780_ );
nor  ( new_n2376_, new_n2375_, new_n2371_ );
and  ( new_n2377_, new_n2376_, new_n2369_ );
and  ( new_n2378_, new_n2377_, new_n2347_ );
not  ( new_n2379_, new_n779_ );
xor  ( new_n2380_, new_n546_, new_n544_ );
and  ( new_n2381_, new_n2380_, new_n2379_ );
not  ( new_n2382_, new_n2381_ );
nor  ( new_n2383_, new_n2380_, new_n2379_ );
nor  ( new_n2384_, new_n2383_, new_n938_ );
and  ( new_n2385_, new_n2384_, new_n2382_ );
not  ( new_n2386_, new_n1588_ );
xor  ( new_n2387_, new_n1356_, new_n1354_ );
and  ( new_n2388_, new_n2387_, new_n2386_ );
not  ( new_n2389_, new_n2388_ );
nor  ( new_n2390_, new_n2387_, new_n2386_ );
nor  ( new_n2391_, new_n2390_, new_n1714_ );
and  ( new_n2392_, new_n2391_, new_n2389_ );
nor  ( new_n2393_, new_n2392_, new_n2385_ );
and  ( new_n2394_, new_n2393_, new_n2378_ );
and  ( new_n2395_, new_n2394_, new_n2345_ );
nor  ( new_n2396_, new_n2395_, new_n2342_ );
not  ( new_n2397_, new_n2396_ );
and  ( new_n2398_, new_n2397_, new_n2178_ );
and  ( new_n2399_, new_n2395_, new_n2342_ );
not  ( new_n2400_, new_n2399_ );
and  ( new_n2401_, new_n2400_, new_n2299_ );
nor  ( new_n2402_, new_n2401_, new_n2398_ );
not  ( new_n2403_, new_n2402_ );
and  ( new_n2404_, new_n255_, new_n1653_ );
and  ( new_n2405_, \d[15] , \c[15]  );
nor  ( new_n2406_, new_n2405_, new_n2294_ );
nor  ( new_n2407_, new_n2406_, new_n2404_ );
xor  ( new_n2408_, new_n2407_, new_n2178_ );
or   ( new_n2409_, new_n2408_, new_n2403_ );
and  ( new_n2410_, new_n2397_, new_n2299_ );
not  ( new_n2411_, new_n2410_ );
or   ( new_n2412_, new_n2411_, new_n2399_ );
and  ( new_n2413_, new_n2412_, new_n2409_ );
nor  ( new_n2414_, new_n2413_, new_n2305_ );
and  ( new_n2415_, new_n2414_, new_n2303_ );
nor  ( new_n2416_, new_n2298_, new_n2232_ );
xor  ( new_n2417_, new_n2407_, new_n2134_ );
nor  ( new_n2418_, new_n2417_, new_n2300_ );
or   ( new_n2419_, new_n2418_, new_n2416_ );
not  ( new_n2420_, new_n2288_ );
and  ( new_n2421_, new_n2420_, new_n2233_ );
xor  ( new_n2422_, new_n2411_, new_n2421_ );
xor  ( new_n2423_, new_n2422_, new_n2419_ );
nand ( new_n2424_, new_n2413_, new_n2305_ );
nor  ( new_n2425_, new_n2424_, new_n2303_ );
nor  ( new_n2426_, new_n2425_, new_n2415_ );
and  ( new_n2427_, new_n2426_, new_n2423_ );
nor  ( new_n2428_, new_n2427_, new_n2415_ );
and  ( new_n2429_, new_n2411_, new_n2421_ );
and  ( new_n2430_, new_n2422_, new_n2419_ );
or   ( new_n2431_, new_n2430_, new_n2429_ );
or   ( new_n2432_, new_n2297_, new_n2134_ );
or   ( new_n2433_, new_n2417_, new_n2232_ );
or   ( new_n2434_, new_n2300_, new_n2134_ );
and  ( new_n2435_, new_n2434_, new_n2433_ );
xor  ( new_n2436_, new_n2435_, new_n2432_ );
xor  ( new_n2437_, new_n2436_, new_n2431_ );
xor  ( new_n2438_, new_n2437_, new_n2428_ );
xor  ( new_n2439_, \d[12] , \c[12]  );
xnor ( new_n2440_, new_n2439_, new_n2282_ );
not  ( new_n2441_, new_n2440_ );
and  ( new_n2442_, new_n2441_, new_n2233_ );
xor  ( new_n2443_, new_n2297_, new_n2299_ );
or   ( new_n2444_, new_n2443_, new_n2403_ );
xor  ( new_n2445_, new_n2395_, new_n2342_ );
not  ( new_n2446_, new_n2445_ );
or   ( new_n2447_, new_n2446_, new_n2408_ );
nand ( new_n2448_, new_n2447_, new_n2444_ );
nand ( new_n2449_, new_n2448_, new_n2442_ );
xnor ( new_n2450_, new_n2448_, new_n2442_ );
or   ( new_n2451_, new_n2100_, new_n2050_ );
or   ( new_n2452_, new_n2076_, new_n352_ );
or   ( new_n2453_, new_n1127_, new_n1038_ );
or   ( new_n2454_, new_n2453_, new_n2058_ );
xor  ( new_n2455_, \d[10] , \b[10]  );
xnor ( new_n2456_, new_n2455_, new_n1831_ );
or   ( new_n2457_, new_n2456_, new_n2061_ );
xor  ( new_n2458_, \d[10] , \c[10]  );
nand ( new_n2459_, new_n2458_, new_n2089_ );
or   ( new_n2460_, new_n1849_, new_n326_ );
or   ( new_n2461_, new_n2067_, new_n1127_ );
or   ( new_n2462_, new_n2065_, new_n1038_ );
and  ( new_n2463_, new_n2462_, new_n2461_ );
and  ( new_n2464_, new_n2463_, new_n2460_ );
and  ( new_n2465_, new_n2464_, new_n2459_ );
and  ( new_n2466_, new_n2465_, new_n2457_ );
and  ( new_n2467_, new_n1038_, new_n352_ );
or   ( new_n2468_, new_n2467_, new_n2056_ );
xor  ( new_n2469_, \c[10] , \a[10]  );
xnor ( new_n2470_, new_n2469_, new_n1767_ );
or   ( new_n2471_, new_n2470_, new_n2062_ );
and  ( new_n2472_, new_n2471_, new_n2468_ );
and  ( new_n2473_, new_n2472_, new_n2466_ );
and  ( new_n2474_, new_n2473_, new_n2454_ );
xor  ( new_n2475_, new_n1396_, new_n1359_ );
not  ( new_n2476_, new_n2475_ );
nor  ( new_n2477_, new_n2476_, new_n1586_ );
and  ( new_n2478_, new_n2476_, new_n1586_ );
or   ( new_n2479_, new_n2478_, new_n1714_ );
or   ( new_n2480_, new_n2479_, new_n2477_ );
xor  ( new_n2481_, new_n586_, new_n549_ );
not  ( new_n2482_, new_n2481_ );
nor  ( new_n2483_, new_n2482_, new_n777_ );
and  ( new_n2484_, new_n2482_, new_n777_ );
or   ( new_n2485_, new_n2484_, new_n938_ );
or   ( new_n2486_, new_n2485_, new_n2483_ );
and  ( new_n2487_, new_n2486_, new_n2480_ );
and  ( new_n2488_, new_n2487_, new_n2474_ );
and  ( new_n2489_, new_n2488_, new_n2452_ );
and  ( new_n2490_, new_n2489_, new_n2451_ );
not  ( new_n2491_, new_n2098_ );
and  ( new_n2492_, new_n2491_, new_n2146_ );
not  ( new_n2493_, new_n2492_ );
and  ( new_n2494_, new_n2075_, \a[9]  );
not  ( new_n2495_, new_n2494_ );
and  ( new_n2496_, \c[9] , \b[9]  );
and  ( new_n2497_, new_n2496_, new_n2084_ );
not  ( new_n2498_, new_n2497_ );
not  ( new_n2499_, new_n775_ );
xor  ( new_n2500_, new_n618_, new_n616_ );
and  ( new_n2501_, new_n2500_, new_n2499_ );
not  ( new_n2502_, new_n2501_ );
nor  ( new_n2503_, new_n2500_, new_n2499_ );
nor  ( new_n2504_, new_n2503_, new_n938_ );
and  ( new_n2505_, new_n2504_, new_n2502_ );
not  ( new_n2506_, new_n2505_ );
xor  ( new_n2507_, \d[9] , \b[9]  );
xnor ( new_n2508_, new_n2507_, new_n1829_ );
not  ( new_n2509_, new_n2508_ );
and  ( new_n2510_, new_n2509_, new_n1844_ );
not  ( new_n2511_, new_n2510_ );
and  ( new_n2512_, new_n1848_, \d[9]  );
not  ( new_n2513_, new_n2512_ );
and  ( new_n2514_, new_n2066_, \c[9]  );
and  ( new_n2515_, new_n2064_, \b[9]  );
nor  ( new_n2516_, new_n2515_, new_n2514_ );
and  ( new_n2517_, new_n2516_, new_n2513_ );
and  ( new_n2518_, new_n2517_, new_n2511_ );
xor  ( new_n2519_, \d[9] , \c[9]  );
and  ( new_n2520_, new_n2519_, new_n2089_ );
xor  ( new_n2521_, \c[9] , \a[9]  );
xnor ( new_n2522_, new_n2521_, new_n1765_ );
not  ( new_n2523_, new_n2522_ );
and  ( new_n2524_, new_n2523_, new_n1780_ );
nor  ( new_n2525_, new_n2524_, new_n2520_ );
and  ( new_n2526_, new_n2525_, new_n2518_ );
and  ( new_n2527_, new_n2526_, new_n2506_ );
and  ( new_n2528_, new_n1296_, new_n137_ );
not  ( new_n2529_, new_n2528_ );
and  ( new_n2530_, new_n2529_, new_n2353_ );
not  ( new_n2531_, new_n1584_ );
xor  ( new_n2532_, new_n1428_, new_n1401_ );
and  ( new_n2533_, new_n2532_, new_n2531_ );
not  ( new_n2534_, new_n2533_ );
nor  ( new_n2535_, new_n2532_, new_n2531_ );
nor  ( new_n2536_, new_n2535_, new_n1714_ );
and  ( new_n2537_, new_n2536_, new_n2534_ );
nor  ( new_n2538_, new_n2537_, new_n2530_ );
and  ( new_n2539_, new_n2538_, new_n2527_ );
and  ( new_n2540_, new_n2539_, new_n2498_ );
and  ( new_n2541_, new_n2540_, new_n2495_ );
and  ( new_n2542_, new_n2541_, new_n2493_ );
nor  ( new_n2543_, new_n2542_, new_n2490_ );
nor  ( new_n2544_, new_n2543_, new_n2395_ );
or   ( new_n2545_, new_n2544_, new_n2450_ );
and  ( new_n2546_, new_n2545_, new_n2449_ );
xor  ( new_n2547_, new_n2413_, new_n2305_ );
xor  ( new_n2548_, new_n2547_, new_n2303_ );
or   ( new_n2549_, new_n2548_, new_n2546_ );
xor  ( new_n2550_, new_n2304_, new_n2233_ );
or   ( new_n2551_, new_n2550_, new_n2232_ );
or   ( new_n2552_, new_n2300_, new_n2289_ );
and  ( new_n2553_, new_n2552_, new_n2551_ );
not  ( new_n2554_, new_n2395_ );
nor  ( new_n2555_, new_n2543_, new_n2554_ );
and  ( new_n2556_, new_n2542_, new_n2490_ );
nor  ( new_n2557_, new_n2556_, new_n2395_ );
nor  ( new_n2558_, new_n2557_, new_n2555_ );
not  ( new_n2559_, new_n2558_ );
xor  ( new_n2560_, new_n2407_, new_n2395_ );
or   ( new_n2561_, new_n2560_, new_n2559_ );
not  ( new_n2562_, new_n2556_ );
nand ( new_n2563_, new_n2562_, new_n2544_ );
and  ( new_n2564_, new_n2563_, new_n2561_ );
nor  ( new_n2565_, new_n2564_, new_n2553_ );
xnor ( new_n2566_, new_n2358_, new_n2280_ );
or   ( new_n2567_, new_n2566_, new_n2134_ );
xor  ( new_n2568_, new_n2288_, new_n2299_ );
or   ( new_n2569_, new_n2568_, new_n2403_ );
or   ( new_n2570_, new_n2446_, new_n2443_ );
and  ( new_n2571_, new_n2570_, new_n2569_ );
nor  ( new_n2572_, new_n2571_, new_n2567_ );
xor  ( new_n2573_, new_n2440_, new_n2233_ );
nor  ( new_n2574_, new_n2573_, new_n2232_ );
nor  ( new_n2575_, new_n2550_, new_n2300_ );
or   ( new_n2576_, new_n2575_, new_n2574_ );
xor  ( new_n2577_, new_n2571_, new_n2567_ );
and  ( new_n2578_, new_n2577_, new_n2576_ );
or   ( new_n2579_, new_n2578_, new_n2572_ );
xor  ( new_n2580_, new_n2564_, new_n2553_ );
and  ( new_n2581_, new_n2580_, new_n2579_ );
nor  ( new_n2582_, new_n2581_, new_n2565_ );
xnor ( new_n2583_, new_n2548_, new_n2546_ );
or   ( new_n2584_, new_n2583_, new_n2582_ );
and  ( new_n2585_, new_n2584_, new_n2549_ );
xnor ( new_n2586_, new_n2426_, new_n2423_ );
or   ( new_n2587_, new_n2586_, new_n2585_ );
and  ( new_n2588_, new_n2586_, new_n2585_ );
xnor ( new_n2589_, new_n2583_, new_n2582_ );
xor  ( new_n2590_, new_n2544_, new_n2450_ );
xor  ( new_n2591_, new_n2580_, new_n2579_ );
nand ( new_n2592_, new_n2591_, new_n2590_ );
nor  ( new_n2593_, new_n2591_, new_n2590_ );
xor  ( new_n2594_, new_n2577_, new_n2576_ );
nand ( new_n2595_, new_n2594_, new_n2564_ );
nor  ( new_n2596_, new_n2594_, new_n2564_ );
xor  ( new_n2597_, new_n2566_, new_n2233_ );
or   ( new_n2598_, new_n2597_, new_n2232_ );
or   ( new_n2599_, new_n2573_, new_n2300_ );
and  ( new_n2600_, new_n2599_, new_n2598_ );
xor  ( new_n2601_, new_n2395_, new_n2297_ );
nand ( new_n2602_, new_n2601_, new_n2558_ );
xor  ( new_n2603_, new_n2542_, new_n2490_ );
not  ( new_n2604_, new_n2603_ );
or   ( new_n2605_, new_n2604_, new_n2560_ );
and  ( new_n2606_, new_n2605_, new_n2602_ );
or   ( new_n2607_, new_n2606_, new_n2600_ );
and  ( new_n2608_, new_n2606_, new_n2600_ );
or   ( new_n2609_, new_n2077_, new_n133_ );
and  ( new_n2610_, new_n2609_, new_n2050_ );
or   ( new_n2611_, new_n2610_, new_n2097_ );
or   ( new_n2612_, new_n2058_, new_n1010_ );
and  ( new_n2613_, new_n2612_, new_n2056_ );
or   ( new_n2614_, new_n2613_, new_n1328_ );
xor  ( new_n2615_, new_n1458_, new_n1456_ );
not  ( new_n2616_, new_n2615_ );
nor  ( new_n2617_, new_n2616_, new_n1582_ );
and  ( new_n2618_, new_n2616_, new_n1582_ );
or   ( new_n2619_, new_n2618_, new_n1714_ );
or   ( new_n2620_, new_n2619_, new_n2617_ );
xor  ( new_n2621_, \c[8] , \a[8]  );
xnor ( new_n2622_, new_n2621_, new_n1763_ );
or   ( new_n2623_, new_n2622_, new_n2062_ );
xor  ( new_n2624_, \d[8] , \b[8]  );
xnor ( new_n2625_, new_n2624_, new_n1827_ );
or   ( new_n2626_, new_n2625_, new_n2061_ );
or   ( new_n2627_, new_n1849_, new_n179_ );
or   ( new_n2628_, new_n2065_, new_n1328_ );
or   ( new_n2629_, new_n2067_, new_n1010_ );
and  ( new_n2630_, new_n2629_, new_n2628_ );
and  ( new_n2631_, new_n2630_, new_n2627_ );
and  ( new_n2632_, new_n2631_, new_n2626_ );
and  ( new_n2633_, new_n2632_, new_n2623_ );
and  ( new_n2634_, new_n2633_, new_n2620_ );
xor  ( new_n2635_, new_n650_, new_n648_ );
not  ( new_n2636_, new_n2635_ );
nor  ( new_n2637_, new_n2636_, new_n773_ );
and  ( new_n2638_, new_n2636_, new_n773_ );
or   ( new_n2639_, new_n2638_, new_n938_ );
or   ( new_n2640_, new_n2639_, new_n2637_ );
xor  ( new_n2641_, \d[8] , \c[8]  );
nand ( new_n2642_, new_n2641_, new_n2089_ );
and  ( new_n2643_, new_n2642_, new_n2640_ );
and  ( new_n2644_, new_n2643_, new_n2634_ );
and  ( new_n2645_, new_n2644_, new_n2614_ );
and  ( new_n2646_, new_n2645_, new_n2611_ );
and  ( new_n2647_, new_n2150_, \a[7]  );
nor  ( new_n2648_, new_n2647_, new_n2146_ );
nor  ( new_n2649_, new_n2648_, new_n2107_ );
not  ( new_n2650_, new_n2649_ );
and  ( new_n2651_, new_n2084_, \c[7]  );
nor  ( new_n2652_, new_n2651_, new_n2353_ );
nor  ( new_n2653_, new_n2652_, new_n1023_ );
not  ( new_n2654_, new_n2653_ );
xor  ( new_n2655_, \d[7] , \c[7]  );
and  ( new_n2656_, new_n2655_, new_n2089_ );
not  ( new_n2657_, new_n2656_ );
not  ( new_n2658_, new_n771_ );
xor  ( new_n2659_, new_n676_, new_n653_ );
and  ( new_n2660_, new_n2659_, new_n2658_ );
not  ( new_n2661_, new_n2660_ );
nor  ( new_n2662_, new_n2659_, new_n2658_ );
nor  ( new_n2663_, new_n2662_, new_n938_ );
and  ( new_n2664_, new_n2663_, new_n2661_ );
not  ( new_n2665_, new_n2664_ );
xor  ( new_n2666_, new_n1484_, new_n1461_ );
xnor ( new_n2667_, new_n2666_, new_n1580_ );
and  ( new_n2668_, new_n2667_, new_n1713_ );
not  ( new_n2669_, new_n2668_ );
xor  ( new_n2670_, \c[7] , \a[7]  );
xnor ( new_n2671_, new_n2670_, new_n1761_ );
not  ( new_n2672_, new_n2671_ );
and  ( new_n2673_, new_n2672_, new_n1780_ );
not  ( new_n2674_, new_n2673_ );
xor  ( new_n2675_, \d[7] , \b[7]  );
xnor ( new_n2676_, new_n2675_, new_n1825_ );
not  ( new_n2677_, new_n2676_ );
and  ( new_n2678_, new_n2677_, new_n1844_ );
not  ( new_n2679_, new_n2678_ );
and  ( new_n2680_, new_n1848_, \d[7]  );
not  ( new_n2681_, new_n2680_ );
and  ( new_n2682_, new_n2064_, \b[7]  );
and  ( new_n2683_, new_n2066_, \c[7]  );
nor  ( new_n2684_, new_n2683_, new_n2682_ );
and  ( new_n2685_, new_n2684_, new_n2681_ );
and  ( new_n2686_, new_n2685_, new_n2679_ );
and  ( new_n2687_, new_n2686_, new_n2674_ );
and  ( new_n2688_, new_n2687_, new_n2669_ );
and  ( new_n2689_, new_n2688_, new_n2665_ );
and  ( new_n2690_, new_n2689_, new_n2657_ );
and  ( new_n2691_, new_n2690_, new_n2654_ );
and  ( new_n2692_, new_n2691_, new_n2650_ );
nor  ( new_n2693_, new_n2692_, new_n2646_ );
nor  ( new_n2694_, new_n2693_, new_n2542_ );
or   ( new_n2695_, new_n2694_, new_n2608_ );
and  ( new_n2696_, new_n2695_, new_n2607_ );
or   ( new_n2697_, new_n2696_, new_n2596_ );
and  ( new_n2698_, new_n2697_, new_n2595_ );
or   ( new_n2699_, new_n2698_, new_n2593_ );
and  ( new_n2700_, new_n2699_, new_n2592_ );
nor  ( new_n2701_, new_n2700_, new_n2589_ );
and  ( new_n2702_, new_n2700_, new_n2589_ );
xor  ( new_n2703_, new_n2591_, new_n2590_ );
xor  ( new_n2704_, new_n2703_, new_n2698_ );
xnor ( new_n2705_, new_n2458_, new_n2278_ );
or   ( new_n2706_, new_n2705_, new_n2134_ );
xor  ( new_n2707_, new_n2304_, new_n2299_ );
or   ( new_n2708_, new_n2707_, new_n2403_ );
or   ( new_n2709_, new_n2568_, new_n2446_ );
and  ( new_n2710_, new_n2709_, new_n2708_ );
or   ( new_n2711_, new_n2710_, new_n2706_ );
xor  ( new_n2712_, new_n2395_, new_n2288_ );
and  ( new_n2713_, new_n2712_, new_n2558_ );
and  ( new_n2714_, new_n2603_, new_n2601_ );
or   ( new_n2715_, new_n2714_, new_n2713_ );
xor  ( new_n2716_, new_n2710_, new_n2706_ );
nand ( new_n2717_, new_n2716_, new_n2715_ );
and  ( new_n2718_, new_n2717_, new_n2711_ );
xor  ( new_n2719_, new_n2594_, new_n2564_ );
xor  ( new_n2720_, new_n2719_, new_n2696_ );
or   ( new_n2721_, new_n2720_, new_n2718_ );
and  ( new_n2722_, new_n2720_, new_n2718_ );
xnor ( new_n2723_, new_n2519_, new_n2276_ );
or   ( new_n2724_, new_n2723_, new_n2134_ );
not  ( new_n2725_, new_n2693_ );
and  ( new_n2726_, new_n2725_, new_n2542_ );
and  ( new_n2727_, new_n2692_, new_n2646_ );
nor  ( new_n2728_, new_n2727_, new_n2542_ );
nor  ( new_n2729_, new_n2728_, new_n2726_ );
not  ( new_n2730_, new_n2729_ );
xor  ( new_n2731_, new_n2542_, new_n2407_ );
or   ( new_n2732_, new_n2731_, new_n2730_ );
not  ( new_n2733_, new_n2694_ );
or   ( new_n2734_, new_n2727_, new_n2733_ );
and  ( new_n2735_, new_n2734_, new_n2732_ );
nor  ( new_n2736_, new_n2735_, new_n2724_ );
xor  ( new_n2737_, new_n2705_, new_n2233_ );
nor  ( new_n2738_, new_n2737_, new_n2232_ );
nor  ( new_n2739_, new_n2597_, new_n2300_ );
or   ( new_n2740_, new_n2739_, new_n2738_ );
xor  ( new_n2741_, new_n2735_, new_n2724_ );
and  ( new_n2742_, new_n2741_, new_n2740_ );
or   ( new_n2743_, new_n2742_, new_n2736_ );
xor  ( new_n2744_, new_n2716_, new_n2715_ );
and  ( new_n2745_, new_n2744_, new_n2743_ );
xor  ( new_n2746_, new_n2744_, new_n2743_ );
xor  ( new_n2747_, new_n2606_, new_n2600_ );
xor  ( new_n2748_, new_n2747_, new_n2733_ );
and  ( new_n2749_, new_n2748_, new_n2746_ );
nor  ( new_n2750_, new_n2749_, new_n2745_ );
or   ( new_n2751_, new_n2750_, new_n2722_ );
and  ( new_n2752_, new_n2751_, new_n2721_ );
nor  ( new_n2753_, new_n2752_, new_n2704_ );
and  ( new_n2754_, new_n2752_, new_n2704_ );
xor  ( new_n2755_, new_n2440_, new_n2178_ );
nand ( new_n2756_, new_n2755_, new_n2402_ );
or   ( new_n2757_, new_n2707_, new_n2446_ );
and  ( new_n2758_, new_n2757_, new_n2756_ );
nor  ( new_n2759_, new_n2758_, new_n2715_ );
xnor ( new_n2760_, new_n2641_, new_n2274_ );
or   ( new_n2761_, new_n2760_, new_n2134_ );
xor  ( new_n2762_, new_n2723_, new_n2233_ );
or   ( new_n2763_, new_n2762_, new_n2232_ );
or   ( new_n2764_, new_n2737_, new_n2300_ );
and  ( new_n2765_, new_n2764_, new_n2763_ );
nor  ( new_n2766_, new_n2765_, new_n2761_ );
xor  ( new_n2767_, new_n2395_, new_n2304_ );
and  ( new_n2768_, new_n2767_, new_n2558_ );
and  ( new_n2769_, new_n2712_, new_n2603_ );
or   ( new_n2770_, new_n2769_, new_n2768_ );
xor  ( new_n2771_, new_n2765_, new_n2761_ );
and  ( new_n2772_, new_n2771_, new_n2770_ );
nor  ( new_n2773_, new_n2772_, new_n2766_ );
and  ( new_n2774_, new_n2758_, new_n2715_ );
nor  ( new_n2775_, new_n2774_, new_n2773_ );
or   ( new_n2776_, new_n2775_, new_n2759_ );
xor  ( new_n2777_, new_n2748_, new_n2746_ );
and  ( new_n2778_, new_n2777_, new_n2776_ );
xor  ( new_n2779_, new_n2542_, new_n2297_ );
nand ( new_n2780_, new_n2779_, new_n2729_ );
xor  ( new_n2781_, new_n2692_, new_n2646_ );
not  ( new_n2782_, new_n2781_ );
or   ( new_n2783_, new_n2782_, new_n2731_ );
and  ( new_n2784_, new_n2783_, new_n2780_ );
or   ( new_n2785_, new_n2077_, new_n212_ );
and  ( new_n2786_, new_n2785_, new_n2050_ );
or   ( new_n2787_, new_n2786_, new_n2108_ );
or   ( new_n2788_, new_n2058_, new_n1373_ );
and  ( new_n2789_, new_n2788_, new_n2056_ );
or   ( new_n2790_, new_n2789_, new_n1019_ );
xor  ( new_n2791_, \d[6] , \c[6]  );
nand ( new_n2792_, new_n2791_, new_n2089_ );
xnor ( new_n2793_, new_n1578_, new_n1508_ );
or   ( new_n2794_, new_n2793_, new_n1714_ );
xnor ( new_n2795_, new_n769_, new_n700_ );
or   ( new_n2796_, new_n2795_, new_n938_ );
xor  ( new_n2797_, \c[6] , \a[6]  );
xnor ( new_n2798_, new_n2797_, new_n1759_ );
or   ( new_n2799_, new_n2798_, new_n2062_ );
xor  ( new_n2800_, \d[6] , \b[6]  );
xnor ( new_n2801_, new_n2800_, new_n1823_ );
or   ( new_n2802_, new_n2801_, new_n2061_ );
or   ( new_n2803_, new_n1849_, new_n563_ );
or   ( new_n2804_, new_n2065_, new_n1019_ );
or   ( new_n2805_, new_n2067_, new_n1373_ );
and  ( new_n2806_, new_n2805_, new_n2804_ );
and  ( new_n2807_, new_n2806_, new_n2803_ );
and  ( new_n2808_, new_n2807_, new_n2802_ );
and  ( new_n2809_, new_n2808_, new_n2799_ );
and  ( new_n2810_, new_n2809_, new_n2796_ );
and  ( new_n2811_, new_n2810_, new_n2794_ );
and  ( new_n2812_, new_n2811_, new_n2792_ );
and  ( new_n2813_, new_n2812_, new_n2790_ );
and  ( new_n2814_, new_n2813_, new_n2787_ );
and  ( new_n2815_, new_n2150_, \a[5]  );
nor  ( new_n2816_, new_n2815_, new_n2146_ );
nor  ( new_n2817_, new_n2816_, new_n2104_ );
not  ( new_n2818_, new_n2817_ );
and  ( new_n2819_, new_n2084_, \c[5]  );
nor  ( new_n2820_, new_n2819_, new_n2353_ );
nor  ( new_n2821_, new_n2820_, new_n847_ );
not  ( new_n2822_, new_n2821_ );
xor  ( new_n2823_, \d[5] , \c[5]  );
and  ( new_n2824_, new_n2823_, new_n2089_ );
not  ( new_n2825_, new_n2824_ );
xor  ( new_n2826_, new_n1524_, new_n1509_ );
xor  ( new_n2827_, new_n2826_, new_n1576_ );
nor  ( new_n2828_, new_n2827_, new_n1714_ );
not  ( new_n2829_, new_n2828_ );
xor  ( new_n2830_, new_n716_, new_n701_ );
xnor ( new_n2831_, new_n2830_, new_n767_ );
and  ( new_n2832_, new_n2831_, new_n937_ );
not  ( new_n2833_, new_n2832_ );
xor  ( new_n2834_, \d[5] , \b[5]  );
xnor ( new_n2835_, new_n2834_, new_n1821_ );
not  ( new_n2836_, new_n2835_ );
and  ( new_n2837_, new_n2836_, new_n1844_ );
not  ( new_n2838_, new_n2837_ );
xor  ( new_n2839_, \c[5] , \a[5]  );
xnor ( new_n2840_, new_n2839_, new_n1757_ );
not  ( new_n2841_, new_n2840_ );
and  ( new_n2842_, new_n2841_, new_n1780_ );
not  ( new_n2843_, new_n2842_ );
and  ( new_n2844_, new_n1848_, \d[5]  );
not  ( new_n2845_, new_n2844_ );
and  ( new_n2846_, new_n2066_, \c[5]  );
and  ( new_n2847_, new_n2064_, \b[5]  );
nor  ( new_n2848_, new_n2847_, new_n2846_ );
and  ( new_n2849_, new_n2848_, new_n2845_ );
and  ( new_n2850_, new_n2849_, new_n2843_ );
and  ( new_n2851_, new_n2850_, new_n2838_ );
and  ( new_n2852_, new_n2851_, new_n2833_ );
and  ( new_n2853_, new_n2852_, new_n2829_ );
and  ( new_n2854_, new_n2853_, new_n2825_ );
and  ( new_n2855_, new_n2854_, new_n2822_ );
and  ( new_n2856_, new_n2855_, new_n2818_ );
nor  ( new_n2857_, new_n2856_, new_n2814_ );
nor  ( new_n2858_, new_n2857_, new_n2692_ );
nor  ( new_n2859_, new_n2858_, new_n2784_ );
xor  ( new_n2860_, new_n2566_, new_n2178_ );
and  ( new_n2861_, new_n2860_, new_n2402_ );
and  ( new_n2862_, new_n2755_, new_n2445_ );
nor  ( new_n2863_, new_n2862_, new_n2861_ );
xnor ( new_n2864_, new_n2858_, new_n2784_ );
nor  ( new_n2865_, new_n2864_, new_n2863_ );
nor  ( new_n2866_, new_n2865_, new_n2859_ );
not  ( new_n2867_, new_n2866_ );
xor  ( new_n2868_, new_n2741_, new_n2740_ );
and  ( new_n2869_, new_n2868_, new_n2867_ );
xor  ( new_n2870_, new_n2868_, new_n2867_ );
not  ( new_n2871_, new_n2870_ );
xor  ( new_n2872_, new_n2758_, new_n2715_ );
xor  ( new_n2873_, new_n2872_, new_n2773_ );
nor  ( new_n2874_, new_n2873_, new_n2871_ );
or   ( new_n2875_, new_n2874_, new_n2869_ );
xor  ( new_n2876_, new_n2777_, new_n2776_ );
and  ( new_n2877_, new_n2876_, new_n2875_ );
or   ( new_n2878_, new_n2877_, new_n2778_ );
xnor ( new_n2879_, new_n2720_, new_n2718_ );
xor  ( new_n2880_, new_n2879_, new_n2750_ );
nor  ( new_n2881_, new_n2880_, new_n2878_ );
and  ( new_n2882_, new_n2880_, new_n2878_ );
xor  ( new_n2883_, new_n2873_, new_n2871_ );
xor  ( new_n2884_, new_n2542_, new_n2288_ );
and  ( new_n2885_, new_n2884_, new_n2729_ );
and  ( new_n2886_, new_n2781_, new_n2779_ );
or   ( new_n2887_, new_n2886_, new_n2885_ );
xor  ( new_n2888_, new_n2771_, new_n2770_ );
nand ( new_n2889_, new_n2888_, new_n2887_ );
nor  ( new_n2890_, new_n2888_, new_n2887_ );
xor  ( new_n2891_, new_n2705_, new_n2178_ );
nand ( new_n2892_, new_n2891_, new_n2402_ );
nand ( new_n2893_, new_n2860_, new_n2445_ );
and  ( new_n2894_, new_n2893_, new_n2892_ );
xor  ( new_n2895_, new_n2760_, new_n2233_ );
or   ( new_n2896_, new_n2895_, new_n2232_ );
or   ( new_n2897_, new_n2762_, new_n2300_ );
and  ( new_n2898_, new_n2897_, new_n2896_ );
or   ( new_n2899_, new_n2898_, new_n2894_ );
and  ( new_n2900_, new_n2898_, new_n2894_ );
not  ( new_n2901_, new_n2692_ );
nor  ( new_n2902_, new_n2857_, new_n2901_ );
and  ( new_n2903_, new_n2856_, new_n2814_ );
nor  ( new_n2904_, new_n2903_, new_n2692_ );
nor  ( new_n2905_, new_n2904_, new_n2902_ );
not  ( new_n2906_, new_n2407_ );
xor  ( new_n2907_, new_n2692_, new_n2906_ );
and  ( new_n2908_, new_n2907_, new_n2905_ );
not  ( new_n2909_, new_n2903_ );
and  ( new_n2910_, new_n2909_, new_n2858_ );
nor  ( new_n2911_, new_n2910_, new_n2908_ );
or   ( new_n2912_, new_n2911_, new_n2900_ );
and  ( new_n2913_, new_n2912_, new_n2899_ );
or   ( new_n2914_, new_n2913_, new_n2890_ );
nand ( new_n2915_, new_n2914_, new_n2889_ );
and  ( new_n2916_, new_n2915_, new_n2883_ );
xnor ( new_n2917_, new_n2915_, new_n2883_ );
xnor ( new_n2918_, new_n2864_, new_n2863_ );
xor  ( new_n2919_, new_n2440_, new_n2395_ );
and  ( new_n2920_, new_n2919_, new_n2558_ );
and  ( new_n2921_, new_n2767_, new_n2603_ );
or   ( new_n2922_, new_n2921_, new_n2920_ );
xnor ( new_n2923_, new_n2655_, new_n2272_ );
not  ( new_n2924_, new_n2923_ );
and  ( new_n2925_, new_n2924_, new_n2233_ );
nand ( new_n2926_, new_n2925_, new_n2922_ );
nor  ( new_n2927_, new_n2925_, new_n2922_ );
or   ( new_n2928_, new_n2927_, new_n2887_ );
and  ( new_n2929_, new_n2928_, new_n2926_ );
or   ( new_n2930_, new_n2929_, new_n2918_ );
and  ( new_n2931_, new_n2929_, new_n2918_ );
xor  ( new_n2932_, new_n2888_, new_n2887_ );
xor  ( new_n2933_, new_n2932_, new_n2913_ );
or   ( new_n2934_, new_n2933_, new_n2931_ );
and  ( new_n2935_, new_n2934_, new_n2930_ );
nor  ( new_n2936_, new_n2935_, new_n2917_ );
or   ( new_n2937_, new_n2936_, new_n2916_ );
xor  ( new_n2938_, new_n2876_, new_n2875_ );
nor  ( new_n2939_, new_n2938_, new_n2937_ );
and  ( new_n2940_, new_n2938_, new_n2937_ );
xor  ( new_n2941_, new_n2898_, new_n2894_ );
xnor ( new_n2942_, new_n2941_, new_n2911_ );
xor  ( new_n2943_, new_n2566_, new_n2554_ );
or   ( new_n2944_, new_n2943_, new_n2559_ );
nand ( new_n2945_, new_n2919_, new_n2603_ );
and  ( new_n2946_, new_n2945_, new_n2944_ );
or   ( new_n2947_, new_n2077_, new_n231_ );
and  ( new_n2948_, new_n2947_, new_n2050_ );
or   ( new_n2949_, new_n2948_, new_n2105_ );
or   ( new_n2950_, new_n2058_, new_n1468_ );
and  ( new_n2951_, new_n2950_, new_n2056_ );
or   ( new_n2952_, new_n2951_, new_n832_ );
xor  ( new_n2953_, \d[4] , \c[4]  );
nand ( new_n2954_, new_n2953_, new_n2089_ );
xor  ( new_n2955_, new_n1542_, new_n1540_ );
xor  ( new_n2956_, new_n2955_, new_n1574_ );
or   ( new_n2957_, new_n2956_, new_n1714_ );
xor  ( new_n2958_, new_n734_, new_n732_ );
xor  ( new_n2959_, new_n2958_, new_n765_ );
or   ( new_n2960_, new_n2959_, new_n938_ );
xor  ( new_n2961_, \d[4] , \b[4]  );
xnor ( new_n2962_, new_n2961_, new_n1819_ );
or   ( new_n2963_, new_n2962_, new_n2061_ );
xor  ( new_n2964_, \c[4] , \a[4]  );
xnor ( new_n2965_, new_n2964_, new_n1755_ );
or   ( new_n2966_, new_n2965_, new_n2062_ );
or   ( new_n2967_, new_n1849_, new_n660_ );
or   ( new_n2968_, new_n2065_, new_n832_ );
or   ( new_n2969_, new_n2067_, new_n1468_ );
and  ( new_n2970_, new_n2969_, new_n2968_ );
and  ( new_n2971_, new_n2970_, new_n2967_ );
and  ( new_n2972_, new_n2971_, new_n2966_ );
and  ( new_n2973_, new_n2972_, new_n2963_ );
and  ( new_n2974_, new_n2973_, new_n2960_ );
and  ( new_n2975_, new_n2974_, new_n2957_ );
and  ( new_n2976_, new_n2975_, new_n2954_ );
and  ( new_n2977_, new_n2976_, new_n2952_ );
and  ( new_n2978_, new_n2977_, new_n2949_ );
not  ( new_n2979_, new_n2092_ );
and  ( new_n2980_, new_n2146_, new_n2979_ );
not  ( new_n2981_, new_n2980_ );
and  ( new_n2982_, new_n2075_, \a[3]  );
not  ( new_n2983_, new_n2982_ );
and  ( new_n2984_, \c[3] , \b[3]  );
and  ( new_n2985_, new_n2084_, new_n2984_ );
not  ( new_n2986_, new_n2985_ );
and  ( new_n2987_, new_n815_, new_n163_ );
not  ( new_n2988_, new_n2987_ );
and  ( new_n2989_, new_n2353_, new_n2988_ );
not  ( new_n2990_, new_n2989_ );
xor  ( new_n2991_, \d[3] , \c[3]  );
and  ( new_n2992_, new_n2991_, new_n2089_ );
not  ( new_n2993_, new_n2992_ );
xor  ( new_n2994_, new_n1553_, new_n1545_ );
xnor ( new_n2995_, new_n2994_, new_n1572_ );
and  ( new_n2996_, new_n2995_, new_n1713_ );
not  ( new_n2997_, new_n2996_ );
xor  ( new_n2998_, new_n745_, new_n737_ );
xnor ( new_n2999_, new_n2998_, new_n763_ );
and  ( new_n3000_, new_n2999_, new_n937_ );
not  ( new_n3001_, new_n3000_ );
xor  ( new_n3002_, \d[3] , \b[3]  );
xnor ( new_n3003_, new_n3002_, new_n1817_ );
not  ( new_n3004_, new_n3003_ );
and  ( new_n3005_, new_n3004_, new_n1844_ );
not  ( new_n3006_, new_n3005_ );
xor  ( new_n3007_, \c[3] , \a[3]  );
xnor ( new_n3008_, new_n3007_, new_n1753_ );
not  ( new_n3009_, new_n3008_ );
and  ( new_n3010_, new_n3009_, new_n1780_ );
not  ( new_n3011_, new_n3010_ );
and  ( new_n3012_, new_n1848_, \d[3]  );
not  ( new_n3013_, new_n3012_ );
and  ( new_n3014_, new_n2064_, \b[3]  );
and  ( new_n3015_, new_n2066_, \c[3]  );
nor  ( new_n3016_, new_n3015_, new_n3014_ );
and  ( new_n3017_, new_n3016_, new_n3013_ );
and  ( new_n3018_, new_n3017_, new_n3011_ );
and  ( new_n3019_, new_n3018_, new_n3006_ );
and  ( new_n3020_, new_n3019_, new_n3001_ );
and  ( new_n3021_, new_n3020_, new_n2997_ );
and  ( new_n3022_, new_n3021_, new_n2993_ );
and  ( new_n3023_, new_n3022_, new_n2990_ );
and  ( new_n3024_, new_n3023_, new_n2986_ );
and  ( new_n3025_, new_n3024_, new_n2983_ );
and  ( new_n3026_, new_n3025_, new_n2981_ );
nor  ( new_n3027_, new_n3026_, new_n2978_ );
nor  ( new_n3028_, new_n3027_, new_n2856_ );
or   ( new_n3029_, new_n3028_, new_n2946_ );
and  ( new_n3030_, new_n3028_, new_n2946_ );
xor  ( new_n3031_, new_n2692_, new_n2297_ );
and  ( new_n3032_, new_n3031_, new_n2905_ );
xor  ( new_n3033_, new_n2856_, new_n2814_ );
and  ( new_n3034_, new_n3033_, new_n2907_ );
nor  ( new_n3035_, new_n3034_, new_n3032_ );
or   ( new_n3036_, new_n3035_, new_n3030_ );
nand ( new_n3037_, new_n3036_, new_n3029_ );
and  ( new_n3038_, new_n3037_, new_n2942_ );
xnor ( new_n3039_, new_n3037_, new_n2942_ );
xor  ( new_n3040_, new_n2723_, new_n2178_ );
and  ( new_n3041_, new_n3040_, new_n2402_ );
and  ( new_n3042_, new_n2891_, new_n2445_ );
nor  ( new_n3043_, new_n3042_, new_n3041_ );
not  ( new_n3044_, new_n3043_ );
xor  ( new_n3045_, new_n2542_, new_n2304_ );
and  ( new_n3046_, new_n3045_, new_n2729_ );
and  ( new_n3047_, new_n2884_, new_n2781_ );
nor  ( new_n3048_, new_n3047_, new_n3046_ );
not  ( new_n3049_, new_n3048_ );
and  ( new_n3050_, new_n3049_, new_n3044_ );
xor  ( new_n3051_, new_n2923_, new_n2233_ );
nor  ( new_n3052_, new_n3051_, new_n2232_ );
nor  ( new_n3053_, new_n2895_, new_n2300_ );
nor  ( new_n3054_, new_n3053_, new_n3052_ );
and  ( new_n3055_, new_n3048_, new_n3043_ );
nor  ( new_n3056_, new_n3055_, new_n3054_ );
nor  ( new_n3057_, new_n3056_, new_n3050_ );
nor  ( new_n3058_, new_n3057_, new_n3039_ );
nor  ( new_n3059_, new_n3058_, new_n3038_ );
xor  ( new_n3060_, new_n2929_, new_n2918_ );
xor  ( new_n3061_, new_n3060_, new_n2933_ );
nor  ( new_n3062_, new_n3061_, new_n3059_ );
xor  ( new_n3063_, new_n3061_, new_n3059_ );
xor  ( new_n3064_, new_n2925_, new_n2922_ );
xnor ( new_n3065_, new_n3064_, new_n2887_ );
xnor ( new_n3066_, new_n2791_, new_n2270_ );
or   ( new_n3067_, new_n3066_, new_n2134_ );
xor  ( new_n3068_, new_n3026_, new_n2978_ );
xnor ( new_n3069_, new_n2978_, new_n2856_ );
nor  ( new_n3070_, new_n3069_, new_n3068_ );
xor  ( new_n3071_, new_n2856_, new_n2906_ );
and  ( new_n3072_, new_n3071_, new_n3070_ );
and  ( new_n3073_, new_n3026_, new_n2978_ );
not  ( new_n3074_, new_n3073_ );
and  ( new_n3075_, new_n3074_, new_n3028_ );
nor  ( new_n3076_, new_n3075_, new_n3072_ );
nand ( new_n3077_, new_n3076_, new_n3067_ );
or   ( new_n3078_, new_n3076_, new_n3067_ );
xor  ( new_n3079_, new_n2760_, new_n2299_ );
or   ( new_n3080_, new_n3079_, new_n2403_ );
nand ( new_n3081_, new_n3040_, new_n2445_ );
and  ( new_n3082_, new_n3081_, new_n3080_ );
xor  ( new_n3083_, new_n2705_, new_n2554_ );
or   ( new_n3084_, new_n3083_, new_n2559_ );
or   ( new_n3085_, new_n2943_, new_n2604_ );
and  ( new_n3086_, new_n3085_, new_n3084_ );
nor  ( new_n3087_, new_n3086_, new_n3082_ );
xor  ( new_n3088_, new_n2692_, new_n2288_ );
and  ( new_n3089_, new_n3088_, new_n2905_ );
and  ( new_n3090_, new_n3033_, new_n3031_ );
nor  ( new_n3091_, new_n3090_, new_n3089_ );
and  ( new_n3092_, new_n3086_, new_n3082_ );
nor  ( new_n3093_, new_n3092_, new_n3091_ );
nor  ( new_n3094_, new_n3093_, new_n3087_ );
nand ( new_n3095_, new_n3094_, new_n3078_ );
and  ( new_n3096_, new_n3095_, new_n3077_ );
nand ( new_n3097_, new_n3096_, new_n3065_ );
nor  ( new_n3098_, new_n3096_, new_n3065_ );
xor  ( new_n3099_, new_n3048_, new_n3044_ );
and  ( new_n3100_, new_n3099_, new_n3054_ );
not  ( new_n3101_, new_n3050_ );
and  ( new_n3102_, new_n3056_, new_n3101_ );
or   ( new_n3103_, new_n3102_, new_n3100_ );
xor  ( new_n3104_, new_n3066_, new_n2233_ );
nor  ( new_n3105_, new_n3104_, new_n2232_ );
nor  ( new_n3106_, new_n3051_, new_n2300_ );
or   ( new_n3107_, new_n3106_, new_n3105_ );
xnor ( new_n3108_, new_n2823_, new_n2268_ );
not  ( new_n3109_, new_n3108_ );
and  ( new_n3110_, new_n3109_, new_n2233_ );
nand ( new_n3111_, new_n3110_, new_n3107_ );
nor  ( new_n3112_, new_n3110_, new_n3107_ );
xor  ( new_n3113_, new_n2542_, new_n2441_ );
or   ( new_n3114_, new_n3113_, new_n2730_ );
nand ( new_n3115_, new_n3045_, new_n2781_ );
and  ( new_n3116_, new_n3115_, new_n3114_ );
or   ( new_n3117_, new_n3116_, new_n3112_ );
and  ( new_n3118_, new_n3117_, new_n3111_ );
nor  ( new_n3119_, new_n3118_, new_n3103_ );
and  ( new_n3120_, new_n3118_, new_n3103_ );
xor  ( new_n3121_, new_n3028_, new_n2946_ );
xnor ( new_n3122_, new_n3121_, new_n3035_ );
not  ( new_n3123_, new_n3122_ );
nor  ( new_n3124_, new_n3123_, new_n3120_ );
nor  ( new_n3125_, new_n3124_, new_n3119_ );
or   ( new_n3126_, new_n3125_, new_n3098_ );
nand ( new_n3127_, new_n3126_, new_n3097_ );
and  ( new_n3128_, new_n3127_, new_n3063_ );
or   ( new_n3129_, new_n3128_, new_n3062_ );
xor  ( new_n3130_, new_n2935_, new_n2917_ );
and  ( new_n3131_, new_n3130_, new_n3129_ );
nor  ( new_n3132_, new_n3130_, new_n3129_ );
xnor ( new_n3133_, new_n3127_, new_n3063_ );
xor  ( new_n3134_, new_n3057_, new_n3039_ );
xnor ( new_n3135_, new_n3096_, new_n3065_ );
xor  ( new_n3136_, new_n3135_, new_n3125_ );
nand ( new_n3137_, new_n3136_, new_n3134_ );
nor  ( new_n3138_, new_n3136_, new_n3134_ );
xor  ( new_n3139_, new_n3076_, new_n3067_ );
xor  ( new_n3140_, new_n3139_, new_n3094_ );
not  ( new_n3141_, new_n3076_ );
not  ( new_n3142_, new_n3070_ );
not  ( new_n3143_, new_n2297_ );
xor  ( new_n3144_, new_n2856_, new_n3143_ );
or   ( new_n3145_, new_n3144_, new_n3142_ );
nand ( new_n3146_, new_n3071_, new_n3068_ );
and  ( new_n3147_, new_n3146_, new_n3145_ );
or   ( new_n3148_, new_n2093_, new_n2050_ );
or   ( new_n3149_, new_n2076_, new_n115_ );
and  ( new_n3150_, \c[2] , \b[2]  );
nand ( new_n3151_, new_n3150_, new_n2084_ );
and  ( new_n3152_, new_n865_, new_n115_ );
or   ( new_n3153_, new_n3152_, new_n2056_ );
xor  ( new_n3154_, \d[2] , \c[2]  );
nand ( new_n3155_, new_n3154_, new_n2089_ );
xor  ( new_n3156_, new_n1563_, new_n1557_ );
xor  ( new_n3157_, new_n3156_, new_n1570_ );
or   ( new_n3158_, new_n3157_, new_n1714_ );
xor  ( new_n3159_, new_n754_, new_n748_ );
xor  ( new_n3160_, new_n3159_, new_n761_ );
or   ( new_n3161_, new_n3160_, new_n938_ );
xor  ( new_n3162_, \d[2] , \b[2]  );
xnor ( new_n3163_, new_n3162_, new_n1815_ );
or   ( new_n3164_, new_n3163_, new_n2061_ );
xor  ( new_n3165_, \c[2] , \a[2]  );
xnor ( new_n3166_, new_n3165_, new_n1751_ );
or   ( new_n3167_, new_n3166_, new_n2062_ );
or   ( new_n3168_, new_n1849_, new_n726_ );
or   ( new_n3169_, new_n2065_, new_n865_ );
or   ( new_n3170_, new_n2067_, new_n1534_ );
and  ( new_n3171_, new_n3170_, new_n3169_ );
and  ( new_n3172_, new_n3171_, new_n3168_ );
and  ( new_n3173_, new_n3172_, new_n3167_ );
and  ( new_n3174_, new_n3173_, new_n3164_ );
and  ( new_n3175_, new_n3174_, new_n3161_ );
and  ( new_n3176_, new_n3175_, new_n3158_ );
and  ( new_n3177_, new_n3176_, new_n3155_ );
and  ( new_n3178_, new_n3177_, new_n3153_ );
and  ( new_n3179_, new_n3178_, new_n3151_ );
and  ( new_n3180_, new_n3179_, new_n3149_ );
and  ( new_n3181_, new_n3180_, new_n3148_ );
and  ( new_n3182_, new_n90_, new_n108_ );
not  ( new_n3183_, new_n3182_ );
and  ( new_n3184_, new_n3183_, new_n2146_ );
not  ( new_n3185_, new_n3184_ );
and  ( new_n3186_, new_n2075_, \a[1]  );
not  ( new_n3187_, new_n3186_ );
and  ( new_n3188_, \c[1] , \b[1]  );
and  ( new_n3189_, new_n3188_, new_n2084_ );
not  ( new_n3190_, new_n3189_ );
and  ( new_n3191_, new_n808_, new_n108_ );
not  ( new_n3192_, new_n3191_ );
and  ( new_n3193_, new_n3192_, new_n2353_ );
not  ( new_n3194_, new_n3193_ );
xor  ( new_n3195_, \d[1] , \c[1]  );
and  ( new_n3196_, new_n3195_, new_n2089_ );
not  ( new_n3197_, new_n3196_ );
and  ( new_n3198_, \c[1] , \b[0]  );
xor  ( new_n3199_, new_n3198_, new_n1566_ );
and  ( new_n3200_, new_n3199_, new_n1713_ );
not  ( new_n3201_, new_n3200_ );
and  ( new_n3202_, \d[1] , \a[0]  );
xor  ( new_n3203_, new_n3202_, new_n757_ );
and  ( new_n3204_, new_n3203_, new_n937_ );
not  ( new_n3205_, new_n3204_ );
xor  ( new_n3206_, \d[1] , \b[1]  );
xnor ( new_n3207_, new_n3206_, new_n1813_ );
not  ( new_n3208_, new_n3207_ );
and  ( new_n3209_, new_n3208_, new_n1844_ );
not  ( new_n3210_, new_n3209_ );
xor  ( new_n3211_, \c[1] , \a[1]  );
xnor ( new_n3212_, new_n3211_, new_n1749_ );
not  ( new_n3213_, new_n3212_ );
and  ( new_n3214_, new_n3213_, new_n1780_ );
not  ( new_n3215_, new_n3214_ );
and  ( new_n3216_, new_n1848_, \d[1]  );
not  ( new_n3217_, new_n3216_ );
and  ( new_n3218_, new_n2064_, \b[1]  );
and  ( new_n3219_, new_n2066_, \c[1]  );
nor  ( new_n3220_, new_n3219_, new_n3218_ );
and  ( new_n3221_, new_n3220_, new_n3217_ );
and  ( new_n3222_, new_n3221_, new_n3215_ );
and  ( new_n3223_, new_n3222_, new_n3210_ );
and  ( new_n3224_, new_n3223_, new_n3205_ );
and  ( new_n3225_, new_n3224_, new_n3201_ );
and  ( new_n3226_, new_n3225_, new_n3197_ );
and  ( new_n3227_, new_n3226_, new_n3194_ );
and  ( new_n3228_, new_n3227_, new_n3190_ );
and  ( new_n3229_, new_n3228_, new_n3187_ );
and  ( new_n3230_, new_n3229_, new_n3185_ );
nor  ( new_n3231_, new_n3230_, new_n3181_ );
nor  ( new_n3232_, new_n3231_, new_n3026_ );
or   ( new_n3233_, new_n3232_, new_n3147_ );
and  ( new_n3234_, new_n3232_, new_n3147_ );
not  ( new_n3235_, new_n2542_ );
xor  ( new_n3236_, new_n2566_, new_n3235_ );
or   ( new_n3237_, new_n3236_, new_n2730_ );
or   ( new_n3238_, new_n3113_, new_n2782_ );
and  ( new_n3239_, new_n3238_, new_n3237_ );
or   ( new_n3240_, new_n3239_, new_n3234_ );
and  ( new_n3241_, new_n3240_, new_n3233_ );
or   ( new_n3242_, new_n3241_, new_n3141_ );
and  ( new_n3243_, new_n3241_, new_n3141_ );
xnor ( new_n3244_, new_n2953_, new_n2266_ );
or   ( new_n3245_, new_n3244_, new_n2134_ );
xor  ( new_n3246_, new_n2723_, new_n2554_ );
or   ( new_n3247_, new_n3246_, new_n2559_ );
or   ( new_n3248_, new_n3083_, new_n2604_ );
and  ( new_n3249_, new_n3248_, new_n3247_ );
nor  ( new_n3250_, new_n3249_, new_n3245_ );
and  ( new_n3251_, new_n3249_, new_n3245_ );
xor  ( new_n3252_, new_n2692_, new_n2304_ );
and  ( new_n3253_, new_n3252_, new_n2905_ );
and  ( new_n3254_, new_n3088_, new_n3033_ );
nor  ( new_n3255_, new_n3254_, new_n3253_ );
nor  ( new_n3256_, new_n3255_, new_n3251_ );
nor  ( new_n3257_, new_n3256_, new_n3250_ );
or   ( new_n3258_, new_n3257_, new_n3243_ );
and  ( new_n3259_, new_n3258_, new_n3242_ );
nor  ( new_n3260_, new_n3259_, new_n3140_ );
and  ( new_n3261_, new_n3259_, new_n3140_ );
xor  ( new_n3262_, new_n3110_, new_n3107_ );
xor  ( new_n3263_, new_n3262_, new_n3116_ );
xor  ( new_n3264_, new_n2923_, new_n2299_ );
or   ( new_n3265_, new_n3264_, new_n2403_ );
or   ( new_n3266_, new_n3079_, new_n2446_ );
and  ( new_n3267_, new_n3266_, new_n3265_ );
not  ( new_n3268_, new_n3231_ );
and  ( new_n3269_, new_n3268_, new_n3026_ );
and  ( new_n3270_, new_n3230_, new_n3181_ );
nor  ( new_n3271_, new_n3270_, new_n3026_ );
nor  ( new_n3272_, new_n3271_, new_n3269_ );
xor  ( new_n3273_, new_n3026_, new_n2906_ );
and  ( new_n3274_, new_n3273_, new_n3272_ );
not  ( new_n3275_, new_n3270_ );
and  ( new_n3276_, new_n3275_, new_n3232_ );
nor  ( new_n3277_, new_n3276_, new_n3274_ );
or   ( new_n3278_, new_n3277_, new_n3267_ );
xor  ( new_n3279_, new_n3108_, new_n2233_ );
nor  ( new_n3280_, new_n3279_, new_n2232_ );
nor  ( new_n3281_, new_n3104_, new_n2300_ );
nor  ( new_n3282_, new_n3281_, new_n3280_ );
and  ( new_n3283_, new_n3277_, new_n3267_ );
or   ( new_n3284_, new_n3283_, new_n3282_ );
and  ( new_n3285_, new_n3284_, new_n3278_ );
and  ( new_n3286_, new_n3285_, new_n3263_ );
xor  ( new_n3287_, new_n3086_, new_n3082_ );
xnor ( new_n3288_, new_n3287_, new_n3091_ );
nor  ( new_n3289_, new_n3285_, new_n3263_ );
nor  ( new_n3290_, new_n3289_, new_n3288_ );
nor  ( new_n3291_, new_n3290_, new_n3286_ );
not  ( new_n3292_, new_n3291_ );
nor  ( new_n3293_, new_n3292_, new_n3261_ );
nor  ( new_n3294_, new_n3293_, new_n3260_ );
or   ( new_n3295_, new_n3294_, new_n3138_ );
and  ( new_n3296_, new_n3295_, new_n3137_ );
nor  ( new_n3297_, new_n3296_, new_n3133_ );
and  ( new_n3298_, new_n3296_, new_n3133_ );
xor  ( new_n3299_, new_n3259_, new_n3140_ );
xor  ( new_n3300_, new_n3299_, new_n3292_ );
xor  ( new_n3301_, new_n3118_, new_n3103_ );
xor  ( new_n3302_, new_n3301_, new_n3123_ );
nand ( new_n3303_, new_n3302_, new_n3300_ );
xor  ( new_n3304_, new_n3232_, new_n3147_ );
xor  ( new_n3305_, new_n3304_, new_n3239_ );
xnor ( new_n3306_, new_n2991_, new_n2264_ );
or   ( new_n3307_, new_n3306_, new_n2134_ );
xor  ( new_n3308_, new_n2856_, new_n2288_ );
nand ( new_n3309_, new_n3308_, new_n3070_ );
not  ( new_n3310_, new_n3068_ );
or   ( new_n3311_, new_n3144_, new_n3310_ );
and  ( new_n3312_, new_n3311_, new_n3309_ );
or   ( new_n3313_, new_n3312_, new_n3307_ );
and  ( new_n3314_, new_n3312_, new_n3307_ );
xor  ( new_n3315_, new_n2705_, new_n2542_ );
nand ( new_n3316_, new_n3315_, new_n2729_ );
or   ( new_n3317_, new_n3236_, new_n2782_ );
and  ( new_n3318_, new_n3317_, new_n3316_ );
or   ( new_n3319_, new_n3318_, new_n3314_ );
and  ( new_n3320_, new_n3319_, new_n3313_ );
nor  ( new_n3321_, new_n3320_, new_n3305_ );
and  ( new_n3322_, new_n3320_, new_n3305_ );
xor  ( new_n3323_, new_n2760_, new_n2395_ );
nand ( new_n3324_, new_n3323_, new_n2558_ );
or   ( new_n3325_, new_n3246_, new_n2604_ );
and  ( new_n3326_, new_n3325_, new_n3324_ );
xor  ( new_n3327_, new_n3066_, new_n2299_ );
or   ( new_n3328_, new_n3327_, new_n2403_ );
or   ( new_n3329_, new_n3264_, new_n2446_ );
and  ( new_n3330_, new_n3329_, new_n3328_ );
nor  ( new_n3331_, new_n3330_, new_n3326_ );
xor  ( new_n3332_, new_n2692_, new_n2440_ );
and  ( new_n3333_, new_n3332_, new_n2905_ );
and  ( new_n3334_, new_n3252_, new_n3033_ );
nor  ( new_n3335_, new_n3334_, new_n3333_ );
and  ( new_n3336_, new_n3330_, new_n3326_ );
nor  ( new_n3337_, new_n3336_, new_n3335_ );
nor  ( new_n3338_, new_n3337_, new_n3331_ );
nor  ( new_n3339_, new_n3338_, new_n3322_ );
nor  ( new_n3340_, new_n3339_, new_n3321_ );
not  ( new_n3341_, new_n3340_ );
xor  ( new_n3342_, new_n3241_, new_n3076_ );
xor  ( new_n3343_, new_n3342_, new_n3257_ );
nor  ( new_n3344_, new_n3343_, new_n3341_ );
xor  ( new_n3345_, new_n3343_, new_n3341_ );
xor  ( new_n3346_, new_n3285_, new_n3263_ );
xnor ( new_n3347_, new_n3346_, new_n3288_ );
and  ( new_n3348_, new_n3347_, new_n3345_ );
or   ( new_n3349_, new_n3348_, new_n3344_ );
xor  ( new_n3350_, new_n3302_, new_n3300_ );
nand ( new_n3351_, new_n3350_, new_n3349_ );
and  ( new_n3352_, new_n3351_, new_n3303_ );
xnor ( new_n3353_, new_n3136_, new_n3134_ );
xor  ( new_n3354_, new_n3353_, new_n3294_ );
nor  ( new_n3355_, new_n3354_, new_n3352_ );
and  ( new_n3356_, new_n3354_, new_n3352_ );
xnor ( new_n3357_, new_n3347_, new_n3345_ );
xnor ( new_n3358_, new_n3249_, new_n3245_ );
xor  ( new_n3359_, new_n3358_, new_n3255_ );
not  ( new_n3360_, new_n3277_ );
xor  ( new_n3361_, new_n3360_, new_n3267_ );
xor  ( new_n3362_, new_n3361_, new_n3282_ );
or   ( new_n3363_, new_n3362_, new_n3359_ );
and  ( new_n3364_, new_n3362_, new_n3359_ );
xor  ( new_n3365_, new_n3244_, new_n2233_ );
or   ( new_n3366_, new_n3365_, new_n2232_ );
or   ( new_n3367_, new_n3279_, new_n2300_ );
and  ( new_n3368_, new_n3367_, new_n3366_ );
and  ( new_n3369_, new_n3368_, new_n3360_ );
nor  ( new_n3370_, new_n3368_, new_n3360_ );
not  ( new_n3371_, new_n3370_ );
xor  ( new_n3372_, new_n3026_, new_n2297_ );
nand ( new_n3373_, new_n3372_, new_n3272_ );
xor  ( new_n3374_, new_n3230_, new_n3181_ );
nand ( new_n3375_, new_n3374_, new_n3273_ );
and  ( new_n3376_, new_n3375_, new_n3373_ );
xor  ( new_n3377_, new_n2692_, new_n2566_ );
nand ( new_n3378_, new_n3377_, new_n2905_ );
nand ( new_n3379_, new_n3332_, new_n3033_ );
and  ( new_n3380_, new_n3379_, new_n3378_ );
and  ( new_n3381_, new_n3380_, new_n3376_ );
and  ( new_n3382_, new_n3381_, new_n3371_ );
nor  ( new_n3383_, new_n3382_, new_n3369_ );
or   ( new_n3384_, new_n3383_, new_n3364_ );
and  ( new_n3385_, new_n3384_, new_n3363_ );
nor  ( new_n3386_, new_n3385_, new_n3357_ );
xor  ( new_n3387_, new_n3385_, new_n3357_ );
xor  ( new_n3388_, new_n2856_, new_n2304_ );
and  ( new_n3389_, new_n3388_, new_n3070_ );
and  ( new_n3390_, new_n3308_, new_n3068_ );
nor  ( new_n3391_, new_n3390_, new_n3389_ );
xor  ( new_n3392_, new_n2923_, new_n2395_ );
and  ( new_n3393_, new_n3392_, new_n2558_ );
and  ( new_n3394_, new_n3323_, new_n2603_ );
nor  ( new_n3395_, new_n3394_, new_n3393_ );
nor  ( new_n3396_, new_n3395_, new_n3391_ );
xor  ( new_n3397_, new_n2723_, new_n2542_ );
and  ( new_n3398_, new_n3397_, new_n2729_ );
and  ( new_n3399_, new_n3315_, new_n2781_ );
nor  ( new_n3400_, new_n3399_, new_n3398_ );
not  ( new_n3401_, new_n3400_ );
and  ( new_n3402_, new_n3395_, new_n3391_ );
not  ( new_n3403_, new_n3402_ );
and  ( new_n3404_, new_n3403_, new_n3401_ );
or   ( new_n3405_, new_n3404_, new_n3396_ );
xnor ( new_n3406_, new_n3154_, new_n2262_ );
not  ( new_n3407_, new_n3406_ );
and  ( new_n3408_, new_n3407_, new_n2233_ );
or   ( new_n3409_, new_n3408_, new_n3230_ );
xor  ( new_n3410_, new_n3306_, new_n2233_ );
nor  ( new_n3411_, new_n3410_, new_n2232_ );
nor  ( new_n3412_, new_n3365_, new_n2300_ );
or   ( new_n3413_, new_n3412_, new_n3411_ );
and  ( new_n3414_, new_n3408_, new_n3230_ );
or   ( new_n3415_, new_n3414_, new_n3413_ );
and  ( new_n3416_, new_n3415_, new_n3409_ );
and  ( new_n3417_, new_n3416_, new_n3405_ );
or   ( new_n3418_, new_n3416_, new_n3405_ );
xor  ( new_n3419_, new_n3330_, new_n3326_ );
xnor ( new_n3420_, new_n3419_, new_n3335_ );
and  ( new_n3421_, new_n3420_, new_n3418_ );
or   ( new_n3422_, new_n3421_, new_n3417_ );
xnor ( new_n3423_, new_n3320_, new_n3305_ );
xor  ( new_n3424_, new_n3423_, new_n3338_ );
nand ( new_n3425_, new_n3424_, new_n3422_ );
nor  ( new_n3426_, new_n3424_, new_n3422_ );
xor  ( new_n3427_, new_n3312_, new_n3307_ );
xor  ( new_n3428_, new_n3427_, new_n3318_ );
xor  ( new_n3429_, new_n3368_, new_n3360_ );
xor  ( new_n3430_, new_n3429_, new_n3381_ );
or   ( new_n3431_, new_n3430_, new_n3428_ );
nand ( new_n3432_, new_n3430_, new_n3428_ );
xor  ( new_n3433_, new_n3380_, new_n3376_ );
xor  ( new_n3434_, new_n3108_, new_n2178_ );
nand ( new_n3435_, new_n3434_, new_n2402_ );
or   ( new_n3436_, new_n3327_, new_n2446_ );
and  ( new_n3437_, new_n3436_, new_n3435_ );
nor  ( new_n3438_, new_n3437_, new_n3433_ );
nand ( new_n3439_, new_n3438_, new_n3432_ );
and  ( new_n3440_, new_n3439_, new_n3431_ );
or   ( new_n3441_, new_n3440_, new_n3426_ );
and  ( new_n3442_, new_n3441_, new_n3425_ );
and  ( new_n3443_, new_n3442_, new_n3387_ );
or   ( new_n3444_, new_n3443_, new_n3386_ );
xor  ( new_n3445_, new_n3350_, new_n3349_ );
and  ( new_n3446_, new_n3445_, new_n3444_ );
nor  ( new_n3447_, new_n3445_, new_n3444_ );
xor  ( new_n3448_, new_n3424_, new_n3422_ );
xor  ( new_n3449_, new_n3448_, new_n3440_ );
xnor ( new_n3450_, new_n3362_, new_n3359_ );
xor  ( new_n3451_, new_n3450_, new_n3383_ );
and  ( new_n3452_, new_n3451_, new_n3449_ );
xnor ( new_n3453_, new_n3416_, new_n3405_ );
xor  ( new_n3454_, new_n3453_, new_n3420_ );
xor  ( new_n3455_, new_n2760_, new_n3235_ );
or   ( new_n3456_, new_n3455_, new_n2730_ );
nand ( new_n3457_, new_n3397_, new_n2781_ );
and  ( new_n3458_, new_n3457_, new_n3456_ );
or   ( new_n3459_, new_n3230_, new_n2407_ );
and  ( new_n3460_, new_n2089_, new_n993_ );
nor  ( new_n3461_, new_n3460_, new_n2052_ );
nor  ( new_n3462_, new_n3461_, new_n86_ );
not  ( new_n3463_, new_n3462_ );
and  ( new_n3464_, new_n2079_, \a[0]  );
not  ( new_n3465_, new_n3464_ );
and  ( new_n3466_, new_n2083_, \b[0]  );
nor  ( new_n3467_, new_n3466_, \c[0]  );
and  ( new_n3468_, new_n2082_, new_n1714_ );
and  ( new_n3469_, new_n3468_, new_n2058_ );
nor  ( new_n3470_, new_n3469_, new_n804_ );
not  ( new_n3471_, new_n3470_ );
and  ( new_n3472_, new_n2089_, new_n86_ );
nor  ( new_n3473_, new_n3472_, new_n2066_ );
and  ( new_n3474_, new_n3473_, new_n3471_ );
nor  ( new_n3475_, new_n3474_, new_n3467_ );
not  ( new_n3476_, new_n3475_ );
and  ( new_n3477_, \d[0] , \a[0]  );
and  ( new_n3478_, new_n3477_, new_n937_ );
not  ( new_n3479_, new_n3478_ );
xor  ( new_n3480_, \d[0] , \b[0]  );
and  ( new_n3481_, new_n3480_, new_n1844_ );
xor  ( new_n3482_, \c[0] , \a[0]  );
and  ( new_n3483_, new_n3482_, new_n1780_ );
nor  ( new_n3484_, new_n3483_, new_n3481_ );
and  ( new_n3485_, new_n3484_, new_n3479_ );
and  ( new_n3486_, new_n3485_, new_n3476_ );
and  ( new_n3487_, new_n3486_, new_n3465_ );
and  ( new_n3488_, new_n3487_, new_n3463_ );
nor  ( new_n3489_, new_n3488_, new_n3230_ );
not  ( new_n3490_, new_n3489_ );
and  ( new_n3491_, new_n3490_, new_n3459_ );
nor  ( new_n3492_, new_n3491_, new_n3458_ );
xor  ( new_n3493_, new_n2856_, new_n2440_ );
and  ( new_n3494_, new_n3493_, new_n3070_ );
and  ( new_n3495_, new_n3388_, new_n3068_ );
or   ( new_n3496_, new_n3495_, new_n3494_ );
xor  ( new_n3497_, new_n3491_, new_n3458_ );
and  ( new_n3498_, new_n3497_, new_n3496_ );
or   ( new_n3499_, new_n3498_, new_n3492_ );
xor  ( new_n3500_, new_n3395_, new_n3391_ );
or   ( new_n3501_, new_n3500_, new_n3401_ );
not  ( new_n3502_, new_n3404_ );
or   ( new_n3503_, new_n3502_, new_n3396_ );
and  ( new_n3504_, new_n3503_, new_n3501_ );
nand ( new_n3505_, new_n3504_, new_n3499_ );
nor  ( new_n3506_, new_n3504_, new_n3499_ );
xnor ( new_n3507_, new_n3195_, new_n2260_ );
or   ( new_n3508_, new_n3507_, new_n2134_ );
xor  ( new_n3509_, new_n3406_, new_n2233_ );
or   ( new_n3510_, new_n3509_, new_n2232_ );
or   ( new_n3511_, new_n3410_, new_n2300_ );
and  ( new_n3512_, new_n3511_, new_n3510_ );
nor  ( new_n3513_, new_n3512_, new_n3508_ );
and  ( new_n3514_, new_n3512_, new_n3508_ );
xor  ( new_n3515_, new_n2705_, new_n2692_ );
and  ( new_n3516_, new_n3515_, new_n2905_ );
and  ( new_n3517_, new_n3377_, new_n3033_ );
nor  ( new_n3518_, new_n3517_, new_n3516_ );
nor  ( new_n3519_, new_n3518_, new_n3514_ );
nor  ( new_n3520_, new_n3519_, new_n3513_ );
or   ( new_n3521_, new_n3520_, new_n3506_ );
and  ( new_n3522_, new_n3521_, new_n3505_ );
nor  ( new_n3523_, new_n3522_, new_n3454_ );
and  ( new_n3524_, new_n3522_, new_n3454_ );
xor  ( new_n3525_, new_n3026_, new_n2288_ );
and  ( new_n3526_, new_n3525_, new_n3272_ );
and  ( new_n3527_, new_n3374_, new_n3372_ );
nor  ( new_n3528_, new_n3527_, new_n3526_ );
not  ( new_n3529_, new_n3528_ );
xor  ( new_n3530_, new_n3244_, new_n2178_ );
and  ( new_n3531_, new_n3530_, new_n2402_ );
and  ( new_n3532_, new_n3434_, new_n2445_ );
nor  ( new_n3533_, new_n3532_, new_n3531_ );
not  ( new_n3534_, new_n3533_ );
and  ( new_n3535_, new_n3534_, new_n3529_ );
xor  ( new_n3536_, new_n3066_, new_n2395_ );
and  ( new_n3537_, new_n3536_, new_n2558_ );
and  ( new_n3538_, new_n3392_, new_n2603_ );
nor  ( new_n3539_, new_n3538_, new_n3537_ );
and  ( new_n3540_, new_n3533_, new_n3528_ );
nor  ( new_n3541_, new_n3540_, new_n3539_ );
or   ( new_n3542_, new_n3541_, new_n3535_ );
xor  ( new_n3543_, new_n3408_, new_n3230_ );
xor  ( new_n3544_, new_n3543_, new_n3413_ );
and  ( new_n3545_, new_n3544_, new_n3542_ );
nor  ( new_n3546_, new_n3544_, new_n3542_ );
xor  ( new_n3547_, \d[0] , \c[0]  );
not  ( new_n3548_, new_n3547_ );
or   ( new_n3549_, new_n3548_, new_n2134_ );
xor  ( new_n3550_, new_n3230_, new_n2407_ );
or   ( new_n3551_, new_n3550_, new_n3488_ );
not  ( new_n3552_, new_n3488_ );
nor  ( new_n3553_, new_n3552_, new_n3230_ );
not  ( new_n3554_, new_n3553_ );
or   ( new_n3555_, new_n3554_, new_n3143_ );
and  ( new_n3556_, new_n3555_, new_n3551_ );
or   ( new_n3557_, new_n3556_, new_n3549_ );
xor  ( new_n3558_, new_n3026_, new_n2304_ );
and  ( new_n3559_, new_n3558_, new_n3272_ );
and  ( new_n3560_, new_n3525_, new_n3374_ );
or   ( new_n3561_, new_n3560_, new_n3559_ );
xor  ( new_n3562_, new_n3556_, new_n3549_ );
nand ( new_n3563_, new_n3562_, new_n3561_ );
and  ( new_n3564_, new_n3563_, new_n3557_ );
xor  ( new_n3565_, new_n3108_, new_n2395_ );
and  ( new_n3566_, new_n3565_, new_n2558_ );
and  ( new_n3567_, new_n3536_, new_n2603_ );
nor  ( new_n3568_, new_n3567_, new_n3566_ );
xor  ( new_n3569_, new_n2856_, new_n2566_ );
and  ( new_n3570_, new_n3569_, new_n3070_ );
and  ( new_n3571_, new_n3493_, new_n3068_ );
nor  ( new_n3572_, new_n3571_, new_n3570_ );
nor  ( new_n3573_, new_n3572_, new_n3568_ );
xor  ( new_n3574_, new_n3306_, new_n2178_ );
and  ( new_n3575_, new_n3574_, new_n2402_ );
and  ( new_n3576_, new_n3530_, new_n2445_ );
nor  ( new_n3577_, new_n3576_, new_n3575_ );
not  ( new_n3578_, new_n3577_ );
and  ( new_n3579_, new_n3572_, new_n3568_ );
not  ( new_n3580_, new_n3579_ );
and  ( new_n3581_, new_n3580_, new_n3578_ );
nor  ( new_n3582_, new_n3581_, new_n3573_ );
nor  ( new_n3583_, new_n3582_, new_n3564_ );
xor  ( new_n3584_, new_n2923_, new_n3235_ );
or   ( new_n3585_, new_n3584_, new_n2730_ );
or   ( new_n3586_, new_n3455_, new_n2782_ );
and  ( new_n3587_, new_n3586_, new_n3585_ );
xor  ( new_n3588_, new_n2723_, new_n2692_ );
nand ( new_n3589_, new_n3588_, new_n2905_ );
nand ( new_n3590_, new_n3515_, new_n3033_ );
and  ( new_n3591_, new_n3590_, new_n3589_ );
nor  ( new_n3592_, new_n3591_, new_n3587_ );
xor  ( new_n3593_, new_n3507_, new_n2233_ );
nor  ( new_n3594_, new_n3593_, new_n2232_ );
nor  ( new_n3595_, new_n3509_, new_n2300_ );
nor  ( new_n3596_, new_n3595_, new_n3594_ );
xnor ( new_n3597_, new_n3591_, new_n3587_ );
nor  ( new_n3598_, new_n3597_, new_n3596_ );
or   ( new_n3599_, new_n3598_, new_n3592_ );
xor  ( new_n3600_, new_n3582_, new_n3564_ );
and  ( new_n3601_, new_n3600_, new_n3599_ );
nor  ( new_n3602_, new_n3601_, new_n3583_ );
nor  ( new_n3603_, new_n3602_, new_n3546_ );
nor  ( new_n3604_, new_n3603_, new_n3545_ );
nor  ( new_n3605_, new_n3604_, new_n3524_ );
nor  ( new_n3606_, new_n3605_, new_n3523_ );
or   ( new_n3607_, new_n3606_, new_n3452_ );
or   ( new_n3608_, new_n3451_, new_n3449_ );
and  ( new_n3609_, new_n3608_, new_n3607_ );
xor  ( new_n3610_, new_n3442_, new_n3387_ );
and  ( new_n3611_, new_n3610_, new_n3609_ );
nor  ( new_n3612_, new_n3610_, new_n3609_ );
xor  ( new_n3613_, new_n3437_, new_n3433_ );
xnor ( new_n3614_, new_n3504_, new_n3499_ );
xor  ( new_n3615_, new_n3614_, new_n3520_ );
nor  ( new_n3616_, new_n3615_, new_n3613_ );
and  ( new_n3617_, new_n3615_, new_n3613_ );
xor  ( new_n3618_, new_n3497_, new_n3496_ );
xnor ( new_n3619_, new_n3512_, new_n3508_ );
xor  ( new_n3620_, new_n3619_, new_n3518_ );
nor  ( new_n3621_, new_n3620_, new_n3618_ );
and  ( new_n3622_, new_n3620_, new_n3618_ );
not  ( new_n3623_, new_n3539_ );
xor  ( new_n3624_, new_n3533_, new_n3528_ );
nor  ( new_n3625_, new_n3624_, new_n3623_ );
not  ( new_n3626_, new_n3535_ );
and  ( new_n3627_, new_n3541_, new_n3626_ );
nor  ( new_n3628_, new_n3627_, new_n3625_ );
nor  ( new_n3629_, new_n3628_, new_n3622_ );
nor  ( new_n3630_, new_n3629_, new_n3621_ );
nor  ( new_n3631_, new_n3630_, new_n3617_ );
nor  ( new_n3632_, new_n3631_, new_n3616_ );
xor  ( new_n3633_, new_n3430_, new_n3428_ );
xor  ( new_n3634_, new_n3633_, new_n3438_ );
or   ( new_n3635_, new_n3634_, new_n3632_ );
xor  ( new_n3636_, new_n3634_, new_n3632_ );
xnor ( new_n3637_, new_n3522_, new_n3454_ );
xnor ( new_n3638_, new_n3637_, new_n3604_ );
nand ( new_n3639_, new_n3638_, new_n3636_ );
and  ( new_n3640_, new_n3639_, new_n3635_ );
xnor ( new_n3641_, new_n3451_, new_n3449_ );
xor  ( new_n3642_, new_n3641_, new_n3606_ );
nor  ( new_n3643_, new_n3642_, new_n3640_ );
and  ( new_n3644_, new_n3642_, new_n3640_ );
xnor ( new_n3645_, new_n3638_, new_n3636_ );
xor  ( new_n3646_, new_n3615_, new_n3613_ );
xor  ( new_n3647_, new_n3646_, new_n3630_ );
xnor ( new_n3648_, new_n3544_, new_n3542_ );
xor  ( new_n3649_, new_n3648_, new_n3602_ );
or   ( new_n3650_, new_n3649_, new_n3647_ );
nand ( new_n3651_, new_n3649_, new_n3647_ );
xor  ( new_n3652_, new_n3026_, new_n2440_ );
and  ( new_n3653_, new_n3652_, new_n3272_ );
and  ( new_n3654_, new_n3558_, new_n3374_ );
or   ( new_n3655_, new_n3654_, new_n3653_ );
and  ( new_n3656_, new_n3547_, new_n2228_ );
or   ( new_n3657_, new_n3656_, new_n2230_ );
nor  ( new_n3658_, new_n3657_, new_n2134_ );
and  ( new_n3659_, new_n3658_, new_n3655_ );
xor  ( new_n3660_, new_n3562_, new_n3561_ );
and  ( new_n3661_, new_n3660_, new_n3659_ );
or   ( new_n3662_, new_n3230_, new_n2420_ );
or   ( new_n3663_, new_n3662_, new_n3552_ );
and  ( new_n3664_, new_n3230_, new_n2297_ );
nor  ( new_n3665_, new_n3230_, new_n2297_ );
or   ( new_n3666_, new_n3665_, new_n3488_ );
or   ( new_n3667_, new_n3666_, new_n3664_ );
and  ( new_n3668_, new_n3667_, new_n3663_ );
or   ( new_n3669_, new_n3593_, new_n2300_ );
nand ( new_n3670_, new_n3548_, new_n2229_ );
nand ( new_n3671_, new_n3547_, new_n2231_ );
and  ( new_n3672_, new_n3671_, new_n3670_ );
and  ( new_n3673_, new_n3672_, new_n3669_ );
nor  ( new_n3674_, new_n3673_, new_n3668_ );
xor  ( new_n3675_, new_n2760_, new_n2692_ );
and  ( new_n3676_, new_n3675_, new_n2905_ );
and  ( new_n3677_, new_n3588_, new_n3033_ );
or   ( new_n3678_, new_n3677_, new_n3676_ );
xor  ( new_n3679_, new_n3673_, new_n3668_ );
and  ( new_n3680_, new_n3679_, new_n3678_ );
or   ( new_n3681_, new_n3680_, new_n3674_ );
xor  ( new_n3682_, new_n3660_, new_n3659_ );
and  ( new_n3683_, new_n3682_, new_n3681_ );
or   ( new_n3684_, new_n3683_, new_n3661_ );
xor  ( new_n3685_, new_n3600_, new_n3599_ );
and  ( new_n3686_, new_n3685_, new_n3684_ );
nor  ( new_n3687_, new_n3685_, new_n3684_ );
xnor ( new_n3688_, new_n3597_, new_n3596_ );
xor  ( new_n3689_, new_n3244_, new_n2395_ );
nand ( new_n3690_, new_n3689_, new_n2558_ );
nand ( new_n3691_, new_n3565_, new_n2603_ );
and  ( new_n3692_, new_n3691_, new_n3690_ );
not  ( new_n3693_, new_n2705_ );
xor  ( new_n3694_, new_n2856_, new_n3693_ );
or   ( new_n3695_, new_n3694_, new_n3142_ );
nand ( new_n3696_, new_n3569_, new_n3068_ );
and  ( new_n3697_, new_n3696_, new_n3695_ );
or   ( new_n3698_, new_n3697_, new_n3692_ );
xor  ( new_n3699_, new_n3066_, new_n3235_ );
or   ( new_n3700_, new_n3699_, new_n2730_ );
or   ( new_n3701_, new_n3584_, new_n2782_ );
and  ( new_n3702_, new_n3701_, new_n3700_ );
and  ( new_n3703_, new_n3697_, new_n3692_ );
or   ( new_n3704_, new_n3703_, new_n3702_ );
and  ( new_n3705_, new_n3704_, new_n3698_ );
nor  ( new_n3706_, new_n3705_, new_n3688_ );
and  ( new_n3707_, new_n3705_, new_n3688_ );
not  ( new_n3708_, new_n3707_ );
xor  ( new_n3709_, new_n3572_, new_n3568_ );
nor  ( new_n3710_, new_n3709_, new_n3578_ );
not  ( new_n3711_, new_n3573_ );
and  ( new_n3712_, new_n3581_, new_n3711_ );
nor  ( new_n3713_, new_n3712_, new_n3710_ );
and  ( new_n3714_, new_n3713_, new_n3708_ );
nor  ( new_n3715_, new_n3714_, new_n3706_ );
nor  ( new_n3716_, new_n3715_, new_n3687_ );
nor  ( new_n3717_, new_n3716_, new_n3686_ );
nand ( new_n3718_, new_n3717_, new_n3651_ );
and  ( new_n3719_, new_n3718_, new_n3650_ );
nor  ( new_n3720_, new_n3719_, new_n3645_ );
and  ( new_n3721_, new_n3719_, new_n3645_ );
xor  ( new_n3722_, new_n3649_, new_n3647_ );
xor  ( new_n3723_, new_n3722_, new_n3717_ );
xor  ( new_n3724_, new_n3406_, new_n2178_ );
and  ( new_n3725_, new_n3724_, new_n2402_ );
and  ( new_n3726_, new_n3574_, new_n2445_ );
or   ( new_n3727_, new_n3726_, new_n3725_ );
xor  ( new_n3728_, new_n3658_, new_n3655_ );
nand ( new_n3729_, new_n3728_, new_n3727_ );
nor  ( new_n3730_, new_n3728_, new_n3727_ );
or   ( new_n3731_, new_n3548_, new_n2300_ );
xnor ( new_n3732_, new_n3230_, new_n2288_ );
or   ( new_n3733_, new_n3732_, new_n3488_ );
not  ( new_n3734_, new_n2304_ );
or   ( new_n3735_, new_n3554_, new_n3734_ );
and  ( new_n3736_, new_n3735_, new_n3733_ );
or   ( new_n3737_, new_n3736_, new_n3731_ );
and  ( new_n3738_, new_n3652_, new_n3374_ );
xor  ( new_n3739_, new_n3026_, new_n2566_ );
and  ( new_n3740_, new_n3739_, new_n3272_ );
nor  ( new_n3741_, new_n3740_, new_n3738_ );
xnor ( new_n3742_, new_n3736_, new_n3731_ );
or   ( new_n3743_, new_n3742_, new_n3741_ );
and  ( new_n3744_, new_n3743_, new_n3737_ );
or   ( new_n3745_, new_n3744_, new_n3730_ );
and  ( new_n3746_, new_n3745_, new_n3729_ );
xor  ( new_n3747_, new_n3697_, new_n3692_ );
xor  ( new_n3748_, new_n3747_, new_n3702_ );
not  ( new_n3749_, new_n2905_ );
xor  ( new_n3750_, new_n2923_, new_n2901_ );
or   ( new_n3751_, new_n3750_, new_n3749_ );
nand ( new_n3752_, new_n3675_, new_n3033_ );
and  ( new_n3753_, new_n3752_, new_n3751_ );
xor  ( new_n3754_, new_n2856_, new_n2723_ );
nand ( new_n3755_, new_n3754_, new_n3070_ );
or   ( new_n3756_, new_n3694_, new_n3310_ );
and  ( new_n3757_, new_n3756_, new_n3755_ );
or   ( new_n3758_, new_n3757_, new_n3753_ );
xor  ( new_n3759_, new_n3108_, new_n2542_ );
nand ( new_n3760_, new_n3759_, new_n2729_ );
or   ( new_n3761_, new_n3699_, new_n2782_ );
and  ( new_n3762_, new_n3761_, new_n3760_ );
and  ( new_n3763_, new_n3757_, new_n3753_ );
or   ( new_n3764_, new_n3763_, new_n3762_ );
and  ( new_n3765_, new_n3764_, new_n3758_ );
or   ( new_n3766_, new_n3765_, new_n3748_ );
and  ( new_n3767_, new_n3765_, new_n3748_ );
and  ( new_n3768_, new_n3739_, new_n3374_ );
xor  ( new_n3769_, new_n3026_, new_n2705_ );
and  ( new_n3770_, new_n3769_, new_n3272_ );
nor  ( new_n3771_, new_n3770_, new_n3768_ );
and  ( new_n3772_, new_n3547_, new_n2400_ );
or   ( new_n3773_, new_n3772_, new_n2411_ );
or   ( new_n3774_, new_n3773_, new_n3771_ );
xor  ( new_n3775_, new_n3507_, new_n2178_ );
nand ( new_n3776_, new_n3775_, new_n2402_ );
nand ( new_n3777_, new_n3724_, new_n2445_ );
and  ( new_n3778_, new_n3777_, new_n3776_ );
nor  ( new_n3779_, new_n3778_, new_n3774_ );
and  ( new_n3780_, new_n3778_, new_n3774_ );
xor  ( new_n3781_, new_n3306_, new_n2395_ );
and  ( new_n3782_, new_n3781_, new_n2558_ );
and  ( new_n3783_, new_n3689_, new_n2603_ );
nor  ( new_n3784_, new_n3783_, new_n3782_ );
nor  ( new_n3785_, new_n3784_, new_n3780_ );
nor  ( new_n3786_, new_n3785_, new_n3779_ );
or   ( new_n3787_, new_n3786_, new_n3767_ );
and  ( new_n3788_, new_n3787_, new_n3766_ );
nor  ( new_n3789_, new_n3788_, new_n3746_ );
nand ( new_n3790_, new_n3788_, new_n3746_ );
xor  ( new_n3791_, new_n3682_, new_n3681_ );
and  ( new_n3792_, new_n3791_, new_n3790_ );
or   ( new_n3793_, new_n3792_, new_n3789_ );
xor  ( new_n3794_, new_n3620_, new_n3618_ );
xor  ( new_n3795_, new_n3794_, new_n3628_ );
nand ( new_n3796_, new_n3795_, new_n3793_ );
nor  ( new_n3797_, new_n3795_, new_n3793_ );
xor  ( new_n3798_, new_n3685_, new_n3684_ );
xor  ( new_n3799_, new_n3798_, new_n3715_ );
or   ( new_n3800_, new_n3799_, new_n3797_ );
and  ( new_n3801_, new_n3800_, new_n3796_ );
nor  ( new_n3802_, new_n3801_, new_n3723_ );
and  ( new_n3803_, new_n3801_, new_n3723_ );
xnor ( new_n3804_, new_n3742_, new_n3741_ );
xor  ( new_n3805_, new_n3066_, new_n2692_ );
nand ( new_n3806_, new_n3805_, new_n2905_ );
xor  ( new_n3807_, new_n2923_, new_n2692_ );
nand ( new_n3808_, new_n3807_, new_n3033_ );
and  ( new_n3809_, new_n3808_, new_n3806_ );
xnor ( new_n3810_, new_n3230_, new_n2304_ );
or   ( new_n3811_, new_n3810_, new_n3488_ );
or   ( new_n3812_, new_n3554_, new_n2441_ );
and  ( new_n3813_, new_n3812_, new_n3811_ );
or   ( new_n3814_, new_n3813_, new_n3809_ );
xor  ( new_n3815_, new_n3244_, new_n2542_ );
and  ( new_n3816_, new_n3815_, new_n2729_ );
and  ( new_n3817_, new_n3759_, new_n2781_ );
nor  ( new_n3818_, new_n3817_, new_n3816_ );
and  ( new_n3819_, new_n3813_, new_n3809_ );
or   ( new_n3820_, new_n3819_, new_n3818_ );
and  ( new_n3821_, new_n3820_, new_n3814_ );
nor  ( new_n3822_, new_n3821_, new_n3804_ );
and  ( new_n3823_, new_n3821_, new_n3804_ );
xor  ( new_n3824_, new_n2856_, new_n2760_ );
and  ( new_n3825_, new_n3824_, new_n3070_ );
and  ( new_n3826_, new_n3754_, new_n3068_ );
nor  ( new_n3827_, new_n3826_, new_n3825_ );
not  ( new_n3828_, new_n3827_ );
and  ( new_n3829_, new_n3775_, new_n2445_ );
xor  ( new_n3830_, new_n3547_, new_n2395_ );
and  ( new_n3831_, new_n3830_, new_n2402_ );
nor  ( new_n3832_, new_n3831_, new_n3829_ );
not  ( new_n3833_, new_n3832_ );
and  ( new_n3834_, new_n3833_, new_n3828_ );
xor  ( new_n3835_, new_n3406_, new_n2395_ );
and  ( new_n3836_, new_n3835_, new_n2558_ );
and  ( new_n3837_, new_n3781_, new_n2603_ );
nor  ( new_n3838_, new_n3837_, new_n3836_ );
and  ( new_n3839_, new_n3832_, new_n3827_ );
nor  ( new_n3840_, new_n3839_, new_n3838_ );
nor  ( new_n3841_, new_n3840_, new_n3834_ );
nor  ( new_n3842_, new_n3841_, new_n3823_ );
nor  ( new_n3843_, new_n3842_, new_n3822_ );
xnor ( new_n3844_, new_n3679_, new_n3678_ );
nor  ( new_n3845_, new_n3844_, new_n3843_ );
xnor ( new_n3846_, new_n3844_, new_n3843_ );
xor  ( new_n3847_, new_n3728_, new_n3727_ );
xor  ( new_n3848_, new_n3847_, new_n3744_ );
nor  ( new_n3849_, new_n3848_, new_n3846_ );
or   ( new_n3850_, new_n3849_, new_n3845_ );
xor  ( new_n3851_, new_n3705_, new_n3688_ );
xor  ( new_n3852_, new_n3851_, new_n3713_ );
nand ( new_n3853_, new_n3852_, new_n3850_ );
xor  ( new_n3854_, new_n3852_, new_n3850_ );
xor  ( new_n3855_, new_n3788_, new_n3746_ );
xor  ( new_n3856_, new_n3855_, new_n3791_ );
nand ( new_n3857_, new_n3856_, new_n3854_ );
and  ( new_n3858_, new_n3857_, new_n3853_ );
xor  ( new_n3859_, new_n3795_, new_n3793_ );
xor  ( new_n3860_, new_n3859_, new_n3799_ );
and  ( new_n3861_, new_n3860_, new_n3858_ );
nor  ( new_n3862_, new_n3860_, new_n3858_ );
xor  ( new_n3863_, new_n3757_, new_n3753_ );
xor  ( new_n3864_, new_n3863_, new_n3762_ );
xor  ( new_n3865_, new_n3778_, new_n3774_ );
xor  ( new_n3866_, new_n3865_, new_n3784_ );
nor  ( new_n3867_, new_n3866_, new_n3864_ );
nand ( new_n3868_, new_n3866_, new_n3864_ );
xnor ( new_n3869_, new_n3773_, new_n3771_ );
xor  ( new_n3870_, new_n3230_, new_n2440_ );
and  ( new_n3871_, new_n3870_, new_n3552_ );
and  ( new_n3872_, new_n3553_, new_n2566_ );
or   ( new_n3873_, new_n3872_, new_n3871_ );
and  ( new_n3874_, new_n3772_, new_n2397_ );
nand ( new_n3875_, new_n3874_, new_n3873_ );
nor  ( new_n3876_, new_n3874_, new_n3873_ );
xor  ( new_n3877_, new_n3026_, new_n2723_ );
and  ( new_n3878_, new_n3877_, new_n3272_ );
and  ( new_n3879_, new_n3769_, new_n3374_ );
nor  ( new_n3880_, new_n3879_, new_n3878_ );
or   ( new_n3881_, new_n3880_, new_n3876_ );
and  ( new_n3882_, new_n3881_, new_n3875_ );
nor  ( new_n3883_, new_n3882_, new_n3869_ );
nand ( new_n3884_, new_n3882_, new_n3869_ );
xor  ( new_n3885_, new_n3306_, new_n2542_ );
and  ( new_n3886_, new_n3885_, new_n2729_ );
and  ( new_n3887_, new_n3815_, new_n2781_ );
nor  ( new_n3888_, new_n3887_, new_n3886_ );
xor  ( new_n3889_, new_n3507_, new_n2395_ );
and  ( new_n3890_, new_n3889_, new_n2558_ );
and  ( new_n3891_, new_n3835_, new_n2603_ );
nor  ( new_n3892_, new_n3891_, new_n3890_ );
nor  ( new_n3893_, new_n3892_, new_n3888_ );
and  ( new_n3894_, new_n3892_, new_n3888_ );
not  ( new_n3895_, new_n3894_ );
xor  ( new_n3896_, new_n3108_, new_n2692_ );
and  ( new_n3897_, new_n3896_, new_n2905_ );
and  ( new_n3898_, new_n3805_, new_n3033_ );
nor  ( new_n3899_, new_n3898_, new_n3897_ );
not  ( new_n3900_, new_n3899_ );
and  ( new_n3901_, new_n3900_, new_n3895_ );
or   ( new_n3902_, new_n3901_, new_n3893_ );
and  ( new_n3903_, new_n3902_, new_n3884_ );
or   ( new_n3904_, new_n3903_, new_n3883_ );
and  ( new_n3905_, new_n3904_, new_n3868_ );
or   ( new_n3906_, new_n3905_, new_n3867_ );
xnor ( new_n3907_, new_n3765_, new_n3748_ );
xor  ( new_n3908_, new_n3907_, new_n3786_ );
and  ( new_n3909_, new_n3908_, new_n3906_ );
xor  ( new_n3910_, new_n3848_, new_n3846_ );
xor  ( new_n3911_, new_n3908_, new_n3906_ );
and  ( new_n3912_, new_n3911_, new_n3910_ );
or   ( new_n3913_, new_n3912_, new_n3909_ );
xor  ( new_n3914_, new_n3856_, new_n3854_ );
nor  ( new_n3915_, new_n3914_, new_n3913_ );
and  ( new_n3916_, new_n3914_, new_n3913_ );
xor  ( new_n3917_, new_n3813_, new_n3809_ );
xnor ( new_n3918_, new_n3917_, new_n3818_ );
not  ( new_n3919_, new_n3918_ );
xor  ( new_n3920_, new_n2923_, new_n2856_ );
and  ( new_n3921_, new_n3920_, new_n3070_ );
and  ( new_n3922_, new_n3824_, new_n3068_ );
or   ( new_n3923_, new_n3922_, new_n3921_ );
and  ( new_n3924_, new_n3877_, new_n3374_ );
xor  ( new_n3925_, new_n3026_, new_n2760_ );
and  ( new_n3926_, new_n3925_, new_n3272_ );
or   ( new_n3927_, new_n3926_, new_n3924_ );
nand ( new_n3928_, new_n3547_, new_n2562_ );
and  ( new_n3929_, new_n3928_, new_n2544_ );
and  ( new_n3930_, new_n3929_, new_n3927_ );
nand ( new_n3931_, new_n3930_, new_n3923_ );
nor  ( new_n3932_, new_n3930_, new_n3923_ );
xor  ( new_n3933_, new_n3244_, new_n2692_ );
and  ( new_n3934_, new_n3933_, new_n2905_ );
and  ( new_n3935_, new_n3896_, new_n3033_ );
nor  ( new_n3936_, new_n3935_, new_n3934_ );
not  ( new_n3937_, new_n3936_ );
nor  ( new_n3938_, new_n3230_, new_n3693_ );
and  ( new_n3939_, new_n3938_, new_n3488_ );
xor  ( new_n3940_, new_n3230_, new_n2566_ );
and  ( new_n3941_, new_n3940_, new_n3552_ );
nor  ( new_n3942_, new_n3941_, new_n3939_ );
not  ( new_n3943_, new_n3942_ );
and  ( new_n3944_, new_n3943_, new_n3937_ );
xor  ( new_n3945_, new_n3406_, new_n2542_ );
and  ( new_n3946_, new_n3945_, new_n2729_ );
and  ( new_n3947_, new_n3885_, new_n2781_ );
nor  ( new_n3948_, new_n3947_, new_n3946_ );
and  ( new_n3949_, new_n3942_, new_n3936_ );
nor  ( new_n3950_, new_n3949_, new_n3948_ );
nor  ( new_n3951_, new_n3950_, new_n3944_ );
or   ( new_n3952_, new_n3951_, new_n3932_ );
and  ( new_n3953_, new_n3952_, new_n3931_ );
and  ( new_n3954_, new_n3953_, new_n3919_ );
xor  ( new_n3955_, new_n3953_, new_n3919_ );
xor  ( new_n3956_, new_n3832_, new_n3828_ );
nand ( new_n3957_, new_n3956_, new_n3838_ );
not  ( new_n3958_, new_n3840_ );
or   ( new_n3959_, new_n3958_, new_n3834_ );
nand ( new_n3960_, new_n3959_, new_n3957_ );
and  ( new_n3961_, new_n3960_, new_n3955_ );
nor  ( new_n3962_, new_n3961_, new_n3954_ );
not  ( new_n3963_, new_n3962_ );
xor  ( new_n3964_, new_n3821_, new_n3804_ );
xor  ( new_n3965_, new_n3964_, new_n3841_ );
nand ( new_n3966_, new_n3965_, new_n3963_ );
xor  ( new_n3967_, new_n3965_, new_n3963_ );
xor  ( new_n3968_, new_n3866_, new_n3864_ );
xnor ( new_n3969_, new_n3968_, new_n3904_ );
nand ( new_n3970_, new_n3969_, new_n3967_ );
and  ( new_n3971_, new_n3970_, new_n3966_ );
xor  ( new_n3972_, new_n3911_, new_n3910_ );
nor  ( new_n3973_, new_n3972_, new_n3971_ );
and  ( new_n3974_, new_n3972_, new_n3971_ );
xnor ( new_n3975_, new_n3969_, new_n3967_ );
xnor ( new_n3976_, new_n3960_, new_n3955_ );
xor  ( new_n3977_, new_n3882_, new_n3869_ );
xor  ( new_n3978_, new_n3977_, new_n3902_ );
or   ( new_n3979_, new_n3978_, new_n3976_ );
and  ( new_n3980_, new_n3978_, new_n3976_ );
xor  ( new_n3981_, new_n3066_, new_n2856_ );
and  ( new_n3982_, new_n3981_, new_n3070_ );
and  ( new_n3983_, new_n3920_, new_n3068_ );
or   ( new_n3984_, new_n3983_, new_n3982_ );
xor  ( new_n3985_, new_n3929_, new_n3927_ );
and  ( new_n3986_, new_n3985_, new_n3984_ );
nor  ( new_n3987_, new_n3830_, new_n2559_ );
and  ( new_n3988_, new_n3889_, new_n2603_ );
nor  ( new_n3989_, new_n3988_, new_n3987_ );
not  ( new_n3990_, new_n3989_ );
xor  ( new_n3991_, new_n3985_, new_n3984_ );
and  ( new_n3992_, new_n3991_, new_n3990_ );
or   ( new_n3993_, new_n3992_, new_n3986_ );
xnor ( new_n3994_, new_n3874_, new_n3873_ );
xor  ( new_n3995_, new_n3994_, new_n3880_ );
or   ( new_n3996_, new_n3995_, new_n3993_ );
and  ( new_n3997_, new_n3995_, new_n3993_ );
xor  ( new_n3998_, new_n3892_, new_n3888_ );
or   ( new_n3999_, new_n3998_, new_n3900_ );
not  ( new_n4000_, new_n3901_ );
or   ( new_n4001_, new_n4000_, new_n3893_ );
and  ( new_n4002_, new_n4001_, new_n3999_ );
or   ( new_n4003_, new_n4002_, new_n3997_ );
and  ( new_n4004_, new_n4003_, new_n3996_ );
or   ( new_n4005_, new_n4004_, new_n3980_ );
and  ( new_n4006_, new_n4005_, new_n3979_ );
nor  ( new_n4007_, new_n4006_, new_n3975_ );
and  ( new_n4008_, new_n4006_, new_n3975_ );
xor  ( new_n4009_, new_n3995_, new_n3993_ );
xor  ( new_n4010_, new_n4009_, new_n4002_ );
xnor ( new_n4011_, new_n3930_, new_n3923_ );
xor  ( new_n4012_, new_n4011_, new_n3951_ );
or   ( new_n4013_, new_n4012_, new_n4010_ );
or   ( new_n4014_, new_n3928_, new_n2543_ );
xnor ( new_n4015_, new_n3230_, new_n2705_ );
or   ( new_n4016_, new_n4015_, new_n3488_ );
not  ( new_n4017_, new_n2723_ );
or   ( new_n4018_, new_n3554_, new_n4017_ );
and  ( new_n4019_, new_n4018_, new_n4016_ );
or   ( new_n4020_, new_n4019_, new_n4014_ );
and  ( new_n4021_, new_n4019_, new_n4014_ );
xor  ( new_n4022_, new_n3026_, new_n2923_ );
and  ( new_n4023_, new_n4022_, new_n3272_ );
and  ( new_n4024_, new_n3925_, new_n3374_ );
nor  ( new_n4025_, new_n4024_, new_n4023_ );
or   ( new_n4026_, new_n4025_, new_n4021_ );
and  ( new_n4027_, new_n4026_, new_n4020_ );
xor  ( new_n4028_, new_n3507_, new_n2542_ );
and  ( new_n4029_, new_n4028_, new_n2729_ );
and  ( new_n4030_, new_n3945_, new_n2781_ );
nor  ( new_n4031_, new_n4030_, new_n4029_ );
not  ( new_n4032_, new_n4031_ );
xor  ( new_n4033_, new_n3306_, new_n2692_ );
and  ( new_n4034_, new_n4033_, new_n2905_ );
and  ( new_n4035_, new_n3933_, new_n3033_ );
nor  ( new_n4036_, new_n4035_, new_n4034_ );
not  ( new_n4037_, new_n4036_ );
and  ( new_n4038_, new_n4037_, new_n4032_ );
and  ( new_n4039_, new_n4036_, new_n4031_ );
xor  ( new_n4040_, new_n3108_, new_n2856_ );
and  ( new_n4041_, new_n4040_, new_n3070_ );
and  ( new_n4042_, new_n3981_, new_n3068_ );
nor  ( new_n4043_, new_n4042_, new_n4041_ );
nor  ( new_n4044_, new_n4043_, new_n4039_ );
nor  ( new_n4045_, new_n4044_, new_n4038_ );
nor  ( new_n4046_, new_n4045_, new_n4027_ );
xor  ( new_n4047_, new_n3991_, new_n3990_ );
xor  ( new_n4048_, new_n4045_, new_n4027_ );
and  ( new_n4049_, new_n4048_, new_n4047_ );
nor  ( new_n4050_, new_n4049_, new_n4046_ );
nand ( new_n4051_, new_n4012_, new_n4010_ );
nand ( new_n4052_, new_n4051_, new_n4050_ );
and  ( new_n4053_, new_n4052_, new_n4013_ );
xor  ( new_n4054_, new_n3978_, new_n3976_ );
xor  ( new_n4055_, new_n4054_, new_n4004_ );
and  ( new_n4056_, new_n4055_, new_n4053_ );
nor  ( new_n4057_, new_n4055_, new_n4053_ );
xor  ( new_n4058_, new_n3942_, new_n3937_ );
and  ( new_n4059_, new_n4058_, new_n3948_ );
not  ( new_n4060_, new_n3944_ );
and  ( new_n4061_, new_n3950_, new_n4060_ );
or   ( new_n4062_, new_n4061_, new_n4059_ );
and  ( new_n4063_, new_n4022_, new_n3374_ );
xor  ( new_n4064_, new_n3066_, new_n3026_ );
and  ( new_n4065_, new_n4064_, new_n3272_ );
or   ( new_n4066_, new_n4065_, new_n4063_ );
nor  ( new_n4067_, new_n3548_, new_n2727_ );
nor  ( new_n4068_, new_n4067_, new_n2733_ );
and  ( new_n4069_, new_n4068_, new_n4066_ );
xnor ( new_n4070_, new_n4019_, new_n4014_ );
xor  ( new_n4071_, new_n4070_, new_n4025_ );
nand ( new_n4072_, new_n4071_, new_n4069_ );
nor  ( new_n4073_, new_n4071_, new_n4069_ );
xor  ( new_n4074_, new_n3406_, new_n2692_ );
nand ( new_n4075_, new_n4074_, new_n2905_ );
nand ( new_n4076_, new_n4033_, new_n3033_ );
and  ( new_n4077_, new_n4076_, new_n4075_ );
nand ( new_n4078_, new_n4028_, new_n2781_ );
xor  ( new_n4079_, new_n3547_, new_n2692_ );
not  ( new_n4080_, new_n4079_ );
or   ( new_n4081_, new_n4080_, new_n2730_ );
and  ( new_n4082_, new_n4081_, new_n4078_ );
or   ( new_n4083_, new_n4082_, new_n4077_ );
and  ( new_n4084_, new_n4082_, new_n4077_ );
not  ( new_n4085_, new_n2760_ );
nor  ( new_n4086_, new_n3230_, new_n4085_ );
and  ( new_n4087_, new_n4086_, new_n3488_ );
xor  ( new_n4088_, new_n3230_, new_n2723_ );
and  ( new_n4089_, new_n4088_, new_n3552_ );
nor  ( new_n4090_, new_n4089_, new_n4087_ );
or   ( new_n4091_, new_n4090_, new_n4084_ );
and  ( new_n4092_, new_n4091_, new_n4083_ );
or   ( new_n4093_, new_n4092_, new_n4073_ );
and  ( new_n4094_, new_n4093_, new_n4072_ );
or   ( new_n4095_, new_n4094_, new_n4062_ );
and  ( new_n4096_, new_n4094_, new_n4062_ );
xnor ( new_n4097_, new_n4048_, new_n4047_ );
or   ( new_n4098_, new_n4097_, new_n4096_ );
and  ( new_n4099_, new_n4098_, new_n4095_ );
xor  ( new_n4100_, new_n4012_, new_n4010_ );
xor  ( new_n4101_, new_n4100_, new_n4050_ );
nor  ( new_n4102_, new_n4101_, new_n4099_ );
and  ( new_n4103_, new_n4101_, new_n4099_ );
xor  ( new_n4104_, new_n4094_, new_n4062_ );
xor  ( new_n4105_, new_n4104_, new_n4097_ );
xor  ( new_n4106_, new_n4036_, new_n4032_ );
and  ( new_n4107_, new_n4106_, new_n4043_ );
not  ( new_n4108_, new_n4038_ );
and  ( new_n4109_, new_n4044_, new_n4108_ );
or   ( new_n4110_, new_n4109_, new_n4107_ );
xor  ( new_n4111_, new_n3244_, new_n2856_ );
and  ( new_n4112_, new_n4111_, new_n3070_ );
and  ( new_n4113_, new_n4040_, new_n3068_ );
or   ( new_n4114_, new_n4113_, new_n4112_ );
xor  ( new_n4115_, new_n4068_, new_n4066_ );
nand ( new_n4116_, new_n4115_, new_n4114_ );
nor  ( new_n4117_, new_n4115_, new_n4114_ );
xor  ( new_n4118_, new_n3108_, new_n3026_ );
and  ( new_n4119_, new_n4118_, new_n3272_ );
and  ( new_n4120_, new_n4064_, new_n3374_ );
or   ( new_n4121_, new_n4120_, new_n4119_ );
and  ( new_n4122_, new_n4067_, new_n2725_ );
and  ( new_n4123_, new_n4122_, new_n4121_ );
nor  ( new_n4124_, new_n4122_, new_n4121_ );
xor  ( new_n4125_, new_n3507_, new_n2692_ );
and  ( new_n4126_, new_n4125_, new_n2905_ );
and  ( new_n4127_, new_n4074_, new_n3033_ );
nor  ( new_n4128_, new_n4127_, new_n4126_ );
nor  ( new_n4129_, new_n4128_, new_n4124_ );
nor  ( new_n4130_, new_n4129_, new_n4123_ );
or   ( new_n4131_, new_n4130_, new_n4117_ );
and  ( new_n4132_, new_n4131_, new_n4116_ );
or   ( new_n4133_, new_n4132_, new_n4110_ );
and  ( new_n4134_, new_n4132_, new_n4110_ );
xor  ( new_n4135_, new_n4071_, new_n4069_ );
xor  ( new_n4136_, new_n4135_, new_n4092_ );
or   ( new_n4137_, new_n4136_, new_n4134_ );
and  ( new_n4138_, new_n4137_, new_n4133_ );
nor  ( new_n4139_, new_n4138_, new_n4105_ );
and  ( new_n4140_, new_n4138_, new_n4105_ );
xor  ( new_n4141_, new_n4082_, new_n4077_ );
xnor ( new_n4142_, new_n4141_, new_n4090_ );
not  ( new_n4143_, new_n2856_ );
xor  ( new_n4144_, new_n3306_, new_n4143_ );
or   ( new_n4145_, new_n4144_, new_n3142_ );
nand ( new_n4146_, new_n4111_, new_n3068_ );
and  ( new_n4147_, new_n4146_, new_n4145_ );
xnor ( new_n4148_, new_n3230_, new_n2760_ );
or   ( new_n4149_, new_n4148_, new_n3488_ );
or   ( new_n4150_, new_n3554_, new_n2924_ );
and  ( new_n4151_, new_n4150_, new_n4149_ );
or   ( new_n4152_, new_n4151_, new_n4147_ );
and  ( new_n4153_, new_n4151_, new_n4147_ );
xor  ( new_n4154_, new_n3244_, new_n3026_ );
and  ( new_n4155_, new_n4154_, new_n3272_ );
and  ( new_n4156_, new_n4118_, new_n3374_ );
or   ( new_n4157_, new_n4156_, new_n4155_ );
nand ( new_n4158_, new_n3547_, new_n2909_ );
and  ( new_n4159_, new_n4158_, new_n2858_ );
nand ( new_n4160_, new_n4159_, new_n4157_ );
or   ( new_n4161_, new_n4160_, new_n4153_ );
nand ( new_n4162_, new_n4161_, new_n4152_ );
nor  ( new_n4163_, new_n4162_, new_n4142_ );
xnor ( new_n4164_, new_n4162_, new_n4142_ );
xnor ( new_n4165_, new_n4115_, new_n4114_ );
xor  ( new_n4166_, new_n4165_, new_n4130_ );
nor  ( new_n4167_, new_n4166_, new_n4164_ );
or   ( new_n4168_, new_n4167_, new_n4163_ );
xor  ( new_n4169_, new_n4132_, new_n4110_ );
xor  ( new_n4170_, new_n4169_, new_n4136_ );
nor  ( new_n4171_, new_n4170_, new_n4168_ );
and  ( new_n4172_, new_n4170_, new_n4168_ );
xor  ( new_n4173_, new_n3406_, new_n2856_ );
nand ( new_n4174_, new_n4173_, new_n3070_ );
or   ( new_n4175_, new_n4144_, new_n3310_ );
and  ( new_n4176_, new_n4175_, new_n4174_ );
not  ( new_n4177_, new_n3066_ );
or   ( new_n4178_, new_n3230_, new_n4177_ );
or   ( new_n4179_, new_n4178_, new_n3552_ );
xnor ( new_n4180_, new_n3230_, new_n2923_ );
or   ( new_n4181_, new_n4180_, new_n3488_ );
and  ( new_n4182_, new_n4181_, new_n4179_ );
nor  ( new_n4183_, new_n4182_, new_n4176_ );
and  ( new_n4184_, new_n4080_, new_n2905_ );
and  ( new_n4185_, new_n4125_, new_n3033_ );
nor  ( new_n4186_, new_n4185_, new_n4184_ );
not  ( new_n4187_, new_n4186_ );
xor  ( new_n4188_, new_n4182_, new_n4176_ );
and  ( new_n4189_, new_n4188_, new_n4187_ );
nor  ( new_n4190_, new_n4189_, new_n4183_ );
xnor ( new_n4191_, new_n4122_, new_n4121_ );
xnor ( new_n4192_, new_n4191_, new_n4128_ );
or   ( new_n4193_, new_n4192_, new_n4190_ );
xnor ( new_n4194_, new_n4192_, new_n4190_ );
xor  ( new_n4195_, new_n4151_, new_n4147_ );
xor  ( new_n4196_, new_n4195_, new_n4160_ );
or   ( new_n4197_, new_n4196_, new_n4194_ );
and  ( new_n4198_, new_n4197_, new_n4193_ );
xor  ( new_n4199_, new_n4166_, new_n4164_ );
nor  ( new_n4200_, new_n4199_, new_n4198_ );
and  ( new_n4201_, new_n4199_, new_n4198_ );
or   ( new_n4202_, new_n4158_, new_n2857_ );
xnor ( new_n4203_, new_n3230_, new_n3066_ );
or   ( new_n4204_, new_n4203_, new_n3488_ );
or   ( new_n4205_, new_n3554_, new_n3109_ );
and  ( new_n4206_, new_n4205_, new_n4204_ );
nor  ( new_n4207_, new_n4206_, new_n4202_ );
xor  ( new_n4208_, new_n3306_, new_n3026_ );
and  ( new_n4209_, new_n4208_, new_n3272_ );
and  ( new_n4210_, new_n4154_, new_n3374_ );
nor  ( new_n4211_, new_n4210_, new_n4209_ );
not  ( new_n4212_, new_n4211_ );
xor  ( new_n4213_, new_n4206_, new_n4202_ );
and  ( new_n4214_, new_n4213_, new_n4212_ );
or   ( new_n4215_, new_n4214_, new_n4207_ );
xor  ( new_n4216_, new_n4159_, new_n4157_ );
and  ( new_n4217_, new_n4216_, new_n4215_ );
xor  ( new_n4218_, new_n4188_, new_n4187_ );
xor  ( new_n4219_, new_n4216_, new_n4215_ );
and  ( new_n4220_, new_n4219_, new_n4218_ );
or   ( new_n4221_, new_n4220_, new_n4217_ );
xor  ( new_n4222_, new_n4196_, new_n4194_ );
and  ( new_n4223_, new_n4222_, new_n4221_ );
nor  ( new_n4224_, new_n4222_, new_n4221_ );
xor  ( new_n4225_, new_n4219_, new_n4218_ );
not  ( new_n4226_, new_n4225_ );
xor  ( new_n4227_, new_n3507_, new_n2856_ );
and  ( new_n4228_, new_n4227_, new_n3070_ );
and  ( new_n4229_, new_n4173_, new_n3068_ );
or   ( new_n4230_, new_n4229_, new_n4228_ );
xor  ( new_n4231_, new_n3406_, new_n3026_ );
and  ( new_n4232_, new_n4231_, new_n3272_ );
and  ( new_n4233_, new_n4208_, new_n3374_ );
or   ( new_n4234_, new_n4233_, new_n4232_ );
not  ( new_n4235_, new_n3028_ );
and  ( new_n4236_, new_n3547_, new_n3074_ );
nor  ( new_n4237_, new_n4236_, new_n4235_ );
and  ( new_n4238_, new_n4237_, new_n4234_ );
nand ( new_n4239_, new_n4238_, new_n4230_ );
or   ( new_n4240_, new_n4238_, new_n4230_ );
xor  ( new_n4241_, new_n4213_, new_n4212_ );
nand ( new_n4242_, new_n4241_, new_n4240_ );
and  ( new_n4243_, new_n4242_, new_n4239_ );
nor  ( new_n4244_, new_n4243_, new_n4226_ );
xor  ( new_n4245_, new_n4243_, new_n4226_ );
not  ( new_n4246_, new_n4245_ );
nand ( new_n4247_, new_n4227_, new_n3068_ );
or   ( new_n4248_, new_n2978_, new_n4143_ );
not  ( new_n4249_, new_n3026_ );
or   ( new_n4250_, new_n3547_, new_n4249_ );
and  ( new_n4251_, new_n4250_, new_n4248_ );
nand ( new_n4252_, new_n2978_, new_n4143_ );
or   ( new_n4253_, new_n3548_, new_n3026_ );
and  ( new_n4254_, new_n4253_, new_n4252_ );
or   ( new_n4255_, new_n4254_, new_n4251_ );
and  ( new_n4256_, new_n4255_, new_n4247_ );
not  ( new_n4257_, new_n3244_ );
or   ( new_n4258_, new_n3554_, new_n4257_ );
xnor ( new_n4259_, new_n3230_, new_n3108_ );
or   ( new_n4260_, new_n4259_, new_n3488_ );
and  ( new_n4261_, new_n4260_, new_n4258_ );
nor  ( new_n4262_, new_n4261_, new_n4256_ );
nand ( new_n4263_, new_n4261_, new_n4256_ );
xor  ( new_n4264_, new_n4237_, new_n4234_ );
and  ( new_n4265_, new_n4264_, new_n4263_ );
or   ( new_n4266_, new_n4265_, new_n4262_ );
xor  ( new_n4267_, new_n4238_, new_n4230_ );
xor  ( new_n4268_, new_n4267_, new_n4241_ );
nand ( new_n4269_, new_n4268_, new_n4266_ );
nor  ( new_n4270_, new_n4268_, new_n4266_ );
not  ( new_n4271_, new_n3027_ );
and  ( new_n4272_, new_n4236_, new_n4271_ );
or   ( new_n4273_, new_n3490_, new_n3244_ );
and  ( new_n4274_, new_n3552_, new_n4257_ );
not  ( new_n4275_, new_n3306_ );
nor  ( new_n4276_, new_n4275_, new_n3230_ );
or   ( new_n4277_, new_n4276_, new_n3489_ );
or   ( new_n4278_, new_n4277_, new_n4274_ );
and  ( new_n4279_, new_n4278_, new_n4273_ );
or   ( new_n4280_, new_n4279_, new_n4272_ );
xor  ( new_n4281_, new_n3507_, new_n3026_ );
and  ( new_n4282_, new_n4281_, new_n3272_ );
and  ( new_n4283_, new_n4231_, new_n3374_ );
or   ( new_n4284_, new_n4283_, new_n4282_ );
and  ( new_n4285_, new_n4279_, new_n4272_ );
or   ( new_n4286_, new_n4285_, new_n4284_ );
and  ( new_n4287_, new_n4286_, new_n4280_ );
xor  ( new_n4288_, new_n4261_, new_n4256_ );
xor  ( new_n4289_, new_n4288_, new_n4264_ );
and  ( new_n4290_, new_n4289_, new_n4287_ );
nor  ( new_n4291_, new_n4289_, new_n4287_ );
and  ( new_n4292_, new_n4281_, new_n3374_ );
xor  ( new_n4293_, new_n3547_, new_n4249_ );
and  ( new_n4294_, new_n4293_, new_n3272_ );
or   ( new_n4295_, new_n4294_, new_n4292_ );
not  ( new_n4296_, new_n3232_ );
and  ( new_n4297_, new_n3547_, new_n3275_ );
nor  ( new_n4298_, new_n4297_, new_n4296_ );
and  ( new_n4299_, new_n4298_, new_n4295_ );
xor  ( new_n4300_, new_n4279_, new_n4272_ );
xor  ( new_n4301_, new_n4300_, new_n4284_ );
and  ( new_n4302_, new_n4301_, new_n4299_ );
nor  ( new_n4303_, new_n4301_, new_n4299_ );
and  ( new_n4304_, new_n3553_, new_n3507_ );
xor  ( new_n4305_, new_n3406_, new_n3230_ );
and  ( new_n4306_, new_n4305_, new_n3552_ );
or   ( new_n4307_, new_n4306_, new_n4304_ );
and  ( new_n4308_, new_n4297_, new_n3268_ );
nor  ( new_n4309_, new_n4308_, new_n4307_ );
and  ( new_n4310_, new_n4308_, new_n4307_ );
not  ( new_n4311_, new_n3507_ );
and  ( new_n4312_, new_n4311_, new_n3552_ );
not  ( new_n4313_, new_n4312_ );
nor  ( new_n4314_, new_n3547_, new_n3230_ );
and  ( new_n4315_, new_n4314_, new_n4313_ );
nor  ( new_n4316_, new_n4315_, new_n4310_ );
nor  ( new_n4317_, new_n4316_, new_n4309_ );
not  ( new_n4318_, new_n4317_ );
xnor ( new_n4319_, new_n3306_, new_n3230_ );
or   ( new_n4320_, new_n4319_, new_n3488_ );
or   ( new_n4321_, new_n3554_, new_n3407_ );
and  ( new_n4322_, new_n4321_, new_n4320_ );
nor  ( new_n4323_, new_n4322_, new_n4318_ );
xor  ( new_n4324_, new_n4322_, new_n4318_ );
xor  ( new_n4325_, new_n4298_, new_n4295_ );
and  ( new_n4326_, new_n4325_, new_n4324_ );
nor  ( new_n4327_, new_n4326_, new_n4323_ );
nor  ( new_n4328_, new_n4327_, new_n4303_ );
nor  ( new_n4329_, new_n4328_, new_n4302_ );
nor  ( new_n4330_, new_n4329_, new_n4291_ );
nor  ( new_n4331_, new_n4330_, new_n4290_ );
or   ( new_n4332_, new_n4331_, new_n4270_ );
and  ( new_n4333_, new_n4332_, new_n4269_ );
nor  ( new_n4334_, new_n4333_, new_n4246_ );
nor  ( new_n4335_, new_n4334_, new_n4244_ );
nor  ( new_n4336_, new_n4335_, new_n4224_ );
nor  ( new_n4337_, new_n4336_, new_n4223_ );
nor  ( new_n4338_, new_n4337_, new_n4201_ );
nor  ( new_n4339_, new_n4338_, new_n4200_ );
nor  ( new_n4340_, new_n4339_, new_n4172_ );
nor  ( new_n4341_, new_n4340_, new_n4171_ );
nor  ( new_n4342_, new_n4341_, new_n4140_ );
nor  ( new_n4343_, new_n4342_, new_n4139_ );
nor  ( new_n4344_, new_n4343_, new_n4103_ );
nor  ( new_n4345_, new_n4344_, new_n4102_ );
nor  ( new_n4346_, new_n4345_, new_n4057_ );
nor  ( new_n4347_, new_n4346_, new_n4056_ );
not  ( new_n4348_, new_n4347_ );
nor  ( new_n4349_, new_n4348_, new_n4008_ );
nor  ( new_n4350_, new_n4349_, new_n4007_ );
nor  ( new_n4351_, new_n4350_, new_n3974_ );
nor  ( new_n4352_, new_n4351_, new_n3973_ );
nor  ( new_n4353_, new_n4352_, new_n3916_ );
nor  ( new_n4354_, new_n4353_, new_n3915_ );
nor  ( new_n4355_, new_n4354_, new_n3862_ );
nor  ( new_n4356_, new_n4355_, new_n3861_ );
not  ( new_n4357_, new_n4356_ );
nor  ( new_n4358_, new_n4357_, new_n3803_ );
nor  ( new_n4359_, new_n4358_, new_n3802_ );
not  ( new_n4360_, new_n4359_ );
nor  ( new_n4361_, new_n4360_, new_n3721_ );
nor  ( new_n4362_, new_n4361_, new_n3720_ );
nor  ( new_n4363_, new_n4362_, new_n3644_ );
nor  ( new_n4364_, new_n4363_, new_n3643_ );
nor  ( new_n4365_, new_n4364_, new_n3612_ );
nor  ( new_n4366_, new_n4365_, new_n3611_ );
nor  ( new_n4367_, new_n4366_, new_n3447_ );
nor  ( new_n4368_, new_n4367_, new_n3446_ );
nor  ( new_n4369_, new_n4368_, new_n3356_ );
nor  ( new_n4370_, new_n4369_, new_n3355_ );
not  ( new_n4371_, new_n4370_ );
nor  ( new_n4372_, new_n4371_, new_n3298_ );
nor  ( new_n4373_, new_n4372_, new_n3297_ );
nor  ( new_n4374_, new_n4373_, new_n3132_ );
nor  ( new_n4375_, new_n4374_, new_n3131_ );
not  ( new_n4376_, new_n4375_ );
nor  ( new_n4377_, new_n4376_, new_n2940_ );
nor  ( new_n4378_, new_n4377_, new_n2939_ );
nor  ( new_n4379_, new_n4378_, new_n2882_ );
nor  ( new_n4380_, new_n4379_, new_n2881_ );
not  ( new_n4381_, new_n4380_ );
nor  ( new_n4382_, new_n4381_, new_n2754_ );
nor  ( new_n4383_, new_n4382_, new_n2753_ );
nor  ( new_n4384_, new_n4383_, new_n2702_ );
nor  ( new_n4385_, new_n4384_, new_n2701_ );
or   ( new_n4386_, new_n4385_, new_n2588_ );
and  ( new_n4387_, new_n4386_, new_n2587_ );
xnor ( new_n4388_, new_n4387_, new_n2438_ );
and  ( new_n4389_, \b[14] , \a[0]  );
and  ( new_n4390_, \b[13] , \a[0]  );
and  ( new_n4391_, \b[12] , \a[0]  );
and  ( new_n4392_, \b[11] , \a[0]  );
and  ( new_n4393_, \b[9] , \a[0]  );
and  ( new_n4394_, \b[8] , \a[0]  );
and  ( new_n4395_, \b[6] , \a[0]  );
and  ( new_n4396_, \b[4] , \a[0]  );
and  ( new_n4397_, new_n2063_, new_n897_ );
and  ( new_n4398_, \b[1] , \a[1]  );
and  ( new_n4399_, \b[0] , \a[2]  );
and  ( new_n4400_, new_n4399_, new_n4398_ );
nand ( new_n4401_, new_n4400_, new_n4397_ );
nor  ( new_n4402_, new_n4399_, new_n4398_ );
or   ( new_n4403_, new_n4400_, new_n4397_ );
or   ( new_n4404_, new_n4403_, new_n4402_ );
and  ( new_n4405_, new_n4404_, new_n4401_ );
nor  ( new_n4406_, new_n4405_, new_n880_ );
and  ( new_n4407_, \b[2] , \a[1]  );
and  ( new_n4408_, \b[0] , \a[3]  );
xor  ( new_n4409_, new_n4408_, new_n891_ );
xor  ( new_n4410_, new_n4409_, new_n4403_ );
xor  ( new_n4411_, new_n4410_, new_n4407_ );
xor  ( new_n4412_, new_n4411_, new_n4406_ );
and  ( new_n4413_, new_n4412_, new_n882_ );
and  ( new_n4414_, \b[3] , \a[1]  );
and  ( new_n4415_, new_n4410_, new_n4407_ );
and  ( new_n4416_, new_n4411_, new_n4406_ );
or   ( new_n4417_, new_n4416_, new_n4415_ );
and  ( new_n4418_, \b[2] , \a[2]  );
and  ( new_n4419_, new_n4408_, new_n891_ );
and  ( new_n4420_, new_n4409_, new_n4403_ );
or   ( new_n4421_, new_n4420_, new_n4419_ );
and  ( new_n4422_, \b[0] , \a[4]  );
xor  ( new_n4423_, new_n4422_, new_n861_ );
xor  ( new_n4424_, new_n4423_, new_n4421_ );
xor  ( new_n4425_, new_n4424_, new_n4418_ );
xor  ( new_n4426_, new_n4425_, new_n4417_ );
xor  ( new_n4427_, new_n4426_, new_n4414_ );
xor  ( new_n4428_, new_n4427_, new_n4413_ );
and  ( new_n4429_, new_n4428_, new_n4396_ );
and  ( new_n4430_, \b[4] , \a[1]  );
and  ( new_n4431_, new_n4426_, new_n4414_ );
and  ( new_n4432_, new_n4427_, new_n4413_ );
or   ( new_n4433_, new_n4432_, new_n4431_ );
and  ( new_n4434_, \b[3] , \a[2]  );
and  ( new_n4435_, new_n4424_, new_n4418_ );
and  ( new_n4436_, new_n4425_, new_n4417_ );
or   ( new_n4437_, new_n4436_, new_n4435_ );
and  ( new_n4438_, \b[2] , \a[3]  );
and  ( new_n4439_, new_n4422_, new_n861_ );
and  ( new_n4440_, new_n4423_, new_n4421_ );
or   ( new_n4441_, new_n4440_, new_n4439_ );
and  ( new_n4442_, \b[0] , \a[5]  );
xor  ( new_n4443_, new_n4442_, new_n810_ );
xor  ( new_n4444_, new_n4443_, new_n4441_ );
xor  ( new_n4445_, new_n4444_, new_n4438_ );
xor  ( new_n4446_, new_n4445_, new_n4437_ );
xor  ( new_n4447_, new_n4446_, new_n4434_ );
xor  ( new_n4448_, new_n4447_, new_n4433_ );
xor  ( new_n4449_, new_n4448_, new_n4430_ );
xor  ( new_n4450_, new_n4449_, new_n4429_ );
and  ( new_n4451_, new_n4450_, new_n1696_ );
and  ( new_n4452_, \b[5] , \a[1]  );
and  ( new_n4453_, new_n4448_, new_n4430_ );
and  ( new_n4454_, new_n4449_, new_n4429_ );
or   ( new_n4455_, new_n4454_, new_n4453_ );
and  ( new_n4456_, \b[4] , \a[2]  );
and  ( new_n4457_, new_n4446_, new_n4434_ );
and  ( new_n4458_, new_n4447_, new_n4433_ );
or   ( new_n4459_, new_n4458_, new_n4457_ );
and  ( new_n4460_, \b[3] , \a[3]  );
and  ( new_n4461_, new_n4444_, new_n4438_ );
and  ( new_n4462_, new_n4445_, new_n4437_ );
or   ( new_n4463_, new_n4462_, new_n4461_ );
and  ( new_n4464_, \b[2] , \a[4]  );
and  ( new_n4465_, new_n4442_, new_n810_ );
and  ( new_n4466_, new_n4443_, new_n4441_ );
or   ( new_n4467_, new_n4466_, new_n4465_ );
and  ( new_n4468_, \b[0] , \a[6]  );
xor  ( new_n4469_, new_n4468_, new_n841_ );
xor  ( new_n4470_, new_n4469_, new_n4467_ );
xor  ( new_n4471_, new_n4470_, new_n4464_ );
xor  ( new_n4472_, new_n4471_, new_n4463_ );
xor  ( new_n4473_, new_n4472_, new_n4460_ );
xor  ( new_n4474_, new_n4473_, new_n4459_ );
xor  ( new_n4475_, new_n4474_, new_n4456_ );
xor  ( new_n4476_, new_n4475_, new_n4455_ );
xor  ( new_n4477_, new_n4476_, new_n4452_ );
xor  ( new_n4478_, new_n4477_, new_n4451_ );
and  ( new_n4479_, new_n4478_, new_n4395_ );
and  ( new_n4480_, \b[6] , \a[1]  );
and  ( new_n4481_, new_n4476_, new_n4452_ );
and  ( new_n4482_, new_n4477_, new_n4451_ );
or   ( new_n4483_, new_n4482_, new_n4481_ );
and  ( new_n4484_, \b[5] , \a[2]  );
and  ( new_n4485_, new_n4474_, new_n4456_ );
and  ( new_n4486_, new_n4475_, new_n4455_ );
or   ( new_n4487_, new_n4486_, new_n4485_ );
and  ( new_n4488_, \b[4] , \a[3]  );
and  ( new_n4489_, new_n4472_, new_n4460_ );
and  ( new_n4490_, new_n4473_, new_n4459_ );
or   ( new_n4491_, new_n4490_, new_n4489_ );
and  ( new_n4492_, \b[3] , \a[4]  );
and  ( new_n4493_, new_n4470_, new_n4464_ );
and  ( new_n4494_, new_n4471_, new_n4463_ );
or   ( new_n4495_, new_n4494_, new_n4493_ );
and  ( new_n4496_, \b[2] , \a[5]  );
and  ( new_n4497_, new_n4468_, new_n841_ );
and  ( new_n4498_, new_n4469_, new_n4467_ );
or   ( new_n4499_, new_n4498_, new_n4497_ );
and  ( new_n4500_, \b[0] , \a[7]  );
xor  ( new_n4501_, new_n4500_, new_n930_ );
xor  ( new_n4502_, new_n4501_, new_n4499_ );
xor  ( new_n4503_, new_n4502_, new_n4496_ );
xor  ( new_n4504_, new_n4503_, new_n4495_ );
xor  ( new_n4505_, new_n4504_, new_n4492_ );
xor  ( new_n4506_, new_n4505_, new_n4491_ );
xor  ( new_n4507_, new_n4506_, new_n4488_ );
xor  ( new_n4508_, new_n4507_, new_n4487_ );
xor  ( new_n4509_, new_n4508_, new_n4484_ );
xor  ( new_n4510_, new_n4509_, new_n4483_ );
xor  ( new_n4511_, new_n4510_, new_n4480_ );
xor  ( new_n4512_, new_n4511_, new_n4479_ );
and  ( new_n4513_, new_n4512_, new_n1896_ );
and  ( new_n4514_, \b[7] , \a[1]  );
and  ( new_n4515_, new_n4510_, new_n4480_ );
and  ( new_n4516_, new_n4511_, new_n4479_ );
or   ( new_n4517_, new_n4516_, new_n4515_ );
and  ( new_n4518_, \b[6] , \a[2]  );
and  ( new_n4519_, new_n4508_, new_n4484_ );
and  ( new_n4520_, new_n4509_, new_n4483_ );
or   ( new_n4521_, new_n4520_, new_n4519_ );
and  ( new_n4522_, \b[5] , \a[3]  );
and  ( new_n4523_, new_n4506_, new_n4488_ );
and  ( new_n4524_, new_n4507_, new_n4487_ );
or   ( new_n4525_, new_n4524_, new_n4523_ );
and  ( new_n4526_, \b[4] , \a[4]  );
and  ( new_n4527_, new_n4504_, new_n4492_ );
and  ( new_n4528_, new_n4505_, new_n4491_ );
or   ( new_n4529_, new_n4528_, new_n4527_ );
and  ( new_n4530_, \b[3] , \a[5]  );
and  ( new_n4531_, new_n4502_, new_n4496_ );
and  ( new_n4532_, new_n4503_, new_n4495_ );
or   ( new_n4533_, new_n4532_, new_n4531_ );
and  ( new_n4534_, \b[2] , \a[6]  );
and  ( new_n4535_, new_n4500_, new_n930_ );
and  ( new_n4536_, new_n4501_, new_n4499_ );
or   ( new_n4537_, new_n4536_, new_n4535_ );
and  ( new_n4538_, \b[0] , \a[8]  );
xor  ( new_n4539_, new_n4538_, new_n1681_ );
xor  ( new_n4540_, new_n4539_, new_n4537_ );
xor  ( new_n4541_, new_n4540_, new_n4534_ );
xor  ( new_n4542_, new_n4541_, new_n4533_ );
xor  ( new_n4543_, new_n4542_, new_n4530_ );
xor  ( new_n4544_, new_n4543_, new_n4529_ );
xor  ( new_n4545_, new_n4544_, new_n4526_ );
xor  ( new_n4546_, new_n4545_, new_n4525_ );
xor  ( new_n4547_, new_n4546_, new_n4522_ );
xor  ( new_n4548_, new_n4547_, new_n4521_ );
xor  ( new_n4549_, new_n4548_, new_n4518_ );
xor  ( new_n4550_, new_n4549_, new_n4517_ );
xor  ( new_n4551_, new_n4550_, new_n4514_ );
xor  ( new_n4552_, new_n4551_, new_n4513_ );
and  ( new_n4553_, new_n4552_, new_n4394_ );
and  ( new_n4554_, \b[8] , \a[1]  );
and  ( new_n4555_, new_n4550_, new_n4514_ );
and  ( new_n4556_, new_n4551_, new_n4513_ );
or   ( new_n4557_, new_n4556_, new_n4555_ );
and  ( new_n4558_, \b[7] , \a[2]  );
and  ( new_n4559_, new_n4548_, new_n4518_ );
and  ( new_n4560_, new_n4549_, new_n4517_ );
or   ( new_n4561_, new_n4560_, new_n4559_ );
and  ( new_n4562_, \b[6] , \a[3]  );
and  ( new_n4563_, new_n4546_, new_n4522_ );
and  ( new_n4564_, new_n4547_, new_n4521_ );
or   ( new_n4565_, new_n4564_, new_n4563_ );
and  ( new_n4566_, \b[5] , \a[4]  );
and  ( new_n4567_, new_n4544_, new_n4526_ );
and  ( new_n4568_, new_n4545_, new_n4525_ );
or   ( new_n4569_, new_n4568_, new_n4567_ );
and  ( new_n4570_, \b[4] , \a[5]  );
and  ( new_n4571_, new_n4542_, new_n4530_ );
and  ( new_n4572_, new_n4543_, new_n4529_ );
or   ( new_n4573_, new_n4572_, new_n4571_ );
and  ( new_n4574_, \b[3] , \a[6]  );
and  ( new_n4575_, new_n4540_, new_n4534_ );
and  ( new_n4576_, new_n4541_, new_n4533_ );
or   ( new_n4577_, new_n4576_, new_n4575_ );
and  ( new_n4578_, \b[2] , \a[7]  );
and  ( new_n4579_, new_n4538_, new_n1681_ );
and  ( new_n4580_, new_n4539_, new_n4537_ );
or   ( new_n4581_, new_n4580_, new_n4579_ );
and  ( new_n4582_, \b[0] , \a[9]  );
xor  ( new_n4583_, new_n4582_, new_n1872_ );
xor  ( new_n4584_, new_n4583_, new_n4581_ );
xor  ( new_n4585_, new_n4584_, new_n4578_ );
xor  ( new_n4586_, new_n4585_, new_n4577_ );
xor  ( new_n4587_, new_n4586_, new_n4574_ );
xor  ( new_n4588_, new_n4587_, new_n4573_ );
xor  ( new_n4589_, new_n4588_, new_n4570_ );
xor  ( new_n4590_, new_n4589_, new_n4569_ );
xor  ( new_n4591_, new_n4590_, new_n4566_ );
xor  ( new_n4592_, new_n4591_, new_n4565_ );
xor  ( new_n4593_, new_n4592_, new_n4562_ );
xor  ( new_n4594_, new_n4593_, new_n4561_ );
xor  ( new_n4595_, new_n4594_, new_n4558_ );
xor  ( new_n4596_, new_n4595_, new_n4557_ );
xor  ( new_n4597_, new_n4596_, new_n4554_ );
xor  ( new_n4598_, new_n4597_, new_n4553_ );
and  ( new_n4599_, new_n4598_, new_n4393_ );
and  ( new_n4600_, \b[9] , \a[1]  );
and  ( new_n4601_, new_n4596_, new_n4554_ );
and  ( new_n4602_, new_n4597_, new_n4553_ );
or   ( new_n4603_, new_n4602_, new_n4601_ );
and  ( new_n4604_, \b[8] , \a[2]  );
and  ( new_n4605_, new_n4594_, new_n4558_ );
and  ( new_n4606_, new_n4595_, new_n4557_ );
or   ( new_n4607_, new_n4606_, new_n4605_ );
and  ( new_n4608_, \b[7] , \a[3]  );
and  ( new_n4609_, new_n4592_, new_n4562_ );
and  ( new_n4610_, new_n4593_, new_n4561_ );
or   ( new_n4611_, new_n4610_, new_n4609_ );
and  ( new_n4612_, \b[6] , \a[4]  );
and  ( new_n4613_, new_n4590_, new_n4566_ );
and  ( new_n4614_, new_n4591_, new_n4565_ );
or   ( new_n4615_, new_n4614_, new_n4613_ );
and  ( new_n4616_, \b[5] , \a[5]  );
and  ( new_n4617_, new_n4588_, new_n4570_ );
and  ( new_n4618_, new_n4589_, new_n4569_ );
or   ( new_n4619_, new_n4618_, new_n4617_ );
and  ( new_n4620_, \b[4] , \a[6]  );
and  ( new_n4621_, new_n4586_, new_n4574_ );
and  ( new_n4622_, new_n4587_, new_n4573_ );
or   ( new_n4623_, new_n4622_, new_n4621_ );
and  ( new_n4624_, \b[3] , \a[7]  );
and  ( new_n4625_, new_n4584_, new_n4578_ );
and  ( new_n4626_, new_n4585_, new_n4577_ );
or   ( new_n4627_, new_n4626_, new_n4625_ );
and  ( new_n4628_, \b[2] , \a[8]  );
and  ( new_n4629_, new_n4582_, new_n1872_ );
and  ( new_n4630_, new_n4583_, new_n4581_ );
or   ( new_n4631_, new_n4630_, new_n4629_ );
and  ( new_n4632_, \b[0] , \a[10]  );
xor  ( new_n4633_, new_n4632_, new_n1862_ );
xor  ( new_n4634_, new_n4633_, new_n4631_ );
xor  ( new_n4635_, new_n4634_, new_n4628_ );
xor  ( new_n4636_, new_n4635_, new_n4627_ );
xor  ( new_n4637_, new_n4636_, new_n4624_ );
xor  ( new_n4638_, new_n4637_, new_n4623_ );
xor  ( new_n4639_, new_n4638_, new_n4620_ );
xor  ( new_n4640_, new_n4639_, new_n4619_ );
xor  ( new_n4641_, new_n4640_, new_n4616_ );
xor  ( new_n4642_, new_n4641_, new_n4615_ );
xor  ( new_n4643_, new_n4642_, new_n4612_ );
xor  ( new_n4644_, new_n4643_, new_n4611_ );
xor  ( new_n4645_, new_n4644_, new_n4608_ );
xor  ( new_n4646_, new_n4645_, new_n4607_ );
xor  ( new_n4647_, new_n4646_, new_n4604_ );
xor  ( new_n4648_, new_n4647_, new_n4603_ );
xor  ( new_n4649_, new_n4648_, new_n4600_ );
xor  ( new_n4650_, new_n4649_, new_n4599_ );
and  ( new_n4651_, new_n4650_, new_n2012_ );
and  ( new_n4652_, \b[10] , \a[1]  );
and  ( new_n4653_, new_n4648_, new_n4600_ );
and  ( new_n4654_, new_n4649_, new_n4599_ );
or   ( new_n4655_, new_n4654_, new_n4653_ );
and  ( new_n4656_, \b[9] , \a[2]  );
and  ( new_n4657_, new_n4646_, new_n4604_ );
and  ( new_n4658_, new_n4647_, new_n4603_ );
or   ( new_n4659_, new_n4658_, new_n4657_ );
and  ( new_n4660_, \b[8] , \a[3]  );
and  ( new_n4661_, new_n4644_, new_n4608_ );
and  ( new_n4662_, new_n4645_, new_n4607_ );
or   ( new_n4663_, new_n4662_, new_n4661_ );
and  ( new_n4664_, \b[7] , \a[4]  );
and  ( new_n4665_, new_n4642_, new_n4612_ );
and  ( new_n4666_, new_n4643_, new_n4611_ );
or   ( new_n4667_, new_n4666_, new_n4665_ );
and  ( new_n4668_, \b[6] , \a[5]  );
and  ( new_n4669_, new_n4640_, new_n4616_ );
and  ( new_n4670_, new_n4641_, new_n4615_ );
or   ( new_n4671_, new_n4670_, new_n4669_ );
and  ( new_n4672_, \b[5] , \a[6]  );
and  ( new_n4673_, new_n4638_, new_n4620_ );
and  ( new_n4674_, new_n4639_, new_n4619_ );
or   ( new_n4675_, new_n4674_, new_n4673_ );
and  ( new_n4676_, \b[4] , \a[7]  );
and  ( new_n4677_, new_n4636_, new_n4624_ );
and  ( new_n4678_, new_n4637_, new_n4623_ );
or   ( new_n4679_, new_n4678_, new_n4677_ );
and  ( new_n4680_, \b[3] , \a[8]  );
and  ( new_n4681_, new_n4634_, new_n4628_ );
and  ( new_n4682_, new_n4635_, new_n4627_ );
or   ( new_n4683_, new_n4682_, new_n4681_ );
and  ( new_n4684_, \b[2] , \a[9]  );
and  ( new_n4685_, new_n4632_, new_n1862_ );
and  ( new_n4686_, new_n4633_, new_n4631_ );
or   ( new_n4687_, new_n4686_, new_n4685_ );
and  ( new_n4688_, \b[0] , \a[11]  );
xor  ( new_n4689_, new_n4688_, new_n1947_ );
xor  ( new_n4690_, new_n4689_, new_n4687_ );
xor  ( new_n4691_, new_n4690_, new_n4684_ );
xor  ( new_n4692_, new_n4691_, new_n4683_ );
xor  ( new_n4693_, new_n4692_, new_n4680_ );
xor  ( new_n4694_, new_n4693_, new_n4679_ );
xor  ( new_n4695_, new_n4694_, new_n4676_ );
xor  ( new_n4696_, new_n4695_, new_n4675_ );
xor  ( new_n4697_, new_n4696_, new_n4672_ );
xor  ( new_n4698_, new_n4697_, new_n4671_ );
xor  ( new_n4699_, new_n4698_, new_n4668_ );
xor  ( new_n4700_, new_n4699_, new_n4667_ );
xor  ( new_n4701_, new_n4700_, new_n4664_ );
xor  ( new_n4702_, new_n4701_, new_n4663_ );
xor  ( new_n4703_, new_n4702_, new_n4660_ );
xor  ( new_n4704_, new_n4703_, new_n4659_ );
xor  ( new_n4705_, new_n4704_, new_n4656_ );
xor  ( new_n4706_, new_n4705_, new_n4655_ );
xor  ( new_n4707_, new_n4706_, new_n4652_ );
xor  ( new_n4708_, new_n4707_, new_n4651_ );
and  ( new_n4709_, new_n4708_, new_n4392_ );
and  ( new_n4710_, \b[11] , \a[1]  );
and  ( new_n4711_, new_n4706_, new_n4652_ );
and  ( new_n4712_, new_n4707_, new_n4651_ );
or   ( new_n4713_, new_n4712_, new_n4711_ );
and  ( new_n4714_, \b[10] , \a[2]  );
and  ( new_n4715_, new_n4704_, new_n4656_ );
and  ( new_n4716_, new_n4705_, new_n4655_ );
or   ( new_n4717_, new_n4716_, new_n4715_ );
and  ( new_n4718_, \b[9] , \a[3]  );
and  ( new_n4719_, new_n4702_, new_n4660_ );
and  ( new_n4720_, new_n4703_, new_n4659_ );
or   ( new_n4721_, new_n4720_, new_n4719_ );
and  ( new_n4722_, \b[8] , \a[4]  );
and  ( new_n4723_, new_n4700_, new_n4664_ );
and  ( new_n4724_, new_n4701_, new_n4663_ );
or   ( new_n4725_, new_n4724_, new_n4723_ );
and  ( new_n4726_, \b[7] , \a[5]  );
and  ( new_n4727_, new_n4698_, new_n4668_ );
and  ( new_n4728_, new_n4699_, new_n4667_ );
or   ( new_n4729_, new_n4728_, new_n4727_ );
and  ( new_n4730_, \b[6] , \a[6]  );
and  ( new_n4731_, new_n4696_, new_n4672_ );
and  ( new_n4732_, new_n4697_, new_n4671_ );
or   ( new_n4733_, new_n4732_, new_n4731_ );
and  ( new_n4734_, \b[5] , \a[7]  );
and  ( new_n4735_, new_n4694_, new_n4676_ );
and  ( new_n4736_, new_n4695_, new_n4675_ );
or   ( new_n4737_, new_n4736_, new_n4735_ );
and  ( new_n4738_, \b[4] , \a[8]  );
and  ( new_n4739_, new_n4692_, new_n4680_ );
and  ( new_n4740_, new_n4693_, new_n4679_ );
or   ( new_n4741_, new_n4740_, new_n4739_ );
and  ( new_n4742_, \b[3] , \a[9]  );
and  ( new_n4743_, new_n4690_, new_n4684_ );
and  ( new_n4744_, new_n4691_, new_n4683_ );
or   ( new_n4745_, new_n4744_, new_n4743_ );
and  ( new_n4746_, \b[2] , \a[10]  );
and  ( new_n4747_, new_n4688_, new_n1947_ );
and  ( new_n4748_, new_n4689_, new_n4687_ );
or   ( new_n4749_, new_n4748_, new_n4747_ );
and  ( new_n4750_, \b[0] , \a[12]  );
xor  ( new_n4751_, new_n4750_, new_n2002_ );
xor  ( new_n4752_, new_n4751_, new_n4749_ );
xor  ( new_n4753_, new_n4752_, new_n4746_ );
xor  ( new_n4754_, new_n4753_, new_n4745_ );
xor  ( new_n4755_, new_n4754_, new_n4742_ );
xor  ( new_n4756_, new_n4755_, new_n4741_ );
xor  ( new_n4757_, new_n4756_, new_n4738_ );
xor  ( new_n4758_, new_n4757_, new_n4737_ );
xor  ( new_n4759_, new_n4758_, new_n4734_ );
xor  ( new_n4760_, new_n4759_, new_n4733_ );
xor  ( new_n4761_, new_n4760_, new_n4730_ );
xor  ( new_n4762_, new_n4761_, new_n4729_ );
xor  ( new_n4763_, new_n4762_, new_n4726_ );
xor  ( new_n4764_, new_n4763_, new_n4725_ );
xor  ( new_n4765_, new_n4764_, new_n4722_ );
xor  ( new_n4766_, new_n4765_, new_n4721_ );
xor  ( new_n4767_, new_n4766_, new_n4718_ );
xor  ( new_n4768_, new_n4767_, new_n4717_ );
xor  ( new_n4769_, new_n4768_, new_n4714_ );
xor  ( new_n4770_, new_n4769_, new_n4713_ );
xor  ( new_n4771_, new_n4770_, new_n4710_ );
xor  ( new_n4772_, new_n4771_, new_n4709_ );
and  ( new_n4773_, new_n4772_, new_n4391_ );
and  ( new_n4774_, \b[12] , \a[1]  );
and  ( new_n4775_, new_n4770_, new_n4710_ );
and  ( new_n4776_, new_n4771_, new_n4709_ );
or   ( new_n4777_, new_n4776_, new_n4775_ );
and  ( new_n4778_, \b[11] , \a[2]  );
and  ( new_n4779_, new_n4768_, new_n4714_ );
and  ( new_n4780_, new_n4769_, new_n4713_ );
or   ( new_n4781_, new_n4780_, new_n4779_ );
and  ( new_n4782_, \b[10] , \a[3]  );
and  ( new_n4783_, new_n4766_, new_n4718_ );
and  ( new_n4784_, new_n4767_, new_n4717_ );
or   ( new_n4785_, new_n4784_, new_n4783_ );
and  ( new_n4786_, \b[9] , \a[4]  );
and  ( new_n4787_, new_n4764_, new_n4722_ );
and  ( new_n4788_, new_n4765_, new_n4721_ );
or   ( new_n4789_, new_n4788_, new_n4787_ );
and  ( new_n4790_, \b[8] , \a[5]  );
and  ( new_n4791_, new_n4762_, new_n4726_ );
and  ( new_n4792_, new_n4763_, new_n4725_ );
or   ( new_n4793_, new_n4792_, new_n4791_ );
and  ( new_n4794_, \b[7] , \a[6]  );
and  ( new_n4795_, new_n4760_, new_n4730_ );
and  ( new_n4796_, new_n4761_, new_n4729_ );
or   ( new_n4797_, new_n4796_, new_n4795_ );
and  ( new_n4798_, \b[6] , \a[7]  );
and  ( new_n4799_, new_n4758_, new_n4734_ );
and  ( new_n4800_, new_n4759_, new_n4733_ );
or   ( new_n4801_, new_n4800_, new_n4799_ );
and  ( new_n4802_, \b[5] , \a[8]  );
and  ( new_n4803_, new_n4756_, new_n4738_ );
and  ( new_n4804_, new_n4757_, new_n4737_ );
or   ( new_n4805_, new_n4804_, new_n4803_ );
and  ( new_n4806_, \b[4] , \a[9]  );
and  ( new_n4807_, new_n4754_, new_n4742_ );
and  ( new_n4808_, new_n4755_, new_n4741_ );
or   ( new_n4809_, new_n4808_, new_n4807_ );
and  ( new_n4810_, \b[3] , \a[10]  );
and  ( new_n4811_, new_n4752_, new_n4746_ );
and  ( new_n4812_, new_n4753_, new_n4745_ );
or   ( new_n4813_, new_n4812_, new_n4811_ );
and  ( new_n4814_, \b[2] , \a[11]  );
and  ( new_n4815_, new_n4750_, new_n2002_ );
and  ( new_n4816_, new_n4751_, new_n4749_ );
or   ( new_n4817_, new_n4816_, new_n4815_ );
and  ( new_n4818_, \b[1] , \a[12]  );
and  ( new_n4819_, \b[0] , \a[13]  );
xor  ( new_n4820_, new_n4819_, new_n4818_ );
xor  ( new_n4821_, new_n4820_, new_n4817_ );
xor  ( new_n4822_, new_n4821_, new_n4814_ );
xor  ( new_n4823_, new_n4822_, new_n4813_ );
xor  ( new_n4824_, new_n4823_, new_n4810_ );
xor  ( new_n4825_, new_n4824_, new_n4809_ );
xor  ( new_n4826_, new_n4825_, new_n4806_ );
xor  ( new_n4827_, new_n4826_, new_n4805_ );
xor  ( new_n4828_, new_n4827_, new_n4802_ );
xor  ( new_n4829_, new_n4828_, new_n4801_ );
xor  ( new_n4830_, new_n4829_, new_n4798_ );
xor  ( new_n4831_, new_n4830_, new_n4797_ );
xor  ( new_n4832_, new_n4831_, new_n4794_ );
xor  ( new_n4833_, new_n4832_, new_n4793_ );
xor  ( new_n4834_, new_n4833_, new_n4790_ );
xor  ( new_n4835_, new_n4834_, new_n4789_ );
xor  ( new_n4836_, new_n4835_, new_n4786_ );
xor  ( new_n4837_, new_n4836_, new_n4785_ );
xor  ( new_n4838_, new_n4837_, new_n4782_ );
xor  ( new_n4839_, new_n4838_, new_n4781_ );
xor  ( new_n4840_, new_n4839_, new_n4778_ );
xor  ( new_n4841_, new_n4840_, new_n4777_ );
xor  ( new_n4842_, new_n4841_, new_n4774_ );
xor  ( new_n4843_, new_n4842_, new_n4773_ );
and  ( new_n4844_, new_n4843_, new_n4390_ );
and  ( new_n4845_, \b[13] , \a[1]  );
and  ( new_n4846_, new_n4841_, new_n4774_ );
and  ( new_n4847_, new_n4842_, new_n4773_ );
or   ( new_n4848_, new_n4847_, new_n4846_ );
and  ( new_n4849_, \b[12] , \a[2]  );
and  ( new_n4850_, new_n4839_, new_n4778_ );
and  ( new_n4851_, new_n4840_, new_n4777_ );
nor  ( new_n4852_, new_n4851_, new_n4850_ );
not  ( new_n4853_, new_n4852_ );
and  ( new_n4854_, \b[11] , \a[3]  );
and  ( new_n4855_, new_n4837_, new_n4782_ );
and  ( new_n4856_, new_n4838_, new_n4781_ );
or   ( new_n4857_, new_n4856_, new_n4855_ );
and  ( new_n4858_, \b[10] , \a[4]  );
and  ( new_n4859_, new_n4835_, new_n4786_ );
and  ( new_n4860_, new_n4836_, new_n4785_ );
or   ( new_n4861_, new_n4860_, new_n4859_ );
and  ( new_n4862_, \b[9] , \a[5]  );
and  ( new_n4863_, new_n4833_, new_n4790_ );
and  ( new_n4864_, new_n4834_, new_n4789_ );
or   ( new_n4865_, new_n4864_, new_n4863_ );
and  ( new_n4866_, \b[8] , \a[6]  );
and  ( new_n4867_, new_n4831_, new_n4794_ );
and  ( new_n4868_, new_n4832_, new_n4793_ );
or   ( new_n4869_, new_n4868_, new_n4867_ );
and  ( new_n4870_, \b[7] , \a[7]  );
and  ( new_n4871_, new_n4829_, new_n4798_ );
and  ( new_n4872_, new_n4830_, new_n4797_ );
or   ( new_n4873_, new_n4872_, new_n4871_ );
and  ( new_n4874_, \b[6] , \a[8]  );
and  ( new_n4875_, new_n4827_, new_n4802_ );
and  ( new_n4876_, new_n4828_, new_n4801_ );
or   ( new_n4877_, new_n4876_, new_n4875_ );
and  ( new_n4878_, \b[5] , \a[9]  );
and  ( new_n4879_, new_n4825_, new_n4806_ );
and  ( new_n4880_, new_n4826_, new_n4805_ );
or   ( new_n4881_, new_n4880_, new_n4879_ );
and  ( new_n4882_, \b[4] , \a[10]  );
and  ( new_n4883_, new_n4823_, new_n4810_ );
and  ( new_n4884_, new_n4824_, new_n4809_ );
or   ( new_n4885_, new_n4884_, new_n4883_ );
and  ( new_n4886_, \b[3] , \a[11]  );
and  ( new_n4887_, new_n4821_, new_n4814_ );
and  ( new_n4888_, new_n4822_, new_n4813_ );
nor  ( new_n4889_, new_n4888_, new_n4887_ );
not  ( new_n4890_, new_n4889_ );
and  ( new_n4891_, \b[2] , \a[12]  );
and  ( new_n4892_, new_n4819_, new_n4818_ );
and  ( new_n4893_, new_n4820_, new_n4817_ );
nor  ( new_n4894_, new_n4893_, new_n4892_ );
not  ( new_n4895_, new_n4894_ );
and  ( new_n4896_, \b[1] , \a[13]  );
and  ( new_n4897_, \b[0] , \a[14]  );
xor  ( new_n4898_, new_n4897_, new_n4896_ );
xor  ( new_n4899_, new_n4898_, new_n4895_ );
xor  ( new_n4900_, new_n4899_, new_n4891_ );
xor  ( new_n4901_, new_n4900_, new_n4890_ );
xor  ( new_n4902_, new_n4901_, new_n4886_ );
xor  ( new_n4903_, new_n4902_, new_n4885_ );
xor  ( new_n4904_, new_n4903_, new_n4882_ );
xor  ( new_n4905_, new_n4904_, new_n4881_ );
xor  ( new_n4906_, new_n4905_, new_n4878_ );
xor  ( new_n4907_, new_n4906_, new_n4877_ );
xor  ( new_n4908_, new_n4907_, new_n4874_ );
xor  ( new_n4909_, new_n4908_, new_n4873_ );
xor  ( new_n4910_, new_n4909_, new_n4870_ );
xor  ( new_n4911_, new_n4910_, new_n4869_ );
xor  ( new_n4912_, new_n4911_, new_n4866_ );
xor  ( new_n4913_, new_n4912_, new_n4865_ );
xor  ( new_n4914_, new_n4913_, new_n4862_ );
xor  ( new_n4915_, new_n4914_, new_n4861_ );
xor  ( new_n4916_, new_n4915_, new_n4858_ );
xor  ( new_n4917_, new_n4916_, new_n4857_ );
xor  ( new_n4918_, new_n4917_, new_n4854_ );
xor  ( new_n4919_, new_n4918_, new_n4853_ );
xor  ( new_n4920_, new_n4919_, new_n4849_ );
xor  ( new_n4921_, new_n4920_, new_n4848_ );
xor  ( new_n4922_, new_n4921_, new_n4845_ );
xor  ( new_n4923_, new_n4922_, new_n4844_ );
and  ( new_n4924_, new_n4923_, new_n4389_ );
and  ( new_n4925_, new_n4921_, new_n4845_ );
and  ( new_n4926_, new_n4922_, new_n4844_ );
nor  ( new_n4927_, new_n4926_, new_n4925_ );
nand ( new_n4928_, new_n4917_, new_n4854_ );
nand ( new_n4929_, new_n4918_, new_n4853_ );
and  ( new_n4930_, new_n4929_, new_n4928_ );
and  ( new_n4931_, new_n4913_, new_n4862_ );
and  ( new_n4932_, new_n4914_, new_n4861_ );
or   ( new_n4933_, new_n4932_, new_n4931_ );
and  ( new_n4934_, new_n4909_, new_n4870_ );
and  ( new_n4935_, new_n4910_, new_n4869_ );
or   ( new_n4936_, new_n4935_, new_n4934_ );
and  ( new_n4937_, new_n4905_, new_n4878_ );
and  ( new_n4938_, new_n4906_, new_n4877_ );
or   ( new_n4939_, new_n4938_, new_n4937_ );
and  ( new_n4940_, new_n4901_, new_n4886_ );
and  ( new_n4941_, new_n4902_, new_n4885_ );
or   ( new_n4942_, new_n4941_, new_n4940_ );
nand ( new_n4943_, new_n4897_, new_n4896_ );
nand ( new_n4944_, new_n4898_, new_n4895_ );
and  ( new_n4945_, new_n4944_, new_n4943_ );
xor  ( new_n4946_, new_n4945_, new_n4942_ );
xor  ( new_n4947_, new_n4946_, new_n4939_ );
xor  ( new_n4948_, new_n4947_, new_n4936_ );
xor  ( new_n4949_, new_n4948_, new_n4933_ );
xor  ( new_n4950_, new_n4949_, new_n4930_ );
and  ( new_n4951_, new_n4919_, new_n4849_ );
and  ( new_n4952_, new_n4920_, new_n4848_ );
or   ( new_n4953_, new_n4952_, new_n4951_ );
and  ( new_n4954_, new_n4915_, new_n4858_ );
and  ( new_n4955_, new_n4916_, new_n4857_ );
or   ( new_n4956_, new_n4955_, new_n4954_ );
and  ( new_n4957_, new_n4911_, new_n4866_ );
and  ( new_n4958_, new_n4912_, new_n4865_ );
or   ( new_n4959_, new_n4958_, new_n4957_ );
and  ( new_n4960_, new_n4907_, new_n4874_ );
and  ( new_n4961_, new_n4908_, new_n4873_ );
or   ( new_n4962_, new_n4961_, new_n4960_ );
and  ( new_n4963_, new_n4903_, new_n4882_ );
and  ( new_n4964_, new_n4904_, new_n4881_ );
or   ( new_n4965_, new_n4964_, new_n4963_ );
nand ( new_n4966_, new_n4899_, new_n4891_ );
nand ( new_n4967_, new_n4900_, new_n4890_ );
and  ( new_n4968_, new_n4967_, new_n4966_ );
xor  ( new_n4969_, new_n4968_, new_n4965_ );
xor  ( new_n4970_, new_n4969_, new_n4962_ );
xor  ( new_n4971_, new_n4970_, new_n4959_ );
xor  ( new_n4972_, new_n4971_, new_n4956_ );
xor  ( new_n4973_, new_n4972_, new_n4953_ );
xor  ( new_n4974_, new_n4973_, new_n4950_ );
xnor ( new_n4975_, new_n4974_, new_n4927_ );
or   ( new_n4976_, new_n2206_, new_n108_ );
or   ( new_n4977_, new_n1053_, new_n163_ );
or   ( new_n4978_, new_n1038_, new_n176_ );
or   ( new_n4979_, new_n1328_, new_n185_ );
or   ( new_n4980_, new_n1019_, new_n137_ );
or   ( new_n4981_, new_n832_, new_n354_ );
and  ( new_n4982_, \b[2] , \a[13]  );
xor  ( new_n4983_, new_n4982_, new_n4981_ );
xor  ( new_n4984_, new_n4983_, new_n4980_ );
xor  ( new_n4985_, new_n4984_, new_n4979_ );
xor  ( new_n4986_, new_n4985_, new_n4978_ );
xor  ( new_n4987_, new_n4986_, new_n4977_ );
xor  ( new_n4988_, new_n4987_, new_n4976_ );
or   ( new_n4989_, new_n1783_, new_n98_ );
or   ( new_n4990_, new_n992_, new_n115_ );
or   ( new_n4991_, new_n1154_, new_n231_ );
or   ( new_n4992_, new_n1296_, new_n212_ );
or   ( new_n4993_, new_n1023_, new_n133_ );
or   ( new_n4994_, new_n847_, new_n352_ );
or   ( new_n4995_, new_n815_, new_n85_ );
or   ( new_n4996_, new_n808_, new_n2116_ );
and  ( new_n4997_, \b[0] , \a[15]  );
xor  ( new_n4998_, new_n4997_, new_n4996_ );
xor  ( new_n4999_, new_n4998_, new_n4995_ );
xor  ( new_n5000_, new_n4999_, new_n4994_ );
xor  ( new_n5001_, new_n5000_, new_n4993_ );
xor  ( new_n5002_, new_n5001_, new_n4992_ );
xor  ( new_n5003_, new_n5002_, new_n4991_ );
xor  ( new_n5004_, new_n5003_, new_n4990_ );
xor  ( new_n5005_, new_n5004_, new_n4989_ );
xor  ( new_n5006_, new_n5005_, new_n4988_ );
xor  ( new_n5007_, new_n5006_, new_n4975_ );
nor  ( new_n5008_, new_n5007_, new_n4924_ );
nor  ( new_n5009_, new_n4923_, new_n4389_ );
not  ( new_n5010_, new_n5009_ );
and  ( new_n5011_, new_n5010_, new_n5007_ );
nor  ( new_n5012_, new_n5011_, new_n5008_ );
xor  ( new_n5013_, new_n4598_, new_n4393_ );
not  ( new_n5014_, new_n5013_ );
xor  ( new_n5015_, new_n4843_, new_n4390_ );
not  ( new_n5016_, new_n5015_ );
xor  ( new_n5017_, new_n4772_, new_n4391_ );
not  ( new_n5018_, new_n5017_ );
xnor ( new_n5019_, new_n4650_, new_n2013_ );
not  ( new_n5020_, new_n5019_ );
xor  ( new_n5021_, new_n4708_, new_n4392_ );
not  ( new_n5022_, new_n5021_ );
and  ( new_n5023_, new_n5022_, new_n5020_ );
and  ( new_n5024_, new_n5023_, new_n5018_ );
and  ( new_n5025_, new_n5024_, new_n5016_ );
and  ( new_n5026_, new_n5025_, new_n5014_ );
and  ( new_n5027_, new_n5026_, new_n5012_ );
xor  ( new_n5028_, new_n4552_, new_n4394_ );
not  ( new_n5029_, new_n5028_ );
xor  ( new_n5030_, new_n4512_, new_n1896_ );
xor  ( new_n5031_, new_n4428_, new_n4396_ );
not  ( new_n5032_, new_n5031_ );
xor  ( new_n5033_, new_n4478_, new_n4395_ );
not  ( new_n5034_, new_n5033_ );
xor  ( new_n5035_, new_n4450_, new_n1696_ );
not  ( new_n5036_, new_n5035_ );
and  ( new_n5037_, new_n5036_, new_n5034_ );
xor  ( new_n5038_, new_n4412_, new_n882_ );
not  ( new_n5039_, new_n5038_ );
nor  ( new_n5040_, new_n2063_, new_n897_ );
and  ( new_n5041_, \b[0] , \a[0]  );
not  ( new_n5042_, new_n5041_ );
xor  ( new_n5043_, new_n4405_, new_n880_ );
not  ( new_n5044_, new_n5043_ );
and  ( new_n5045_, new_n5044_, new_n5042_ );
and  ( new_n5046_, new_n5045_, new_n5040_ );
and  ( new_n5047_, new_n5046_, new_n5039_ );
and  ( new_n5048_, new_n5047_, new_n5037_ );
and  ( new_n5049_, new_n5048_, new_n5032_ );
and  ( new_n5050_, new_n5049_, new_n5030_ );
and  ( new_n5051_, new_n5050_, new_n5029_ );
and  ( new_n5052_, new_n5051_, new_n5027_ );
not  ( new_n5053_, new_n5030_ );
and  ( new_n5054_, new_n5049_, new_n5053_ );
and  ( new_n5055_, new_n5054_, new_n5028_ );
and  ( new_n5056_, new_n5055_, new_n5027_ );
and  ( new_n5057_, new_n5053_, new_n5029_ );
and  ( new_n5058_, new_n5057_, new_n5049_ );
and  ( new_n5059_, new_n5058_, new_n5014_ );
and  ( new_n5060_, new_n5059_, new_n5018_ );
and  ( new_n5061_, new_n5060_, new_n5012_ );
and  ( new_n5062_, new_n5022_, new_n5019_ );
and  ( new_n5063_, new_n5062_, new_n5016_ );
and  ( new_n5064_, new_n5063_, new_n5061_ );
or   ( new_n5065_, new_n5064_, new_n5056_ );
or   ( new_n5066_, new_n5065_, new_n5052_ );
and  ( new_n5067_, new_n5057_, new_n5034_ );
and  ( new_n5068_, new_n5046_, new_n5038_ );
and  ( new_n5069_, new_n5068_, new_n5032_ );
and  ( new_n5070_, new_n5069_, new_n5036_ );
and  ( new_n5071_, new_n5070_, new_n5067_ );
and  ( new_n5072_, new_n5071_, new_n5027_ );
and  ( new_n5073_, new_n5047_, new_n5032_ );
and  ( new_n5074_, new_n5073_, new_n5035_ );
and  ( new_n5075_, new_n5074_, new_n5067_ );
and  ( new_n5076_, new_n5075_, new_n5027_ );
or   ( new_n5077_, new_n5076_, new_n5072_ );
and  ( new_n5078_, new_n5048_, new_n5031_ );
and  ( new_n5079_, new_n5078_, new_n5057_ );
and  ( new_n5080_, new_n5079_, new_n5027_ );
and  ( new_n5081_, new_n5021_, new_n5020_ );
and  ( new_n5082_, new_n5081_, new_n5016_ );
and  ( new_n5083_, new_n5082_, new_n5061_ );
or   ( new_n5084_, new_n5083_, new_n5080_ );
or   ( new_n5085_, new_n5084_, new_n5077_ );
and  ( new_n5086_, new_n5039_, new_n5032_ );
and  ( new_n5087_, new_n5042_, new_n5040_ );
and  ( new_n5088_, new_n5087_, new_n5043_ );
and  ( new_n5089_, new_n5088_, new_n5086_ );
and  ( new_n5090_, new_n5089_, new_n5036_ );
and  ( new_n5091_, new_n5090_, new_n5067_ );
and  ( new_n5092_, new_n5091_, new_n5027_ );
and  ( new_n5093_, new_n5073_, new_n5036_ );
and  ( new_n5094_, new_n5093_, new_n5033_ );
and  ( new_n5095_, new_n5094_, new_n5057_ );
and  ( new_n5096_, new_n5095_, new_n5014_ );
and  ( new_n5097_, new_n5096_, new_n5025_ );
and  ( new_n5098_, new_n5097_, new_n5012_ );
and  ( new_n5099_, new_n5054_, new_n5029_ );
and  ( new_n5100_, new_n5099_, new_n5013_ );
and  ( new_n5101_, new_n5100_, new_n5025_ );
and  ( new_n5102_, new_n5101_, new_n5012_ );
or   ( new_n5103_, new_n5102_, new_n5098_ );
or   ( new_n5104_, new_n5103_, new_n5092_ );
and  ( new_n5105_, new_n5041_, new_n2065_ );
and  ( new_n5106_, new_n5105_, new_n5044_ );
and  ( new_n5107_, new_n5106_, new_n5086_ );
and  ( new_n5108_, new_n5107_, new_n5037_ );
and  ( new_n5109_, new_n5108_, new_n5057_ );
and  ( new_n5110_, new_n5109_, new_n5027_ );
not  ( new_n5111_, new_n5040_ );
and  ( new_n5112_, new_n5045_, new_n5111_ );
and  ( new_n5113_, new_n5112_, new_n5086_ );
and  ( new_n5114_, new_n5113_, new_n5037_ );
and  ( new_n5115_, new_n5114_, new_n5057_ );
and  ( new_n5116_, new_n5115_, new_n5027_ );
or   ( new_n5117_, new_n5116_, new_n5110_ );
or   ( new_n5118_, new_n5117_, new_n5104_ );
or   ( new_n5119_, new_n5118_, new_n5085_ );
or   ( new_n5120_, new_n5119_, new_n5066_ );
and  ( new_n5121_, new_n5083_, new_n2203_ );
not  ( new_n5122_, new_n5121_ );
and  ( new_n5123_, \d[8] , \a[0]  );
and  ( new_n5124_, new_n3202_, new_n757_ );
and  ( new_n5125_, \d[1] , \a[1]  );
and  ( new_n5126_, \d[0] , \a[2]  );
and  ( new_n5127_, new_n5126_, new_n5125_ );
xnor ( new_n5128_, new_n5127_, new_n5124_ );
or   ( new_n5129_, new_n5126_, new_n5125_ );
and  ( new_n5130_, new_n5129_, new_n5128_ );
and  ( new_n5131_, new_n5130_, new_n740_ );
and  ( new_n5132_, \d[2] , \a[1]  );
or   ( new_n5133_, new_n5127_, new_n5124_ );
and  ( new_n5134_, \d[0] , \a[3]  );
xor  ( new_n5135_, new_n5134_, new_n751_ );
xor  ( new_n5136_, new_n5135_, new_n5133_ );
xor  ( new_n5137_, new_n5136_, new_n5132_ );
xor  ( new_n5138_, new_n5137_, new_n5131_ );
and  ( new_n5139_, new_n5138_, new_n742_ );
and  ( new_n5140_, \d[3] , \a[1]  );
and  ( new_n5141_, new_n5136_, new_n5132_ );
and  ( new_n5142_, new_n5137_, new_n5131_ );
or   ( new_n5143_, new_n5142_, new_n5141_ );
and  ( new_n5144_, \d[2] , \a[2]  );
and  ( new_n5145_, new_n5134_, new_n751_ );
and  ( new_n5146_, new_n5135_, new_n5133_ );
or   ( new_n5147_, new_n5146_, new_n5145_ );
and  ( new_n5148_, \d[0] , \a[4]  );
xor  ( new_n5149_, new_n5148_, new_n722_ );
xor  ( new_n5150_, new_n5149_, new_n5147_ );
xor  ( new_n5151_, new_n5150_, new_n5144_ );
xor  ( new_n5152_, new_n5151_, new_n5143_ );
xor  ( new_n5153_, new_n5152_, new_n5140_ );
xor  ( new_n5154_, new_n5153_, new_n5139_ );
and  ( new_n5155_, new_n5154_, new_n685_ );
and  ( new_n5156_, \d[4] , \a[1]  );
and  ( new_n5157_, new_n5152_, new_n5140_ );
and  ( new_n5158_, new_n5153_, new_n5139_ );
or   ( new_n5159_, new_n5158_, new_n5157_ );
and  ( new_n5160_, \d[3] , \a[2]  );
and  ( new_n5161_, new_n5150_, new_n5144_ );
and  ( new_n5162_, new_n5151_, new_n5143_ );
or   ( new_n5163_, new_n5162_, new_n5161_ );
and  ( new_n5164_, \d[2] , \a[3]  );
and  ( new_n5165_, new_n5148_, new_n722_ );
and  ( new_n5166_, new_n5149_, new_n5147_ );
or   ( new_n5167_, new_n5166_, new_n5165_ );
and  ( new_n5168_, \d[0] , \a[5]  );
xor  ( new_n5169_, new_n5168_, new_n705_ );
xor  ( new_n5170_, new_n5169_, new_n5167_ );
xor  ( new_n5171_, new_n5170_, new_n5164_ );
xor  ( new_n5172_, new_n5171_, new_n5163_ );
xor  ( new_n5173_, new_n5172_, new_n5160_ );
xor  ( new_n5174_, new_n5173_, new_n5159_ );
xor  ( new_n5175_, new_n5174_, new_n5156_ );
xor  ( new_n5176_, new_n5175_, new_n5155_ );
and  ( new_n5177_, new_n5176_, new_n687_ );
and  ( new_n5178_, \d[5] , \a[1]  );
and  ( new_n5179_, new_n5174_, new_n5156_ );
and  ( new_n5180_, new_n5175_, new_n5155_ );
or   ( new_n5181_, new_n5180_, new_n5179_ );
and  ( new_n5182_, \d[4] , \a[2]  );
and  ( new_n5183_, new_n5172_, new_n5160_ );
and  ( new_n5184_, new_n5173_, new_n5159_ );
or   ( new_n5185_, new_n5184_, new_n5183_ );
and  ( new_n5186_, \d[3] , \a[3]  );
and  ( new_n5187_, new_n5170_, new_n5164_ );
and  ( new_n5188_, new_n5171_, new_n5163_ );
or   ( new_n5189_, new_n5188_, new_n5187_ );
and  ( new_n5190_, \d[2] , \a[4]  );
and  ( new_n5191_, new_n5168_, new_n705_ );
and  ( new_n5192_, new_n5169_, new_n5167_ );
or   ( new_n5193_, new_n5192_, new_n5191_ );
and  ( new_n5194_, \d[0] , \a[6]  );
xor  ( new_n5195_, new_n5194_, new_n656_ );
xor  ( new_n5196_, new_n5195_, new_n5193_ );
xor  ( new_n5197_, new_n5196_, new_n5190_ );
xor  ( new_n5198_, new_n5197_, new_n5189_ );
xor  ( new_n5199_, new_n5198_, new_n5186_ );
xor  ( new_n5200_, new_n5199_, new_n5185_ );
xor  ( new_n5201_, new_n5200_, new_n5182_ );
xor  ( new_n5202_, new_n5201_, new_n5181_ );
xor  ( new_n5203_, new_n5202_, new_n5178_ );
xor  ( new_n5204_, new_n5203_, new_n5177_ );
and  ( new_n5205_, new_n5204_, new_n602_ );
and  ( new_n5206_, \d[6] , \a[1]  );
and  ( new_n5207_, new_n5202_, new_n5178_ );
and  ( new_n5208_, new_n5203_, new_n5177_ );
or   ( new_n5209_, new_n5208_, new_n5207_ );
and  ( new_n5210_, \d[5] , \a[2]  );
and  ( new_n5211_, new_n5200_, new_n5182_ );
and  ( new_n5212_, new_n5201_, new_n5181_ );
or   ( new_n5213_, new_n5212_, new_n5211_ );
and  ( new_n5214_, \d[4] , \a[3]  );
and  ( new_n5215_, new_n5198_, new_n5186_ );
and  ( new_n5216_, new_n5199_, new_n5185_ );
or   ( new_n5217_, new_n5216_, new_n5215_ );
and  ( new_n5218_, \d[3] , \a[4]  );
and  ( new_n5219_, new_n5196_, new_n5190_ );
and  ( new_n5220_, new_n5197_, new_n5189_ );
or   ( new_n5221_, new_n5220_, new_n5219_ );
and  ( new_n5222_, \d[2] , \a[5]  );
and  ( new_n5223_, new_n5194_, new_n656_ );
and  ( new_n5224_, new_n5195_, new_n5193_ );
or   ( new_n5225_, new_n5224_, new_n5223_ );
and  ( new_n5226_, \d[0] , \a[7]  );
xor  ( new_n5227_, new_n5226_, new_n626_ );
xor  ( new_n5228_, new_n5227_, new_n5225_ );
xor  ( new_n5229_, new_n5228_, new_n5222_ );
xor  ( new_n5230_, new_n5229_, new_n5221_ );
xor  ( new_n5231_, new_n5230_, new_n5218_ );
xor  ( new_n5232_, new_n5231_, new_n5217_ );
xor  ( new_n5233_, new_n5232_, new_n5214_ );
xor  ( new_n5234_, new_n5233_, new_n5213_ );
xor  ( new_n5235_, new_n5234_, new_n5210_ );
xor  ( new_n5236_, new_n5235_, new_n5209_ );
xor  ( new_n5237_, new_n5236_, new_n5206_ );
xor  ( new_n5238_, new_n5237_, new_n5205_ );
and  ( new_n5239_, new_n5238_, new_n472_ );
and  ( new_n5240_, \d[7] , \a[1]  );
and  ( new_n5241_, new_n5236_, new_n5206_ );
and  ( new_n5242_, new_n5237_, new_n5205_ );
or   ( new_n5243_, new_n5242_, new_n5241_ );
and  ( new_n5244_, \d[6] , \a[2]  );
and  ( new_n5245_, new_n5234_, new_n5210_ );
and  ( new_n5246_, new_n5235_, new_n5209_ );
or   ( new_n5247_, new_n5246_, new_n5245_ );
and  ( new_n5248_, \d[5] , \a[3]  );
and  ( new_n5249_, new_n5232_, new_n5214_ );
and  ( new_n5250_, new_n5233_, new_n5213_ );
or   ( new_n5251_, new_n5250_, new_n5249_ );
and  ( new_n5252_, \d[4] , \a[4]  );
and  ( new_n5253_, new_n5230_, new_n5218_ );
and  ( new_n5254_, new_n5231_, new_n5217_ );
or   ( new_n5255_, new_n5254_, new_n5253_ );
and  ( new_n5256_, \d[3] , \a[5]  );
and  ( new_n5257_, new_n5228_, new_n5222_ );
and  ( new_n5258_, new_n5229_, new_n5221_ );
or   ( new_n5259_, new_n5258_, new_n5257_ );
and  ( new_n5260_, \d[2] , \a[6]  );
and  ( new_n5261_, new_n5226_, new_n626_ );
and  ( new_n5262_, new_n5227_, new_n5225_ );
or   ( new_n5263_, new_n5262_, new_n5261_ );
and  ( new_n5264_, \d[0] , \a[8]  );
xor  ( new_n5265_, new_n5264_, new_n558_ );
xor  ( new_n5266_, new_n5265_, new_n5263_ );
xor  ( new_n5267_, new_n5266_, new_n5260_ );
xor  ( new_n5268_, new_n5267_, new_n5259_ );
xor  ( new_n5269_, new_n5268_, new_n5256_ );
xor  ( new_n5270_, new_n5269_, new_n5255_ );
xor  ( new_n5271_, new_n5270_, new_n5252_ );
xor  ( new_n5272_, new_n5271_, new_n5251_ );
xor  ( new_n5273_, new_n5272_, new_n5248_ );
xor  ( new_n5274_, new_n5273_, new_n5247_ );
xor  ( new_n5275_, new_n5274_, new_n5244_ );
xor  ( new_n5276_, new_n5275_, new_n5243_ );
xor  ( new_n5277_, new_n5276_, new_n5240_ );
xor  ( new_n5278_, new_n5277_, new_n5239_ );
and  ( new_n5279_, new_n5278_, new_n5123_ );
and  ( new_n5280_, \d[8] , \a[1]  );
and  ( new_n5281_, new_n5276_, new_n5240_ );
and  ( new_n5282_, new_n5277_, new_n5239_ );
or   ( new_n5283_, new_n5282_, new_n5281_ );
and  ( new_n5284_, \d[7] , \a[2]  );
and  ( new_n5285_, new_n5274_, new_n5244_ );
and  ( new_n5286_, new_n5275_, new_n5243_ );
or   ( new_n5287_, new_n5286_, new_n5285_ );
and  ( new_n5288_, \d[6] , \a[3]  );
and  ( new_n5289_, new_n5272_, new_n5248_ );
and  ( new_n5290_, new_n5273_, new_n5247_ );
or   ( new_n5291_, new_n5290_, new_n5289_ );
and  ( new_n5292_, \d[5] , \a[4]  );
and  ( new_n5293_, new_n5270_, new_n5252_ );
and  ( new_n5294_, new_n5271_, new_n5251_ );
or   ( new_n5295_, new_n5294_, new_n5293_ );
and  ( new_n5296_, \d[4] , \a[5]  );
and  ( new_n5297_, new_n5268_, new_n5256_ );
and  ( new_n5298_, new_n5269_, new_n5255_ );
or   ( new_n5299_, new_n5298_, new_n5297_ );
and  ( new_n5300_, \d[3] , \a[6]  );
and  ( new_n5301_, new_n5266_, new_n5260_ );
and  ( new_n5302_, new_n5267_, new_n5259_ );
or   ( new_n5303_, new_n5302_, new_n5301_ );
and  ( new_n5304_, \d[2] , \a[7]  );
and  ( new_n5305_, new_n5264_, new_n558_ );
and  ( new_n5306_, new_n5265_, new_n5263_ );
or   ( new_n5307_, new_n5306_, new_n5305_ );
and  ( new_n5308_, \d[0] , \a[9]  );
xor  ( new_n5309_, new_n5308_, new_n518_ );
xor  ( new_n5310_, new_n5309_, new_n5307_ );
xor  ( new_n5311_, new_n5310_, new_n5304_ );
xor  ( new_n5312_, new_n5311_, new_n5303_ );
xor  ( new_n5313_, new_n5312_, new_n5300_ );
xor  ( new_n5314_, new_n5313_, new_n5299_ );
xor  ( new_n5315_, new_n5314_, new_n5296_ );
xor  ( new_n5316_, new_n5315_, new_n5295_ );
xor  ( new_n5317_, new_n5316_, new_n5292_ );
xor  ( new_n5318_, new_n5317_, new_n5291_ );
xor  ( new_n5319_, new_n5318_, new_n5288_ );
xor  ( new_n5320_, new_n5319_, new_n5287_ );
xor  ( new_n5321_, new_n5320_, new_n5284_ );
xor  ( new_n5322_, new_n5321_, new_n5283_ );
xor  ( new_n5323_, new_n5322_, new_n5280_ );
xor  ( new_n5324_, new_n5323_, new_n5279_ );
and  ( new_n5325_, new_n5324_, new_n329_ );
and  ( new_n5326_, \d[9] , \a[1]  );
and  ( new_n5327_, new_n5322_, new_n5280_ );
and  ( new_n5328_, new_n5323_, new_n5279_ );
or   ( new_n5329_, new_n5328_, new_n5327_ );
and  ( new_n5330_, \d[8] , \a[2]  );
and  ( new_n5331_, new_n5320_, new_n5284_ );
and  ( new_n5332_, new_n5321_, new_n5283_ );
or   ( new_n5333_, new_n5332_, new_n5331_ );
and  ( new_n5334_, \d[7] , \a[3]  );
and  ( new_n5335_, new_n5318_, new_n5288_ );
and  ( new_n5336_, new_n5319_, new_n5287_ );
or   ( new_n5337_, new_n5336_, new_n5335_ );
and  ( new_n5338_, \d[6] , \a[4]  );
and  ( new_n5339_, new_n5316_, new_n5292_ );
and  ( new_n5340_, new_n5317_, new_n5291_ );
or   ( new_n5341_, new_n5340_, new_n5339_ );
and  ( new_n5342_, \d[5] , \a[5]  );
and  ( new_n5343_, new_n5314_, new_n5296_ );
and  ( new_n5344_, new_n5315_, new_n5295_ );
or   ( new_n5345_, new_n5344_, new_n5343_ );
and  ( new_n5346_, \d[4] , \a[6]  );
and  ( new_n5347_, new_n5312_, new_n5300_ );
and  ( new_n5348_, new_n5313_, new_n5299_ );
or   ( new_n5349_, new_n5348_, new_n5347_ );
and  ( new_n5350_, \d[3] , \a[7]  );
and  ( new_n5351_, new_n5310_, new_n5304_ );
and  ( new_n5352_, new_n5311_, new_n5303_ );
or   ( new_n5353_, new_n5352_, new_n5351_ );
and  ( new_n5354_, \d[2] , \a[8]  );
and  ( new_n5355_, new_n5308_, new_n518_ );
and  ( new_n5356_, new_n5309_, new_n5307_ );
or   ( new_n5357_, new_n5356_, new_n5355_ );
and  ( new_n5358_, \d[0] , \a[10]  );
xor  ( new_n5359_, new_n5358_, new_n487_ );
xor  ( new_n5360_, new_n5359_, new_n5357_ );
xor  ( new_n5361_, new_n5360_, new_n5354_ );
xor  ( new_n5362_, new_n5361_, new_n5353_ );
xor  ( new_n5363_, new_n5362_, new_n5350_ );
xor  ( new_n5364_, new_n5363_, new_n5349_ );
xor  ( new_n5365_, new_n5364_, new_n5346_ );
xor  ( new_n5366_, new_n5365_, new_n5345_ );
xor  ( new_n5367_, new_n5366_, new_n5342_ );
xor  ( new_n5368_, new_n5367_, new_n5341_ );
xor  ( new_n5369_, new_n5368_, new_n5338_ );
xor  ( new_n5370_, new_n5369_, new_n5337_ );
xor  ( new_n5371_, new_n5370_, new_n5334_ );
xor  ( new_n5372_, new_n5371_, new_n5333_ );
xor  ( new_n5373_, new_n5372_, new_n5330_ );
xor  ( new_n5374_, new_n5373_, new_n5329_ );
xor  ( new_n5375_, new_n5374_, new_n5326_ );
xor  ( new_n5376_, new_n5375_, new_n5325_ );
and  ( new_n5377_, new_n5376_, new_n387_ );
and  ( new_n5378_, \d[10] , \a[1]  );
and  ( new_n5379_, new_n5374_, new_n5326_ );
and  ( new_n5380_, new_n5375_, new_n5325_ );
or   ( new_n5381_, new_n5380_, new_n5379_ );
and  ( new_n5382_, \d[9] , \a[2]  );
and  ( new_n5383_, new_n5372_, new_n5330_ );
and  ( new_n5384_, new_n5373_, new_n5329_ );
or   ( new_n5385_, new_n5384_, new_n5383_ );
and  ( new_n5386_, \d[8] , \a[3]  );
and  ( new_n5387_, new_n5370_, new_n5334_ );
and  ( new_n5388_, new_n5371_, new_n5333_ );
or   ( new_n5389_, new_n5388_, new_n5387_ );
and  ( new_n5390_, \d[7] , \a[4]  );
and  ( new_n5391_, new_n5368_, new_n5338_ );
and  ( new_n5392_, new_n5369_, new_n5337_ );
or   ( new_n5393_, new_n5392_, new_n5391_ );
and  ( new_n5394_, \d[6] , \a[5]  );
and  ( new_n5395_, new_n5366_, new_n5342_ );
and  ( new_n5396_, new_n5367_, new_n5341_ );
or   ( new_n5397_, new_n5396_, new_n5395_ );
and  ( new_n5398_, \d[5] , \a[6]  );
and  ( new_n5399_, new_n5364_, new_n5346_ );
and  ( new_n5400_, new_n5365_, new_n5345_ );
or   ( new_n5401_, new_n5400_, new_n5399_ );
and  ( new_n5402_, \d[4] , \a[7]  );
and  ( new_n5403_, new_n5362_, new_n5350_ );
and  ( new_n5404_, new_n5363_, new_n5349_ );
or   ( new_n5405_, new_n5404_, new_n5403_ );
and  ( new_n5406_, \d[3] , \a[8]  );
and  ( new_n5407_, new_n5360_, new_n5354_ );
and  ( new_n5408_, new_n5361_, new_n5353_ );
or   ( new_n5409_, new_n5408_, new_n5407_ );
and  ( new_n5410_, \d[2] , \a[9]  );
and  ( new_n5411_, new_n5358_, new_n487_ );
and  ( new_n5412_, new_n5359_, new_n5357_ );
or   ( new_n5413_, new_n5412_, new_n5411_ );
and  ( new_n5414_, \d[0] , \a[11]  );
xor  ( new_n5415_, new_n5414_, new_n422_ );
xor  ( new_n5416_, new_n5415_, new_n5413_ );
xor  ( new_n5417_, new_n5416_, new_n5410_ );
xor  ( new_n5418_, new_n5417_, new_n5409_ );
xor  ( new_n5419_, new_n5418_, new_n5406_ );
xor  ( new_n5420_, new_n5419_, new_n5405_ );
xor  ( new_n5421_, new_n5420_, new_n5402_ );
xor  ( new_n5422_, new_n5421_, new_n5401_ );
xor  ( new_n5423_, new_n5422_, new_n5398_ );
xor  ( new_n5424_, new_n5423_, new_n5397_ );
xor  ( new_n5425_, new_n5424_, new_n5394_ );
xor  ( new_n5426_, new_n5425_, new_n5393_ );
xor  ( new_n5427_, new_n5426_, new_n5390_ );
xor  ( new_n5428_, new_n5427_, new_n5389_ );
xor  ( new_n5429_, new_n5428_, new_n5386_ );
xor  ( new_n5430_, new_n5429_, new_n5385_ );
xor  ( new_n5431_, new_n5430_, new_n5382_ );
xor  ( new_n5432_, new_n5431_, new_n5381_ );
xor  ( new_n5433_, new_n5432_, new_n5378_ );
xor  ( new_n5434_, new_n5433_, new_n5377_ );
and  ( new_n5435_, new_n5434_, new_n389_ );
and  ( new_n5436_, \d[11] , \a[1]  );
and  ( new_n5437_, new_n5432_, new_n5378_ );
and  ( new_n5438_, new_n5433_, new_n5377_ );
or   ( new_n5439_, new_n5438_, new_n5437_ );
and  ( new_n5440_, \d[10] , \a[2]  );
and  ( new_n5441_, new_n5430_, new_n5382_ );
and  ( new_n5442_, new_n5431_, new_n5381_ );
or   ( new_n5443_, new_n5442_, new_n5441_ );
and  ( new_n5444_, \d[9] , \a[3]  );
and  ( new_n5445_, new_n5428_, new_n5386_ );
and  ( new_n5446_, new_n5429_, new_n5385_ );
or   ( new_n5447_, new_n5446_, new_n5445_ );
and  ( new_n5448_, \d[8] , \a[4]  );
and  ( new_n5449_, new_n5426_, new_n5390_ );
and  ( new_n5450_, new_n5427_, new_n5389_ );
or   ( new_n5451_, new_n5450_, new_n5449_ );
and  ( new_n5452_, \d[7] , \a[5]  );
and  ( new_n5453_, new_n5424_, new_n5394_ );
and  ( new_n5454_, new_n5425_, new_n5393_ );
or   ( new_n5455_, new_n5454_, new_n5453_ );
and  ( new_n5456_, \d[6] , \a[6]  );
and  ( new_n5457_, new_n5422_, new_n5398_ );
and  ( new_n5458_, new_n5423_, new_n5397_ );
or   ( new_n5459_, new_n5458_, new_n5457_ );
and  ( new_n5460_, \d[5] , \a[7]  );
and  ( new_n5461_, new_n5420_, new_n5402_ );
and  ( new_n5462_, new_n5421_, new_n5401_ );
or   ( new_n5463_, new_n5462_, new_n5461_ );
and  ( new_n5464_, \d[4] , \a[8]  );
and  ( new_n5465_, new_n5418_, new_n5406_ );
and  ( new_n5466_, new_n5419_, new_n5405_ );
or   ( new_n5467_, new_n5466_, new_n5465_ );
and  ( new_n5468_, \d[3] , \a[9]  );
and  ( new_n5469_, new_n5416_, new_n5410_ );
and  ( new_n5470_, new_n5417_, new_n5409_ );
or   ( new_n5471_, new_n5470_, new_n5469_ );
and  ( new_n5472_, \d[2] , \a[10]  );
and  ( new_n5473_, new_n5414_, new_n422_ );
and  ( new_n5474_, new_n5415_, new_n5413_ );
or   ( new_n5475_, new_n5474_, new_n5473_ );
and  ( new_n5476_, \d[0] , \a[12]  );
xor  ( new_n5477_, new_n5476_, new_n357_ );
xor  ( new_n5478_, new_n5477_, new_n5475_ );
xor  ( new_n5479_, new_n5478_, new_n5472_ );
xor  ( new_n5480_, new_n5479_, new_n5471_ );
xor  ( new_n5481_, new_n5480_, new_n5468_ );
xor  ( new_n5482_, new_n5481_, new_n5467_ );
xor  ( new_n5483_, new_n5482_, new_n5464_ );
xor  ( new_n5484_, new_n5483_, new_n5463_ );
xor  ( new_n5485_, new_n5484_, new_n5460_ );
xor  ( new_n5486_, new_n5485_, new_n5459_ );
xor  ( new_n5487_, new_n5486_, new_n5456_ );
xor  ( new_n5488_, new_n5487_, new_n5455_ );
xor  ( new_n5489_, new_n5488_, new_n5452_ );
xor  ( new_n5490_, new_n5489_, new_n5451_ );
xor  ( new_n5491_, new_n5490_, new_n5448_ );
xor  ( new_n5492_, new_n5491_, new_n5447_ );
xor  ( new_n5493_, new_n5492_, new_n5444_ );
xor  ( new_n5494_, new_n5493_, new_n5443_ );
xor  ( new_n5495_, new_n5494_, new_n5440_ );
xor  ( new_n5496_, new_n5495_, new_n5439_ );
xor  ( new_n5497_, new_n5496_, new_n5436_ );
xor  ( new_n5498_, new_n5497_, new_n5435_ );
and  ( new_n5499_, new_n5498_, new_n275_ );
and  ( new_n5500_, \d[12] , \a[1]  );
and  ( new_n5501_, new_n5496_, new_n5436_ );
and  ( new_n5502_, new_n5497_, new_n5435_ );
or   ( new_n5503_, new_n5502_, new_n5501_ );
and  ( new_n5504_, \d[11] , \a[2]  );
and  ( new_n5505_, new_n5494_, new_n5440_ );
and  ( new_n5506_, new_n5495_, new_n5439_ );
or   ( new_n5507_, new_n5506_, new_n5505_ );
and  ( new_n5508_, \d[10] , \a[3]  );
and  ( new_n5509_, new_n5492_, new_n5444_ );
and  ( new_n5510_, new_n5493_, new_n5443_ );
or   ( new_n5511_, new_n5510_, new_n5509_ );
and  ( new_n5512_, \d[9] , \a[4]  );
and  ( new_n5513_, new_n5490_, new_n5448_ );
and  ( new_n5514_, new_n5491_, new_n5447_ );
or   ( new_n5515_, new_n5514_, new_n5513_ );
and  ( new_n5516_, \d[8] , \a[5]  );
and  ( new_n5517_, new_n5488_, new_n5452_ );
and  ( new_n5518_, new_n5489_, new_n5451_ );
or   ( new_n5519_, new_n5518_, new_n5517_ );
and  ( new_n5520_, \d[7] , \a[6]  );
and  ( new_n5521_, new_n5486_, new_n5456_ );
and  ( new_n5522_, new_n5487_, new_n5455_ );
or   ( new_n5523_, new_n5522_, new_n5521_ );
and  ( new_n5524_, \d[6] , \a[7]  );
and  ( new_n5525_, new_n5484_, new_n5460_ );
and  ( new_n5526_, new_n5485_, new_n5459_ );
or   ( new_n5527_, new_n5526_, new_n5525_ );
and  ( new_n5528_, \d[5] , \a[8]  );
and  ( new_n5529_, new_n5482_, new_n5464_ );
and  ( new_n5530_, new_n5483_, new_n5463_ );
or   ( new_n5531_, new_n5530_, new_n5529_ );
and  ( new_n5532_, \d[4] , \a[9]  );
and  ( new_n5533_, new_n5480_, new_n5468_ );
and  ( new_n5534_, new_n5481_, new_n5467_ );
or   ( new_n5535_, new_n5534_, new_n5533_ );
and  ( new_n5536_, \d[3] , \a[10]  );
and  ( new_n5537_, new_n5478_, new_n5472_ );
and  ( new_n5538_, new_n5479_, new_n5471_ );
or   ( new_n5539_, new_n5538_, new_n5537_ );
and  ( new_n5540_, \d[2] , \a[11]  );
and  ( new_n5541_, new_n5476_, new_n357_ );
and  ( new_n5542_, new_n5477_, new_n5475_ );
or   ( new_n5543_, new_n5542_, new_n5541_ );
and  ( new_n5544_, \d[0] , \a[13]  );
xor  ( new_n5545_, new_n5544_, new_n238_ );
xor  ( new_n5546_, new_n5545_, new_n5543_ );
xor  ( new_n5547_, new_n5546_, new_n5540_ );
xor  ( new_n5548_, new_n5547_, new_n5539_ );
xor  ( new_n5549_, new_n5548_, new_n5536_ );
xor  ( new_n5550_, new_n5549_, new_n5535_ );
xor  ( new_n5551_, new_n5550_, new_n5532_ );
xor  ( new_n5552_, new_n5551_, new_n5531_ );
xor  ( new_n5553_, new_n5552_, new_n5528_ );
xor  ( new_n5554_, new_n5553_, new_n5527_ );
xor  ( new_n5555_, new_n5554_, new_n5524_ );
xor  ( new_n5556_, new_n5555_, new_n5523_ );
xor  ( new_n5557_, new_n5556_, new_n5520_ );
xor  ( new_n5558_, new_n5557_, new_n5519_ );
xor  ( new_n5559_, new_n5558_, new_n5516_ );
xor  ( new_n5560_, new_n5559_, new_n5515_ );
xor  ( new_n5561_, new_n5560_, new_n5512_ );
xor  ( new_n5562_, new_n5561_, new_n5511_ );
xor  ( new_n5563_, new_n5562_, new_n5508_ );
xor  ( new_n5564_, new_n5563_, new_n5507_ );
xor  ( new_n5565_, new_n5564_, new_n5504_ );
xor  ( new_n5566_, new_n5565_, new_n5503_ );
xor  ( new_n5567_, new_n5566_, new_n5500_ );
xor  ( new_n5568_, new_n5567_, new_n5499_ );
and  ( new_n5569_, new_n5568_, new_n277_ );
and  ( new_n5570_, \d[13] , \a[1]  );
and  ( new_n5571_, new_n5566_, new_n5500_ );
and  ( new_n5572_, new_n5567_, new_n5499_ );
or   ( new_n5573_, new_n5572_, new_n5571_ );
and  ( new_n5574_, \d[12] , \a[2]  );
and  ( new_n5575_, new_n5564_, new_n5504_ );
and  ( new_n5576_, new_n5565_, new_n5503_ );
or   ( new_n5577_, new_n5576_, new_n5575_ );
and  ( new_n5578_, \d[11] , \a[3]  );
and  ( new_n5579_, new_n5562_, new_n5508_ );
and  ( new_n5580_, new_n5563_, new_n5507_ );
or   ( new_n5581_, new_n5580_, new_n5579_ );
and  ( new_n5582_, \d[10] , \a[4]  );
and  ( new_n5583_, new_n5560_, new_n5512_ );
and  ( new_n5584_, new_n5561_, new_n5511_ );
or   ( new_n5585_, new_n5584_, new_n5583_ );
and  ( new_n5586_, \d[9] , \a[5]  );
and  ( new_n5587_, new_n5558_, new_n5516_ );
and  ( new_n5588_, new_n5559_, new_n5515_ );
or   ( new_n5589_, new_n5588_, new_n5587_ );
and  ( new_n5590_, \d[8] , \a[6]  );
and  ( new_n5591_, new_n5556_, new_n5520_ );
and  ( new_n5592_, new_n5557_, new_n5519_ );
or   ( new_n5593_, new_n5592_, new_n5591_ );
and  ( new_n5594_, \d[7] , \a[7]  );
and  ( new_n5595_, new_n5554_, new_n5524_ );
and  ( new_n5596_, new_n5555_, new_n5523_ );
or   ( new_n5597_, new_n5596_, new_n5595_ );
and  ( new_n5598_, \d[6] , \a[8]  );
and  ( new_n5599_, new_n5552_, new_n5528_ );
and  ( new_n5600_, new_n5553_, new_n5527_ );
or   ( new_n5601_, new_n5600_, new_n5599_ );
and  ( new_n5602_, \d[5] , \a[9]  );
and  ( new_n5603_, new_n5550_, new_n5532_ );
and  ( new_n5604_, new_n5551_, new_n5531_ );
or   ( new_n5605_, new_n5604_, new_n5603_ );
and  ( new_n5606_, \d[4] , \a[10]  );
and  ( new_n5607_, new_n5548_, new_n5536_ );
and  ( new_n5608_, new_n5549_, new_n5535_ );
or   ( new_n5609_, new_n5608_, new_n5607_ );
and  ( new_n5610_, \d[3] , \a[11]  );
and  ( new_n5611_, new_n5546_, new_n5540_ );
and  ( new_n5612_, new_n5547_, new_n5539_ );
nor  ( new_n5613_, new_n5612_, new_n5611_ );
not  ( new_n5614_, new_n5613_ );
and  ( new_n5615_, \d[2] , \a[12]  );
and  ( new_n5616_, new_n5544_, new_n238_ );
and  ( new_n5617_, new_n5545_, new_n5543_ );
nor  ( new_n5618_, new_n5617_, new_n5616_ );
not  ( new_n5619_, new_n5618_ );
and  ( new_n5620_, \d[0] , \a[14]  );
xor  ( new_n5621_, new_n5620_, new_n93_ );
xor  ( new_n5622_, new_n5621_, new_n5619_ );
xor  ( new_n5623_, new_n5622_, new_n5615_ );
xor  ( new_n5624_, new_n5623_, new_n5614_ );
xor  ( new_n5625_, new_n5624_, new_n5610_ );
xor  ( new_n5626_, new_n5625_, new_n5609_ );
xor  ( new_n5627_, new_n5626_, new_n5606_ );
xor  ( new_n5628_, new_n5627_, new_n5605_ );
xor  ( new_n5629_, new_n5628_, new_n5602_ );
xor  ( new_n5630_, new_n5629_, new_n5601_ );
xor  ( new_n5631_, new_n5630_, new_n5598_ );
xor  ( new_n5632_, new_n5631_, new_n5597_ );
xor  ( new_n5633_, new_n5632_, new_n5594_ );
xor  ( new_n5634_, new_n5633_, new_n5593_ );
xor  ( new_n5635_, new_n5634_, new_n5590_ );
xor  ( new_n5636_, new_n5635_, new_n5589_ );
xor  ( new_n5637_, new_n5636_, new_n5586_ );
xor  ( new_n5638_, new_n5637_, new_n5585_ );
xor  ( new_n5639_, new_n5638_, new_n5582_ );
xor  ( new_n5640_, new_n5639_, new_n5581_ );
xor  ( new_n5641_, new_n5640_, new_n5578_ );
xor  ( new_n5642_, new_n5641_, new_n5577_ );
xor  ( new_n5643_, new_n5642_, new_n5574_ );
xor  ( new_n5644_, new_n5643_, new_n5573_ );
xor  ( new_n5645_, new_n5644_, new_n5570_ );
xor  ( new_n5646_, new_n5645_, new_n5569_ );
xnor ( new_n5647_, new_n5646_, new_n260_ );
and  ( new_n5648_, new_n5647_, new_n5098_ );
or   ( new_n5649_, \b[14] , \a[14]  );
and  ( new_n5650_, new_n5649_, new_n5102_ );
nor  ( new_n5651_, new_n5650_, new_n5648_ );
and  ( new_n5652_, new_n5651_, new_n5122_ );
and  ( new_n5653_, new_n5110_, \a[14]  );
and  ( new_n5654_, new_n5092_, \c[14]  );
nor  ( new_n5655_, new_n5654_, new_n5653_ );
and  ( new_n5656_, new_n5076_, new_n2200_ );
and  ( new_n5657_, new_n5080_, new_n2195_ );
nor  ( new_n5658_, new_n5657_, new_n5656_ );
and  ( new_n5659_, new_n5658_, new_n5655_ );
and  ( new_n5660_, new_n5659_, new_n5652_ );
and  ( new_n5661_, new_n5064_, \c[14]  );
nor  ( new_n5662_, new_n5661_, new_n5116_ );
nor  ( new_n5663_, new_n5662_, new_n2206_ );
not  ( new_n5664_, new_n5663_ );
and  ( new_n5665_, \c[8] , \b[0]  );
and  ( new_n5666_, new_n3198_, new_n1566_ );
and  ( new_n5667_, \c[0] , \b[2]  );
and  ( new_n5668_, new_n5667_, new_n3188_ );
xnor ( new_n5669_, new_n5668_, new_n5666_ );
or   ( new_n5670_, new_n5667_, new_n3188_ );
and  ( new_n5671_, new_n5670_, new_n5669_ );
and  ( new_n5672_, new_n5671_, new_n1548_ );
and  ( new_n5673_, \c[2] , \b[1]  );
or   ( new_n5674_, new_n5668_, new_n5666_ );
and  ( new_n5675_, \c[0] , \b[3]  );
xor  ( new_n5676_, new_n5675_, new_n1560_ );
xor  ( new_n5677_, new_n5676_, new_n5674_ );
xor  ( new_n5678_, new_n5677_, new_n5673_ );
xor  ( new_n5679_, new_n5678_, new_n5672_ );
and  ( new_n5680_, new_n5679_, new_n1550_ );
and  ( new_n5681_, \c[3] , \b[1]  );
and  ( new_n5682_, new_n5677_, new_n5673_ );
and  ( new_n5683_, new_n5678_, new_n5672_ );
or   ( new_n5684_, new_n5683_, new_n5682_ );
and  ( new_n5685_, new_n5675_, new_n1560_ );
and  ( new_n5686_, new_n5676_, new_n5674_ );
or   ( new_n5687_, new_n5686_, new_n5685_ );
and  ( new_n5688_, \c[0] , \b[4]  );
xor  ( new_n5689_, new_n5688_, new_n1530_ );
xor  ( new_n5690_, new_n5689_, new_n5687_ );
xor  ( new_n5691_, new_n5690_, new_n3150_ );
xor  ( new_n5692_, new_n5691_, new_n5684_ );
xor  ( new_n5693_, new_n5692_, new_n5681_ );
xor  ( new_n5694_, new_n5693_, new_n5680_ );
and  ( new_n5695_, new_n5694_, new_n1493_ );
and  ( new_n5696_, \c[4] , \b[1]  );
and  ( new_n5697_, new_n5692_, new_n5681_ );
and  ( new_n5698_, new_n5693_, new_n5680_ );
or   ( new_n5699_, new_n5698_, new_n5697_ );
and  ( new_n5700_, \c[3] , \b[2]  );
and  ( new_n5701_, new_n5690_, new_n3150_ );
and  ( new_n5702_, new_n5691_, new_n5684_ );
or   ( new_n5703_, new_n5702_, new_n5701_ );
and  ( new_n5704_, \c[2] , \b[3]  );
and  ( new_n5705_, new_n5688_, new_n1530_ );
and  ( new_n5706_, new_n5689_, new_n5687_ );
or   ( new_n5707_, new_n5706_, new_n5705_ );
and  ( new_n5708_, \c[0] , \b[5]  );
xor  ( new_n5709_, new_n5708_, new_n1513_ );
xor  ( new_n5710_, new_n5709_, new_n5707_ );
xor  ( new_n5711_, new_n5710_, new_n5704_ );
xor  ( new_n5712_, new_n5711_, new_n5703_ );
xor  ( new_n5713_, new_n5712_, new_n5700_ );
xor  ( new_n5714_, new_n5713_, new_n5699_ );
xor  ( new_n5715_, new_n5714_, new_n5696_ );
xor  ( new_n5716_, new_n5715_, new_n5695_ );
and  ( new_n5717_, new_n5716_, new_n1495_ );
and  ( new_n5718_, \c[5] , \b[1]  );
and  ( new_n5719_, new_n5714_, new_n5696_ );
and  ( new_n5720_, new_n5715_, new_n5695_ );
or   ( new_n5721_, new_n5720_, new_n5719_ );
and  ( new_n5722_, \c[4] , \b[2]  );
and  ( new_n5723_, new_n5712_, new_n5700_ );
and  ( new_n5724_, new_n5713_, new_n5699_ );
or   ( new_n5725_, new_n5724_, new_n5723_ );
and  ( new_n5726_, new_n5710_, new_n5704_ );
and  ( new_n5727_, new_n5711_, new_n5703_ );
or   ( new_n5728_, new_n5727_, new_n5726_ );
and  ( new_n5729_, \c[2] , \b[4]  );
and  ( new_n5730_, new_n5708_, new_n1513_ );
and  ( new_n5731_, new_n5709_, new_n5707_ );
or   ( new_n5732_, new_n5731_, new_n5730_ );
and  ( new_n5733_, \c[0] , \b[6]  );
xor  ( new_n5734_, new_n5733_, new_n1464_ );
xor  ( new_n5735_, new_n5734_, new_n5732_ );
xor  ( new_n5736_, new_n5735_, new_n5729_ );
xor  ( new_n5737_, new_n5736_, new_n5728_ );
xor  ( new_n5738_, new_n5737_, new_n2984_ );
xor  ( new_n5739_, new_n5738_, new_n5725_ );
xor  ( new_n5740_, new_n5739_, new_n5722_ );
xor  ( new_n5741_, new_n5740_, new_n5721_ );
xor  ( new_n5742_, new_n5741_, new_n5718_ );
xor  ( new_n5743_, new_n5742_, new_n5717_ );
and  ( new_n5744_, new_n5743_, new_n1415_ );
and  ( new_n5745_, \c[6] , \b[1]  );
and  ( new_n5746_, new_n5741_, new_n5718_ );
and  ( new_n5747_, new_n5742_, new_n5717_ );
or   ( new_n5748_, new_n5747_, new_n5746_ );
and  ( new_n5749_, \c[5] , \b[2]  );
and  ( new_n5750_, new_n5739_, new_n5722_ );
and  ( new_n5751_, new_n5740_, new_n5721_ );
or   ( new_n5752_, new_n5751_, new_n5750_ );
and  ( new_n5753_, \c[4] , \b[3]  );
and  ( new_n5754_, new_n5737_, new_n2984_ );
and  ( new_n5755_, new_n5738_, new_n5725_ );
or   ( new_n5756_, new_n5755_, new_n5754_ );
and  ( new_n5757_, \c[3] , \b[4]  );
and  ( new_n5758_, new_n5735_, new_n5729_ );
and  ( new_n5759_, new_n5736_, new_n5728_ );
or   ( new_n5760_, new_n5759_, new_n5758_ );
and  ( new_n5761_, \c[2] , \b[5]  );
and  ( new_n5762_, new_n5733_, new_n1464_ );
and  ( new_n5763_, new_n5734_, new_n5732_ );
or   ( new_n5764_, new_n5763_, new_n5762_ );
and  ( new_n5765_, \c[0] , \b[7]  );
xor  ( new_n5766_, new_n5765_, new_n1435_ );
xor  ( new_n5767_, new_n5766_, new_n5764_ );
xor  ( new_n5768_, new_n5767_, new_n5761_ );
xor  ( new_n5769_, new_n5768_, new_n5760_ );
xor  ( new_n5770_, new_n5769_, new_n5757_ );
xor  ( new_n5771_, new_n5770_, new_n5756_ );
xor  ( new_n5772_, new_n5771_, new_n5753_ );
xor  ( new_n5773_, new_n5772_, new_n5752_ );
xor  ( new_n5774_, new_n5773_, new_n5749_ );
xor  ( new_n5775_, new_n5774_, new_n5748_ );
xor  ( new_n5776_, new_n5775_, new_n5745_ );
xor  ( new_n5777_, new_n5776_, new_n5744_ );
and  ( new_n5778_, new_n5777_, new_n1282_ );
and  ( new_n5779_, \c[7] , \b[1]  );
and  ( new_n5780_, new_n5775_, new_n5745_ );
and  ( new_n5781_, new_n5776_, new_n5744_ );
or   ( new_n5782_, new_n5781_, new_n5780_ );
and  ( new_n5783_, \c[6] , \b[2]  );
and  ( new_n5784_, new_n5773_, new_n5749_ );
and  ( new_n5785_, new_n5774_, new_n5748_ );
or   ( new_n5786_, new_n5785_, new_n5784_ );
and  ( new_n5787_, \c[5] , \b[3]  );
and  ( new_n5788_, new_n5771_, new_n5753_ );
and  ( new_n5789_, new_n5772_, new_n5752_ );
or   ( new_n5790_, new_n5789_, new_n5788_ );
and  ( new_n5791_, \c[4] , \b[4]  );
and  ( new_n5792_, new_n5769_, new_n5757_ );
and  ( new_n5793_, new_n5770_, new_n5756_ );
or   ( new_n5794_, new_n5793_, new_n5792_ );
and  ( new_n5795_, \c[3] , \b[5]  );
and  ( new_n5796_, new_n5767_, new_n5761_ );
and  ( new_n5797_, new_n5768_, new_n5760_ );
or   ( new_n5798_, new_n5797_, new_n5796_ );
and  ( new_n5799_, \c[2] , \b[6]  );
and  ( new_n5800_, new_n5765_, new_n1435_ );
and  ( new_n5801_, new_n5766_, new_n5764_ );
or   ( new_n5802_, new_n5801_, new_n5800_ );
and  ( new_n5803_, \c[0] , \b[8]  );
xor  ( new_n5804_, new_n5803_, new_n1368_ );
xor  ( new_n5805_, new_n5804_, new_n5802_ );
xor  ( new_n5806_, new_n5805_, new_n5799_ );
xor  ( new_n5807_, new_n5806_, new_n5798_ );
xor  ( new_n5808_, new_n5807_, new_n5795_ );
xor  ( new_n5809_, new_n5808_, new_n5794_ );
xor  ( new_n5810_, new_n5809_, new_n5791_ );
xor  ( new_n5811_, new_n5810_, new_n5790_ );
xor  ( new_n5812_, new_n5811_, new_n5787_ );
xor  ( new_n5813_, new_n5812_, new_n5786_ );
xor  ( new_n5814_, new_n5813_, new_n5783_ );
xor  ( new_n5815_, new_n5814_, new_n5782_ );
xor  ( new_n5816_, new_n5815_, new_n5779_ );
xor  ( new_n5817_, new_n5816_, new_n5778_ );
and  ( new_n5818_, new_n5817_, new_n5665_ );
and  ( new_n5819_, \c[8] , \b[1]  );
and  ( new_n5820_, new_n5815_, new_n5779_ );
and  ( new_n5821_, new_n5816_, new_n5778_ );
or   ( new_n5822_, new_n5821_, new_n5820_ );
and  ( new_n5823_, \c[7] , \b[2]  );
and  ( new_n5824_, new_n5813_, new_n5783_ );
and  ( new_n5825_, new_n5814_, new_n5782_ );
or   ( new_n5826_, new_n5825_, new_n5824_ );
and  ( new_n5827_, \c[6] , \b[3]  );
and  ( new_n5828_, new_n5811_, new_n5787_ );
and  ( new_n5829_, new_n5812_, new_n5786_ );
or   ( new_n5830_, new_n5829_, new_n5828_ );
and  ( new_n5831_, \c[5] , \b[4]  );
and  ( new_n5832_, new_n5809_, new_n5791_ );
and  ( new_n5833_, new_n5810_, new_n5790_ );
or   ( new_n5834_, new_n5833_, new_n5832_ );
and  ( new_n5835_, \c[4] , \b[5]  );
and  ( new_n5836_, new_n5807_, new_n5795_ );
and  ( new_n5837_, new_n5808_, new_n5794_ );
or   ( new_n5838_, new_n5837_, new_n5836_ );
and  ( new_n5839_, \c[3] , \b[6]  );
and  ( new_n5840_, new_n5805_, new_n5799_ );
and  ( new_n5841_, new_n5806_, new_n5798_ );
or   ( new_n5842_, new_n5841_, new_n5840_ );
and  ( new_n5843_, \c[2] , \b[7]  );
and  ( new_n5844_, new_n5803_, new_n1368_ );
and  ( new_n5845_, new_n5804_, new_n5802_ );
or   ( new_n5846_, new_n5845_, new_n5844_ );
and  ( new_n5847_, \c[0] , \b[9]  );
xor  ( new_n5848_, new_n5847_, new_n1330_ );
xor  ( new_n5849_, new_n5848_, new_n5846_ );
xor  ( new_n5850_, new_n5849_, new_n5843_ );
xor  ( new_n5851_, new_n5850_, new_n5842_ );
xor  ( new_n5852_, new_n5851_, new_n5839_ );
xor  ( new_n5853_, new_n5852_, new_n5838_ );
xor  ( new_n5854_, new_n5853_, new_n5835_ );
xor  ( new_n5855_, new_n5854_, new_n5834_ );
xor  ( new_n5856_, new_n5855_, new_n5831_ );
xor  ( new_n5857_, new_n5856_, new_n5830_ );
xor  ( new_n5858_, new_n5857_, new_n5827_ );
xor  ( new_n5859_, new_n5858_, new_n5826_ );
xor  ( new_n5860_, new_n5859_, new_n5823_ );
xor  ( new_n5861_, new_n5860_, new_n5822_ );
xor  ( new_n5862_, new_n5861_, new_n5819_ );
xor  ( new_n5863_, new_n5862_, new_n5818_ );
and  ( new_n5864_, new_n5863_, new_n1130_ );
and  ( new_n5865_, \c[9] , \b[1]  );
and  ( new_n5866_, new_n5861_, new_n5819_ );
and  ( new_n5867_, new_n5862_, new_n5818_ );
or   ( new_n5868_, new_n5867_, new_n5866_ );
and  ( new_n5869_, \c[8] , \b[2]  );
and  ( new_n5870_, new_n5859_, new_n5823_ );
and  ( new_n5871_, new_n5860_, new_n5822_ );
or   ( new_n5872_, new_n5871_, new_n5870_ );
and  ( new_n5873_, \c[7] , \b[3]  );
and  ( new_n5874_, new_n5857_, new_n5827_ );
and  ( new_n5875_, new_n5858_, new_n5826_ );
or   ( new_n5876_, new_n5875_, new_n5874_ );
and  ( new_n5877_, \c[6] , \b[4]  );
and  ( new_n5878_, new_n5855_, new_n5831_ );
and  ( new_n5879_, new_n5856_, new_n5830_ );
or   ( new_n5880_, new_n5879_, new_n5878_ );
and  ( new_n5881_, \c[5] , \b[5]  );
and  ( new_n5882_, new_n5853_, new_n5835_ );
and  ( new_n5883_, new_n5854_, new_n5834_ );
or   ( new_n5884_, new_n5883_, new_n5882_ );
and  ( new_n5885_, \c[4] , \b[6]  );
and  ( new_n5886_, new_n5851_, new_n5839_ );
and  ( new_n5887_, new_n5852_, new_n5838_ );
or   ( new_n5888_, new_n5887_, new_n5886_ );
and  ( new_n5889_, \c[3] , \b[7]  );
and  ( new_n5890_, new_n5849_, new_n5843_ );
and  ( new_n5891_, new_n5850_, new_n5842_ );
or   ( new_n5892_, new_n5891_, new_n5890_ );
and  ( new_n5893_, \c[2] , \b[8]  );
and  ( new_n5894_, new_n5847_, new_n1330_ );
and  ( new_n5895_, new_n5848_, new_n5846_ );
or   ( new_n5896_, new_n5895_, new_n5894_ );
and  ( new_n5897_, \c[0] , \b[10]  );
xor  ( new_n5898_, new_n5897_, new_n1298_ );
xor  ( new_n5899_, new_n5898_, new_n5896_ );
xor  ( new_n5900_, new_n5899_, new_n5893_ );
xor  ( new_n5901_, new_n5900_, new_n5892_ );
xor  ( new_n5902_, new_n5901_, new_n5889_ );
xor  ( new_n5903_, new_n5902_, new_n5888_ );
xor  ( new_n5904_, new_n5903_, new_n5885_ );
xor  ( new_n5905_, new_n5904_, new_n5884_ );
xor  ( new_n5906_, new_n5905_, new_n5881_ );
xor  ( new_n5907_, new_n5906_, new_n5880_ );
xor  ( new_n5908_, new_n5907_, new_n5877_ );
xor  ( new_n5909_, new_n5908_, new_n5876_ );
xor  ( new_n5910_, new_n5909_, new_n5873_ );
xor  ( new_n5911_, new_n5910_, new_n5872_ );
xor  ( new_n5912_, new_n5911_, new_n5869_ );
xor  ( new_n5913_, new_n5912_, new_n5868_ );
xor  ( new_n5914_, new_n5913_, new_n5865_ );
xor  ( new_n5915_, new_n5914_, new_n5864_ );
and  ( new_n5916_, new_n5915_, new_n1204_ );
and  ( new_n5917_, \c[10] , \b[1]  );
and  ( new_n5918_, new_n5913_, new_n5865_ );
and  ( new_n5919_, new_n5914_, new_n5864_ );
or   ( new_n5920_, new_n5919_, new_n5918_ );
and  ( new_n5921_, \c[9] , \b[2]  );
and  ( new_n5922_, new_n5911_, new_n5869_ );
and  ( new_n5923_, new_n5912_, new_n5868_ );
or   ( new_n5924_, new_n5923_, new_n5922_ );
and  ( new_n5925_, \c[8] , \b[3]  );
and  ( new_n5926_, new_n5909_, new_n5873_ );
and  ( new_n5927_, new_n5910_, new_n5872_ );
or   ( new_n5928_, new_n5927_, new_n5926_ );
and  ( new_n5929_, \c[7] , \b[4]  );
and  ( new_n5930_, new_n5907_, new_n5877_ );
and  ( new_n5931_, new_n5908_, new_n5876_ );
or   ( new_n5932_, new_n5931_, new_n5930_ );
and  ( new_n5933_, \c[6] , \b[5]  );
and  ( new_n5934_, new_n5905_, new_n5881_ );
and  ( new_n5935_, new_n5906_, new_n5880_ );
or   ( new_n5936_, new_n5935_, new_n5934_ );
and  ( new_n5937_, \c[5] , \b[6]  );
and  ( new_n5938_, new_n5903_, new_n5885_ );
and  ( new_n5939_, new_n5904_, new_n5884_ );
or   ( new_n5940_, new_n5939_, new_n5938_ );
and  ( new_n5941_, \c[4] , \b[7]  );
and  ( new_n5942_, new_n5901_, new_n5889_ );
and  ( new_n5943_, new_n5902_, new_n5888_ );
or   ( new_n5944_, new_n5943_, new_n5942_ );
and  ( new_n5945_, \c[3] , \b[8]  );
and  ( new_n5946_, new_n5899_, new_n5893_ );
and  ( new_n5947_, new_n5900_, new_n5892_ );
or   ( new_n5948_, new_n5947_, new_n5946_ );
and  ( new_n5949_, \c[2] , \b[9]  );
and  ( new_n5950_, new_n5897_, new_n1298_ );
and  ( new_n5951_, new_n5898_, new_n5896_ );
or   ( new_n5952_, new_n5951_, new_n5950_ );
and  ( new_n5953_, \c[0] , \b[11]  );
xor  ( new_n5954_, new_n5953_, new_n1235_ );
xor  ( new_n5955_, new_n5954_, new_n5952_ );
xor  ( new_n5956_, new_n5955_, new_n5949_ );
xor  ( new_n5957_, new_n5956_, new_n5948_ );
xor  ( new_n5958_, new_n5957_, new_n5945_ );
xor  ( new_n5959_, new_n5958_, new_n5944_ );
xor  ( new_n5960_, new_n5959_, new_n5941_ );
xor  ( new_n5961_, new_n5960_, new_n5940_ );
xor  ( new_n5962_, new_n5961_, new_n5937_ );
xor  ( new_n5963_, new_n5962_, new_n5936_ );
xor  ( new_n5964_, new_n5963_, new_n5933_ );
xor  ( new_n5965_, new_n5964_, new_n5932_ );
xor  ( new_n5966_, new_n5965_, new_n5929_ );
xor  ( new_n5967_, new_n5966_, new_n5928_ );
xor  ( new_n5968_, new_n5967_, new_n5925_ );
xor  ( new_n5969_, new_n5968_, new_n5924_ );
xor  ( new_n5970_, new_n5969_, new_n5921_ );
xor  ( new_n5971_, new_n5970_, new_n5920_ );
xor  ( new_n5972_, new_n5971_, new_n5917_ );
xor  ( new_n5973_, new_n5972_, new_n5916_ );
and  ( new_n5974_, new_n5973_, new_n1206_ );
and  ( new_n5975_, \c[11] , \b[1]  );
and  ( new_n5976_, new_n5971_, new_n5917_ );
and  ( new_n5977_, new_n5972_, new_n5916_ );
or   ( new_n5978_, new_n5977_, new_n5976_ );
and  ( new_n5979_, \c[10] , \b[2]  );
and  ( new_n5980_, new_n5969_, new_n5921_ );
and  ( new_n5981_, new_n5970_, new_n5920_ );
or   ( new_n5982_, new_n5981_, new_n5980_ );
and  ( new_n5983_, \c[9] , \b[3]  );
and  ( new_n5984_, new_n5967_, new_n5925_ );
and  ( new_n5985_, new_n5968_, new_n5924_ );
or   ( new_n5986_, new_n5985_, new_n5984_ );
and  ( new_n5987_, \c[8] , \b[4]  );
and  ( new_n5988_, new_n5965_, new_n5929_ );
and  ( new_n5989_, new_n5966_, new_n5928_ );
or   ( new_n5990_, new_n5989_, new_n5988_ );
and  ( new_n5991_, \c[7] , \b[5]  );
and  ( new_n5992_, new_n5963_, new_n5933_ );
and  ( new_n5993_, new_n5964_, new_n5932_ );
or   ( new_n5994_, new_n5993_, new_n5992_ );
and  ( new_n5995_, \c[6] , \b[6]  );
and  ( new_n5996_, new_n5961_, new_n5937_ );
and  ( new_n5997_, new_n5962_, new_n5936_ );
or   ( new_n5998_, new_n5997_, new_n5996_ );
and  ( new_n5999_, \c[5] , \b[7]  );
and  ( new_n6000_, new_n5959_, new_n5941_ );
and  ( new_n6001_, new_n5960_, new_n5940_ );
or   ( new_n6002_, new_n6001_, new_n6000_ );
and  ( new_n6003_, \c[4] , \b[8]  );
and  ( new_n6004_, new_n5957_, new_n5945_ );
and  ( new_n6005_, new_n5958_, new_n5944_ );
or   ( new_n6006_, new_n6005_, new_n6004_ );
and  ( new_n6007_, \c[3] , \b[9]  );
and  ( new_n6008_, new_n5955_, new_n5949_ );
and  ( new_n6009_, new_n5956_, new_n5948_ );
or   ( new_n6010_, new_n6009_, new_n6008_ );
and  ( new_n6011_, \c[2] , \b[10]  );
and  ( new_n6012_, new_n5953_, new_n1235_ );
and  ( new_n6013_, new_n5954_, new_n5952_ );
or   ( new_n6014_, new_n6013_, new_n6012_ );
and  ( new_n6015_, \c[0] , \b[12]  );
xor  ( new_n6016_, new_n6015_, new_n1157_ );
xor  ( new_n6017_, new_n6016_, new_n6014_ );
xor  ( new_n6018_, new_n6017_, new_n6011_ );
xor  ( new_n6019_, new_n6018_, new_n6010_ );
xor  ( new_n6020_, new_n6019_, new_n6007_ );
xor  ( new_n6021_, new_n6020_, new_n6006_ );
xor  ( new_n6022_, new_n6021_, new_n6003_ );
xor  ( new_n6023_, new_n6022_, new_n6002_ );
xor  ( new_n6024_, new_n6023_, new_n5999_ );
xor  ( new_n6025_, new_n6024_, new_n5998_ );
xor  ( new_n6026_, new_n6025_, new_n5995_ );
xor  ( new_n6027_, new_n6026_, new_n5994_ );
xor  ( new_n6028_, new_n6027_, new_n5991_ );
xor  ( new_n6029_, new_n6028_, new_n5990_ );
xor  ( new_n6030_, new_n6029_, new_n5987_ );
xor  ( new_n6031_, new_n6030_, new_n5986_ );
xor  ( new_n6032_, new_n6031_, new_n5983_ );
xor  ( new_n6033_, new_n6032_, new_n5982_ );
xor  ( new_n6034_, new_n6033_, new_n5979_ );
xor  ( new_n6035_, new_n6034_, new_n5978_ );
xor  ( new_n6036_, new_n6035_, new_n5975_ );
xor  ( new_n6037_, new_n6036_, new_n5974_ );
and  ( new_n6038_, new_n6037_, new_n968_ );
and  ( new_n6039_, \c[12] , \b[1]  );
and  ( new_n6040_, new_n6035_, new_n5975_ );
and  ( new_n6041_, new_n6036_, new_n5974_ );
or   ( new_n6042_, new_n6041_, new_n6040_ );
and  ( new_n6043_, \c[11] , \b[2]  );
and  ( new_n6044_, new_n6033_, new_n5979_ );
and  ( new_n6045_, new_n6034_, new_n5978_ );
or   ( new_n6046_, new_n6045_, new_n6044_ );
and  ( new_n6047_, \c[10] , \b[3]  );
and  ( new_n6048_, new_n6031_, new_n5983_ );
and  ( new_n6049_, new_n6032_, new_n5982_ );
or   ( new_n6050_, new_n6049_, new_n6048_ );
and  ( new_n6051_, \c[9] , \b[4]  );
and  ( new_n6052_, new_n6029_, new_n5987_ );
and  ( new_n6053_, new_n6030_, new_n5986_ );
or   ( new_n6054_, new_n6053_, new_n6052_ );
and  ( new_n6055_, \c[8] , \b[5]  );
and  ( new_n6056_, new_n6027_, new_n5991_ );
and  ( new_n6057_, new_n6028_, new_n5990_ );
or   ( new_n6058_, new_n6057_, new_n6056_ );
and  ( new_n6059_, \c[7] , \b[6]  );
and  ( new_n6060_, new_n6025_, new_n5995_ );
and  ( new_n6061_, new_n6026_, new_n5994_ );
or   ( new_n6062_, new_n6061_, new_n6060_ );
and  ( new_n6063_, \c[6] , \b[7]  );
and  ( new_n6064_, new_n6023_, new_n5999_ );
and  ( new_n6065_, new_n6024_, new_n5998_ );
or   ( new_n6066_, new_n6065_, new_n6064_ );
and  ( new_n6067_, \c[5] , \b[8]  );
and  ( new_n6068_, new_n6021_, new_n6003_ );
and  ( new_n6069_, new_n6022_, new_n6002_ );
or   ( new_n6070_, new_n6069_, new_n6068_ );
and  ( new_n6071_, \c[4] , \b[9]  );
and  ( new_n6072_, new_n6019_, new_n6007_ );
and  ( new_n6073_, new_n6020_, new_n6006_ );
or   ( new_n6074_, new_n6073_, new_n6072_ );
and  ( new_n6075_, \c[3] , \b[10]  );
and  ( new_n6076_, new_n6017_, new_n6011_ );
and  ( new_n6077_, new_n6018_, new_n6010_ );
or   ( new_n6078_, new_n6077_, new_n6076_ );
and  ( new_n6079_, \c[2] , \b[11]  );
and  ( new_n6080_, new_n6015_, new_n1157_ );
and  ( new_n6081_, new_n6016_, new_n6014_ );
or   ( new_n6082_, new_n6081_, new_n6080_ );
and  ( new_n6083_, \c[0] , \b[13]  );
xor  ( new_n6084_, new_n6083_, new_n1106_ );
xor  ( new_n6085_, new_n6084_, new_n6082_ );
xor  ( new_n6086_, new_n6085_, new_n6079_ );
xor  ( new_n6087_, new_n6086_, new_n6078_ );
xor  ( new_n6088_, new_n6087_, new_n6075_ );
xor  ( new_n6089_, new_n6088_, new_n6074_ );
xor  ( new_n6090_, new_n6089_, new_n6071_ );
xor  ( new_n6091_, new_n6090_, new_n6070_ );
xor  ( new_n6092_, new_n6091_, new_n6067_ );
xor  ( new_n6093_, new_n6092_, new_n6066_ );
xor  ( new_n6094_, new_n6093_, new_n6063_ );
xor  ( new_n6095_, new_n6094_, new_n6062_ );
xor  ( new_n6096_, new_n6095_, new_n6059_ );
xor  ( new_n6097_, new_n6096_, new_n6058_ );
xor  ( new_n6098_, new_n6097_, new_n6055_ );
xor  ( new_n6099_, new_n6098_, new_n6054_ );
xor  ( new_n6100_, new_n6099_, new_n6051_ );
xor  ( new_n6101_, new_n6100_, new_n6050_ );
xor  ( new_n6102_, new_n6101_, new_n6047_ );
xor  ( new_n6103_, new_n6102_, new_n6046_ );
xor  ( new_n6104_, new_n6103_, new_n6043_ );
xor  ( new_n6105_, new_n6104_, new_n6042_ );
xor  ( new_n6106_, new_n6105_, new_n6039_ );
xor  ( new_n6107_, new_n6106_, new_n6038_ );
and  ( new_n6108_, new_n6107_, new_n972_ );
and  ( new_n6109_, \c[13] , \b[1]  );
and  ( new_n6110_, new_n6105_, new_n6039_ );
and  ( new_n6111_, new_n6106_, new_n6038_ );
or   ( new_n6112_, new_n6111_, new_n6110_ );
and  ( new_n6113_, \c[12] , \b[2]  );
and  ( new_n6114_, new_n6103_, new_n6043_ );
and  ( new_n6115_, new_n6104_, new_n6042_ );
or   ( new_n6116_, new_n6115_, new_n6114_ );
and  ( new_n6117_, \c[11] , \b[3]  );
and  ( new_n6118_, new_n6101_, new_n6047_ );
and  ( new_n6119_, new_n6102_, new_n6046_ );
or   ( new_n6120_, new_n6119_, new_n6118_ );
and  ( new_n6121_, \c[10] , \b[4]  );
and  ( new_n6122_, new_n6099_, new_n6051_ );
and  ( new_n6123_, new_n6100_, new_n6050_ );
or   ( new_n6124_, new_n6123_, new_n6122_ );
and  ( new_n6125_, \c[9] , \b[5]  );
and  ( new_n6126_, new_n6097_, new_n6055_ );
and  ( new_n6127_, new_n6098_, new_n6054_ );
or   ( new_n6128_, new_n6127_, new_n6126_ );
and  ( new_n6129_, \c[8] , \b[6]  );
and  ( new_n6130_, new_n6095_, new_n6059_ );
and  ( new_n6131_, new_n6096_, new_n6058_ );
or   ( new_n6132_, new_n6131_, new_n6130_ );
and  ( new_n6133_, \c[7] , \b[7]  );
and  ( new_n6134_, new_n6093_, new_n6063_ );
and  ( new_n6135_, new_n6094_, new_n6062_ );
or   ( new_n6136_, new_n6135_, new_n6134_ );
and  ( new_n6137_, \c[6] , \b[8]  );
and  ( new_n6138_, new_n6091_, new_n6067_ );
and  ( new_n6139_, new_n6092_, new_n6066_ );
or   ( new_n6140_, new_n6139_, new_n6138_ );
and  ( new_n6141_, \c[5] , \b[9]  );
and  ( new_n6142_, new_n6089_, new_n6071_ );
and  ( new_n6143_, new_n6090_, new_n6070_ );
or   ( new_n6144_, new_n6143_, new_n6142_ );
and  ( new_n6145_, \c[4] , \b[10]  );
and  ( new_n6146_, new_n6087_, new_n6075_ );
and  ( new_n6147_, new_n6088_, new_n6074_ );
or   ( new_n6148_, new_n6147_, new_n6146_ );
and  ( new_n6149_, \c[3] , \b[11]  );
and  ( new_n6150_, new_n6085_, new_n6079_ );
and  ( new_n6151_, new_n6086_, new_n6078_ );
nor  ( new_n6152_, new_n6151_, new_n6150_ );
not  ( new_n6153_, new_n6152_ );
and  ( new_n6154_, \c[2] , \b[12]  );
and  ( new_n6155_, new_n6083_, new_n1106_ );
and  ( new_n6156_, new_n6084_, new_n6082_ );
nor  ( new_n6157_, new_n6156_, new_n6155_ );
not  ( new_n6158_, new_n6157_ );
and  ( new_n6159_, \c[0] , \b[14]  );
xor  ( new_n6160_, new_n6159_, new_n1056_ );
xor  ( new_n6161_, new_n6160_, new_n6158_ );
xor  ( new_n6162_, new_n6161_, new_n6154_ );
xor  ( new_n6163_, new_n6162_, new_n6153_ );
xor  ( new_n6164_, new_n6163_, new_n6149_ );
xor  ( new_n6165_, new_n6164_, new_n6148_ );
xor  ( new_n6166_, new_n6165_, new_n6145_ );
xor  ( new_n6167_, new_n6166_, new_n6144_ );
xor  ( new_n6168_, new_n6167_, new_n6141_ );
xor  ( new_n6169_, new_n6168_, new_n6140_ );
xor  ( new_n6170_, new_n6169_, new_n6137_ );
xor  ( new_n6171_, new_n6170_, new_n6136_ );
xor  ( new_n6172_, new_n6171_, new_n6133_ );
xor  ( new_n6173_, new_n6172_, new_n6132_ );
xor  ( new_n6174_, new_n6173_, new_n6129_ );
xor  ( new_n6175_, new_n6174_, new_n6128_ );
xor  ( new_n6176_, new_n6175_, new_n6125_ );
xor  ( new_n6177_, new_n6176_, new_n6124_ );
xor  ( new_n6178_, new_n6177_, new_n6121_ );
xor  ( new_n6179_, new_n6178_, new_n6120_ );
xor  ( new_n6180_, new_n6179_, new_n6117_ );
xor  ( new_n6181_, new_n6180_, new_n6116_ );
xor  ( new_n6182_, new_n6181_, new_n6113_ );
xor  ( new_n6183_, new_n6182_, new_n6112_ );
xor  ( new_n6184_, new_n6183_, new_n6109_ );
xor  ( new_n6185_, new_n6184_, new_n6108_ );
xnor ( new_n6186_, new_n6185_, new_n1628_ );
and  ( new_n6187_, new_n6186_, new_n5052_ );
not  ( new_n6188_, new_n6187_ );
and  ( new_n6189_, new_n5072_, \d[14]  );
and  ( new_n6190_, new_n5056_, new_n2213_ );
nor  ( new_n6191_, new_n6190_, new_n6189_ );
and  ( new_n6192_, new_n6191_, new_n6188_ );
and  ( new_n6193_, new_n6192_, new_n5664_ );
and  ( new_n6194_, new_n6193_, new_n5660_ );
and  ( new_n6195_, new_n6194_, new_n5120_ );
or   ( new_n6196_, new_n6195_, new_n2906_ );
and  ( new_n6197_, new_n5056_, new_n3195_ );
not  ( new_n6198_, new_n6197_ );
and  ( new_n6199_, new_n5052_, new_n3199_ );
and  ( new_n6200_, new_n5083_, new_n3183_ );
nor  ( new_n6201_, new_n6200_, new_n6199_ );
and  ( new_n6202_, new_n6201_, new_n6198_ );
and  ( new_n6203_, new_n5064_, new_n3188_ );
and  ( new_n6204_, new_n5072_, \d[1]  );
nor  ( new_n6205_, new_n6204_, new_n6203_ );
and  ( new_n6206_, new_n5110_, \a[1]  );
and  ( new_n6207_, new_n5116_, \b[1]  );
nor  ( new_n6208_, new_n6207_, new_n6206_ );
and  ( new_n6209_, new_n6208_, new_n6205_ );
and  ( new_n6210_, new_n5092_, \c[1]  );
not  ( new_n6211_, new_n6210_ );
and  ( new_n6212_, new_n5098_, new_n3203_ );
and  ( new_n6213_, new_n5102_, new_n3192_ );
nor  ( new_n6214_, new_n6213_, new_n6212_ );
and  ( new_n6215_, new_n6214_, new_n6211_ );
and  ( new_n6216_, new_n5076_, new_n3208_ );
and  ( new_n6217_, new_n5080_, new_n3213_ );
nor  ( new_n6218_, new_n6217_, new_n6216_ );
and  ( new_n6219_, new_n6218_, new_n6215_ );
and  ( new_n6220_, new_n6219_, new_n6209_ );
and  ( new_n6221_, new_n6220_, new_n6202_ );
not  ( new_n6222_, new_n6221_ );
and  ( new_n6223_, new_n6222_, new_n2407_ );
and  ( new_n6224_, new_n6221_, new_n5120_ );
or   ( new_n6225_, new_n6224_, new_n3507_ );
and  ( new_n6226_, \c[0] , \b[0]  );
and  ( new_n6227_, new_n6226_, new_n5064_ );
not  ( new_n6228_, new_n6227_ );
and  ( new_n6229_, new_n5116_, \b[0]  );
and  ( new_n6230_, new_n5056_, new_n3547_ );
nor  ( new_n6231_, new_n6230_, new_n6229_ );
and  ( new_n6232_, new_n6231_, new_n6228_ );
and  ( new_n6233_, new_n5076_, new_n3480_ );
and  ( new_n6234_, new_n86_, new_n98_ );
not  ( new_n6235_, new_n6234_ );
and  ( new_n6236_, new_n5083_, new_n6235_ );
nor  ( new_n6237_, new_n6236_, new_n6233_ );
and  ( new_n6238_, new_n5072_, \d[0]  );
and  ( new_n6239_, new_n5110_, \a[0]  );
nor  ( new_n6240_, new_n6239_, new_n6238_ );
and  ( new_n6241_, new_n6240_, new_n6237_ );
and  ( new_n6242_, new_n5092_, \c[0]  );
not  ( new_n6243_, new_n6242_ );
or   ( new_n6244_, \b[0] , \a[0]  );
and  ( new_n6245_, new_n6244_, new_n5102_ );
and  ( new_n6246_, new_n5098_, new_n3477_ );
nor  ( new_n6247_, new_n6246_, new_n6245_ );
and  ( new_n6248_, new_n6247_, new_n6243_ );
and  ( new_n6249_, new_n6226_, new_n5052_ );
and  ( new_n6250_, new_n5080_, new_n3482_ );
nor  ( new_n6251_, new_n6250_, new_n6249_ );
and  ( new_n6252_, new_n6251_, new_n6248_ );
and  ( new_n6253_, new_n6252_, new_n6241_ );
and  ( new_n6254_, new_n6253_, new_n6232_ );
and  ( new_n6255_, new_n6254_, new_n5120_ );
or   ( new_n6256_, new_n6255_, new_n3406_ );
and  ( new_n6257_, new_n6256_, new_n6225_ );
not  ( new_n6258_, new_n6254_ );
and  ( new_n6259_, new_n6258_, new_n3407_ );
and  ( new_n6260_, new_n6222_, new_n4311_ );
and  ( new_n6261_, new_n6260_, new_n6259_ );
or   ( new_n6262_, new_n6261_, new_n6257_ );
or   ( new_n6263_, new_n3548_, new_n3507_ );
or   ( new_n6264_, new_n6263_, new_n6224_ );
or   ( new_n6265_, new_n6264_, new_n6255_ );
or   ( new_n6266_, new_n6265_, new_n6262_ );
or   ( new_n6267_, new_n6256_, new_n6225_ );
and  ( new_n6268_, new_n6267_, new_n6266_ );
and  ( new_n6269_, new_n6222_, new_n3407_ );
and  ( new_n6270_, new_n6258_, new_n4275_ );
and  ( new_n6271_, new_n6270_, new_n6269_ );
or   ( new_n6272_, new_n6224_, new_n3406_ );
or   ( new_n6273_, new_n6255_, new_n3306_ );
and  ( new_n6274_, new_n6273_, new_n6272_ );
or   ( new_n6275_, new_n6274_, new_n6271_ );
or   ( new_n6276_, new_n6275_, new_n6268_ );
or   ( new_n6277_, new_n6273_, new_n6272_ );
and  ( new_n6278_, new_n6277_, new_n6276_ );
or   ( new_n6279_, new_n6224_, new_n3306_ );
or   ( new_n6280_, new_n6255_, new_n3244_ );
and  ( new_n6281_, new_n6280_, new_n6279_ );
and  ( new_n6282_, new_n6222_, new_n4257_ );
and  ( new_n6283_, new_n6282_, new_n6270_ );
or   ( new_n6284_, new_n6283_, new_n6281_ );
or   ( new_n6285_, new_n6284_, new_n6278_ );
or   ( new_n6286_, new_n6280_, new_n6279_ );
and  ( new_n6287_, new_n6286_, new_n6285_ );
and  ( new_n6288_, new_n6258_, new_n3109_ );
and  ( new_n6289_, new_n6288_, new_n6282_ );
or   ( new_n6290_, new_n6224_, new_n3244_ );
or   ( new_n6291_, new_n6255_, new_n3108_ );
and  ( new_n6292_, new_n6291_, new_n6290_ );
or   ( new_n6293_, new_n6292_, new_n6289_ );
or   ( new_n6294_, new_n6293_, new_n6287_ );
or   ( new_n6295_, new_n6291_, new_n6290_ );
and  ( new_n6296_, new_n6295_, new_n6294_ );
or   ( new_n6297_, new_n6224_, new_n3108_ );
or   ( new_n6298_, new_n6255_, new_n3066_ );
and  ( new_n6299_, new_n6298_, new_n6297_ );
and  ( new_n6300_, new_n6222_, new_n4177_ );
and  ( new_n6301_, new_n6300_, new_n6288_ );
or   ( new_n6302_, new_n6301_, new_n6299_ );
or   ( new_n6303_, new_n6302_, new_n6296_ );
or   ( new_n6304_, new_n6298_, new_n6297_ );
and  ( new_n6305_, new_n6304_, new_n6303_ );
and  ( new_n6306_, new_n6258_, new_n2924_ );
and  ( new_n6307_, new_n6306_, new_n6300_ );
or   ( new_n6308_, new_n6224_, new_n3066_ );
or   ( new_n6309_, new_n6255_, new_n2923_ );
and  ( new_n6310_, new_n6309_, new_n6308_ );
or   ( new_n6311_, new_n6310_, new_n6307_ );
or   ( new_n6312_, new_n6311_, new_n6305_ );
or   ( new_n6313_, new_n6309_, new_n6308_ );
and  ( new_n6314_, new_n6313_, new_n6312_ );
or   ( new_n6315_, new_n6224_, new_n2923_ );
or   ( new_n6316_, new_n6255_, new_n2760_ );
and  ( new_n6317_, new_n6316_, new_n6315_ );
and  ( new_n6318_, new_n6222_, new_n4085_ );
and  ( new_n6319_, new_n6318_, new_n6306_ );
or   ( new_n6320_, new_n6319_, new_n6317_ );
or   ( new_n6321_, new_n6320_, new_n6314_ );
or   ( new_n6322_, new_n6316_, new_n6315_ );
and  ( new_n6323_, new_n6322_, new_n6321_ );
and  ( new_n6324_, new_n6258_, new_n4017_ );
and  ( new_n6325_, new_n6324_, new_n6318_ );
or   ( new_n6326_, new_n6224_, new_n2760_ );
or   ( new_n6327_, new_n6255_, new_n2723_ );
and  ( new_n6328_, new_n6327_, new_n6326_ );
or   ( new_n6329_, new_n6328_, new_n6325_ );
or   ( new_n6330_, new_n6329_, new_n6323_ );
or   ( new_n6331_, new_n6327_, new_n6326_ );
and  ( new_n6332_, new_n6331_, new_n6330_ );
or   ( new_n6333_, new_n6224_, new_n2723_ );
or   ( new_n6334_, new_n6255_, new_n2705_ );
and  ( new_n6335_, new_n6334_, new_n6333_ );
and  ( new_n6336_, new_n6222_, new_n3693_ );
and  ( new_n6337_, new_n6336_, new_n6324_ );
or   ( new_n6338_, new_n6337_, new_n6335_ );
or   ( new_n6339_, new_n6338_, new_n6332_ );
or   ( new_n6340_, new_n6334_, new_n6333_ );
and  ( new_n6341_, new_n6340_, new_n6339_ );
not  ( new_n6342_, new_n2566_ );
and  ( new_n6343_, new_n6258_, new_n6342_ );
and  ( new_n6344_, new_n6343_, new_n6336_ );
or   ( new_n6345_, new_n6224_, new_n2705_ );
or   ( new_n6346_, new_n6255_, new_n2566_ );
and  ( new_n6347_, new_n6346_, new_n6345_ );
or   ( new_n6348_, new_n6347_, new_n6344_ );
or   ( new_n6349_, new_n6348_, new_n6341_ );
or   ( new_n6350_, new_n6346_, new_n6345_ );
and  ( new_n6351_, new_n6350_, new_n6349_ );
or   ( new_n6352_, new_n6224_, new_n2566_ );
or   ( new_n6353_, new_n6255_, new_n2440_ );
and  ( new_n6354_, new_n6353_, new_n6352_ );
and  ( new_n6355_, new_n6222_, new_n2441_ );
and  ( new_n6356_, new_n6355_, new_n6343_ );
or   ( new_n6357_, new_n6356_, new_n6354_ );
or   ( new_n6358_, new_n6357_, new_n6351_ );
or   ( new_n6359_, new_n6353_, new_n6352_ );
and  ( new_n6360_, new_n6359_, new_n6358_ );
and  ( new_n6361_, new_n6258_, new_n3734_ );
and  ( new_n6362_, new_n6361_, new_n6355_ );
or   ( new_n6363_, new_n6224_, new_n2440_ );
or   ( new_n6364_, new_n6255_, new_n2304_ );
and  ( new_n6365_, new_n6364_, new_n6363_ );
or   ( new_n6366_, new_n6365_, new_n6362_ );
or   ( new_n6367_, new_n6366_, new_n6360_ );
or   ( new_n6368_, new_n6364_, new_n6363_ );
and  ( new_n6369_, new_n6368_, new_n6367_ );
or   ( new_n6370_, new_n6224_, new_n2304_ );
or   ( new_n6371_, new_n6255_, new_n2288_ );
and  ( new_n6372_, new_n6371_, new_n6370_ );
and  ( new_n6373_, new_n6222_, new_n2420_ );
and  ( new_n6374_, new_n6373_, new_n6361_ );
or   ( new_n6375_, new_n6374_, new_n6372_ );
or   ( new_n6376_, new_n6375_, new_n6369_ );
or   ( new_n6377_, new_n6371_, new_n6370_ );
and  ( new_n6378_, new_n6377_, new_n6376_ );
and  ( new_n6379_, new_n6258_, new_n3143_ );
and  ( new_n6380_, new_n6379_, new_n6373_ );
or   ( new_n6381_, new_n6224_, new_n2288_ );
or   ( new_n6382_, new_n6255_, new_n2297_ );
and  ( new_n6383_, new_n6382_, new_n6381_ );
or   ( new_n6384_, new_n6383_, new_n6380_ );
or   ( new_n6385_, new_n6384_, new_n6378_ );
or   ( new_n6386_, new_n6382_, new_n6381_ );
and  ( new_n6387_, new_n6386_, new_n6385_ );
or   ( new_n6388_, new_n6224_, new_n2297_ );
or   ( new_n6389_, new_n6255_, new_n2906_ );
and  ( new_n6390_, new_n6389_, new_n6388_ );
and  ( new_n6391_, new_n6379_, new_n6223_ );
or   ( new_n6392_, new_n6391_, new_n6390_ );
or   ( new_n6393_, new_n6392_, new_n6387_ );
or   ( new_n6394_, new_n6389_, new_n6388_ );
and  ( new_n6395_, new_n6394_, new_n6393_ );
and  ( new_n6396_, new_n6395_, new_n6223_ );
or   ( new_n6397_, new_n6224_, new_n2906_ );
and  ( new_n6398_, new_n6381_, new_n6379_ );
and  ( new_n6399_, new_n6382_, new_n6373_ );
or   ( new_n6400_, new_n6399_, new_n6398_ );
and  ( new_n6401_, new_n6363_, new_n6361_ );
and  ( new_n6402_, new_n6364_, new_n6355_ );
or   ( new_n6403_, new_n6402_, new_n6401_ );
and  ( new_n6404_, new_n6345_, new_n6343_ );
and  ( new_n6405_, new_n6346_, new_n6336_ );
or   ( new_n6406_, new_n6405_, new_n6404_ );
and  ( new_n6407_, new_n6326_, new_n6324_ );
and  ( new_n6408_, new_n6327_, new_n6318_ );
or   ( new_n6409_, new_n6408_, new_n6407_ );
and  ( new_n6410_, new_n6308_, new_n6306_ );
and  ( new_n6411_, new_n6309_, new_n6300_ );
or   ( new_n6412_, new_n6411_, new_n6410_ );
and  ( new_n6413_, new_n6290_, new_n6288_ );
and  ( new_n6414_, new_n6291_, new_n6282_ );
or   ( new_n6415_, new_n6414_, new_n6413_ );
and  ( new_n6416_, new_n6272_, new_n6270_ );
and  ( new_n6417_, new_n6273_, new_n6269_ );
or   ( new_n6418_, new_n6417_, new_n6416_ );
and  ( new_n6419_, new_n6259_, new_n6225_ );
and  ( new_n6420_, new_n6260_, new_n6256_ );
or   ( new_n6421_, new_n6420_, new_n6419_ );
and  ( new_n6422_, new_n6258_, new_n3547_ );
and  ( new_n6423_, new_n6422_, new_n6260_ );
and  ( new_n6424_, new_n6423_, new_n6421_ );
or   ( new_n6425_, new_n6424_, new_n6261_ );
and  ( new_n6426_, new_n6425_, new_n6418_ );
or   ( new_n6427_, new_n6426_, new_n6271_ );
and  ( new_n6428_, new_n6258_, new_n4257_ );
and  ( new_n6429_, new_n6428_, new_n6279_ );
and  ( new_n6430_, new_n6222_, new_n4275_ );
and  ( new_n6431_, new_n6430_, new_n6280_ );
or   ( new_n6432_, new_n6431_, new_n6429_ );
and  ( new_n6433_, new_n6432_, new_n6427_ );
or   ( new_n6434_, new_n6433_, new_n6283_ );
and  ( new_n6435_, new_n6434_, new_n6415_ );
or   ( new_n6436_, new_n6435_, new_n6289_ );
and  ( new_n6437_, new_n6258_, new_n4177_ );
and  ( new_n6438_, new_n6437_, new_n6297_ );
and  ( new_n6439_, new_n6222_, new_n3109_ );
and  ( new_n6440_, new_n6439_, new_n6298_ );
or   ( new_n6441_, new_n6440_, new_n6438_ );
and  ( new_n6442_, new_n6441_, new_n6436_ );
or   ( new_n6443_, new_n6442_, new_n6301_ );
and  ( new_n6444_, new_n6443_, new_n6412_ );
or   ( new_n6445_, new_n6444_, new_n6307_ );
and  ( new_n6446_, new_n6258_, new_n4085_ );
and  ( new_n6447_, new_n6446_, new_n6315_ );
and  ( new_n6448_, new_n6222_, new_n2924_ );
and  ( new_n6449_, new_n6448_, new_n6316_ );
or   ( new_n6450_, new_n6449_, new_n6447_ );
and  ( new_n6451_, new_n6450_, new_n6445_ );
or   ( new_n6452_, new_n6451_, new_n6319_ );
and  ( new_n6453_, new_n6452_, new_n6409_ );
or   ( new_n6454_, new_n6453_, new_n6325_ );
and  ( new_n6455_, new_n6258_, new_n3693_ );
and  ( new_n6456_, new_n6455_, new_n6333_ );
and  ( new_n6457_, new_n6222_, new_n4017_ );
and  ( new_n6458_, new_n6457_, new_n6334_ );
or   ( new_n6459_, new_n6458_, new_n6456_ );
and  ( new_n6460_, new_n6459_, new_n6454_ );
or   ( new_n6461_, new_n6460_, new_n6337_ );
and  ( new_n6462_, new_n6461_, new_n6406_ );
or   ( new_n6463_, new_n6462_, new_n6344_ );
and  ( new_n6464_, new_n6258_, new_n2441_ );
and  ( new_n6465_, new_n6464_, new_n6352_ );
and  ( new_n6466_, new_n6222_, new_n6342_ );
and  ( new_n6467_, new_n6466_, new_n6353_ );
or   ( new_n6468_, new_n6467_, new_n6465_ );
and  ( new_n6469_, new_n6468_, new_n6463_ );
or   ( new_n6470_, new_n6469_, new_n6356_ );
and  ( new_n6471_, new_n6470_, new_n6403_ );
or   ( new_n6472_, new_n6471_, new_n6362_ );
and  ( new_n6473_, new_n6258_, new_n2420_ );
and  ( new_n6474_, new_n6473_, new_n6370_ );
and  ( new_n6475_, new_n6222_, new_n3734_ );
and  ( new_n6476_, new_n6475_, new_n6371_ );
or   ( new_n6477_, new_n6476_, new_n6474_ );
and  ( new_n6478_, new_n6477_, new_n6472_ );
or   ( new_n6479_, new_n6478_, new_n6374_ );
and  ( new_n6480_, new_n6479_, new_n6400_ );
or   ( new_n6481_, new_n6480_, new_n6380_ );
and  ( new_n6482_, new_n6222_, new_n3143_ );
and  ( new_n6483_, new_n6482_, new_n6389_ );
and  ( new_n6484_, new_n6258_, new_n2407_ );
and  ( new_n6485_, new_n6484_, new_n6388_ );
or   ( new_n6486_, new_n6485_, new_n6483_ );
and  ( new_n6487_, new_n6486_, new_n6481_ );
or   ( new_n6488_, new_n6487_, new_n6391_ );
and  ( new_n6489_, new_n6488_, new_n6397_ );
or   ( new_n6490_, new_n6489_, new_n6396_ );
and  ( new_n6491_, new_n5110_, \a[2]  );
not  ( new_n6492_, new_n6491_ );
xor  ( new_n6493_, new_n5130_, new_n740_ );
and  ( new_n6494_, new_n6493_, new_n5098_ );
not  ( new_n6495_, new_n3152_ );
and  ( new_n6496_, new_n5102_, new_n6495_ );
nor  ( new_n6497_, new_n6496_, new_n6494_ );
and  ( new_n6498_, new_n6497_, new_n6492_ );
and  ( new_n6499_, new_n5092_, \c[2]  );
nand ( new_n6500_, new_n5075_, new_n5027_ );
nor  ( new_n6501_, new_n6500_, new_n3163_ );
nor  ( new_n6502_, new_n6501_, new_n6499_ );
nand ( new_n6503_, new_n5079_, new_n5027_ );
nor  ( new_n6504_, new_n6503_, new_n3166_ );
and  ( new_n6505_, new_n5056_, new_n3154_ );
nor  ( new_n6506_, new_n6505_, new_n6504_ );
and  ( new_n6507_, new_n6506_, new_n6502_ );
and  ( new_n6508_, new_n6507_, new_n6498_ );
and  ( new_n6509_, new_n5064_, \c[2]  );
nor  ( new_n6510_, new_n6509_, new_n5116_ );
nor  ( new_n6511_, new_n6510_, new_n865_ );
not  ( new_n6512_, new_n6511_ );
not  ( new_n6513_, new_n2093_ );
and  ( new_n6514_, new_n5083_, new_n6513_ );
not  ( new_n6515_, new_n6514_ );
xor  ( new_n6516_, new_n5671_, new_n1548_ );
and  ( new_n6517_, new_n6516_, new_n5052_ );
and  ( new_n6518_, new_n5072_, \d[2]  );
nor  ( new_n6519_, new_n6518_, new_n6517_ );
and  ( new_n6520_, new_n6519_, new_n6515_ );
and  ( new_n6521_, new_n6520_, new_n6512_ );
and  ( new_n6522_, new_n6521_, new_n6508_ );
not  ( new_n6523_, new_n6522_ );
and  ( new_n6524_, new_n6523_, new_n3143_ );
and  ( new_n6525_, new_n6524_, new_n6490_ );
and  ( new_n6526_, new_n6522_, new_n5120_ );
or   ( new_n6527_, new_n6526_, new_n2297_ );
and  ( new_n6528_, new_n6527_, new_n6490_ );
and  ( new_n6529_, new_n6488_, new_n6223_ );
and  ( new_n6530_, new_n6397_, new_n6393_ );
or   ( new_n6531_, new_n6530_, new_n6529_ );
and  ( new_n6532_, new_n6531_, new_n6524_ );
or   ( new_n6533_, new_n6532_, new_n6528_ );
and  ( new_n6534_, new_n6486_, new_n6387_ );
and  ( new_n6535_, new_n6481_, new_n6392_ );
or   ( new_n6536_, new_n6535_, new_n6534_ );
and  ( new_n6537_, new_n6523_, new_n2420_ );
and  ( new_n6538_, new_n6537_, new_n6536_ );
or   ( new_n6539_, new_n6526_, new_n2288_ );
and  ( new_n6540_, new_n6539_, new_n6536_ );
and  ( new_n6541_, new_n6392_, new_n6387_ );
or   ( new_n6542_, new_n6541_, new_n6487_ );
and  ( new_n6543_, new_n6542_, new_n6537_ );
or   ( new_n6544_, new_n6543_, new_n6540_ );
and  ( new_n6545_, new_n6400_, new_n6378_ );
and  ( new_n6546_, new_n6479_, new_n6384_ );
or   ( new_n6547_, new_n6546_, new_n6545_ );
and  ( new_n6548_, new_n6523_, new_n3734_ );
and  ( new_n6549_, new_n6548_, new_n6547_ );
or   ( new_n6550_, new_n6526_, new_n2304_ );
and  ( new_n6551_, new_n6550_, new_n6547_ );
and  ( new_n6552_, new_n6384_, new_n6378_ );
or   ( new_n6553_, new_n6552_, new_n6480_ );
and  ( new_n6554_, new_n6553_, new_n6548_ );
or   ( new_n6555_, new_n6554_, new_n6551_ );
and  ( new_n6556_, new_n6477_, new_n6369_ );
and  ( new_n6557_, new_n6472_, new_n6375_ );
or   ( new_n6558_, new_n6557_, new_n6556_ );
and  ( new_n6559_, new_n6523_, new_n2441_ );
and  ( new_n6560_, new_n6559_, new_n6558_ );
or   ( new_n6561_, new_n6526_, new_n2440_ );
and  ( new_n6562_, new_n6561_, new_n6558_ );
and  ( new_n6563_, new_n6375_, new_n6369_ );
or   ( new_n6564_, new_n6563_, new_n6478_ );
and  ( new_n6565_, new_n6564_, new_n6559_ );
or   ( new_n6566_, new_n6565_, new_n6562_ );
and  ( new_n6567_, new_n6403_, new_n6360_ );
and  ( new_n6568_, new_n6470_, new_n6366_ );
or   ( new_n6569_, new_n6568_, new_n6567_ );
and  ( new_n6570_, new_n6523_, new_n6342_ );
and  ( new_n6571_, new_n6570_, new_n6569_ );
or   ( new_n6572_, new_n6526_, new_n2566_ );
and  ( new_n6573_, new_n6572_, new_n6569_ );
and  ( new_n6574_, new_n6366_, new_n6360_ );
or   ( new_n6575_, new_n6574_, new_n6471_ );
and  ( new_n6576_, new_n6575_, new_n6570_ );
or   ( new_n6577_, new_n6576_, new_n6573_ );
and  ( new_n6578_, new_n6468_, new_n6351_ );
and  ( new_n6579_, new_n6463_, new_n6357_ );
or   ( new_n6580_, new_n6579_, new_n6578_ );
and  ( new_n6581_, new_n6523_, new_n3693_ );
and  ( new_n6582_, new_n6581_, new_n6580_ );
or   ( new_n6583_, new_n6526_, new_n2705_ );
and  ( new_n6584_, new_n6583_, new_n6580_ );
and  ( new_n6585_, new_n6357_, new_n6351_ );
or   ( new_n6586_, new_n6585_, new_n6469_ );
and  ( new_n6587_, new_n6586_, new_n6581_ );
or   ( new_n6588_, new_n6587_, new_n6584_ );
and  ( new_n6589_, new_n6406_, new_n6341_ );
and  ( new_n6590_, new_n6461_, new_n6348_ );
or   ( new_n6591_, new_n6590_, new_n6589_ );
and  ( new_n6592_, new_n6523_, new_n4017_ );
and  ( new_n6593_, new_n6592_, new_n6591_ );
or   ( new_n6594_, new_n6526_, new_n2723_ );
and  ( new_n6595_, new_n6594_, new_n6591_ );
and  ( new_n6596_, new_n6348_, new_n6341_ );
or   ( new_n6597_, new_n6596_, new_n6462_ );
and  ( new_n6598_, new_n6597_, new_n6592_ );
or   ( new_n6599_, new_n6598_, new_n6595_ );
and  ( new_n6600_, new_n6459_, new_n6332_ );
and  ( new_n6601_, new_n6454_, new_n6338_ );
or   ( new_n6602_, new_n6601_, new_n6600_ );
and  ( new_n6603_, new_n6523_, new_n4085_ );
and  ( new_n6604_, new_n6603_, new_n6602_ );
or   ( new_n6605_, new_n6526_, new_n2760_ );
and  ( new_n6606_, new_n6605_, new_n6602_ );
and  ( new_n6607_, new_n6338_, new_n6332_ );
or   ( new_n6608_, new_n6607_, new_n6460_ );
and  ( new_n6609_, new_n6608_, new_n6603_ );
or   ( new_n6610_, new_n6609_, new_n6606_ );
and  ( new_n6611_, new_n6409_, new_n6323_ );
and  ( new_n6612_, new_n6452_, new_n6329_ );
or   ( new_n6613_, new_n6612_, new_n6611_ );
and  ( new_n6614_, new_n6523_, new_n2924_ );
and  ( new_n6615_, new_n6614_, new_n6613_ );
or   ( new_n6616_, new_n6526_, new_n2923_ );
and  ( new_n6617_, new_n6616_, new_n6613_ );
and  ( new_n6618_, new_n6329_, new_n6323_ );
or   ( new_n6619_, new_n6618_, new_n6453_ );
and  ( new_n6620_, new_n6619_, new_n6614_ );
or   ( new_n6621_, new_n6620_, new_n6617_ );
and  ( new_n6622_, new_n6450_, new_n6314_ );
and  ( new_n6623_, new_n6445_, new_n6320_ );
or   ( new_n6624_, new_n6623_, new_n6622_ );
and  ( new_n6625_, new_n6523_, new_n4177_ );
and  ( new_n6626_, new_n6625_, new_n6624_ );
or   ( new_n6627_, new_n6526_, new_n3066_ );
and  ( new_n6628_, new_n6627_, new_n6624_ );
and  ( new_n6629_, new_n6320_, new_n6314_ );
or   ( new_n6630_, new_n6629_, new_n6451_ );
and  ( new_n6631_, new_n6630_, new_n6625_ );
or   ( new_n6632_, new_n6631_, new_n6628_ );
and  ( new_n6633_, new_n6412_, new_n6305_ );
and  ( new_n6634_, new_n6443_, new_n6311_ );
or   ( new_n6635_, new_n6634_, new_n6633_ );
and  ( new_n6636_, new_n6523_, new_n3109_ );
and  ( new_n6637_, new_n6636_, new_n6635_ );
or   ( new_n6638_, new_n6526_, new_n3108_ );
and  ( new_n6639_, new_n6638_, new_n6635_ );
and  ( new_n6640_, new_n6311_, new_n6305_ );
or   ( new_n6641_, new_n6640_, new_n6444_ );
and  ( new_n6642_, new_n6641_, new_n6636_ );
or   ( new_n6643_, new_n6642_, new_n6639_ );
and  ( new_n6644_, new_n6441_, new_n6296_ );
and  ( new_n6645_, new_n6436_, new_n6302_ );
or   ( new_n6646_, new_n6645_, new_n6644_ );
and  ( new_n6647_, new_n6523_, new_n4257_ );
and  ( new_n6648_, new_n6647_, new_n6646_ );
or   ( new_n6649_, new_n6526_, new_n3244_ );
and  ( new_n6650_, new_n6649_, new_n6646_ );
and  ( new_n6651_, new_n6302_, new_n6296_ );
or   ( new_n6652_, new_n6651_, new_n6442_ );
and  ( new_n6653_, new_n6652_, new_n6647_ );
or   ( new_n6654_, new_n6653_, new_n6650_ );
and  ( new_n6655_, new_n6415_, new_n6287_ );
and  ( new_n6656_, new_n6434_, new_n6293_ );
or   ( new_n6657_, new_n6656_, new_n6655_ );
and  ( new_n6658_, new_n6523_, new_n4275_ );
and  ( new_n6659_, new_n6658_, new_n6657_ );
or   ( new_n6660_, new_n6526_, new_n3306_ );
and  ( new_n6661_, new_n6660_, new_n6657_ );
and  ( new_n6662_, new_n6293_, new_n6287_ );
or   ( new_n6663_, new_n6662_, new_n6435_ );
and  ( new_n6664_, new_n6663_, new_n6658_ );
or   ( new_n6665_, new_n6664_, new_n6661_ );
and  ( new_n6666_, new_n6432_, new_n6278_ );
and  ( new_n6667_, new_n6427_, new_n6284_ );
or   ( new_n6668_, new_n6667_, new_n6666_ );
and  ( new_n6669_, new_n6523_, new_n3407_ );
and  ( new_n6670_, new_n6669_, new_n6668_ );
or   ( new_n6671_, new_n6526_, new_n3406_ );
and  ( new_n6672_, new_n6671_, new_n6668_ );
and  ( new_n6673_, new_n6284_, new_n6278_ );
or   ( new_n6674_, new_n6673_, new_n6433_ );
and  ( new_n6675_, new_n6674_, new_n6669_ );
or   ( new_n6676_, new_n6675_, new_n6672_ );
and  ( new_n6677_, new_n6418_, new_n6268_ );
and  ( new_n6678_, new_n6425_, new_n6275_ );
or   ( new_n6679_, new_n6678_, new_n6677_ );
and  ( new_n6680_, new_n6523_, new_n4311_ );
and  ( new_n6681_, new_n6680_, new_n6679_ );
and  ( new_n6682_, new_n6421_, new_n6265_ );
and  ( new_n6683_, new_n6423_, new_n6262_ );
or   ( new_n6684_, new_n6683_, new_n6682_ );
and  ( new_n6685_, new_n6523_, new_n3547_ );
and  ( new_n6686_, new_n6685_, new_n6684_ );
or   ( new_n6687_, new_n6526_, new_n3507_ );
and  ( new_n6688_, new_n6687_, new_n6679_ );
and  ( new_n6689_, new_n6275_, new_n6268_ );
or   ( new_n6690_, new_n6689_, new_n6426_ );
and  ( new_n6691_, new_n6690_, new_n6680_ );
or   ( new_n6692_, new_n6691_, new_n6688_ );
and  ( new_n6693_, new_n6692_, new_n6686_ );
or   ( new_n6694_, new_n6693_, new_n6681_ );
and  ( new_n6695_, new_n6694_, new_n6676_ );
or   ( new_n6696_, new_n6695_, new_n6670_ );
and  ( new_n6697_, new_n6696_, new_n6665_ );
or   ( new_n6698_, new_n6697_, new_n6659_ );
and  ( new_n6699_, new_n6698_, new_n6654_ );
or   ( new_n6700_, new_n6699_, new_n6648_ );
and  ( new_n6701_, new_n6700_, new_n6643_ );
or   ( new_n6702_, new_n6701_, new_n6637_ );
and  ( new_n6703_, new_n6702_, new_n6632_ );
or   ( new_n6704_, new_n6703_, new_n6626_ );
and  ( new_n6705_, new_n6704_, new_n6621_ );
or   ( new_n6706_, new_n6705_, new_n6615_ );
and  ( new_n6707_, new_n6706_, new_n6610_ );
or   ( new_n6708_, new_n6707_, new_n6604_ );
and  ( new_n6709_, new_n6708_, new_n6599_ );
or   ( new_n6710_, new_n6709_, new_n6593_ );
and  ( new_n6711_, new_n6710_, new_n6588_ );
or   ( new_n6712_, new_n6711_, new_n6582_ );
and  ( new_n6713_, new_n6712_, new_n6577_ );
or   ( new_n6714_, new_n6713_, new_n6571_ );
and  ( new_n6715_, new_n6714_, new_n6566_ );
or   ( new_n6716_, new_n6715_, new_n6560_ );
and  ( new_n6717_, new_n6716_, new_n6555_ );
or   ( new_n6718_, new_n6717_, new_n6549_ );
and  ( new_n6719_, new_n6718_, new_n6544_ );
or   ( new_n6720_, new_n6719_, new_n6538_ );
and  ( new_n6721_, new_n6720_, new_n6533_ );
or   ( new_n6722_, new_n6721_, new_n6525_ );
and  ( new_n6723_, new_n6529_, new_n6526_ );
or   ( new_n6724_, new_n6397_, new_n6395_ );
and  ( new_n6725_, new_n6523_, new_n2407_ );
and  ( new_n6726_, new_n6725_, new_n6724_ );
or   ( new_n6727_, new_n6726_, new_n6723_ );
and  ( new_n6728_, new_n6727_, new_n6722_ );
and  ( new_n6729_, new_n6529_, new_n6523_ );
or   ( new_n6730_, new_n6729_, new_n6728_ );
and  ( new_n6731_, new_n5083_, new_n2979_ );
not  ( new_n6732_, new_n6731_ );
xor  ( new_n6733_, new_n5138_, new_n742_ );
and  ( new_n6734_, new_n6733_, new_n5098_ );
and  ( new_n6735_, new_n5102_, new_n2988_ );
nor  ( new_n6736_, new_n6735_, new_n6734_ );
and  ( new_n6737_, new_n6736_, new_n6732_ );
and  ( new_n6738_, new_n5110_, \a[3]  );
and  ( new_n6739_, new_n5092_, \c[3]  );
nor  ( new_n6740_, new_n6739_, new_n6738_ );
and  ( new_n6741_, new_n5076_, new_n3004_ );
and  ( new_n6742_, new_n5080_, new_n3009_ );
nor  ( new_n6743_, new_n6742_, new_n6741_ );
and  ( new_n6744_, new_n6743_, new_n6740_ );
and  ( new_n6745_, new_n6744_, new_n6737_ );
and  ( new_n6746_, new_n5064_, \c[3]  );
nor  ( new_n6747_, new_n6746_, new_n5116_ );
nor  ( new_n6748_, new_n6747_, new_n815_ );
not  ( new_n6749_, new_n6748_ );
xor  ( new_n6750_, new_n5679_, new_n1550_ );
and  ( new_n6751_, new_n6750_, new_n5052_ );
not  ( new_n6752_, new_n6751_ );
and  ( new_n6753_, new_n5072_, \d[3]  );
and  ( new_n6754_, new_n5056_, new_n2991_ );
nor  ( new_n6755_, new_n6754_, new_n6753_ );
and  ( new_n6756_, new_n6755_, new_n6752_ );
and  ( new_n6757_, new_n6756_, new_n6749_ );
and  ( new_n6758_, new_n6757_, new_n6745_ );
not  ( new_n6759_, new_n6758_ );
and  ( new_n6760_, new_n6759_, new_n2407_ );
and  ( new_n6761_, new_n6760_, new_n6730_ );
and  ( new_n6762_, new_n6758_, new_n5120_ );
or   ( new_n6763_, new_n6762_, new_n2906_ );
and  ( new_n6764_, new_n6763_, new_n6730_ );
or   ( new_n6765_, new_n6531_, new_n6527_ );
or   ( new_n6766_, new_n6542_, new_n6539_ );
or   ( new_n6767_, new_n6553_, new_n6550_ );
or   ( new_n6768_, new_n6564_, new_n6561_ );
or   ( new_n6769_, new_n6575_, new_n6572_ );
or   ( new_n6770_, new_n6586_, new_n6583_ );
or   ( new_n6771_, new_n6597_, new_n6594_ );
or   ( new_n6772_, new_n6608_, new_n6605_ );
or   ( new_n6773_, new_n6619_, new_n6616_ );
or   ( new_n6774_, new_n6630_, new_n6627_ );
or   ( new_n6775_, new_n6641_, new_n6638_ );
or   ( new_n6776_, new_n6652_, new_n6649_ );
or   ( new_n6777_, new_n6663_, new_n6660_ );
or   ( new_n6778_, new_n6674_, new_n6671_ );
or   ( new_n6779_, new_n6690_, new_n6687_ );
and  ( new_n6780_, new_n6265_, new_n6262_ );
or   ( new_n6781_, new_n6780_, new_n6424_ );
or   ( new_n6782_, new_n6526_, new_n3548_ );
or   ( new_n6783_, new_n6782_, new_n6781_ );
and  ( new_n6784_, new_n6690_, new_n6687_ );
or   ( new_n6785_, new_n6784_, new_n6681_ );
or   ( new_n6786_, new_n6785_, new_n6783_ );
and  ( new_n6787_, new_n6786_, new_n6779_ );
and  ( new_n6788_, new_n6674_, new_n6671_ );
or   ( new_n6789_, new_n6788_, new_n6670_ );
or   ( new_n6790_, new_n6789_, new_n6787_ );
and  ( new_n6791_, new_n6790_, new_n6778_ );
and  ( new_n6792_, new_n6663_, new_n6660_ );
or   ( new_n6793_, new_n6792_, new_n6659_ );
or   ( new_n6794_, new_n6793_, new_n6791_ );
and  ( new_n6795_, new_n6794_, new_n6777_ );
and  ( new_n6796_, new_n6652_, new_n6649_ );
or   ( new_n6797_, new_n6796_, new_n6648_ );
or   ( new_n6798_, new_n6797_, new_n6795_ );
and  ( new_n6799_, new_n6798_, new_n6776_ );
and  ( new_n6800_, new_n6641_, new_n6638_ );
or   ( new_n6801_, new_n6800_, new_n6637_ );
or   ( new_n6802_, new_n6801_, new_n6799_ );
and  ( new_n6803_, new_n6802_, new_n6775_ );
and  ( new_n6804_, new_n6630_, new_n6627_ );
or   ( new_n6805_, new_n6804_, new_n6626_ );
or   ( new_n6806_, new_n6805_, new_n6803_ );
and  ( new_n6807_, new_n6806_, new_n6774_ );
and  ( new_n6808_, new_n6619_, new_n6616_ );
or   ( new_n6809_, new_n6808_, new_n6615_ );
or   ( new_n6810_, new_n6809_, new_n6807_ );
and  ( new_n6811_, new_n6810_, new_n6773_ );
and  ( new_n6812_, new_n6608_, new_n6605_ );
or   ( new_n6813_, new_n6812_, new_n6604_ );
or   ( new_n6814_, new_n6813_, new_n6811_ );
and  ( new_n6815_, new_n6814_, new_n6772_ );
and  ( new_n6816_, new_n6597_, new_n6594_ );
or   ( new_n6817_, new_n6816_, new_n6593_ );
or   ( new_n6818_, new_n6817_, new_n6815_ );
and  ( new_n6819_, new_n6818_, new_n6771_ );
and  ( new_n6820_, new_n6586_, new_n6583_ );
or   ( new_n6821_, new_n6820_, new_n6582_ );
or   ( new_n6822_, new_n6821_, new_n6819_ );
and  ( new_n6823_, new_n6822_, new_n6770_ );
and  ( new_n6824_, new_n6575_, new_n6572_ );
or   ( new_n6825_, new_n6824_, new_n6571_ );
or   ( new_n6826_, new_n6825_, new_n6823_ );
and  ( new_n6827_, new_n6826_, new_n6769_ );
and  ( new_n6828_, new_n6564_, new_n6561_ );
or   ( new_n6829_, new_n6828_, new_n6560_ );
or   ( new_n6830_, new_n6829_, new_n6827_ );
and  ( new_n6831_, new_n6830_, new_n6768_ );
and  ( new_n6832_, new_n6553_, new_n6550_ );
or   ( new_n6833_, new_n6832_, new_n6549_ );
or   ( new_n6834_, new_n6833_, new_n6831_ );
and  ( new_n6835_, new_n6834_, new_n6767_ );
and  ( new_n6836_, new_n6542_, new_n6539_ );
or   ( new_n6837_, new_n6836_, new_n6538_ );
or   ( new_n6838_, new_n6837_, new_n6835_ );
and  ( new_n6839_, new_n6838_, new_n6766_ );
and  ( new_n6840_, new_n6531_, new_n6527_ );
or   ( new_n6841_, new_n6840_, new_n6525_ );
or   ( new_n6842_, new_n6841_, new_n6839_ );
and  ( new_n6843_, new_n6842_, new_n6765_ );
or   ( new_n6844_, new_n6526_, new_n2906_ );
and  ( new_n6845_, new_n6844_, new_n6724_ );
or   ( new_n6846_, new_n6845_, new_n6729_ );
or   ( new_n6847_, new_n6846_, new_n6843_ );
or   ( new_n6848_, new_n6724_, new_n6526_ );
and  ( new_n6849_, new_n6848_, new_n6847_ );
and  ( new_n6850_, new_n6849_, new_n6760_ );
or   ( new_n6851_, new_n6850_, new_n6764_ );
and  ( new_n6852_, new_n6843_, new_n6727_ );
and  ( new_n6853_, new_n6846_, new_n6722_ );
or   ( new_n6854_, new_n6853_, new_n6852_ );
and  ( new_n6855_, new_n6759_, new_n3143_ );
and  ( new_n6856_, new_n6855_, new_n6854_ );
or   ( new_n6857_, new_n6762_, new_n2297_ );
and  ( new_n6858_, new_n6857_, new_n6854_ );
and  ( new_n6859_, new_n6846_, new_n6843_ );
or   ( new_n6860_, new_n6859_, new_n6728_ );
and  ( new_n6861_, new_n6860_, new_n6855_ );
or   ( new_n6862_, new_n6861_, new_n6858_ );
and  ( new_n6863_, new_n6839_, new_n6533_ );
and  ( new_n6864_, new_n6841_, new_n6720_ );
or   ( new_n6865_, new_n6864_, new_n6863_ );
and  ( new_n6866_, new_n6759_, new_n2420_ );
and  ( new_n6867_, new_n6866_, new_n6865_ );
or   ( new_n6868_, new_n6762_, new_n2288_ );
and  ( new_n6869_, new_n6868_, new_n6865_ );
and  ( new_n6870_, new_n6841_, new_n6839_ );
or   ( new_n6871_, new_n6870_, new_n6721_ );
and  ( new_n6872_, new_n6871_, new_n6866_ );
or   ( new_n6873_, new_n6872_, new_n6869_ );
and  ( new_n6874_, new_n6835_, new_n6544_ );
and  ( new_n6875_, new_n6837_, new_n6718_ );
or   ( new_n6876_, new_n6875_, new_n6874_ );
and  ( new_n6877_, new_n6759_, new_n3734_ );
and  ( new_n6878_, new_n6877_, new_n6876_ );
or   ( new_n6879_, new_n6762_, new_n2304_ );
and  ( new_n6880_, new_n6879_, new_n6876_ );
and  ( new_n6881_, new_n6837_, new_n6835_ );
or   ( new_n6882_, new_n6881_, new_n6719_ );
and  ( new_n6883_, new_n6882_, new_n6877_ );
or   ( new_n6884_, new_n6883_, new_n6880_ );
and  ( new_n6885_, new_n6831_, new_n6555_ );
and  ( new_n6886_, new_n6833_, new_n6716_ );
or   ( new_n6887_, new_n6886_, new_n6885_ );
and  ( new_n6888_, new_n6759_, new_n2441_ );
and  ( new_n6889_, new_n6888_, new_n6887_ );
or   ( new_n6890_, new_n6762_, new_n2440_ );
and  ( new_n6891_, new_n6890_, new_n6887_ );
and  ( new_n6892_, new_n6833_, new_n6831_ );
or   ( new_n6893_, new_n6892_, new_n6717_ );
and  ( new_n6894_, new_n6893_, new_n6888_ );
or   ( new_n6895_, new_n6894_, new_n6891_ );
and  ( new_n6896_, new_n6827_, new_n6566_ );
and  ( new_n6897_, new_n6829_, new_n6714_ );
or   ( new_n6898_, new_n6897_, new_n6896_ );
and  ( new_n6899_, new_n6759_, new_n6342_ );
and  ( new_n6900_, new_n6899_, new_n6898_ );
or   ( new_n6901_, new_n6762_, new_n2566_ );
and  ( new_n6902_, new_n6901_, new_n6898_ );
and  ( new_n6903_, new_n6829_, new_n6827_ );
or   ( new_n6904_, new_n6903_, new_n6715_ );
and  ( new_n6905_, new_n6904_, new_n6899_ );
or   ( new_n6906_, new_n6905_, new_n6902_ );
and  ( new_n6907_, new_n6823_, new_n6577_ );
and  ( new_n6908_, new_n6825_, new_n6712_ );
or   ( new_n6909_, new_n6908_, new_n6907_ );
and  ( new_n6910_, new_n6759_, new_n3693_ );
and  ( new_n6911_, new_n6910_, new_n6909_ );
or   ( new_n6912_, new_n6762_, new_n2705_ );
and  ( new_n6913_, new_n6912_, new_n6909_ );
and  ( new_n6914_, new_n6825_, new_n6823_ );
or   ( new_n6915_, new_n6914_, new_n6713_ );
and  ( new_n6916_, new_n6915_, new_n6910_ );
or   ( new_n6917_, new_n6916_, new_n6913_ );
and  ( new_n6918_, new_n6819_, new_n6588_ );
and  ( new_n6919_, new_n6821_, new_n6710_ );
or   ( new_n6920_, new_n6919_, new_n6918_ );
and  ( new_n6921_, new_n6759_, new_n4017_ );
and  ( new_n6922_, new_n6921_, new_n6920_ );
or   ( new_n6923_, new_n6762_, new_n2723_ );
and  ( new_n6924_, new_n6923_, new_n6920_ );
and  ( new_n6925_, new_n6821_, new_n6819_ );
or   ( new_n6926_, new_n6925_, new_n6711_ );
and  ( new_n6927_, new_n6926_, new_n6921_ );
or   ( new_n6928_, new_n6927_, new_n6924_ );
and  ( new_n6929_, new_n6815_, new_n6599_ );
and  ( new_n6930_, new_n6817_, new_n6708_ );
or   ( new_n6931_, new_n6930_, new_n6929_ );
and  ( new_n6932_, new_n6759_, new_n4085_ );
and  ( new_n6933_, new_n6932_, new_n6931_ );
or   ( new_n6934_, new_n6762_, new_n2760_ );
and  ( new_n6935_, new_n6934_, new_n6931_ );
and  ( new_n6936_, new_n6817_, new_n6815_ );
or   ( new_n6937_, new_n6936_, new_n6709_ );
and  ( new_n6938_, new_n6937_, new_n6932_ );
or   ( new_n6939_, new_n6938_, new_n6935_ );
and  ( new_n6940_, new_n6811_, new_n6610_ );
and  ( new_n6941_, new_n6813_, new_n6706_ );
or   ( new_n6942_, new_n6941_, new_n6940_ );
and  ( new_n6943_, new_n6759_, new_n2924_ );
and  ( new_n6944_, new_n6943_, new_n6942_ );
or   ( new_n6945_, new_n6762_, new_n2923_ );
and  ( new_n6946_, new_n6945_, new_n6942_ );
and  ( new_n6947_, new_n6813_, new_n6811_ );
or   ( new_n6948_, new_n6947_, new_n6707_ );
and  ( new_n6949_, new_n6948_, new_n6943_ );
or   ( new_n6950_, new_n6949_, new_n6946_ );
and  ( new_n6951_, new_n6807_, new_n6621_ );
and  ( new_n6952_, new_n6809_, new_n6704_ );
or   ( new_n6953_, new_n6952_, new_n6951_ );
and  ( new_n6954_, new_n6759_, new_n4177_ );
and  ( new_n6955_, new_n6954_, new_n6953_ );
or   ( new_n6956_, new_n6762_, new_n3066_ );
and  ( new_n6957_, new_n6956_, new_n6953_ );
and  ( new_n6958_, new_n6809_, new_n6807_ );
or   ( new_n6959_, new_n6958_, new_n6705_ );
and  ( new_n6960_, new_n6959_, new_n6954_ );
or   ( new_n6961_, new_n6960_, new_n6957_ );
and  ( new_n6962_, new_n6803_, new_n6632_ );
and  ( new_n6963_, new_n6805_, new_n6702_ );
or   ( new_n6964_, new_n6963_, new_n6962_ );
and  ( new_n6965_, new_n6759_, new_n3109_ );
and  ( new_n6966_, new_n6965_, new_n6964_ );
or   ( new_n6967_, new_n6762_, new_n3108_ );
and  ( new_n6968_, new_n6967_, new_n6964_ );
and  ( new_n6969_, new_n6805_, new_n6803_ );
or   ( new_n6970_, new_n6969_, new_n6703_ );
and  ( new_n6971_, new_n6970_, new_n6965_ );
or   ( new_n6972_, new_n6971_, new_n6968_ );
and  ( new_n6973_, new_n6799_, new_n6643_ );
and  ( new_n6974_, new_n6801_, new_n6700_ );
or   ( new_n6975_, new_n6974_, new_n6973_ );
and  ( new_n6976_, new_n6759_, new_n4257_ );
and  ( new_n6977_, new_n6976_, new_n6975_ );
or   ( new_n6978_, new_n6762_, new_n3244_ );
and  ( new_n6979_, new_n6978_, new_n6975_ );
and  ( new_n6980_, new_n6801_, new_n6799_ );
or   ( new_n6981_, new_n6980_, new_n6701_ );
and  ( new_n6982_, new_n6981_, new_n6976_ );
or   ( new_n6983_, new_n6982_, new_n6979_ );
and  ( new_n6984_, new_n6795_, new_n6654_ );
and  ( new_n6985_, new_n6797_, new_n6698_ );
or   ( new_n6986_, new_n6985_, new_n6984_ );
and  ( new_n6987_, new_n6759_, new_n4275_ );
and  ( new_n6988_, new_n6987_, new_n6986_ );
or   ( new_n6989_, new_n6762_, new_n3306_ );
and  ( new_n6990_, new_n6989_, new_n6986_ );
and  ( new_n6991_, new_n6797_, new_n6795_ );
or   ( new_n6992_, new_n6991_, new_n6699_ );
and  ( new_n6993_, new_n6992_, new_n6987_ );
or   ( new_n6994_, new_n6993_, new_n6990_ );
and  ( new_n6995_, new_n6791_, new_n6665_ );
and  ( new_n6996_, new_n6793_, new_n6696_ );
or   ( new_n6997_, new_n6996_, new_n6995_ );
and  ( new_n6998_, new_n6759_, new_n3407_ );
and  ( new_n6999_, new_n6998_, new_n6997_ );
or   ( new_n7000_, new_n6762_, new_n3406_ );
and  ( new_n7001_, new_n7000_, new_n6997_ );
and  ( new_n7002_, new_n6793_, new_n6791_ );
or   ( new_n7003_, new_n7002_, new_n6697_ );
and  ( new_n7004_, new_n7003_, new_n6998_ );
or   ( new_n7005_, new_n7004_, new_n7001_ );
and  ( new_n7006_, new_n6787_, new_n6676_ );
and  ( new_n7007_, new_n6789_, new_n6694_ );
or   ( new_n7008_, new_n7007_, new_n7006_ );
and  ( new_n7009_, new_n6759_, new_n4311_ );
and  ( new_n7010_, new_n7009_, new_n7008_ );
and  ( new_n7011_, new_n6783_, new_n6692_ );
and  ( new_n7012_, new_n6785_, new_n6686_ );
or   ( new_n7013_, new_n7012_, new_n7011_ );
and  ( new_n7014_, new_n6759_, new_n3547_ );
and  ( new_n7015_, new_n7014_, new_n7013_ );
or   ( new_n7016_, new_n6762_, new_n3507_ );
and  ( new_n7017_, new_n7016_, new_n7008_ );
and  ( new_n7018_, new_n6789_, new_n6787_ );
or   ( new_n7019_, new_n7018_, new_n6695_ );
and  ( new_n7020_, new_n7019_, new_n7009_ );
or   ( new_n7021_, new_n7020_, new_n7017_ );
and  ( new_n7022_, new_n7021_, new_n7015_ );
or   ( new_n7023_, new_n7022_, new_n7010_ );
and  ( new_n7024_, new_n7023_, new_n7005_ );
or   ( new_n7025_, new_n7024_, new_n6999_ );
and  ( new_n7026_, new_n7025_, new_n6994_ );
or   ( new_n7027_, new_n7026_, new_n6988_ );
and  ( new_n7028_, new_n7027_, new_n6983_ );
or   ( new_n7029_, new_n7028_, new_n6977_ );
and  ( new_n7030_, new_n7029_, new_n6972_ );
or   ( new_n7031_, new_n7030_, new_n6966_ );
and  ( new_n7032_, new_n7031_, new_n6961_ );
or   ( new_n7033_, new_n7032_, new_n6955_ );
and  ( new_n7034_, new_n7033_, new_n6950_ );
or   ( new_n7035_, new_n7034_, new_n6944_ );
and  ( new_n7036_, new_n7035_, new_n6939_ );
or   ( new_n7037_, new_n7036_, new_n6933_ );
and  ( new_n7038_, new_n7037_, new_n6928_ );
or   ( new_n7039_, new_n7038_, new_n6922_ );
and  ( new_n7040_, new_n7039_, new_n6917_ );
or   ( new_n7041_, new_n7040_, new_n6911_ );
and  ( new_n7042_, new_n7041_, new_n6906_ );
or   ( new_n7043_, new_n7042_, new_n6900_ );
and  ( new_n7044_, new_n7043_, new_n6895_ );
or   ( new_n7045_, new_n7044_, new_n6889_ );
and  ( new_n7046_, new_n7045_, new_n6884_ );
or   ( new_n7047_, new_n7046_, new_n6878_ );
and  ( new_n7048_, new_n7047_, new_n6873_ );
or   ( new_n7049_, new_n7048_, new_n6867_ );
and  ( new_n7050_, new_n7049_, new_n6862_ );
or   ( new_n7051_, new_n7050_, new_n6856_ );
and  ( new_n7052_, new_n7051_, new_n6851_ );
or   ( new_n7053_, new_n7052_, new_n6761_ );
not  ( new_n7054_, new_n2105_ );
and  ( new_n7055_, new_n5083_, new_n7054_ );
not  ( new_n7056_, new_n7055_ );
xor  ( new_n7057_, new_n5154_, new_n685_ );
and  ( new_n7058_, new_n7057_, new_n5098_ );
or   ( new_n7059_, \b[4] , \a[4]  );
and  ( new_n7060_, new_n7059_, new_n5102_ );
nor  ( new_n7061_, new_n7060_, new_n7058_ );
and  ( new_n7062_, new_n7061_, new_n7056_ );
and  ( new_n7063_, new_n5110_, \a[4]  );
and  ( new_n7064_, new_n5092_, \c[4]  );
nor  ( new_n7065_, new_n7064_, new_n7063_ );
nor  ( new_n7066_, new_n6500_, new_n2962_ );
nor  ( new_n7067_, new_n6503_, new_n2965_ );
nor  ( new_n7068_, new_n7067_, new_n7066_ );
and  ( new_n7069_, new_n7068_, new_n7065_ );
and  ( new_n7070_, new_n7069_, new_n7062_ );
and  ( new_n7071_, new_n5064_, \c[4]  );
nor  ( new_n7072_, new_n7071_, new_n5116_ );
nor  ( new_n7073_, new_n7072_, new_n832_ );
not  ( new_n7074_, new_n7073_ );
xor  ( new_n7075_, new_n5694_, new_n1493_ );
and  ( new_n7076_, new_n7075_, new_n5052_ );
not  ( new_n7077_, new_n7076_ );
and  ( new_n7078_, new_n5072_, \d[4]  );
and  ( new_n7079_, new_n5056_, new_n2953_ );
nor  ( new_n7080_, new_n7079_, new_n7078_ );
and  ( new_n7081_, new_n7080_, new_n7077_ );
and  ( new_n7082_, new_n7081_, new_n7074_ );
and  ( new_n7083_, new_n7082_, new_n7070_ );
not  ( new_n7084_, new_n7083_ );
and  ( new_n7085_, new_n7084_, new_n2407_ );
and  ( new_n7086_, new_n7085_, new_n7053_ );
and  ( new_n7087_, new_n7083_, new_n5120_ );
or   ( new_n7088_, new_n7087_, new_n2906_ );
and  ( new_n7089_, new_n7088_, new_n7053_ );
or   ( new_n7090_, new_n6849_, new_n6763_ );
or   ( new_n7091_, new_n6860_, new_n6857_ );
or   ( new_n7092_, new_n6871_, new_n6868_ );
or   ( new_n7093_, new_n6882_, new_n6879_ );
or   ( new_n7094_, new_n6893_, new_n6890_ );
or   ( new_n7095_, new_n6904_, new_n6901_ );
or   ( new_n7096_, new_n6915_, new_n6912_ );
or   ( new_n7097_, new_n6926_, new_n6923_ );
or   ( new_n7098_, new_n6937_, new_n6934_ );
or   ( new_n7099_, new_n6948_, new_n6945_ );
or   ( new_n7100_, new_n6959_, new_n6956_ );
or   ( new_n7101_, new_n6970_, new_n6967_ );
or   ( new_n7102_, new_n6981_, new_n6978_ );
or   ( new_n7103_, new_n6992_, new_n6989_ );
or   ( new_n7104_, new_n7003_, new_n7000_ );
or   ( new_n7105_, new_n7019_, new_n7016_ );
and  ( new_n7106_, new_n6785_, new_n6783_ );
or   ( new_n7107_, new_n7106_, new_n6693_ );
or   ( new_n7108_, new_n6762_, new_n3548_ );
or   ( new_n7109_, new_n7108_, new_n7107_ );
and  ( new_n7110_, new_n7019_, new_n7016_ );
or   ( new_n7111_, new_n7110_, new_n7010_ );
or   ( new_n7112_, new_n7111_, new_n7109_ );
and  ( new_n7113_, new_n7112_, new_n7105_ );
and  ( new_n7114_, new_n7003_, new_n7000_ );
or   ( new_n7115_, new_n7114_, new_n6999_ );
or   ( new_n7116_, new_n7115_, new_n7113_ );
and  ( new_n7117_, new_n7116_, new_n7104_ );
and  ( new_n7118_, new_n6992_, new_n6989_ );
or   ( new_n7119_, new_n7118_, new_n6988_ );
or   ( new_n7120_, new_n7119_, new_n7117_ );
and  ( new_n7121_, new_n7120_, new_n7103_ );
and  ( new_n7122_, new_n6981_, new_n6978_ );
or   ( new_n7123_, new_n7122_, new_n6977_ );
or   ( new_n7124_, new_n7123_, new_n7121_ );
and  ( new_n7125_, new_n7124_, new_n7102_ );
and  ( new_n7126_, new_n6970_, new_n6967_ );
or   ( new_n7127_, new_n7126_, new_n6966_ );
or   ( new_n7128_, new_n7127_, new_n7125_ );
and  ( new_n7129_, new_n7128_, new_n7101_ );
and  ( new_n7130_, new_n6959_, new_n6956_ );
or   ( new_n7131_, new_n7130_, new_n6955_ );
or   ( new_n7132_, new_n7131_, new_n7129_ );
and  ( new_n7133_, new_n7132_, new_n7100_ );
and  ( new_n7134_, new_n6948_, new_n6945_ );
or   ( new_n7135_, new_n7134_, new_n6944_ );
or   ( new_n7136_, new_n7135_, new_n7133_ );
and  ( new_n7137_, new_n7136_, new_n7099_ );
and  ( new_n7138_, new_n6937_, new_n6934_ );
or   ( new_n7139_, new_n7138_, new_n6933_ );
or   ( new_n7140_, new_n7139_, new_n7137_ );
and  ( new_n7141_, new_n7140_, new_n7098_ );
and  ( new_n7142_, new_n6926_, new_n6923_ );
or   ( new_n7143_, new_n7142_, new_n6922_ );
or   ( new_n7144_, new_n7143_, new_n7141_ );
and  ( new_n7145_, new_n7144_, new_n7097_ );
and  ( new_n7146_, new_n6915_, new_n6912_ );
or   ( new_n7147_, new_n7146_, new_n6911_ );
or   ( new_n7148_, new_n7147_, new_n7145_ );
and  ( new_n7149_, new_n7148_, new_n7096_ );
and  ( new_n7150_, new_n6904_, new_n6901_ );
or   ( new_n7151_, new_n7150_, new_n6900_ );
or   ( new_n7152_, new_n7151_, new_n7149_ );
and  ( new_n7153_, new_n7152_, new_n7095_ );
and  ( new_n7154_, new_n6893_, new_n6890_ );
or   ( new_n7155_, new_n7154_, new_n6889_ );
or   ( new_n7156_, new_n7155_, new_n7153_ );
and  ( new_n7157_, new_n7156_, new_n7094_ );
and  ( new_n7158_, new_n6882_, new_n6879_ );
or   ( new_n7159_, new_n7158_, new_n6878_ );
or   ( new_n7160_, new_n7159_, new_n7157_ );
and  ( new_n7161_, new_n7160_, new_n7093_ );
and  ( new_n7162_, new_n6871_, new_n6868_ );
or   ( new_n7163_, new_n7162_, new_n6867_ );
or   ( new_n7164_, new_n7163_, new_n7161_ );
and  ( new_n7165_, new_n7164_, new_n7092_ );
and  ( new_n7166_, new_n6860_, new_n6857_ );
or   ( new_n7167_, new_n7166_, new_n6856_ );
or   ( new_n7168_, new_n7167_, new_n7165_ );
and  ( new_n7169_, new_n7168_, new_n7091_ );
and  ( new_n7170_, new_n6849_, new_n6763_ );
or   ( new_n7171_, new_n7170_, new_n6761_ );
or   ( new_n7172_, new_n7171_, new_n7169_ );
and  ( new_n7173_, new_n7172_, new_n7090_ );
and  ( new_n7174_, new_n7173_, new_n7085_ );
or   ( new_n7175_, new_n7174_, new_n7089_ );
and  ( new_n7176_, new_n7169_, new_n6851_ );
and  ( new_n7177_, new_n7171_, new_n7051_ );
or   ( new_n7178_, new_n7177_, new_n7176_ );
and  ( new_n7179_, new_n7084_, new_n3143_ );
and  ( new_n7180_, new_n7179_, new_n7178_ );
or   ( new_n7181_, new_n7087_, new_n2297_ );
and  ( new_n7182_, new_n7181_, new_n7178_ );
and  ( new_n7183_, new_n7171_, new_n7169_ );
or   ( new_n7184_, new_n7183_, new_n7052_ );
and  ( new_n7185_, new_n7184_, new_n7179_ );
or   ( new_n7186_, new_n7185_, new_n7182_ );
and  ( new_n7187_, new_n7165_, new_n6862_ );
and  ( new_n7188_, new_n7167_, new_n7049_ );
or   ( new_n7189_, new_n7188_, new_n7187_ );
and  ( new_n7190_, new_n7084_, new_n2420_ );
and  ( new_n7191_, new_n7190_, new_n7189_ );
or   ( new_n7192_, new_n7087_, new_n2288_ );
and  ( new_n7193_, new_n7192_, new_n7189_ );
and  ( new_n7194_, new_n7167_, new_n7165_ );
or   ( new_n7195_, new_n7194_, new_n7050_ );
and  ( new_n7196_, new_n7195_, new_n7190_ );
or   ( new_n7197_, new_n7196_, new_n7193_ );
and  ( new_n7198_, new_n7161_, new_n6873_ );
and  ( new_n7199_, new_n7163_, new_n7047_ );
or   ( new_n7200_, new_n7199_, new_n7198_ );
and  ( new_n7201_, new_n7084_, new_n3734_ );
and  ( new_n7202_, new_n7201_, new_n7200_ );
or   ( new_n7203_, new_n7087_, new_n2304_ );
and  ( new_n7204_, new_n7203_, new_n7200_ );
and  ( new_n7205_, new_n7163_, new_n7161_ );
or   ( new_n7206_, new_n7205_, new_n7048_ );
and  ( new_n7207_, new_n7206_, new_n7201_ );
or   ( new_n7208_, new_n7207_, new_n7204_ );
and  ( new_n7209_, new_n7157_, new_n6884_ );
and  ( new_n7210_, new_n7159_, new_n7045_ );
or   ( new_n7211_, new_n7210_, new_n7209_ );
and  ( new_n7212_, new_n7084_, new_n2441_ );
and  ( new_n7213_, new_n7212_, new_n7211_ );
or   ( new_n7214_, new_n7087_, new_n2440_ );
and  ( new_n7215_, new_n7214_, new_n7211_ );
and  ( new_n7216_, new_n7159_, new_n7157_ );
or   ( new_n7217_, new_n7216_, new_n7046_ );
and  ( new_n7218_, new_n7217_, new_n7212_ );
or   ( new_n7219_, new_n7218_, new_n7215_ );
and  ( new_n7220_, new_n7153_, new_n6895_ );
and  ( new_n7221_, new_n7155_, new_n7043_ );
or   ( new_n7222_, new_n7221_, new_n7220_ );
and  ( new_n7223_, new_n7084_, new_n6342_ );
and  ( new_n7224_, new_n7223_, new_n7222_ );
or   ( new_n7225_, new_n7087_, new_n2566_ );
and  ( new_n7226_, new_n7225_, new_n7222_ );
and  ( new_n7227_, new_n7155_, new_n7153_ );
or   ( new_n7228_, new_n7227_, new_n7044_ );
and  ( new_n7229_, new_n7228_, new_n7223_ );
or   ( new_n7230_, new_n7229_, new_n7226_ );
and  ( new_n7231_, new_n7149_, new_n6906_ );
and  ( new_n7232_, new_n7151_, new_n7041_ );
or   ( new_n7233_, new_n7232_, new_n7231_ );
and  ( new_n7234_, new_n7084_, new_n3693_ );
and  ( new_n7235_, new_n7234_, new_n7233_ );
or   ( new_n7236_, new_n7087_, new_n2705_ );
and  ( new_n7237_, new_n7236_, new_n7233_ );
and  ( new_n7238_, new_n7151_, new_n7149_ );
or   ( new_n7239_, new_n7238_, new_n7042_ );
and  ( new_n7240_, new_n7239_, new_n7234_ );
or   ( new_n7241_, new_n7240_, new_n7237_ );
and  ( new_n7242_, new_n7145_, new_n6917_ );
and  ( new_n7243_, new_n7147_, new_n7039_ );
or   ( new_n7244_, new_n7243_, new_n7242_ );
and  ( new_n7245_, new_n7084_, new_n4017_ );
and  ( new_n7246_, new_n7245_, new_n7244_ );
or   ( new_n7247_, new_n7087_, new_n2723_ );
and  ( new_n7248_, new_n7247_, new_n7244_ );
and  ( new_n7249_, new_n7147_, new_n7145_ );
or   ( new_n7250_, new_n7249_, new_n7040_ );
and  ( new_n7251_, new_n7250_, new_n7245_ );
or   ( new_n7252_, new_n7251_, new_n7248_ );
and  ( new_n7253_, new_n7141_, new_n6928_ );
and  ( new_n7254_, new_n7143_, new_n7037_ );
or   ( new_n7255_, new_n7254_, new_n7253_ );
and  ( new_n7256_, new_n7084_, new_n4085_ );
and  ( new_n7257_, new_n7256_, new_n7255_ );
or   ( new_n7258_, new_n7087_, new_n2760_ );
and  ( new_n7259_, new_n7258_, new_n7255_ );
and  ( new_n7260_, new_n7143_, new_n7141_ );
or   ( new_n7261_, new_n7260_, new_n7038_ );
and  ( new_n7262_, new_n7261_, new_n7256_ );
or   ( new_n7263_, new_n7262_, new_n7259_ );
and  ( new_n7264_, new_n7137_, new_n6939_ );
and  ( new_n7265_, new_n7139_, new_n7035_ );
or   ( new_n7266_, new_n7265_, new_n7264_ );
and  ( new_n7267_, new_n7084_, new_n2924_ );
and  ( new_n7268_, new_n7267_, new_n7266_ );
or   ( new_n7269_, new_n7087_, new_n2923_ );
and  ( new_n7270_, new_n7269_, new_n7266_ );
and  ( new_n7271_, new_n7139_, new_n7137_ );
or   ( new_n7272_, new_n7271_, new_n7036_ );
and  ( new_n7273_, new_n7272_, new_n7267_ );
or   ( new_n7274_, new_n7273_, new_n7270_ );
and  ( new_n7275_, new_n7133_, new_n6950_ );
and  ( new_n7276_, new_n7135_, new_n7033_ );
or   ( new_n7277_, new_n7276_, new_n7275_ );
and  ( new_n7278_, new_n7084_, new_n4177_ );
and  ( new_n7279_, new_n7278_, new_n7277_ );
or   ( new_n7280_, new_n7087_, new_n3066_ );
and  ( new_n7281_, new_n7280_, new_n7277_ );
and  ( new_n7282_, new_n7135_, new_n7133_ );
or   ( new_n7283_, new_n7282_, new_n7034_ );
and  ( new_n7284_, new_n7283_, new_n7278_ );
or   ( new_n7285_, new_n7284_, new_n7281_ );
and  ( new_n7286_, new_n7129_, new_n6961_ );
and  ( new_n7287_, new_n7131_, new_n7031_ );
or   ( new_n7288_, new_n7287_, new_n7286_ );
and  ( new_n7289_, new_n7084_, new_n3109_ );
and  ( new_n7290_, new_n7289_, new_n7288_ );
or   ( new_n7291_, new_n7087_, new_n3108_ );
and  ( new_n7292_, new_n7291_, new_n7288_ );
and  ( new_n7293_, new_n7131_, new_n7129_ );
or   ( new_n7294_, new_n7293_, new_n7032_ );
and  ( new_n7295_, new_n7294_, new_n7289_ );
or   ( new_n7296_, new_n7295_, new_n7292_ );
and  ( new_n7297_, new_n7125_, new_n6972_ );
and  ( new_n7298_, new_n7127_, new_n7029_ );
or   ( new_n7299_, new_n7298_, new_n7297_ );
and  ( new_n7300_, new_n7084_, new_n4257_ );
and  ( new_n7301_, new_n7300_, new_n7299_ );
or   ( new_n7302_, new_n7087_, new_n3244_ );
and  ( new_n7303_, new_n7302_, new_n7299_ );
and  ( new_n7304_, new_n7127_, new_n7125_ );
or   ( new_n7305_, new_n7304_, new_n7030_ );
and  ( new_n7306_, new_n7305_, new_n7300_ );
or   ( new_n7307_, new_n7306_, new_n7303_ );
and  ( new_n7308_, new_n7121_, new_n6983_ );
and  ( new_n7309_, new_n7123_, new_n7027_ );
or   ( new_n7310_, new_n7309_, new_n7308_ );
and  ( new_n7311_, new_n7084_, new_n4275_ );
and  ( new_n7312_, new_n7311_, new_n7310_ );
or   ( new_n7313_, new_n7087_, new_n3306_ );
and  ( new_n7314_, new_n7313_, new_n7310_ );
and  ( new_n7315_, new_n7123_, new_n7121_ );
or   ( new_n7316_, new_n7315_, new_n7028_ );
and  ( new_n7317_, new_n7316_, new_n7311_ );
or   ( new_n7318_, new_n7317_, new_n7314_ );
and  ( new_n7319_, new_n7117_, new_n6994_ );
and  ( new_n7320_, new_n7119_, new_n7025_ );
or   ( new_n7321_, new_n7320_, new_n7319_ );
and  ( new_n7322_, new_n7084_, new_n3407_ );
and  ( new_n7323_, new_n7322_, new_n7321_ );
or   ( new_n7324_, new_n7087_, new_n3406_ );
and  ( new_n7325_, new_n7324_, new_n7321_ );
and  ( new_n7326_, new_n7119_, new_n7117_ );
or   ( new_n7327_, new_n7326_, new_n7026_ );
and  ( new_n7328_, new_n7327_, new_n7322_ );
or   ( new_n7329_, new_n7328_, new_n7325_ );
and  ( new_n7330_, new_n7113_, new_n7005_ );
and  ( new_n7331_, new_n7115_, new_n7023_ );
or   ( new_n7332_, new_n7331_, new_n7330_ );
and  ( new_n7333_, new_n7084_, new_n4311_ );
and  ( new_n7334_, new_n7333_, new_n7332_ );
and  ( new_n7335_, new_n7109_, new_n7021_ );
and  ( new_n7336_, new_n7111_, new_n7015_ );
or   ( new_n7337_, new_n7336_, new_n7335_ );
and  ( new_n7338_, new_n7084_, new_n3547_ );
and  ( new_n7339_, new_n7338_, new_n7337_ );
or   ( new_n7340_, new_n7087_, new_n3507_ );
and  ( new_n7341_, new_n7340_, new_n7332_ );
and  ( new_n7342_, new_n7115_, new_n7113_ );
or   ( new_n7343_, new_n7342_, new_n7024_ );
and  ( new_n7344_, new_n7343_, new_n7333_ );
or   ( new_n7345_, new_n7344_, new_n7341_ );
and  ( new_n7346_, new_n7345_, new_n7339_ );
or   ( new_n7347_, new_n7346_, new_n7334_ );
and  ( new_n7348_, new_n7347_, new_n7329_ );
or   ( new_n7349_, new_n7348_, new_n7323_ );
and  ( new_n7350_, new_n7349_, new_n7318_ );
or   ( new_n7351_, new_n7350_, new_n7312_ );
and  ( new_n7352_, new_n7351_, new_n7307_ );
or   ( new_n7353_, new_n7352_, new_n7301_ );
and  ( new_n7354_, new_n7353_, new_n7296_ );
or   ( new_n7355_, new_n7354_, new_n7290_ );
and  ( new_n7356_, new_n7355_, new_n7285_ );
or   ( new_n7357_, new_n7356_, new_n7279_ );
and  ( new_n7358_, new_n7357_, new_n7274_ );
or   ( new_n7359_, new_n7358_, new_n7268_ );
and  ( new_n7360_, new_n7359_, new_n7263_ );
or   ( new_n7361_, new_n7360_, new_n7257_ );
and  ( new_n7362_, new_n7361_, new_n7252_ );
or   ( new_n7363_, new_n7362_, new_n7246_ );
and  ( new_n7364_, new_n7363_, new_n7241_ );
or   ( new_n7365_, new_n7364_, new_n7235_ );
and  ( new_n7366_, new_n7365_, new_n7230_ );
or   ( new_n7367_, new_n7366_, new_n7224_ );
and  ( new_n7368_, new_n7367_, new_n7219_ );
or   ( new_n7369_, new_n7368_, new_n7213_ );
and  ( new_n7370_, new_n7369_, new_n7208_ );
or   ( new_n7371_, new_n7370_, new_n7202_ );
and  ( new_n7372_, new_n7371_, new_n7197_ );
or   ( new_n7373_, new_n7372_, new_n7191_ );
and  ( new_n7374_, new_n7373_, new_n7186_ );
or   ( new_n7375_, new_n7374_, new_n7180_ );
and  ( new_n7376_, new_n7375_, new_n7175_ );
or   ( new_n7377_, new_n7376_, new_n7086_ );
not  ( new_n7378_, new_n2104_ );
and  ( new_n7379_, new_n5083_, new_n7378_ );
not  ( new_n7380_, new_n7379_ );
xor  ( new_n7381_, new_n5176_, new_n687_ );
and  ( new_n7382_, new_n7381_, new_n5098_ );
and  ( new_n7383_, new_n847_, new_n176_ );
not  ( new_n7384_, new_n7383_ );
and  ( new_n7385_, new_n5102_, new_n7384_ );
nor  ( new_n7386_, new_n7385_, new_n7382_ );
and  ( new_n7387_, new_n7386_, new_n7380_ );
and  ( new_n7388_, new_n5110_, \a[5]  );
and  ( new_n7389_, new_n5092_, \c[5]  );
nor  ( new_n7390_, new_n7389_, new_n7388_ );
and  ( new_n7391_, new_n5076_, new_n2836_ );
and  ( new_n7392_, new_n5080_, new_n2841_ );
nor  ( new_n7393_, new_n7392_, new_n7391_ );
and  ( new_n7394_, new_n7393_, new_n7390_ );
and  ( new_n7395_, new_n7394_, new_n7387_ );
and  ( new_n7396_, new_n5064_, \c[5]  );
nor  ( new_n7397_, new_n7396_, new_n5116_ );
nor  ( new_n7398_, new_n7397_, new_n847_ );
not  ( new_n7399_, new_n7398_ );
xor  ( new_n7400_, new_n5716_, new_n1495_ );
and  ( new_n7401_, new_n7400_, new_n5052_ );
not  ( new_n7402_, new_n7401_ );
and  ( new_n7403_, new_n5072_, \d[5]  );
and  ( new_n7404_, new_n5056_, new_n2823_ );
nor  ( new_n7405_, new_n7404_, new_n7403_ );
and  ( new_n7406_, new_n7405_, new_n7402_ );
and  ( new_n7407_, new_n7406_, new_n7399_ );
and  ( new_n7408_, new_n7407_, new_n7395_ );
not  ( new_n7409_, new_n7408_ );
and  ( new_n7410_, new_n7409_, new_n2407_ );
and  ( new_n7411_, new_n7410_, new_n7377_ );
and  ( new_n7412_, new_n7408_, new_n5120_ );
or   ( new_n7413_, new_n7412_, new_n2906_ );
and  ( new_n7414_, new_n7413_, new_n7377_ );
or   ( new_n7415_, new_n7173_, new_n7088_ );
or   ( new_n7416_, new_n7184_, new_n7181_ );
or   ( new_n7417_, new_n7195_, new_n7192_ );
or   ( new_n7418_, new_n7206_, new_n7203_ );
or   ( new_n7419_, new_n7217_, new_n7214_ );
or   ( new_n7420_, new_n7228_, new_n7225_ );
or   ( new_n7421_, new_n7239_, new_n7236_ );
or   ( new_n7422_, new_n7250_, new_n7247_ );
or   ( new_n7423_, new_n7261_, new_n7258_ );
or   ( new_n7424_, new_n7272_, new_n7269_ );
or   ( new_n7425_, new_n7283_, new_n7280_ );
or   ( new_n7426_, new_n7294_, new_n7291_ );
or   ( new_n7427_, new_n7305_, new_n7302_ );
or   ( new_n7428_, new_n7316_, new_n7313_ );
or   ( new_n7429_, new_n7327_, new_n7324_ );
or   ( new_n7430_, new_n7343_, new_n7340_ );
and  ( new_n7431_, new_n7111_, new_n7109_ );
or   ( new_n7432_, new_n7431_, new_n7022_ );
or   ( new_n7433_, new_n7087_, new_n3548_ );
or   ( new_n7434_, new_n7433_, new_n7432_ );
and  ( new_n7435_, new_n7343_, new_n7340_ );
or   ( new_n7436_, new_n7435_, new_n7334_ );
or   ( new_n7437_, new_n7436_, new_n7434_ );
and  ( new_n7438_, new_n7437_, new_n7430_ );
and  ( new_n7439_, new_n7327_, new_n7324_ );
or   ( new_n7440_, new_n7439_, new_n7323_ );
or   ( new_n7441_, new_n7440_, new_n7438_ );
and  ( new_n7442_, new_n7441_, new_n7429_ );
and  ( new_n7443_, new_n7316_, new_n7313_ );
or   ( new_n7444_, new_n7443_, new_n7312_ );
or   ( new_n7445_, new_n7444_, new_n7442_ );
and  ( new_n7446_, new_n7445_, new_n7428_ );
and  ( new_n7447_, new_n7305_, new_n7302_ );
or   ( new_n7448_, new_n7447_, new_n7301_ );
or   ( new_n7449_, new_n7448_, new_n7446_ );
and  ( new_n7450_, new_n7449_, new_n7427_ );
and  ( new_n7451_, new_n7294_, new_n7291_ );
or   ( new_n7452_, new_n7451_, new_n7290_ );
or   ( new_n7453_, new_n7452_, new_n7450_ );
and  ( new_n7454_, new_n7453_, new_n7426_ );
and  ( new_n7455_, new_n7283_, new_n7280_ );
or   ( new_n7456_, new_n7455_, new_n7279_ );
or   ( new_n7457_, new_n7456_, new_n7454_ );
and  ( new_n7458_, new_n7457_, new_n7425_ );
and  ( new_n7459_, new_n7272_, new_n7269_ );
or   ( new_n7460_, new_n7459_, new_n7268_ );
or   ( new_n7461_, new_n7460_, new_n7458_ );
and  ( new_n7462_, new_n7461_, new_n7424_ );
and  ( new_n7463_, new_n7261_, new_n7258_ );
or   ( new_n7464_, new_n7463_, new_n7257_ );
or   ( new_n7465_, new_n7464_, new_n7462_ );
and  ( new_n7466_, new_n7465_, new_n7423_ );
and  ( new_n7467_, new_n7250_, new_n7247_ );
or   ( new_n7468_, new_n7467_, new_n7246_ );
or   ( new_n7469_, new_n7468_, new_n7466_ );
and  ( new_n7470_, new_n7469_, new_n7422_ );
and  ( new_n7471_, new_n7239_, new_n7236_ );
or   ( new_n7472_, new_n7471_, new_n7235_ );
or   ( new_n7473_, new_n7472_, new_n7470_ );
and  ( new_n7474_, new_n7473_, new_n7421_ );
and  ( new_n7475_, new_n7228_, new_n7225_ );
or   ( new_n7476_, new_n7475_, new_n7224_ );
or   ( new_n7477_, new_n7476_, new_n7474_ );
and  ( new_n7478_, new_n7477_, new_n7420_ );
and  ( new_n7479_, new_n7217_, new_n7214_ );
or   ( new_n7480_, new_n7479_, new_n7213_ );
or   ( new_n7481_, new_n7480_, new_n7478_ );
and  ( new_n7482_, new_n7481_, new_n7419_ );
and  ( new_n7483_, new_n7206_, new_n7203_ );
or   ( new_n7484_, new_n7483_, new_n7202_ );
or   ( new_n7485_, new_n7484_, new_n7482_ );
and  ( new_n7486_, new_n7485_, new_n7418_ );
and  ( new_n7487_, new_n7195_, new_n7192_ );
or   ( new_n7488_, new_n7487_, new_n7191_ );
or   ( new_n7489_, new_n7488_, new_n7486_ );
and  ( new_n7490_, new_n7489_, new_n7417_ );
and  ( new_n7491_, new_n7184_, new_n7181_ );
or   ( new_n7492_, new_n7491_, new_n7180_ );
or   ( new_n7493_, new_n7492_, new_n7490_ );
and  ( new_n7494_, new_n7493_, new_n7416_ );
and  ( new_n7495_, new_n7173_, new_n7088_ );
or   ( new_n7496_, new_n7495_, new_n7086_ );
or   ( new_n7497_, new_n7496_, new_n7494_ );
and  ( new_n7498_, new_n7497_, new_n7415_ );
and  ( new_n7499_, new_n7498_, new_n7410_ );
or   ( new_n7500_, new_n7499_, new_n7414_ );
and  ( new_n7501_, new_n7494_, new_n7175_ );
and  ( new_n7502_, new_n7496_, new_n7375_ );
or   ( new_n7503_, new_n7502_, new_n7501_ );
and  ( new_n7504_, new_n7409_, new_n3143_ );
and  ( new_n7505_, new_n7504_, new_n7503_ );
or   ( new_n7506_, new_n7412_, new_n2297_ );
and  ( new_n7507_, new_n7506_, new_n7503_ );
and  ( new_n7508_, new_n7496_, new_n7494_ );
or   ( new_n7509_, new_n7508_, new_n7376_ );
and  ( new_n7510_, new_n7509_, new_n7504_ );
or   ( new_n7511_, new_n7510_, new_n7507_ );
and  ( new_n7512_, new_n7490_, new_n7186_ );
and  ( new_n7513_, new_n7492_, new_n7373_ );
or   ( new_n7514_, new_n7513_, new_n7512_ );
and  ( new_n7515_, new_n7409_, new_n2420_ );
and  ( new_n7516_, new_n7515_, new_n7514_ );
or   ( new_n7517_, new_n7412_, new_n2288_ );
and  ( new_n7518_, new_n7517_, new_n7514_ );
and  ( new_n7519_, new_n7492_, new_n7490_ );
or   ( new_n7520_, new_n7519_, new_n7374_ );
and  ( new_n7521_, new_n7520_, new_n7515_ );
or   ( new_n7522_, new_n7521_, new_n7518_ );
and  ( new_n7523_, new_n7486_, new_n7197_ );
and  ( new_n7524_, new_n7488_, new_n7371_ );
or   ( new_n7525_, new_n7524_, new_n7523_ );
and  ( new_n7526_, new_n7409_, new_n3734_ );
and  ( new_n7527_, new_n7526_, new_n7525_ );
or   ( new_n7528_, new_n7412_, new_n2304_ );
and  ( new_n7529_, new_n7528_, new_n7525_ );
and  ( new_n7530_, new_n7488_, new_n7486_ );
or   ( new_n7531_, new_n7530_, new_n7372_ );
and  ( new_n7532_, new_n7531_, new_n7526_ );
or   ( new_n7533_, new_n7532_, new_n7529_ );
and  ( new_n7534_, new_n7482_, new_n7208_ );
and  ( new_n7535_, new_n7484_, new_n7369_ );
or   ( new_n7536_, new_n7535_, new_n7534_ );
and  ( new_n7537_, new_n7409_, new_n2441_ );
and  ( new_n7538_, new_n7537_, new_n7536_ );
or   ( new_n7539_, new_n7412_, new_n2440_ );
and  ( new_n7540_, new_n7539_, new_n7536_ );
and  ( new_n7541_, new_n7484_, new_n7482_ );
or   ( new_n7542_, new_n7541_, new_n7370_ );
and  ( new_n7543_, new_n7542_, new_n7537_ );
or   ( new_n7544_, new_n7543_, new_n7540_ );
and  ( new_n7545_, new_n7478_, new_n7219_ );
and  ( new_n7546_, new_n7480_, new_n7367_ );
or   ( new_n7547_, new_n7546_, new_n7545_ );
and  ( new_n7548_, new_n7409_, new_n6342_ );
and  ( new_n7549_, new_n7548_, new_n7547_ );
or   ( new_n7550_, new_n7412_, new_n2566_ );
and  ( new_n7551_, new_n7550_, new_n7547_ );
and  ( new_n7552_, new_n7480_, new_n7478_ );
or   ( new_n7553_, new_n7552_, new_n7368_ );
and  ( new_n7554_, new_n7553_, new_n7548_ );
or   ( new_n7555_, new_n7554_, new_n7551_ );
and  ( new_n7556_, new_n7474_, new_n7230_ );
and  ( new_n7557_, new_n7476_, new_n7365_ );
or   ( new_n7558_, new_n7557_, new_n7556_ );
and  ( new_n7559_, new_n7409_, new_n3693_ );
and  ( new_n7560_, new_n7559_, new_n7558_ );
or   ( new_n7561_, new_n7412_, new_n2705_ );
and  ( new_n7562_, new_n7561_, new_n7558_ );
and  ( new_n7563_, new_n7476_, new_n7474_ );
or   ( new_n7564_, new_n7563_, new_n7366_ );
and  ( new_n7565_, new_n7564_, new_n7559_ );
or   ( new_n7566_, new_n7565_, new_n7562_ );
and  ( new_n7567_, new_n7470_, new_n7241_ );
and  ( new_n7568_, new_n7472_, new_n7363_ );
or   ( new_n7569_, new_n7568_, new_n7567_ );
and  ( new_n7570_, new_n7409_, new_n4017_ );
and  ( new_n7571_, new_n7570_, new_n7569_ );
or   ( new_n7572_, new_n7412_, new_n2723_ );
and  ( new_n7573_, new_n7572_, new_n7569_ );
and  ( new_n7574_, new_n7472_, new_n7470_ );
or   ( new_n7575_, new_n7574_, new_n7364_ );
and  ( new_n7576_, new_n7575_, new_n7570_ );
or   ( new_n7577_, new_n7576_, new_n7573_ );
and  ( new_n7578_, new_n7466_, new_n7252_ );
and  ( new_n7579_, new_n7468_, new_n7361_ );
or   ( new_n7580_, new_n7579_, new_n7578_ );
and  ( new_n7581_, new_n7409_, new_n4085_ );
and  ( new_n7582_, new_n7581_, new_n7580_ );
or   ( new_n7583_, new_n7412_, new_n2760_ );
and  ( new_n7584_, new_n7583_, new_n7580_ );
and  ( new_n7585_, new_n7468_, new_n7466_ );
or   ( new_n7586_, new_n7585_, new_n7362_ );
and  ( new_n7587_, new_n7586_, new_n7581_ );
or   ( new_n7588_, new_n7587_, new_n7584_ );
and  ( new_n7589_, new_n7462_, new_n7263_ );
and  ( new_n7590_, new_n7464_, new_n7359_ );
or   ( new_n7591_, new_n7590_, new_n7589_ );
and  ( new_n7592_, new_n7409_, new_n2924_ );
and  ( new_n7593_, new_n7592_, new_n7591_ );
or   ( new_n7594_, new_n7412_, new_n2923_ );
and  ( new_n7595_, new_n7594_, new_n7591_ );
and  ( new_n7596_, new_n7464_, new_n7462_ );
or   ( new_n7597_, new_n7596_, new_n7360_ );
and  ( new_n7598_, new_n7597_, new_n7592_ );
or   ( new_n7599_, new_n7598_, new_n7595_ );
and  ( new_n7600_, new_n7458_, new_n7274_ );
and  ( new_n7601_, new_n7460_, new_n7357_ );
or   ( new_n7602_, new_n7601_, new_n7600_ );
and  ( new_n7603_, new_n7409_, new_n4177_ );
and  ( new_n7604_, new_n7603_, new_n7602_ );
or   ( new_n7605_, new_n7412_, new_n3066_ );
and  ( new_n7606_, new_n7605_, new_n7602_ );
and  ( new_n7607_, new_n7460_, new_n7458_ );
or   ( new_n7608_, new_n7607_, new_n7358_ );
and  ( new_n7609_, new_n7608_, new_n7603_ );
or   ( new_n7610_, new_n7609_, new_n7606_ );
and  ( new_n7611_, new_n7454_, new_n7285_ );
and  ( new_n7612_, new_n7456_, new_n7355_ );
or   ( new_n7613_, new_n7612_, new_n7611_ );
and  ( new_n7614_, new_n7409_, new_n3109_ );
and  ( new_n7615_, new_n7614_, new_n7613_ );
or   ( new_n7616_, new_n7412_, new_n3108_ );
and  ( new_n7617_, new_n7616_, new_n7613_ );
and  ( new_n7618_, new_n7456_, new_n7454_ );
or   ( new_n7619_, new_n7618_, new_n7356_ );
and  ( new_n7620_, new_n7619_, new_n7614_ );
or   ( new_n7621_, new_n7620_, new_n7617_ );
and  ( new_n7622_, new_n7450_, new_n7296_ );
and  ( new_n7623_, new_n7452_, new_n7353_ );
or   ( new_n7624_, new_n7623_, new_n7622_ );
and  ( new_n7625_, new_n7409_, new_n4257_ );
and  ( new_n7626_, new_n7625_, new_n7624_ );
or   ( new_n7627_, new_n7412_, new_n3244_ );
and  ( new_n7628_, new_n7627_, new_n7624_ );
and  ( new_n7629_, new_n7452_, new_n7450_ );
or   ( new_n7630_, new_n7629_, new_n7354_ );
and  ( new_n7631_, new_n7630_, new_n7625_ );
or   ( new_n7632_, new_n7631_, new_n7628_ );
and  ( new_n7633_, new_n7446_, new_n7307_ );
and  ( new_n7634_, new_n7448_, new_n7351_ );
or   ( new_n7635_, new_n7634_, new_n7633_ );
and  ( new_n7636_, new_n7409_, new_n4275_ );
and  ( new_n7637_, new_n7636_, new_n7635_ );
or   ( new_n7638_, new_n7412_, new_n3306_ );
and  ( new_n7639_, new_n7638_, new_n7635_ );
and  ( new_n7640_, new_n7448_, new_n7446_ );
or   ( new_n7641_, new_n7640_, new_n7352_ );
and  ( new_n7642_, new_n7641_, new_n7636_ );
or   ( new_n7643_, new_n7642_, new_n7639_ );
and  ( new_n7644_, new_n7442_, new_n7318_ );
and  ( new_n7645_, new_n7444_, new_n7349_ );
or   ( new_n7646_, new_n7645_, new_n7644_ );
and  ( new_n7647_, new_n7409_, new_n3407_ );
and  ( new_n7648_, new_n7647_, new_n7646_ );
or   ( new_n7649_, new_n7412_, new_n3406_ );
and  ( new_n7650_, new_n7649_, new_n7646_ );
and  ( new_n7651_, new_n7444_, new_n7442_ );
or   ( new_n7652_, new_n7651_, new_n7350_ );
and  ( new_n7653_, new_n7652_, new_n7647_ );
or   ( new_n7654_, new_n7653_, new_n7650_ );
and  ( new_n7655_, new_n7438_, new_n7329_ );
and  ( new_n7656_, new_n7440_, new_n7347_ );
or   ( new_n7657_, new_n7656_, new_n7655_ );
and  ( new_n7658_, new_n7409_, new_n4311_ );
and  ( new_n7659_, new_n7658_, new_n7657_ );
and  ( new_n7660_, new_n7434_, new_n7345_ );
and  ( new_n7661_, new_n7436_, new_n7339_ );
or   ( new_n7662_, new_n7661_, new_n7660_ );
and  ( new_n7663_, new_n7409_, new_n3547_ );
and  ( new_n7664_, new_n7663_, new_n7662_ );
or   ( new_n7665_, new_n7412_, new_n3507_ );
and  ( new_n7666_, new_n7665_, new_n7657_ );
and  ( new_n7667_, new_n7440_, new_n7438_ );
or   ( new_n7668_, new_n7667_, new_n7348_ );
and  ( new_n7669_, new_n7668_, new_n7658_ );
or   ( new_n7670_, new_n7669_, new_n7666_ );
and  ( new_n7671_, new_n7670_, new_n7664_ );
or   ( new_n7672_, new_n7671_, new_n7659_ );
and  ( new_n7673_, new_n7672_, new_n7654_ );
or   ( new_n7674_, new_n7673_, new_n7648_ );
and  ( new_n7675_, new_n7674_, new_n7643_ );
or   ( new_n7676_, new_n7675_, new_n7637_ );
and  ( new_n7677_, new_n7676_, new_n7632_ );
or   ( new_n7678_, new_n7677_, new_n7626_ );
and  ( new_n7679_, new_n7678_, new_n7621_ );
or   ( new_n7680_, new_n7679_, new_n7615_ );
and  ( new_n7681_, new_n7680_, new_n7610_ );
or   ( new_n7682_, new_n7681_, new_n7604_ );
and  ( new_n7683_, new_n7682_, new_n7599_ );
or   ( new_n7684_, new_n7683_, new_n7593_ );
and  ( new_n7685_, new_n7684_, new_n7588_ );
or   ( new_n7686_, new_n7685_, new_n7582_ );
and  ( new_n7687_, new_n7686_, new_n7577_ );
or   ( new_n7688_, new_n7687_, new_n7571_ );
and  ( new_n7689_, new_n7688_, new_n7566_ );
or   ( new_n7690_, new_n7689_, new_n7560_ );
and  ( new_n7691_, new_n7690_, new_n7555_ );
or   ( new_n7692_, new_n7691_, new_n7549_ );
and  ( new_n7693_, new_n7692_, new_n7544_ );
or   ( new_n7694_, new_n7693_, new_n7538_ );
and  ( new_n7695_, new_n7694_, new_n7533_ );
or   ( new_n7696_, new_n7695_, new_n7527_ );
and  ( new_n7697_, new_n7696_, new_n7522_ );
or   ( new_n7698_, new_n7697_, new_n7516_ );
and  ( new_n7699_, new_n7698_, new_n7511_ );
or   ( new_n7700_, new_n7699_, new_n7505_ );
and  ( new_n7701_, new_n7700_, new_n7500_ );
or   ( new_n7702_, new_n7701_, new_n7411_ );
not  ( new_n7703_, new_n2108_ );
and  ( new_n7704_, new_n5083_, new_n7703_ );
not  ( new_n7705_, new_n7704_ );
xor  ( new_n7706_, new_n5204_, new_n602_ );
and  ( new_n7707_, new_n7706_, new_n5098_ );
or   ( new_n7708_, \b[6] , \a[6]  );
and  ( new_n7709_, new_n7708_, new_n5102_ );
nor  ( new_n7710_, new_n7709_, new_n7707_ );
and  ( new_n7711_, new_n7710_, new_n7705_ );
and  ( new_n7712_, new_n5110_, \a[6]  );
and  ( new_n7713_, new_n5092_, \c[6]  );
nor  ( new_n7714_, new_n7713_, new_n7712_ );
nor  ( new_n7715_, new_n6500_, new_n2801_ );
nor  ( new_n7716_, new_n6503_, new_n2798_ );
nor  ( new_n7717_, new_n7716_, new_n7715_ );
and  ( new_n7718_, new_n7717_, new_n7714_ );
and  ( new_n7719_, new_n7718_, new_n7711_ );
and  ( new_n7720_, new_n5064_, \c[6]  );
nor  ( new_n7721_, new_n7720_, new_n5116_ );
nor  ( new_n7722_, new_n7721_, new_n1019_ );
not  ( new_n7723_, new_n7722_ );
xor  ( new_n7724_, new_n5743_, new_n1415_ );
and  ( new_n7725_, new_n7724_, new_n5052_ );
not  ( new_n7726_, new_n7725_ );
and  ( new_n7727_, new_n5072_, \d[6]  );
and  ( new_n7728_, new_n5056_, new_n2791_ );
nor  ( new_n7729_, new_n7728_, new_n7727_ );
and  ( new_n7730_, new_n7729_, new_n7726_ );
and  ( new_n7731_, new_n7730_, new_n7723_ );
and  ( new_n7732_, new_n7731_, new_n7719_ );
not  ( new_n7733_, new_n7732_ );
and  ( new_n7734_, new_n7733_, new_n2407_ );
and  ( new_n7735_, new_n7734_, new_n7702_ );
and  ( new_n7736_, new_n7732_, new_n5120_ );
or   ( new_n7737_, new_n7736_, new_n2906_ );
and  ( new_n7738_, new_n7737_, new_n7702_ );
or   ( new_n7739_, new_n7498_, new_n7413_ );
or   ( new_n7740_, new_n7509_, new_n7506_ );
or   ( new_n7741_, new_n7520_, new_n7517_ );
or   ( new_n7742_, new_n7531_, new_n7528_ );
or   ( new_n7743_, new_n7542_, new_n7539_ );
or   ( new_n7744_, new_n7553_, new_n7550_ );
or   ( new_n7745_, new_n7564_, new_n7561_ );
or   ( new_n7746_, new_n7575_, new_n7572_ );
or   ( new_n7747_, new_n7586_, new_n7583_ );
or   ( new_n7748_, new_n7597_, new_n7594_ );
or   ( new_n7749_, new_n7608_, new_n7605_ );
or   ( new_n7750_, new_n7619_, new_n7616_ );
or   ( new_n7751_, new_n7630_, new_n7627_ );
or   ( new_n7752_, new_n7641_, new_n7638_ );
or   ( new_n7753_, new_n7652_, new_n7649_ );
or   ( new_n7754_, new_n7668_, new_n7665_ );
and  ( new_n7755_, new_n7436_, new_n7434_ );
or   ( new_n7756_, new_n7755_, new_n7346_ );
or   ( new_n7757_, new_n7412_, new_n3548_ );
or   ( new_n7758_, new_n7757_, new_n7756_ );
and  ( new_n7759_, new_n7668_, new_n7665_ );
or   ( new_n7760_, new_n7759_, new_n7659_ );
or   ( new_n7761_, new_n7760_, new_n7758_ );
and  ( new_n7762_, new_n7761_, new_n7754_ );
and  ( new_n7763_, new_n7652_, new_n7649_ );
or   ( new_n7764_, new_n7763_, new_n7648_ );
or   ( new_n7765_, new_n7764_, new_n7762_ );
and  ( new_n7766_, new_n7765_, new_n7753_ );
and  ( new_n7767_, new_n7641_, new_n7638_ );
or   ( new_n7768_, new_n7767_, new_n7637_ );
or   ( new_n7769_, new_n7768_, new_n7766_ );
and  ( new_n7770_, new_n7769_, new_n7752_ );
and  ( new_n7771_, new_n7630_, new_n7627_ );
or   ( new_n7772_, new_n7771_, new_n7626_ );
or   ( new_n7773_, new_n7772_, new_n7770_ );
and  ( new_n7774_, new_n7773_, new_n7751_ );
and  ( new_n7775_, new_n7619_, new_n7616_ );
or   ( new_n7776_, new_n7775_, new_n7615_ );
or   ( new_n7777_, new_n7776_, new_n7774_ );
and  ( new_n7778_, new_n7777_, new_n7750_ );
and  ( new_n7779_, new_n7608_, new_n7605_ );
or   ( new_n7780_, new_n7779_, new_n7604_ );
or   ( new_n7781_, new_n7780_, new_n7778_ );
and  ( new_n7782_, new_n7781_, new_n7749_ );
and  ( new_n7783_, new_n7597_, new_n7594_ );
or   ( new_n7784_, new_n7783_, new_n7593_ );
or   ( new_n7785_, new_n7784_, new_n7782_ );
and  ( new_n7786_, new_n7785_, new_n7748_ );
and  ( new_n7787_, new_n7586_, new_n7583_ );
or   ( new_n7788_, new_n7787_, new_n7582_ );
or   ( new_n7789_, new_n7788_, new_n7786_ );
and  ( new_n7790_, new_n7789_, new_n7747_ );
and  ( new_n7791_, new_n7575_, new_n7572_ );
or   ( new_n7792_, new_n7791_, new_n7571_ );
or   ( new_n7793_, new_n7792_, new_n7790_ );
and  ( new_n7794_, new_n7793_, new_n7746_ );
and  ( new_n7795_, new_n7564_, new_n7561_ );
or   ( new_n7796_, new_n7795_, new_n7560_ );
or   ( new_n7797_, new_n7796_, new_n7794_ );
and  ( new_n7798_, new_n7797_, new_n7745_ );
and  ( new_n7799_, new_n7553_, new_n7550_ );
or   ( new_n7800_, new_n7799_, new_n7549_ );
or   ( new_n7801_, new_n7800_, new_n7798_ );
and  ( new_n7802_, new_n7801_, new_n7744_ );
and  ( new_n7803_, new_n7542_, new_n7539_ );
or   ( new_n7804_, new_n7803_, new_n7538_ );
or   ( new_n7805_, new_n7804_, new_n7802_ );
and  ( new_n7806_, new_n7805_, new_n7743_ );
and  ( new_n7807_, new_n7531_, new_n7528_ );
or   ( new_n7808_, new_n7807_, new_n7527_ );
or   ( new_n7809_, new_n7808_, new_n7806_ );
and  ( new_n7810_, new_n7809_, new_n7742_ );
and  ( new_n7811_, new_n7520_, new_n7517_ );
or   ( new_n7812_, new_n7811_, new_n7516_ );
or   ( new_n7813_, new_n7812_, new_n7810_ );
and  ( new_n7814_, new_n7813_, new_n7741_ );
and  ( new_n7815_, new_n7509_, new_n7506_ );
or   ( new_n7816_, new_n7815_, new_n7505_ );
or   ( new_n7817_, new_n7816_, new_n7814_ );
and  ( new_n7818_, new_n7817_, new_n7740_ );
and  ( new_n7819_, new_n7498_, new_n7413_ );
or   ( new_n7820_, new_n7819_, new_n7411_ );
or   ( new_n7821_, new_n7820_, new_n7818_ );
and  ( new_n7822_, new_n7821_, new_n7739_ );
and  ( new_n7823_, new_n7822_, new_n7734_ );
or   ( new_n7824_, new_n7823_, new_n7738_ );
and  ( new_n7825_, new_n7818_, new_n7500_ );
and  ( new_n7826_, new_n7820_, new_n7700_ );
or   ( new_n7827_, new_n7826_, new_n7825_ );
and  ( new_n7828_, new_n7733_, new_n3143_ );
and  ( new_n7829_, new_n7828_, new_n7827_ );
or   ( new_n7830_, new_n7736_, new_n2297_ );
and  ( new_n7831_, new_n7830_, new_n7827_ );
and  ( new_n7832_, new_n7820_, new_n7818_ );
or   ( new_n7833_, new_n7832_, new_n7701_ );
and  ( new_n7834_, new_n7833_, new_n7828_ );
or   ( new_n7835_, new_n7834_, new_n7831_ );
and  ( new_n7836_, new_n7814_, new_n7511_ );
and  ( new_n7837_, new_n7816_, new_n7698_ );
or   ( new_n7838_, new_n7837_, new_n7836_ );
and  ( new_n7839_, new_n7733_, new_n2420_ );
and  ( new_n7840_, new_n7839_, new_n7838_ );
or   ( new_n7841_, new_n7736_, new_n2288_ );
and  ( new_n7842_, new_n7841_, new_n7838_ );
and  ( new_n7843_, new_n7816_, new_n7814_ );
or   ( new_n7844_, new_n7843_, new_n7699_ );
and  ( new_n7845_, new_n7844_, new_n7839_ );
or   ( new_n7846_, new_n7845_, new_n7842_ );
and  ( new_n7847_, new_n7810_, new_n7522_ );
and  ( new_n7848_, new_n7812_, new_n7696_ );
or   ( new_n7849_, new_n7848_, new_n7847_ );
and  ( new_n7850_, new_n7733_, new_n3734_ );
and  ( new_n7851_, new_n7850_, new_n7849_ );
or   ( new_n7852_, new_n7736_, new_n2304_ );
and  ( new_n7853_, new_n7852_, new_n7849_ );
and  ( new_n7854_, new_n7812_, new_n7810_ );
or   ( new_n7855_, new_n7854_, new_n7697_ );
and  ( new_n7856_, new_n7855_, new_n7850_ );
or   ( new_n7857_, new_n7856_, new_n7853_ );
and  ( new_n7858_, new_n7806_, new_n7533_ );
and  ( new_n7859_, new_n7808_, new_n7694_ );
or   ( new_n7860_, new_n7859_, new_n7858_ );
and  ( new_n7861_, new_n7733_, new_n2441_ );
and  ( new_n7862_, new_n7861_, new_n7860_ );
or   ( new_n7863_, new_n7736_, new_n2440_ );
and  ( new_n7864_, new_n7863_, new_n7860_ );
and  ( new_n7865_, new_n7808_, new_n7806_ );
or   ( new_n7866_, new_n7865_, new_n7695_ );
and  ( new_n7867_, new_n7866_, new_n7861_ );
or   ( new_n7868_, new_n7867_, new_n7864_ );
and  ( new_n7869_, new_n7802_, new_n7544_ );
and  ( new_n7870_, new_n7804_, new_n7692_ );
or   ( new_n7871_, new_n7870_, new_n7869_ );
and  ( new_n7872_, new_n7733_, new_n6342_ );
and  ( new_n7873_, new_n7872_, new_n7871_ );
or   ( new_n7874_, new_n7736_, new_n2566_ );
and  ( new_n7875_, new_n7874_, new_n7871_ );
and  ( new_n7876_, new_n7804_, new_n7802_ );
or   ( new_n7877_, new_n7876_, new_n7693_ );
and  ( new_n7878_, new_n7877_, new_n7872_ );
or   ( new_n7879_, new_n7878_, new_n7875_ );
and  ( new_n7880_, new_n7798_, new_n7555_ );
and  ( new_n7881_, new_n7800_, new_n7690_ );
or   ( new_n7882_, new_n7881_, new_n7880_ );
and  ( new_n7883_, new_n7733_, new_n3693_ );
and  ( new_n7884_, new_n7883_, new_n7882_ );
or   ( new_n7885_, new_n7736_, new_n2705_ );
and  ( new_n7886_, new_n7885_, new_n7882_ );
and  ( new_n7887_, new_n7800_, new_n7798_ );
or   ( new_n7888_, new_n7887_, new_n7691_ );
and  ( new_n7889_, new_n7888_, new_n7883_ );
or   ( new_n7890_, new_n7889_, new_n7886_ );
and  ( new_n7891_, new_n7794_, new_n7566_ );
and  ( new_n7892_, new_n7796_, new_n7688_ );
or   ( new_n7893_, new_n7892_, new_n7891_ );
and  ( new_n7894_, new_n7733_, new_n4017_ );
and  ( new_n7895_, new_n7894_, new_n7893_ );
or   ( new_n7896_, new_n7736_, new_n2723_ );
and  ( new_n7897_, new_n7896_, new_n7893_ );
and  ( new_n7898_, new_n7796_, new_n7794_ );
or   ( new_n7899_, new_n7898_, new_n7689_ );
and  ( new_n7900_, new_n7899_, new_n7894_ );
or   ( new_n7901_, new_n7900_, new_n7897_ );
and  ( new_n7902_, new_n7790_, new_n7577_ );
and  ( new_n7903_, new_n7792_, new_n7686_ );
or   ( new_n7904_, new_n7903_, new_n7902_ );
and  ( new_n7905_, new_n7733_, new_n4085_ );
and  ( new_n7906_, new_n7905_, new_n7904_ );
or   ( new_n7907_, new_n7736_, new_n2760_ );
and  ( new_n7908_, new_n7907_, new_n7904_ );
and  ( new_n7909_, new_n7792_, new_n7790_ );
or   ( new_n7910_, new_n7909_, new_n7687_ );
and  ( new_n7911_, new_n7910_, new_n7905_ );
or   ( new_n7912_, new_n7911_, new_n7908_ );
and  ( new_n7913_, new_n7786_, new_n7588_ );
and  ( new_n7914_, new_n7788_, new_n7684_ );
or   ( new_n7915_, new_n7914_, new_n7913_ );
and  ( new_n7916_, new_n7733_, new_n2924_ );
and  ( new_n7917_, new_n7916_, new_n7915_ );
or   ( new_n7918_, new_n7736_, new_n2923_ );
and  ( new_n7919_, new_n7918_, new_n7915_ );
and  ( new_n7920_, new_n7788_, new_n7786_ );
or   ( new_n7921_, new_n7920_, new_n7685_ );
and  ( new_n7922_, new_n7921_, new_n7916_ );
or   ( new_n7923_, new_n7922_, new_n7919_ );
and  ( new_n7924_, new_n7782_, new_n7599_ );
and  ( new_n7925_, new_n7784_, new_n7682_ );
or   ( new_n7926_, new_n7925_, new_n7924_ );
and  ( new_n7927_, new_n7733_, new_n4177_ );
and  ( new_n7928_, new_n7927_, new_n7926_ );
or   ( new_n7929_, new_n7736_, new_n3066_ );
and  ( new_n7930_, new_n7929_, new_n7926_ );
and  ( new_n7931_, new_n7784_, new_n7782_ );
or   ( new_n7932_, new_n7931_, new_n7683_ );
and  ( new_n7933_, new_n7932_, new_n7927_ );
or   ( new_n7934_, new_n7933_, new_n7930_ );
and  ( new_n7935_, new_n7778_, new_n7610_ );
and  ( new_n7936_, new_n7780_, new_n7680_ );
or   ( new_n7937_, new_n7936_, new_n7935_ );
and  ( new_n7938_, new_n7733_, new_n3109_ );
and  ( new_n7939_, new_n7938_, new_n7937_ );
or   ( new_n7940_, new_n7736_, new_n3108_ );
and  ( new_n7941_, new_n7940_, new_n7937_ );
and  ( new_n7942_, new_n7780_, new_n7778_ );
or   ( new_n7943_, new_n7942_, new_n7681_ );
and  ( new_n7944_, new_n7943_, new_n7938_ );
or   ( new_n7945_, new_n7944_, new_n7941_ );
and  ( new_n7946_, new_n7774_, new_n7621_ );
and  ( new_n7947_, new_n7776_, new_n7678_ );
or   ( new_n7948_, new_n7947_, new_n7946_ );
and  ( new_n7949_, new_n7733_, new_n4257_ );
and  ( new_n7950_, new_n7949_, new_n7948_ );
or   ( new_n7951_, new_n7736_, new_n3244_ );
and  ( new_n7952_, new_n7951_, new_n7948_ );
and  ( new_n7953_, new_n7776_, new_n7774_ );
or   ( new_n7954_, new_n7953_, new_n7679_ );
and  ( new_n7955_, new_n7954_, new_n7949_ );
or   ( new_n7956_, new_n7955_, new_n7952_ );
and  ( new_n7957_, new_n7770_, new_n7632_ );
and  ( new_n7958_, new_n7772_, new_n7676_ );
or   ( new_n7959_, new_n7958_, new_n7957_ );
and  ( new_n7960_, new_n7733_, new_n4275_ );
and  ( new_n7961_, new_n7960_, new_n7959_ );
or   ( new_n7962_, new_n7736_, new_n3306_ );
and  ( new_n7963_, new_n7962_, new_n7959_ );
and  ( new_n7964_, new_n7772_, new_n7770_ );
or   ( new_n7965_, new_n7964_, new_n7677_ );
and  ( new_n7966_, new_n7965_, new_n7960_ );
or   ( new_n7967_, new_n7966_, new_n7963_ );
and  ( new_n7968_, new_n7766_, new_n7643_ );
and  ( new_n7969_, new_n7768_, new_n7674_ );
or   ( new_n7970_, new_n7969_, new_n7968_ );
and  ( new_n7971_, new_n7733_, new_n3407_ );
and  ( new_n7972_, new_n7971_, new_n7970_ );
or   ( new_n7973_, new_n7736_, new_n3406_ );
and  ( new_n7974_, new_n7973_, new_n7970_ );
and  ( new_n7975_, new_n7768_, new_n7766_ );
or   ( new_n7976_, new_n7975_, new_n7675_ );
and  ( new_n7977_, new_n7976_, new_n7971_ );
or   ( new_n7978_, new_n7977_, new_n7974_ );
and  ( new_n7979_, new_n7762_, new_n7654_ );
and  ( new_n7980_, new_n7764_, new_n7672_ );
or   ( new_n7981_, new_n7980_, new_n7979_ );
and  ( new_n7982_, new_n7733_, new_n4311_ );
and  ( new_n7983_, new_n7982_, new_n7981_ );
and  ( new_n7984_, new_n7758_, new_n7670_ );
and  ( new_n7985_, new_n7760_, new_n7664_ );
or   ( new_n7986_, new_n7985_, new_n7984_ );
and  ( new_n7987_, new_n7733_, new_n3547_ );
and  ( new_n7988_, new_n7987_, new_n7986_ );
or   ( new_n7989_, new_n7736_, new_n3507_ );
and  ( new_n7990_, new_n7989_, new_n7981_ );
and  ( new_n7991_, new_n7764_, new_n7762_ );
or   ( new_n7992_, new_n7991_, new_n7673_ );
and  ( new_n7993_, new_n7992_, new_n7982_ );
or   ( new_n7994_, new_n7993_, new_n7990_ );
and  ( new_n7995_, new_n7994_, new_n7988_ );
or   ( new_n7996_, new_n7995_, new_n7983_ );
and  ( new_n7997_, new_n7996_, new_n7978_ );
or   ( new_n7998_, new_n7997_, new_n7972_ );
and  ( new_n7999_, new_n7998_, new_n7967_ );
or   ( new_n8000_, new_n7999_, new_n7961_ );
and  ( new_n8001_, new_n8000_, new_n7956_ );
or   ( new_n8002_, new_n8001_, new_n7950_ );
and  ( new_n8003_, new_n8002_, new_n7945_ );
or   ( new_n8004_, new_n8003_, new_n7939_ );
and  ( new_n8005_, new_n8004_, new_n7934_ );
or   ( new_n8006_, new_n8005_, new_n7928_ );
and  ( new_n8007_, new_n8006_, new_n7923_ );
or   ( new_n8008_, new_n8007_, new_n7917_ );
and  ( new_n8009_, new_n8008_, new_n7912_ );
or   ( new_n8010_, new_n8009_, new_n7906_ );
and  ( new_n8011_, new_n8010_, new_n7901_ );
or   ( new_n8012_, new_n8011_, new_n7895_ );
and  ( new_n8013_, new_n8012_, new_n7890_ );
or   ( new_n8014_, new_n8013_, new_n7884_ );
and  ( new_n8015_, new_n8014_, new_n7879_ );
or   ( new_n8016_, new_n8015_, new_n7873_ );
and  ( new_n8017_, new_n8016_, new_n7868_ );
or   ( new_n8018_, new_n8017_, new_n7862_ );
and  ( new_n8019_, new_n8018_, new_n7857_ );
or   ( new_n8020_, new_n8019_, new_n7851_ );
and  ( new_n8021_, new_n8020_, new_n7846_ );
or   ( new_n8022_, new_n8021_, new_n7840_ );
and  ( new_n8023_, new_n8022_, new_n7835_ );
or   ( new_n8024_, new_n8023_, new_n7829_ );
and  ( new_n8025_, new_n8024_, new_n7824_ );
or   ( new_n8026_, new_n8025_, new_n7735_ );
not  ( new_n8027_, new_n2107_ );
and  ( new_n8028_, new_n5083_, new_n8027_ );
not  ( new_n8029_, new_n8028_ );
xor  ( new_n8030_, new_n5238_, new_n472_ );
and  ( new_n8031_, new_n8030_, new_n5098_ );
or   ( new_n8032_, \b[7] , \a[7]  );
and  ( new_n8033_, new_n8032_, new_n5102_ );
nor  ( new_n8034_, new_n8033_, new_n8031_ );
and  ( new_n8035_, new_n8034_, new_n8029_ );
and  ( new_n8036_, new_n5110_, \a[7]  );
and  ( new_n8037_, new_n5092_, \c[7]  );
nor  ( new_n8038_, new_n8037_, new_n8036_ );
and  ( new_n8039_, new_n5076_, new_n2677_ );
and  ( new_n8040_, new_n5080_, new_n2672_ );
nor  ( new_n8041_, new_n8040_, new_n8039_ );
and  ( new_n8042_, new_n8041_, new_n8038_ );
and  ( new_n8043_, new_n8042_, new_n8035_ );
and  ( new_n8044_, new_n5064_, \c[7]  );
nor  ( new_n8045_, new_n8044_, new_n5116_ );
nor  ( new_n8046_, new_n8045_, new_n1023_ );
not  ( new_n8047_, new_n8046_ );
xor  ( new_n8048_, new_n5777_, new_n1282_ );
and  ( new_n8049_, new_n8048_, new_n5052_ );
not  ( new_n8050_, new_n8049_ );
and  ( new_n8051_, new_n5072_, \d[7]  );
and  ( new_n8052_, new_n5056_, new_n2655_ );
nor  ( new_n8053_, new_n8052_, new_n8051_ );
and  ( new_n8054_, new_n8053_, new_n8050_ );
and  ( new_n8055_, new_n8054_, new_n8047_ );
and  ( new_n8056_, new_n8055_, new_n8043_ );
not  ( new_n8057_, new_n8056_ );
and  ( new_n8058_, new_n8057_, new_n2407_ );
and  ( new_n8059_, new_n8058_, new_n8026_ );
and  ( new_n8060_, new_n8056_, new_n5120_ );
or   ( new_n8061_, new_n8060_, new_n2906_ );
and  ( new_n8062_, new_n8061_, new_n8026_ );
or   ( new_n8063_, new_n7822_, new_n7737_ );
or   ( new_n8064_, new_n7833_, new_n7830_ );
or   ( new_n8065_, new_n7844_, new_n7841_ );
or   ( new_n8066_, new_n7855_, new_n7852_ );
or   ( new_n8067_, new_n7866_, new_n7863_ );
or   ( new_n8068_, new_n7877_, new_n7874_ );
or   ( new_n8069_, new_n7888_, new_n7885_ );
or   ( new_n8070_, new_n7899_, new_n7896_ );
or   ( new_n8071_, new_n7910_, new_n7907_ );
or   ( new_n8072_, new_n7921_, new_n7918_ );
or   ( new_n8073_, new_n7932_, new_n7929_ );
or   ( new_n8074_, new_n7943_, new_n7940_ );
or   ( new_n8075_, new_n7954_, new_n7951_ );
or   ( new_n8076_, new_n7965_, new_n7962_ );
or   ( new_n8077_, new_n7976_, new_n7973_ );
or   ( new_n8078_, new_n7992_, new_n7989_ );
and  ( new_n8079_, new_n7760_, new_n7758_ );
or   ( new_n8080_, new_n8079_, new_n7671_ );
or   ( new_n8081_, new_n7736_, new_n3548_ );
or   ( new_n8082_, new_n8081_, new_n8080_ );
and  ( new_n8083_, new_n7992_, new_n7989_ );
or   ( new_n8084_, new_n8083_, new_n7983_ );
or   ( new_n8085_, new_n8084_, new_n8082_ );
and  ( new_n8086_, new_n8085_, new_n8078_ );
and  ( new_n8087_, new_n7976_, new_n7973_ );
or   ( new_n8088_, new_n8087_, new_n7972_ );
or   ( new_n8089_, new_n8088_, new_n8086_ );
and  ( new_n8090_, new_n8089_, new_n8077_ );
and  ( new_n8091_, new_n7965_, new_n7962_ );
or   ( new_n8092_, new_n8091_, new_n7961_ );
or   ( new_n8093_, new_n8092_, new_n8090_ );
and  ( new_n8094_, new_n8093_, new_n8076_ );
and  ( new_n8095_, new_n7954_, new_n7951_ );
or   ( new_n8096_, new_n8095_, new_n7950_ );
or   ( new_n8097_, new_n8096_, new_n8094_ );
and  ( new_n8098_, new_n8097_, new_n8075_ );
and  ( new_n8099_, new_n7943_, new_n7940_ );
or   ( new_n8100_, new_n8099_, new_n7939_ );
or   ( new_n8101_, new_n8100_, new_n8098_ );
and  ( new_n8102_, new_n8101_, new_n8074_ );
and  ( new_n8103_, new_n7932_, new_n7929_ );
or   ( new_n8104_, new_n8103_, new_n7928_ );
or   ( new_n8105_, new_n8104_, new_n8102_ );
and  ( new_n8106_, new_n8105_, new_n8073_ );
and  ( new_n8107_, new_n7921_, new_n7918_ );
or   ( new_n8108_, new_n8107_, new_n7917_ );
or   ( new_n8109_, new_n8108_, new_n8106_ );
and  ( new_n8110_, new_n8109_, new_n8072_ );
and  ( new_n8111_, new_n7910_, new_n7907_ );
or   ( new_n8112_, new_n8111_, new_n7906_ );
or   ( new_n8113_, new_n8112_, new_n8110_ );
and  ( new_n8114_, new_n8113_, new_n8071_ );
and  ( new_n8115_, new_n7899_, new_n7896_ );
or   ( new_n8116_, new_n8115_, new_n7895_ );
or   ( new_n8117_, new_n8116_, new_n8114_ );
and  ( new_n8118_, new_n8117_, new_n8070_ );
and  ( new_n8119_, new_n7888_, new_n7885_ );
or   ( new_n8120_, new_n8119_, new_n7884_ );
or   ( new_n8121_, new_n8120_, new_n8118_ );
and  ( new_n8122_, new_n8121_, new_n8069_ );
and  ( new_n8123_, new_n7877_, new_n7874_ );
or   ( new_n8124_, new_n8123_, new_n7873_ );
or   ( new_n8125_, new_n8124_, new_n8122_ );
and  ( new_n8126_, new_n8125_, new_n8068_ );
and  ( new_n8127_, new_n7866_, new_n7863_ );
or   ( new_n8128_, new_n8127_, new_n7862_ );
or   ( new_n8129_, new_n8128_, new_n8126_ );
and  ( new_n8130_, new_n8129_, new_n8067_ );
and  ( new_n8131_, new_n7855_, new_n7852_ );
or   ( new_n8132_, new_n8131_, new_n7851_ );
or   ( new_n8133_, new_n8132_, new_n8130_ );
and  ( new_n8134_, new_n8133_, new_n8066_ );
and  ( new_n8135_, new_n7844_, new_n7841_ );
or   ( new_n8136_, new_n8135_, new_n7840_ );
or   ( new_n8137_, new_n8136_, new_n8134_ );
and  ( new_n8138_, new_n8137_, new_n8065_ );
and  ( new_n8139_, new_n7833_, new_n7830_ );
or   ( new_n8140_, new_n8139_, new_n7829_ );
or   ( new_n8141_, new_n8140_, new_n8138_ );
and  ( new_n8142_, new_n8141_, new_n8064_ );
and  ( new_n8143_, new_n7822_, new_n7737_ );
or   ( new_n8144_, new_n8143_, new_n7735_ );
or   ( new_n8145_, new_n8144_, new_n8142_ );
and  ( new_n8146_, new_n8145_, new_n8063_ );
and  ( new_n8147_, new_n8146_, new_n8058_ );
or   ( new_n8148_, new_n8147_, new_n8062_ );
and  ( new_n8149_, new_n8142_, new_n7824_ );
and  ( new_n8150_, new_n8144_, new_n8024_ );
or   ( new_n8151_, new_n8150_, new_n8149_ );
and  ( new_n8152_, new_n8057_, new_n3143_ );
and  ( new_n8153_, new_n8152_, new_n8151_ );
or   ( new_n8154_, new_n8060_, new_n2297_ );
and  ( new_n8155_, new_n8154_, new_n8151_ );
and  ( new_n8156_, new_n8144_, new_n8142_ );
or   ( new_n8157_, new_n8156_, new_n8025_ );
and  ( new_n8158_, new_n8157_, new_n8152_ );
or   ( new_n8159_, new_n8158_, new_n8155_ );
and  ( new_n8160_, new_n8138_, new_n7835_ );
and  ( new_n8161_, new_n8140_, new_n8022_ );
or   ( new_n8162_, new_n8161_, new_n8160_ );
and  ( new_n8163_, new_n8057_, new_n2420_ );
and  ( new_n8164_, new_n8163_, new_n8162_ );
or   ( new_n8165_, new_n8060_, new_n2288_ );
and  ( new_n8166_, new_n8165_, new_n8162_ );
and  ( new_n8167_, new_n8140_, new_n8138_ );
or   ( new_n8168_, new_n8167_, new_n8023_ );
and  ( new_n8169_, new_n8168_, new_n8163_ );
or   ( new_n8170_, new_n8169_, new_n8166_ );
and  ( new_n8171_, new_n8134_, new_n7846_ );
and  ( new_n8172_, new_n8136_, new_n8020_ );
or   ( new_n8173_, new_n8172_, new_n8171_ );
and  ( new_n8174_, new_n8057_, new_n3734_ );
and  ( new_n8175_, new_n8174_, new_n8173_ );
or   ( new_n8176_, new_n8060_, new_n2304_ );
and  ( new_n8177_, new_n8176_, new_n8173_ );
and  ( new_n8178_, new_n8136_, new_n8134_ );
or   ( new_n8179_, new_n8178_, new_n8021_ );
and  ( new_n8180_, new_n8179_, new_n8174_ );
or   ( new_n8181_, new_n8180_, new_n8177_ );
and  ( new_n8182_, new_n8130_, new_n7857_ );
and  ( new_n8183_, new_n8132_, new_n8018_ );
or   ( new_n8184_, new_n8183_, new_n8182_ );
and  ( new_n8185_, new_n8057_, new_n2441_ );
and  ( new_n8186_, new_n8185_, new_n8184_ );
or   ( new_n8187_, new_n8060_, new_n2440_ );
and  ( new_n8188_, new_n8187_, new_n8184_ );
and  ( new_n8189_, new_n8132_, new_n8130_ );
or   ( new_n8190_, new_n8189_, new_n8019_ );
and  ( new_n8191_, new_n8190_, new_n8185_ );
or   ( new_n8192_, new_n8191_, new_n8188_ );
and  ( new_n8193_, new_n8126_, new_n7868_ );
and  ( new_n8194_, new_n8128_, new_n8016_ );
or   ( new_n8195_, new_n8194_, new_n8193_ );
and  ( new_n8196_, new_n8057_, new_n6342_ );
and  ( new_n8197_, new_n8196_, new_n8195_ );
or   ( new_n8198_, new_n8060_, new_n2566_ );
and  ( new_n8199_, new_n8198_, new_n8195_ );
and  ( new_n8200_, new_n8128_, new_n8126_ );
or   ( new_n8201_, new_n8200_, new_n8017_ );
and  ( new_n8202_, new_n8201_, new_n8196_ );
or   ( new_n8203_, new_n8202_, new_n8199_ );
and  ( new_n8204_, new_n8122_, new_n7879_ );
and  ( new_n8205_, new_n8124_, new_n8014_ );
or   ( new_n8206_, new_n8205_, new_n8204_ );
and  ( new_n8207_, new_n8057_, new_n3693_ );
and  ( new_n8208_, new_n8207_, new_n8206_ );
or   ( new_n8209_, new_n8060_, new_n2705_ );
and  ( new_n8210_, new_n8209_, new_n8206_ );
and  ( new_n8211_, new_n8124_, new_n8122_ );
or   ( new_n8212_, new_n8211_, new_n8015_ );
and  ( new_n8213_, new_n8212_, new_n8207_ );
or   ( new_n8214_, new_n8213_, new_n8210_ );
and  ( new_n8215_, new_n8118_, new_n7890_ );
and  ( new_n8216_, new_n8120_, new_n8012_ );
or   ( new_n8217_, new_n8216_, new_n8215_ );
and  ( new_n8218_, new_n8057_, new_n4017_ );
and  ( new_n8219_, new_n8218_, new_n8217_ );
or   ( new_n8220_, new_n8060_, new_n2723_ );
and  ( new_n8221_, new_n8220_, new_n8217_ );
and  ( new_n8222_, new_n8120_, new_n8118_ );
or   ( new_n8223_, new_n8222_, new_n8013_ );
and  ( new_n8224_, new_n8223_, new_n8218_ );
or   ( new_n8225_, new_n8224_, new_n8221_ );
and  ( new_n8226_, new_n8114_, new_n7901_ );
and  ( new_n8227_, new_n8116_, new_n8010_ );
or   ( new_n8228_, new_n8227_, new_n8226_ );
and  ( new_n8229_, new_n8057_, new_n4085_ );
and  ( new_n8230_, new_n8229_, new_n8228_ );
or   ( new_n8231_, new_n8060_, new_n2760_ );
and  ( new_n8232_, new_n8231_, new_n8228_ );
and  ( new_n8233_, new_n8116_, new_n8114_ );
or   ( new_n8234_, new_n8233_, new_n8011_ );
and  ( new_n8235_, new_n8234_, new_n8229_ );
or   ( new_n8236_, new_n8235_, new_n8232_ );
and  ( new_n8237_, new_n8110_, new_n7912_ );
and  ( new_n8238_, new_n8112_, new_n8008_ );
or   ( new_n8239_, new_n8238_, new_n8237_ );
and  ( new_n8240_, new_n8057_, new_n2924_ );
and  ( new_n8241_, new_n8240_, new_n8239_ );
or   ( new_n8242_, new_n8060_, new_n2923_ );
and  ( new_n8243_, new_n8242_, new_n8239_ );
and  ( new_n8244_, new_n8112_, new_n8110_ );
or   ( new_n8245_, new_n8244_, new_n8009_ );
and  ( new_n8246_, new_n8245_, new_n8240_ );
or   ( new_n8247_, new_n8246_, new_n8243_ );
and  ( new_n8248_, new_n8106_, new_n7923_ );
and  ( new_n8249_, new_n8108_, new_n8006_ );
or   ( new_n8250_, new_n8249_, new_n8248_ );
and  ( new_n8251_, new_n8057_, new_n4177_ );
and  ( new_n8252_, new_n8251_, new_n8250_ );
or   ( new_n8253_, new_n8060_, new_n3066_ );
and  ( new_n8254_, new_n8253_, new_n8250_ );
and  ( new_n8255_, new_n8108_, new_n8106_ );
or   ( new_n8256_, new_n8255_, new_n8007_ );
and  ( new_n8257_, new_n8256_, new_n8251_ );
or   ( new_n8258_, new_n8257_, new_n8254_ );
and  ( new_n8259_, new_n8102_, new_n7934_ );
and  ( new_n8260_, new_n8104_, new_n8004_ );
or   ( new_n8261_, new_n8260_, new_n8259_ );
and  ( new_n8262_, new_n8057_, new_n3109_ );
and  ( new_n8263_, new_n8262_, new_n8261_ );
or   ( new_n8264_, new_n8060_, new_n3108_ );
and  ( new_n8265_, new_n8264_, new_n8261_ );
and  ( new_n8266_, new_n8104_, new_n8102_ );
or   ( new_n8267_, new_n8266_, new_n8005_ );
and  ( new_n8268_, new_n8267_, new_n8262_ );
or   ( new_n8269_, new_n8268_, new_n8265_ );
and  ( new_n8270_, new_n8098_, new_n7945_ );
and  ( new_n8271_, new_n8100_, new_n8002_ );
or   ( new_n8272_, new_n8271_, new_n8270_ );
and  ( new_n8273_, new_n8057_, new_n4257_ );
and  ( new_n8274_, new_n8273_, new_n8272_ );
or   ( new_n8275_, new_n8060_, new_n3244_ );
and  ( new_n8276_, new_n8275_, new_n8272_ );
and  ( new_n8277_, new_n8100_, new_n8098_ );
or   ( new_n8278_, new_n8277_, new_n8003_ );
and  ( new_n8279_, new_n8278_, new_n8273_ );
or   ( new_n8280_, new_n8279_, new_n8276_ );
and  ( new_n8281_, new_n8094_, new_n7956_ );
and  ( new_n8282_, new_n8096_, new_n8000_ );
or   ( new_n8283_, new_n8282_, new_n8281_ );
and  ( new_n8284_, new_n8057_, new_n4275_ );
and  ( new_n8285_, new_n8284_, new_n8283_ );
or   ( new_n8286_, new_n8060_, new_n3306_ );
and  ( new_n8287_, new_n8286_, new_n8283_ );
and  ( new_n8288_, new_n8096_, new_n8094_ );
or   ( new_n8289_, new_n8288_, new_n8001_ );
and  ( new_n8290_, new_n8289_, new_n8284_ );
or   ( new_n8291_, new_n8290_, new_n8287_ );
and  ( new_n8292_, new_n8090_, new_n7967_ );
and  ( new_n8293_, new_n8092_, new_n7998_ );
or   ( new_n8294_, new_n8293_, new_n8292_ );
and  ( new_n8295_, new_n8057_, new_n3407_ );
and  ( new_n8296_, new_n8295_, new_n8294_ );
or   ( new_n8297_, new_n8060_, new_n3406_ );
and  ( new_n8298_, new_n8297_, new_n8294_ );
and  ( new_n8299_, new_n8092_, new_n8090_ );
or   ( new_n8300_, new_n8299_, new_n7999_ );
and  ( new_n8301_, new_n8300_, new_n8295_ );
or   ( new_n8302_, new_n8301_, new_n8298_ );
and  ( new_n8303_, new_n8086_, new_n7978_ );
and  ( new_n8304_, new_n8088_, new_n7996_ );
or   ( new_n8305_, new_n8304_, new_n8303_ );
and  ( new_n8306_, new_n8057_, new_n4311_ );
and  ( new_n8307_, new_n8306_, new_n8305_ );
and  ( new_n8308_, new_n8082_, new_n7994_ );
and  ( new_n8309_, new_n8084_, new_n7988_ );
or   ( new_n8310_, new_n8309_, new_n8308_ );
and  ( new_n8311_, new_n8057_, new_n3547_ );
and  ( new_n8312_, new_n8311_, new_n8310_ );
or   ( new_n8313_, new_n8060_, new_n3507_ );
and  ( new_n8314_, new_n8313_, new_n8305_ );
and  ( new_n8315_, new_n8088_, new_n8086_ );
or   ( new_n8316_, new_n8315_, new_n7997_ );
and  ( new_n8317_, new_n8316_, new_n8306_ );
or   ( new_n8318_, new_n8317_, new_n8314_ );
and  ( new_n8319_, new_n8318_, new_n8312_ );
or   ( new_n8320_, new_n8319_, new_n8307_ );
and  ( new_n8321_, new_n8320_, new_n8302_ );
or   ( new_n8322_, new_n8321_, new_n8296_ );
and  ( new_n8323_, new_n8322_, new_n8291_ );
or   ( new_n8324_, new_n8323_, new_n8285_ );
and  ( new_n8325_, new_n8324_, new_n8280_ );
or   ( new_n8326_, new_n8325_, new_n8274_ );
and  ( new_n8327_, new_n8326_, new_n8269_ );
or   ( new_n8328_, new_n8327_, new_n8263_ );
and  ( new_n8329_, new_n8328_, new_n8258_ );
or   ( new_n8330_, new_n8329_, new_n8252_ );
and  ( new_n8331_, new_n8330_, new_n8247_ );
or   ( new_n8332_, new_n8331_, new_n8241_ );
and  ( new_n8333_, new_n8332_, new_n8236_ );
or   ( new_n8334_, new_n8333_, new_n8230_ );
and  ( new_n8335_, new_n8334_, new_n8225_ );
or   ( new_n8336_, new_n8335_, new_n8219_ );
and  ( new_n8337_, new_n8336_, new_n8214_ );
or   ( new_n8338_, new_n8337_, new_n8208_ );
and  ( new_n8339_, new_n8338_, new_n8203_ );
or   ( new_n8340_, new_n8339_, new_n8197_ );
and  ( new_n8341_, new_n8340_, new_n8192_ );
or   ( new_n8342_, new_n8341_, new_n8186_ );
and  ( new_n8343_, new_n8342_, new_n8181_ );
or   ( new_n8344_, new_n8343_, new_n8175_ );
and  ( new_n8345_, new_n8344_, new_n8170_ );
or   ( new_n8346_, new_n8345_, new_n8164_ );
and  ( new_n8347_, new_n8346_, new_n8159_ );
or   ( new_n8348_, new_n8347_, new_n8153_ );
and  ( new_n8349_, new_n8348_, new_n8148_ );
or   ( new_n8350_, new_n8349_, new_n8059_ );
xor  ( new_n8351_, new_n5817_, new_n5665_ );
and  ( new_n8352_, new_n8351_, new_n5052_ );
not  ( new_n8353_, new_n8352_ );
and  ( new_n8354_, new_n5116_, \b[8]  );
not  ( new_n8355_, new_n2097_ );
and  ( new_n8356_, new_n5083_, new_n8355_ );
nor  ( new_n8357_, new_n8356_, new_n8354_ );
and  ( new_n8358_, new_n8357_, new_n8353_ );
nor  ( new_n8359_, new_n6500_, new_n2625_ );
nor  ( new_n8360_, new_n6503_, new_n2622_ );
nor  ( new_n8361_, new_n8360_, new_n8359_ );
and  ( new_n8362_, \c[8] , \b[8]  );
and  ( new_n8363_, new_n8362_, new_n5064_ );
and  ( new_n8364_, new_n5110_, \a[8]  );
nor  ( new_n8365_, new_n8364_, new_n8363_ );
and  ( new_n8366_, new_n8365_, new_n8361_ );
and  ( new_n8367_, new_n5056_, new_n2641_ );
not  ( new_n8368_, new_n8367_ );
xor  ( new_n8369_, new_n5278_, new_n5123_ );
and  ( new_n8370_, new_n8369_, new_n5098_ );
or   ( new_n8371_, \b[8] , \a[8]  );
and  ( new_n8372_, new_n8371_, new_n5102_ );
nor  ( new_n8373_, new_n8372_, new_n8370_ );
and  ( new_n8374_, new_n8373_, new_n8368_ );
and  ( new_n8375_, new_n5072_, \d[8]  );
and  ( new_n8376_, new_n5092_, \c[8]  );
nor  ( new_n8377_, new_n8376_, new_n8375_ );
and  ( new_n8378_, new_n8377_, new_n8374_ );
and  ( new_n8379_, new_n8378_, new_n8366_ );
and  ( new_n8380_, new_n8379_, new_n8358_ );
not  ( new_n8381_, new_n8380_ );
and  ( new_n8382_, new_n8381_, new_n2407_ );
and  ( new_n8383_, new_n8382_, new_n8350_ );
and  ( new_n8384_, new_n8380_, new_n5120_ );
or   ( new_n8385_, new_n8384_, new_n2906_ );
and  ( new_n8386_, new_n8385_, new_n8350_ );
or   ( new_n8387_, new_n8146_, new_n8061_ );
or   ( new_n8388_, new_n8157_, new_n8154_ );
or   ( new_n8389_, new_n8168_, new_n8165_ );
or   ( new_n8390_, new_n8179_, new_n8176_ );
or   ( new_n8391_, new_n8190_, new_n8187_ );
or   ( new_n8392_, new_n8201_, new_n8198_ );
or   ( new_n8393_, new_n8212_, new_n8209_ );
or   ( new_n8394_, new_n8223_, new_n8220_ );
or   ( new_n8395_, new_n8234_, new_n8231_ );
or   ( new_n8396_, new_n8245_, new_n8242_ );
or   ( new_n8397_, new_n8256_, new_n8253_ );
or   ( new_n8398_, new_n8267_, new_n8264_ );
or   ( new_n8399_, new_n8278_, new_n8275_ );
or   ( new_n8400_, new_n8289_, new_n8286_ );
or   ( new_n8401_, new_n8300_, new_n8297_ );
or   ( new_n8402_, new_n8316_, new_n8313_ );
and  ( new_n8403_, new_n8084_, new_n8082_ );
or   ( new_n8404_, new_n8403_, new_n7995_ );
or   ( new_n8405_, new_n8060_, new_n3548_ );
or   ( new_n8406_, new_n8405_, new_n8404_ );
and  ( new_n8407_, new_n8316_, new_n8313_ );
or   ( new_n8408_, new_n8407_, new_n8307_ );
or   ( new_n8409_, new_n8408_, new_n8406_ );
and  ( new_n8410_, new_n8409_, new_n8402_ );
and  ( new_n8411_, new_n8300_, new_n8297_ );
or   ( new_n8412_, new_n8411_, new_n8296_ );
or   ( new_n8413_, new_n8412_, new_n8410_ );
and  ( new_n8414_, new_n8413_, new_n8401_ );
and  ( new_n8415_, new_n8289_, new_n8286_ );
or   ( new_n8416_, new_n8415_, new_n8285_ );
or   ( new_n8417_, new_n8416_, new_n8414_ );
and  ( new_n8418_, new_n8417_, new_n8400_ );
and  ( new_n8419_, new_n8278_, new_n8275_ );
or   ( new_n8420_, new_n8419_, new_n8274_ );
or   ( new_n8421_, new_n8420_, new_n8418_ );
and  ( new_n8422_, new_n8421_, new_n8399_ );
and  ( new_n8423_, new_n8267_, new_n8264_ );
or   ( new_n8424_, new_n8423_, new_n8263_ );
or   ( new_n8425_, new_n8424_, new_n8422_ );
and  ( new_n8426_, new_n8425_, new_n8398_ );
and  ( new_n8427_, new_n8256_, new_n8253_ );
or   ( new_n8428_, new_n8427_, new_n8252_ );
or   ( new_n8429_, new_n8428_, new_n8426_ );
and  ( new_n8430_, new_n8429_, new_n8397_ );
and  ( new_n8431_, new_n8245_, new_n8242_ );
or   ( new_n8432_, new_n8431_, new_n8241_ );
or   ( new_n8433_, new_n8432_, new_n8430_ );
and  ( new_n8434_, new_n8433_, new_n8396_ );
and  ( new_n8435_, new_n8234_, new_n8231_ );
or   ( new_n8436_, new_n8435_, new_n8230_ );
or   ( new_n8437_, new_n8436_, new_n8434_ );
and  ( new_n8438_, new_n8437_, new_n8395_ );
and  ( new_n8439_, new_n8223_, new_n8220_ );
or   ( new_n8440_, new_n8439_, new_n8219_ );
or   ( new_n8441_, new_n8440_, new_n8438_ );
and  ( new_n8442_, new_n8441_, new_n8394_ );
and  ( new_n8443_, new_n8212_, new_n8209_ );
or   ( new_n8444_, new_n8443_, new_n8208_ );
or   ( new_n8445_, new_n8444_, new_n8442_ );
and  ( new_n8446_, new_n8445_, new_n8393_ );
and  ( new_n8447_, new_n8201_, new_n8198_ );
or   ( new_n8448_, new_n8447_, new_n8197_ );
or   ( new_n8449_, new_n8448_, new_n8446_ );
and  ( new_n8450_, new_n8449_, new_n8392_ );
and  ( new_n8451_, new_n8190_, new_n8187_ );
or   ( new_n8452_, new_n8451_, new_n8186_ );
or   ( new_n8453_, new_n8452_, new_n8450_ );
and  ( new_n8454_, new_n8453_, new_n8391_ );
and  ( new_n8455_, new_n8179_, new_n8176_ );
or   ( new_n8456_, new_n8455_, new_n8175_ );
or   ( new_n8457_, new_n8456_, new_n8454_ );
and  ( new_n8458_, new_n8457_, new_n8390_ );
and  ( new_n8459_, new_n8168_, new_n8165_ );
or   ( new_n8460_, new_n8459_, new_n8164_ );
or   ( new_n8461_, new_n8460_, new_n8458_ );
and  ( new_n8462_, new_n8461_, new_n8389_ );
and  ( new_n8463_, new_n8157_, new_n8154_ );
or   ( new_n8464_, new_n8463_, new_n8153_ );
or   ( new_n8465_, new_n8464_, new_n8462_ );
and  ( new_n8466_, new_n8465_, new_n8388_ );
and  ( new_n8467_, new_n8146_, new_n8061_ );
or   ( new_n8468_, new_n8467_, new_n8059_ );
or   ( new_n8469_, new_n8468_, new_n8466_ );
and  ( new_n8470_, new_n8469_, new_n8387_ );
and  ( new_n8471_, new_n8470_, new_n8382_ );
or   ( new_n8472_, new_n8471_, new_n8386_ );
and  ( new_n8473_, new_n8466_, new_n8148_ );
and  ( new_n8474_, new_n8468_, new_n8348_ );
or   ( new_n8475_, new_n8474_, new_n8473_ );
and  ( new_n8476_, new_n8381_, new_n3143_ );
and  ( new_n8477_, new_n8476_, new_n8475_ );
or   ( new_n8478_, new_n8384_, new_n2297_ );
and  ( new_n8479_, new_n8478_, new_n8475_ );
and  ( new_n8480_, new_n8468_, new_n8466_ );
or   ( new_n8481_, new_n8480_, new_n8349_ );
and  ( new_n8482_, new_n8481_, new_n8476_ );
or   ( new_n8483_, new_n8482_, new_n8479_ );
and  ( new_n8484_, new_n8462_, new_n8159_ );
and  ( new_n8485_, new_n8464_, new_n8346_ );
or   ( new_n8486_, new_n8485_, new_n8484_ );
and  ( new_n8487_, new_n8381_, new_n2420_ );
and  ( new_n8488_, new_n8487_, new_n8486_ );
or   ( new_n8489_, new_n8384_, new_n2288_ );
and  ( new_n8490_, new_n8489_, new_n8486_ );
and  ( new_n8491_, new_n8464_, new_n8462_ );
or   ( new_n8492_, new_n8491_, new_n8347_ );
and  ( new_n8493_, new_n8492_, new_n8487_ );
or   ( new_n8494_, new_n8493_, new_n8490_ );
and  ( new_n8495_, new_n8458_, new_n8170_ );
and  ( new_n8496_, new_n8460_, new_n8344_ );
or   ( new_n8497_, new_n8496_, new_n8495_ );
and  ( new_n8498_, new_n8381_, new_n3734_ );
and  ( new_n8499_, new_n8498_, new_n8497_ );
or   ( new_n8500_, new_n8384_, new_n2304_ );
and  ( new_n8501_, new_n8500_, new_n8497_ );
and  ( new_n8502_, new_n8460_, new_n8458_ );
or   ( new_n8503_, new_n8502_, new_n8345_ );
and  ( new_n8504_, new_n8503_, new_n8498_ );
or   ( new_n8505_, new_n8504_, new_n8501_ );
and  ( new_n8506_, new_n8454_, new_n8181_ );
and  ( new_n8507_, new_n8456_, new_n8342_ );
or   ( new_n8508_, new_n8507_, new_n8506_ );
and  ( new_n8509_, new_n8381_, new_n2441_ );
and  ( new_n8510_, new_n8509_, new_n8508_ );
or   ( new_n8511_, new_n8384_, new_n2440_ );
and  ( new_n8512_, new_n8511_, new_n8508_ );
and  ( new_n8513_, new_n8456_, new_n8454_ );
or   ( new_n8514_, new_n8513_, new_n8343_ );
and  ( new_n8515_, new_n8514_, new_n8509_ );
or   ( new_n8516_, new_n8515_, new_n8512_ );
and  ( new_n8517_, new_n8450_, new_n8192_ );
and  ( new_n8518_, new_n8452_, new_n8340_ );
or   ( new_n8519_, new_n8518_, new_n8517_ );
and  ( new_n8520_, new_n8381_, new_n6342_ );
and  ( new_n8521_, new_n8520_, new_n8519_ );
or   ( new_n8522_, new_n8384_, new_n2566_ );
and  ( new_n8523_, new_n8522_, new_n8519_ );
and  ( new_n8524_, new_n8452_, new_n8450_ );
or   ( new_n8525_, new_n8524_, new_n8341_ );
and  ( new_n8526_, new_n8525_, new_n8520_ );
or   ( new_n8527_, new_n8526_, new_n8523_ );
and  ( new_n8528_, new_n8446_, new_n8203_ );
and  ( new_n8529_, new_n8448_, new_n8338_ );
or   ( new_n8530_, new_n8529_, new_n8528_ );
and  ( new_n8531_, new_n8381_, new_n3693_ );
and  ( new_n8532_, new_n8531_, new_n8530_ );
or   ( new_n8533_, new_n8384_, new_n2705_ );
and  ( new_n8534_, new_n8533_, new_n8530_ );
and  ( new_n8535_, new_n8448_, new_n8446_ );
or   ( new_n8536_, new_n8535_, new_n8339_ );
and  ( new_n8537_, new_n8536_, new_n8531_ );
or   ( new_n8538_, new_n8537_, new_n8534_ );
and  ( new_n8539_, new_n8442_, new_n8214_ );
and  ( new_n8540_, new_n8444_, new_n8336_ );
or   ( new_n8541_, new_n8540_, new_n8539_ );
and  ( new_n8542_, new_n8381_, new_n4017_ );
and  ( new_n8543_, new_n8542_, new_n8541_ );
or   ( new_n8544_, new_n8384_, new_n2723_ );
and  ( new_n8545_, new_n8544_, new_n8541_ );
and  ( new_n8546_, new_n8444_, new_n8442_ );
or   ( new_n8547_, new_n8546_, new_n8337_ );
and  ( new_n8548_, new_n8547_, new_n8542_ );
or   ( new_n8549_, new_n8548_, new_n8545_ );
and  ( new_n8550_, new_n8438_, new_n8225_ );
and  ( new_n8551_, new_n8440_, new_n8334_ );
or   ( new_n8552_, new_n8551_, new_n8550_ );
and  ( new_n8553_, new_n8381_, new_n4085_ );
and  ( new_n8554_, new_n8553_, new_n8552_ );
or   ( new_n8555_, new_n8384_, new_n2760_ );
and  ( new_n8556_, new_n8555_, new_n8552_ );
and  ( new_n8557_, new_n8440_, new_n8438_ );
or   ( new_n8558_, new_n8557_, new_n8335_ );
and  ( new_n8559_, new_n8558_, new_n8553_ );
or   ( new_n8560_, new_n8559_, new_n8556_ );
and  ( new_n8561_, new_n8434_, new_n8236_ );
and  ( new_n8562_, new_n8436_, new_n8332_ );
or   ( new_n8563_, new_n8562_, new_n8561_ );
and  ( new_n8564_, new_n8381_, new_n2924_ );
and  ( new_n8565_, new_n8564_, new_n8563_ );
or   ( new_n8566_, new_n8384_, new_n2923_ );
and  ( new_n8567_, new_n8566_, new_n8563_ );
and  ( new_n8568_, new_n8436_, new_n8434_ );
or   ( new_n8569_, new_n8568_, new_n8333_ );
and  ( new_n8570_, new_n8569_, new_n8564_ );
or   ( new_n8571_, new_n8570_, new_n8567_ );
and  ( new_n8572_, new_n8430_, new_n8247_ );
and  ( new_n8573_, new_n8432_, new_n8330_ );
or   ( new_n8574_, new_n8573_, new_n8572_ );
and  ( new_n8575_, new_n8381_, new_n4177_ );
and  ( new_n8576_, new_n8575_, new_n8574_ );
or   ( new_n8577_, new_n8384_, new_n3066_ );
and  ( new_n8578_, new_n8577_, new_n8574_ );
and  ( new_n8579_, new_n8432_, new_n8430_ );
or   ( new_n8580_, new_n8579_, new_n8331_ );
and  ( new_n8581_, new_n8580_, new_n8575_ );
or   ( new_n8582_, new_n8581_, new_n8578_ );
and  ( new_n8583_, new_n8426_, new_n8258_ );
and  ( new_n8584_, new_n8428_, new_n8328_ );
or   ( new_n8585_, new_n8584_, new_n8583_ );
and  ( new_n8586_, new_n8381_, new_n3109_ );
and  ( new_n8587_, new_n8586_, new_n8585_ );
or   ( new_n8588_, new_n8384_, new_n3108_ );
and  ( new_n8589_, new_n8588_, new_n8585_ );
and  ( new_n8590_, new_n8428_, new_n8426_ );
or   ( new_n8591_, new_n8590_, new_n8329_ );
and  ( new_n8592_, new_n8591_, new_n8586_ );
or   ( new_n8593_, new_n8592_, new_n8589_ );
and  ( new_n8594_, new_n8422_, new_n8269_ );
and  ( new_n8595_, new_n8424_, new_n8326_ );
or   ( new_n8596_, new_n8595_, new_n8594_ );
and  ( new_n8597_, new_n8381_, new_n4257_ );
and  ( new_n8598_, new_n8597_, new_n8596_ );
or   ( new_n8599_, new_n8384_, new_n3244_ );
and  ( new_n8600_, new_n8599_, new_n8596_ );
and  ( new_n8601_, new_n8424_, new_n8422_ );
or   ( new_n8602_, new_n8601_, new_n8327_ );
and  ( new_n8603_, new_n8602_, new_n8597_ );
or   ( new_n8604_, new_n8603_, new_n8600_ );
and  ( new_n8605_, new_n8418_, new_n8280_ );
and  ( new_n8606_, new_n8420_, new_n8324_ );
or   ( new_n8607_, new_n8606_, new_n8605_ );
and  ( new_n8608_, new_n8381_, new_n4275_ );
and  ( new_n8609_, new_n8608_, new_n8607_ );
or   ( new_n8610_, new_n8384_, new_n3306_ );
and  ( new_n8611_, new_n8610_, new_n8607_ );
and  ( new_n8612_, new_n8420_, new_n8418_ );
or   ( new_n8613_, new_n8612_, new_n8325_ );
and  ( new_n8614_, new_n8613_, new_n8608_ );
or   ( new_n8615_, new_n8614_, new_n8611_ );
and  ( new_n8616_, new_n8414_, new_n8291_ );
and  ( new_n8617_, new_n8416_, new_n8322_ );
or   ( new_n8618_, new_n8617_, new_n8616_ );
and  ( new_n8619_, new_n8381_, new_n3407_ );
and  ( new_n8620_, new_n8619_, new_n8618_ );
or   ( new_n8621_, new_n8384_, new_n3406_ );
and  ( new_n8622_, new_n8621_, new_n8618_ );
and  ( new_n8623_, new_n8416_, new_n8414_ );
or   ( new_n8624_, new_n8623_, new_n8323_ );
and  ( new_n8625_, new_n8624_, new_n8619_ );
or   ( new_n8626_, new_n8625_, new_n8622_ );
and  ( new_n8627_, new_n8410_, new_n8302_ );
and  ( new_n8628_, new_n8412_, new_n8320_ );
or   ( new_n8629_, new_n8628_, new_n8627_ );
and  ( new_n8630_, new_n8381_, new_n4311_ );
and  ( new_n8631_, new_n8630_, new_n8629_ );
and  ( new_n8632_, new_n8406_, new_n8318_ );
and  ( new_n8633_, new_n8408_, new_n8312_ );
or   ( new_n8634_, new_n8633_, new_n8632_ );
and  ( new_n8635_, new_n8381_, new_n3547_ );
and  ( new_n8636_, new_n8635_, new_n8634_ );
or   ( new_n8637_, new_n8384_, new_n3507_ );
and  ( new_n8638_, new_n8637_, new_n8629_ );
and  ( new_n8639_, new_n8412_, new_n8410_ );
or   ( new_n8640_, new_n8639_, new_n8321_ );
and  ( new_n8641_, new_n8640_, new_n8630_ );
or   ( new_n8642_, new_n8641_, new_n8638_ );
and  ( new_n8643_, new_n8642_, new_n8636_ );
or   ( new_n8644_, new_n8643_, new_n8631_ );
and  ( new_n8645_, new_n8644_, new_n8626_ );
or   ( new_n8646_, new_n8645_, new_n8620_ );
and  ( new_n8647_, new_n8646_, new_n8615_ );
or   ( new_n8648_, new_n8647_, new_n8609_ );
and  ( new_n8649_, new_n8648_, new_n8604_ );
or   ( new_n8650_, new_n8649_, new_n8598_ );
and  ( new_n8651_, new_n8650_, new_n8593_ );
or   ( new_n8652_, new_n8651_, new_n8587_ );
and  ( new_n8653_, new_n8652_, new_n8582_ );
or   ( new_n8654_, new_n8653_, new_n8576_ );
and  ( new_n8655_, new_n8654_, new_n8571_ );
or   ( new_n8656_, new_n8655_, new_n8565_ );
and  ( new_n8657_, new_n8656_, new_n8560_ );
or   ( new_n8658_, new_n8657_, new_n8554_ );
and  ( new_n8659_, new_n8658_, new_n8549_ );
or   ( new_n8660_, new_n8659_, new_n8543_ );
and  ( new_n8661_, new_n8660_, new_n8538_ );
or   ( new_n8662_, new_n8661_, new_n8532_ );
and  ( new_n8663_, new_n8662_, new_n8527_ );
or   ( new_n8664_, new_n8663_, new_n8521_ );
and  ( new_n8665_, new_n8664_, new_n8516_ );
or   ( new_n8666_, new_n8665_, new_n8510_ );
and  ( new_n8667_, new_n8666_, new_n8505_ );
or   ( new_n8668_, new_n8667_, new_n8499_ );
and  ( new_n8669_, new_n8668_, new_n8494_ );
or   ( new_n8670_, new_n8669_, new_n8488_ );
and  ( new_n8671_, new_n8670_, new_n8483_ );
or   ( new_n8672_, new_n8671_, new_n8477_ );
and  ( new_n8673_, new_n8672_, new_n8472_ );
or   ( new_n8674_, new_n8673_, new_n8383_ );
and  ( new_n8675_, new_n5083_, new_n2491_ );
not  ( new_n8676_, new_n8675_ );
xor  ( new_n8677_, new_n5324_, new_n329_ );
and  ( new_n8678_, new_n8677_, new_n5098_ );
and  ( new_n8679_, new_n5102_, new_n2529_ );
nor  ( new_n8680_, new_n8679_, new_n8678_ );
and  ( new_n8681_, new_n8680_, new_n8676_ );
and  ( new_n8682_, new_n5110_, \a[9]  );
and  ( new_n8683_, new_n5092_, \c[9]  );
nor  ( new_n8684_, new_n8683_, new_n8682_ );
and  ( new_n8685_, new_n5076_, new_n2509_ );
and  ( new_n8686_, new_n5080_, new_n2523_ );
nor  ( new_n8687_, new_n8686_, new_n8685_ );
and  ( new_n8688_, new_n8687_, new_n8684_ );
and  ( new_n8689_, new_n8688_, new_n8681_ );
and  ( new_n8690_, new_n5064_, \c[9]  );
nor  ( new_n8691_, new_n8690_, new_n5116_ );
nor  ( new_n8692_, new_n8691_, new_n1296_ );
not  ( new_n8693_, new_n8692_ );
xor  ( new_n8694_, new_n5863_, new_n1130_ );
and  ( new_n8695_, new_n8694_, new_n5052_ );
not  ( new_n8696_, new_n8695_ );
and  ( new_n8697_, new_n5072_, \d[9]  );
and  ( new_n8698_, new_n5056_, new_n2519_ );
nor  ( new_n8699_, new_n8698_, new_n8697_ );
and  ( new_n8700_, new_n8699_, new_n8696_ );
and  ( new_n8701_, new_n8700_, new_n8693_ );
and  ( new_n8702_, new_n8701_, new_n8689_ );
not  ( new_n8703_, new_n8702_ );
and  ( new_n8704_, new_n8703_, new_n2407_ );
and  ( new_n8705_, new_n8704_, new_n8674_ );
and  ( new_n8706_, new_n8702_, new_n5120_ );
or   ( new_n8707_, new_n8706_, new_n2906_ );
and  ( new_n8708_, new_n8707_, new_n8674_ );
or   ( new_n8709_, new_n8470_, new_n8385_ );
or   ( new_n8710_, new_n8481_, new_n8478_ );
or   ( new_n8711_, new_n8492_, new_n8489_ );
or   ( new_n8712_, new_n8503_, new_n8500_ );
or   ( new_n8713_, new_n8514_, new_n8511_ );
or   ( new_n8714_, new_n8525_, new_n8522_ );
or   ( new_n8715_, new_n8536_, new_n8533_ );
or   ( new_n8716_, new_n8547_, new_n8544_ );
or   ( new_n8717_, new_n8558_, new_n8555_ );
or   ( new_n8718_, new_n8569_, new_n8566_ );
or   ( new_n8719_, new_n8580_, new_n8577_ );
or   ( new_n8720_, new_n8591_, new_n8588_ );
or   ( new_n8721_, new_n8602_, new_n8599_ );
or   ( new_n8722_, new_n8613_, new_n8610_ );
or   ( new_n8723_, new_n8624_, new_n8621_ );
or   ( new_n8724_, new_n8640_, new_n8637_ );
and  ( new_n8725_, new_n8408_, new_n8406_ );
or   ( new_n8726_, new_n8725_, new_n8319_ );
or   ( new_n8727_, new_n8384_, new_n3548_ );
or   ( new_n8728_, new_n8727_, new_n8726_ );
and  ( new_n8729_, new_n8640_, new_n8637_ );
or   ( new_n8730_, new_n8729_, new_n8631_ );
or   ( new_n8731_, new_n8730_, new_n8728_ );
and  ( new_n8732_, new_n8731_, new_n8724_ );
and  ( new_n8733_, new_n8624_, new_n8621_ );
or   ( new_n8734_, new_n8733_, new_n8620_ );
or   ( new_n8735_, new_n8734_, new_n8732_ );
and  ( new_n8736_, new_n8735_, new_n8723_ );
and  ( new_n8737_, new_n8613_, new_n8610_ );
or   ( new_n8738_, new_n8737_, new_n8609_ );
or   ( new_n8739_, new_n8738_, new_n8736_ );
and  ( new_n8740_, new_n8739_, new_n8722_ );
and  ( new_n8741_, new_n8602_, new_n8599_ );
or   ( new_n8742_, new_n8741_, new_n8598_ );
or   ( new_n8743_, new_n8742_, new_n8740_ );
and  ( new_n8744_, new_n8743_, new_n8721_ );
and  ( new_n8745_, new_n8591_, new_n8588_ );
or   ( new_n8746_, new_n8745_, new_n8587_ );
or   ( new_n8747_, new_n8746_, new_n8744_ );
and  ( new_n8748_, new_n8747_, new_n8720_ );
and  ( new_n8749_, new_n8580_, new_n8577_ );
or   ( new_n8750_, new_n8749_, new_n8576_ );
or   ( new_n8751_, new_n8750_, new_n8748_ );
and  ( new_n8752_, new_n8751_, new_n8719_ );
and  ( new_n8753_, new_n8569_, new_n8566_ );
or   ( new_n8754_, new_n8753_, new_n8565_ );
or   ( new_n8755_, new_n8754_, new_n8752_ );
and  ( new_n8756_, new_n8755_, new_n8718_ );
and  ( new_n8757_, new_n8558_, new_n8555_ );
or   ( new_n8758_, new_n8757_, new_n8554_ );
or   ( new_n8759_, new_n8758_, new_n8756_ );
and  ( new_n8760_, new_n8759_, new_n8717_ );
and  ( new_n8761_, new_n8547_, new_n8544_ );
or   ( new_n8762_, new_n8761_, new_n8543_ );
or   ( new_n8763_, new_n8762_, new_n8760_ );
and  ( new_n8764_, new_n8763_, new_n8716_ );
and  ( new_n8765_, new_n8536_, new_n8533_ );
or   ( new_n8766_, new_n8765_, new_n8532_ );
or   ( new_n8767_, new_n8766_, new_n8764_ );
and  ( new_n8768_, new_n8767_, new_n8715_ );
and  ( new_n8769_, new_n8525_, new_n8522_ );
or   ( new_n8770_, new_n8769_, new_n8521_ );
or   ( new_n8771_, new_n8770_, new_n8768_ );
and  ( new_n8772_, new_n8771_, new_n8714_ );
and  ( new_n8773_, new_n8514_, new_n8511_ );
or   ( new_n8774_, new_n8773_, new_n8510_ );
or   ( new_n8775_, new_n8774_, new_n8772_ );
and  ( new_n8776_, new_n8775_, new_n8713_ );
and  ( new_n8777_, new_n8503_, new_n8500_ );
or   ( new_n8778_, new_n8777_, new_n8499_ );
or   ( new_n8779_, new_n8778_, new_n8776_ );
and  ( new_n8780_, new_n8779_, new_n8712_ );
and  ( new_n8781_, new_n8492_, new_n8489_ );
or   ( new_n8782_, new_n8781_, new_n8488_ );
or   ( new_n8783_, new_n8782_, new_n8780_ );
and  ( new_n8784_, new_n8783_, new_n8711_ );
and  ( new_n8785_, new_n8481_, new_n8478_ );
or   ( new_n8786_, new_n8785_, new_n8477_ );
or   ( new_n8787_, new_n8786_, new_n8784_ );
and  ( new_n8788_, new_n8787_, new_n8710_ );
and  ( new_n8789_, new_n8470_, new_n8385_ );
or   ( new_n8790_, new_n8789_, new_n8383_ );
or   ( new_n8791_, new_n8790_, new_n8788_ );
and  ( new_n8792_, new_n8791_, new_n8709_ );
and  ( new_n8793_, new_n8792_, new_n8704_ );
or   ( new_n8794_, new_n8793_, new_n8708_ );
and  ( new_n8795_, new_n8788_, new_n8472_ );
and  ( new_n8796_, new_n8790_, new_n8672_ );
or   ( new_n8797_, new_n8796_, new_n8795_ );
and  ( new_n8798_, new_n8703_, new_n3143_ );
and  ( new_n8799_, new_n8798_, new_n8797_ );
or   ( new_n8800_, new_n8706_, new_n2297_ );
and  ( new_n8801_, new_n8800_, new_n8797_ );
and  ( new_n8802_, new_n8790_, new_n8788_ );
or   ( new_n8803_, new_n8802_, new_n8673_ );
and  ( new_n8804_, new_n8803_, new_n8798_ );
or   ( new_n8805_, new_n8804_, new_n8801_ );
and  ( new_n8806_, new_n8784_, new_n8483_ );
and  ( new_n8807_, new_n8786_, new_n8670_ );
or   ( new_n8808_, new_n8807_, new_n8806_ );
and  ( new_n8809_, new_n8703_, new_n2420_ );
and  ( new_n8810_, new_n8809_, new_n8808_ );
or   ( new_n8811_, new_n8706_, new_n2288_ );
and  ( new_n8812_, new_n8811_, new_n8808_ );
and  ( new_n8813_, new_n8786_, new_n8784_ );
or   ( new_n8814_, new_n8813_, new_n8671_ );
and  ( new_n8815_, new_n8814_, new_n8809_ );
or   ( new_n8816_, new_n8815_, new_n8812_ );
and  ( new_n8817_, new_n8780_, new_n8494_ );
and  ( new_n8818_, new_n8782_, new_n8668_ );
or   ( new_n8819_, new_n8818_, new_n8817_ );
and  ( new_n8820_, new_n8703_, new_n3734_ );
and  ( new_n8821_, new_n8820_, new_n8819_ );
or   ( new_n8822_, new_n8706_, new_n2304_ );
and  ( new_n8823_, new_n8822_, new_n8819_ );
and  ( new_n8824_, new_n8782_, new_n8780_ );
or   ( new_n8825_, new_n8824_, new_n8669_ );
and  ( new_n8826_, new_n8825_, new_n8820_ );
or   ( new_n8827_, new_n8826_, new_n8823_ );
and  ( new_n8828_, new_n8776_, new_n8505_ );
and  ( new_n8829_, new_n8778_, new_n8666_ );
or   ( new_n8830_, new_n8829_, new_n8828_ );
and  ( new_n8831_, new_n8703_, new_n2441_ );
and  ( new_n8832_, new_n8831_, new_n8830_ );
or   ( new_n8833_, new_n8706_, new_n2440_ );
and  ( new_n8834_, new_n8833_, new_n8830_ );
and  ( new_n8835_, new_n8778_, new_n8776_ );
or   ( new_n8836_, new_n8835_, new_n8667_ );
and  ( new_n8837_, new_n8836_, new_n8831_ );
or   ( new_n8838_, new_n8837_, new_n8834_ );
and  ( new_n8839_, new_n8772_, new_n8516_ );
and  ( new_n8840_, new_n8774_, new_n8664_ );
or   ( new_n8841_, new_n8840_, new_n8839_ );
and  ( new_n8842_, new_n8703_, new_n6342_ );
and  ( new_n8843_, new_n8842_, new_n8841_ );
or   ( new_n8844_, new_n8706_, new_n2566_ );
and  ( new_n8845_, new_n8844_, new_n8841_ );
and  ( new_n8846_, new_n8774_, new_n8772_ );
or   ( new_n8847_, new_n8846_, new_n8665_ );
and  ( new_n8848_, new_n8847_, new_n8842_ );
or   ( new_n8849_, new_n8848_, new_n8845_ );
and  ( new_n8850_, new_n8768_, new_n8527_ );
and  ( new_n8851_, new_n8770_, new_n8662_ );
or   ( new_n8852_, new_n8851_, new_n8850_ );
and  ( new_n8853_, new_n8703_, new_n3693_ );
and  ( new_n8854_, new_n8853_, new_n8852_ );
or   ( new_n8855_, new_n8706_, new_n2705_ );
and  ( new_n8856_, new_n8855_, new_n8852_ );
and  ( new_n8857_, new_n8770_, new_n8768_ );
or   ( new_n8858_, new_n8857_, new_n8663_ );
and  ( new_n8859_, new_n8858_, new_n8853_ );
or   ( new_n8860_, new_n8859_, new_n8856_ );
and  ( new_n8861_, new_n8764_, new_n8538_ );
and  ( new_n8862_, new_n8766_, new_n8660_ );
or   ( new_n8863_, new_n8862_, new_n8861_ );
and  ( new_n8864_, new_n8703_, new_n4017_ );
and  ( new_n8865_, new_n8864_, new_n8863_ );
or   ( new_n8866_, new_n8706_, new_n2723_ );
and  ( new_n8867_, new_n8866_, new_n8863_ );
and  ( new_n8868_, new_n8766_, new_n8764_ );
or   ( new_n8869_, new_n8868_, new_n8661_ );
and  ( new_n8870_, new_n8869_, new_n8864_ );
or   ( new_n8871_, new_n8870_, new_n8867_ );
and  ( new_n8872_, new_n8760_, new_n8549_ );
and  ( new_n8873_, new_n8762_, new_n8658_ );
or   ( new_n8874_, new_n8873_, new_n8872_ );
and  ( new_n8875_, new_n8703_, new_n4085_ );
and  ( new_n8876_, new_n8875_, new_n8874_ );
or   ( new_n8877_, new_n8706_, new_n2760_ );
and  ( new_n8878_, new_n8877_, new_n8874_ );
and  ( new_n8879_, new_n8762_, new_n8760_ );
or   ( new_n8880_, new_n8879_, new_n8659_ );
and  ( new_n8881_, new_n8880_, new_n8875_ );
or   ( new_n8882_, new_n8881_, new_n8878_ );
and  ( new_n8883_, new_n8756_, new_n8560_ );
and  ( new_n8884_, new_n8758_, new_n8656_ );
or   ( new_n8885_, new_n8884_, new_n8883_ );
and  ( new_n8886_, new_n8703_, new_n2924_ );
and  ( new_n8887_, new_n8886_, new_n8885_ );
or   ( new_n8888_, new_n8706_, new_n2923_ );
and  ( new_n8889_, new_n8888_, new_n8885_ );
and  ( new_n8890_, new_n8758_, new_n8756_ );
or   ( new_n8891_, new_n8890_, new_n8657_ );
and  ( new_n8892_, new_n8891_, new_n8886_ );
or   ( new_n8893_, new_n8892_, new_n8889_ );
and  ( new_n8894_, new_n8752_, new_n8571_ );
and  ( new_n8895_, new_n8754_, new_n8654_ );
or   ( new_n8896_, new_n8895_, new_n8894_ );
and  ( new_n8897_, new_n8703_, new_n4177_ );
and  ( new_n8898_, new_n8897_, new_n8896_ );
or   ( new_n8899_, new_n8706_, new_n3066_ );
and  ( new_n8900_, new_n8899_, new_n8896_ );
and  ( new_n8901_, new_n8754_, new_n8752_ );
or   ( new_n8902_, new_n8901_, new_n8655_ );
and  ( new_n8903_, new_n8902_, new_n8897_ );
or   ( new_n8904_, new_n8903_, new_n8900_ );
and  ( new_n8905_, new_n8748_, new_n8582_ );
and  ( new_n8906_, new_n8750_, new_n8652_ );
or   ( new_n8907_, new_n8906_, new_n8905_ );
and  ( new_n8908_, new_n8703_, new_n3109_ );
and  ( new_n8909_, new_n8908_, new_n8907_ );
or   ( new_n8910_, new_n8706_, new_n3108_ );
and  ( new_n8911_, new_n8910_, new_n8907_ );
and  ( new_n8912_, new_n8750_, new_n8748_ );
or   ( new_n8913_, new_n8912_, new_n8653_ );
and  ( new_n8914_, new_n8913_, new_n8908_ );
or   ( new_n8915_, new_n8914_, new_n8911_ );
and  ( new_n8916_, new_n8744_, new_n8593_ );
and  ( new_n8917_, new_n8746_, new_n8650_ );
or   ( new_n8918_, new_n8917_, new_n8916_ );
and  ( new_n8919_, new_n8703_, new_n4257_ );
and  ( new_n8920_, new_n8919_, new_n8918_ );
or   ( new_n8921_, new_n8706_, new_n3244_ );
and  ( new_n8922_, new_n8921_, new_n8918_ );
and  ( new_n8923_, new_n8746_, new_n8744_ );
or   ( new_n8924_, new_n8923_, new_n8651_ );
and  ( new_n8925_, new_n8924_, new_n8919_ );
or   ( new_n8926_, new_n8925_, new_n8922_ );
and  ( new_n8927_, new_n8740_, new_n8604_ );
and  ( new_n8928_, new_n8742_, new_n8648_ );
or   ( new_n8929_, new_n8928_, new_n8927_ );
and  ( new_n8930_, new_n8703_, new_n4275_ );
and  ( new_n8931_, new_n8930_, new_n8929_ );
or   ( new_n8932_, new_n8706_, new_n3306_ );
and  ( new_n8933_, new_n8932_, new_n8929_ );
and  ( new_n8934_, new_n8742_, new_n8740_ );
or   ( new_n8935_, new_n8934_, new_n8649_ );
and  ( new_n8936_, new_n8935_, new_n8930_ );
or   ( new_n8937_, new_n8936_, new_n8933_ );
and  ( new_n8938_, new_n8736_, new_n8615_ );
and  ( new_n8939_, new_n8738_, new_n8646_ );
or   ( new_n8940_, new_n8939_, new_n8938_ );
and  ( new_n8941_, new_n8703_, new_n3407_ );
and  ( new_n8942_, new_n8941_, new_n8940_ );
or   ( new_n8943_, new_n8706_, new_n3406_ );
and  ( new_n8944_, new_n8943_, new_n8940_ );
and  ( new_n8945_, new_n8738_, new_n8736_ );
or   ( new_n8946_, new_n8945_, new_n8647_ );
and  ( new_n8947_, new_n8946_, new_n8941_ );
or   ( new_n8948_, new_n8947_, new_n8944_ );
and  ( new_n8949_, new_n8732_, new_n8626_ );
and  ( new_n8950_, new_n8734_, new_n8644_ );
or   ( new_n8951_, new_n8950_, new_n8949_ );
and  ( new_n8952_, new_n8703_, new_n4311_ );
and  ( new_n8953_, new_n8952_, new_n8951_ );
and  ( new_n8954_, new_n8728_, new_n8642_ );
and  ( new_n8955_, new_n8730_, new_n8636_ );
or   ( new_n8956_, new_n8955_, new_n8954_ );
and  ( new_n8957_, new_n8703_, new_n3547_ );
and  ( new_n8958_, new_n8957_, new_n8956_ );
or   ( new_n8959_, new_n8706_, new_n3507_ );
and  ( new_n8960_, new_n8959_, new_n8951_ );
and  ( new_n8961_, new_n8734_, new_n8732_ );
or   ( new_n8962_, new_n8961_, new_n8645_ );
and  ( new_n8963_, new_n8962_, new_n8952_ );
or   ( new_n8964_, new_n8963_, new_n8960_ );
and  ( new_n8965_, new_n8964_, new_n8958_ );
or   ( new_n8966_, new_n8965_, new_n8953_ );
and  ( new_n8967_, new_n8966_, new_n8948_ );
or   ( new_n8968_, new_n8967_, new_n8942_ );
and  ( new_n8969_, new_n8968_, new_n8937_ );
or   ( new_n8970_, new_n8969_, new_n8931_ );
and  ( new_n8971_, new_n8970_, new_n8926_ );
or   ( new_n8972_, new_n8971_, new_n8920_ );
and  ( new_n8973_, new_n8972_, new_n8915_ );
or   ( new_n8974_, new_n8973_, new_n8909_ );
and  ( new_n8975_, new_n8974_, new_n8904_ );
or   ( new_n8976_, new_n8975_, new_n8898_ );
and  ( new_n8977_, new_n8976_, new_n8893_ );
or   ( new_n8978_, new_n8977_, new_n8887_ );
and  ( new_n8979_, new_n8978_, new_n8882_ );
or   ( new_n8980_, new_n8979_, new_n8876_ );
and  ( new_n8981_, new_n8980_, new_n8871_ );
or   ( new_n8982_, new_n8981_, new_n8865_ );
and  ( new_n8983_, new_n8982_, new_n8860_ );
or   ( new_n8984_, new_n8983_, new_n8854_ );
and  ( new_n8985_, new_n8984_, new_n8849_ );
or   ( new_n8986_, new_n8985_, new_n8843_ );
and  ( new_n8987_, new_n8986_, new_n8838_ );
or   ( new_n8988_, new_n8987_, new_n8832_ );
and  ( new_n8989_, new_n8988_, new_n8827_ );
or   ( new_n8990_, new_n8989_, new_n8821_ );
and  ( new_n8991_, new_n8990_, new_n8816_ );
or   ( new_n8992_, new_n8991_, new_n8810_ );
and  ( new_n8993_, new_n8992_, new_n8805_ );
or   ( new_n8994_, new_n8993_, new_n8799_ );
and  ( new_n8995_, new_n8994_, new_n8794_ );
or   ( new_n8996_, new_n8995_, new_n8705_ );
not  ( new_n8997_, new_n2100_ );
and  ( new_n8998_, new_n5083_, new_n8997_ );
not  ( new_n8999_, new_n8998_ );
xor  ( new_n9000_, new_n5376_, new_n387_ );
and  ( new_n9001_, new_n9000_, new_n5098_ );
not  ( new_n9002_, new_n2467_ );
and  ( new_n9003_, new_n5102_, new_n9002_ );
nor  ( new_n9004_, new_n9003_, new_n9001_ );
and  ( new_n9005_, new_n9004_, new_n8999_ );
and  ( new_n9006_, new_n5110_, \a[10]  );
and  ( new_n9007_, new_n5092_, \c[10]  );
nor  ( new_n9008_, new_n9007_, new_n9006_ );
nor  ( new_n9009_, new_n6500_, new_n2456_ );
nor  ( new_n9010_, new_n6503_, new_n2470_ );
nor  ( new_n9011_, new_n9010_, new_n9009_ );
and  ( new_n9012_, new_n9011_, new_n9008_ );
and  ( new_n9013_, new_n9012_, new_n9005_ );
and  ( new_n9014_, new_n5064_, \c[10]  );
nor  ( new_n9015_, new_n9014_, new_n5116_ );
nor  ( new_n9016_, new_n9015_, new_n1038_ );
not  ( new_n9017_, new_n9016_ );
xor  ( new_n9018_, new_n5915_, new_n1204_ );
and  ( new_n9019_, new_n9018_, new_n5052_ );
not  ( new_n9020_, new_n9019_ );
and  ( new_n9021_, new_n5072_, \d[10]  );
and  ( new_n9022_, new_n5056_, new_n2458_ );
nor  ( new_n9023_, new_n9022_, new_n9021_ );
and  ( new_n9024_, new_n9023_, new_n9020_ );
and  ( new_n9025_, new_n9024_, new_n9017_ );
and  ( new_n9026_, new_n9025_, new_n9013_ );
not  ( new_n9027_, new_n9026_ );
and  ( new_n9028_, new_n9027_, new_n2407_ );
and  ( new_n9029_, new_n9028_, new_n8996_ );
and  ( new_n9030_, new_n9026_, new_n5120_ );
or   ( new_n9031_, new_n9030_, new_n2906_ );
and  ( new_n9032_, new_n9031_, new_n8996_ );
or   ( new_n9033_, new_n8792_, new_n8707_ );
or   ( new_n9034_, new_n8803_, new_n8800_ );
or   ( new_n9035_, new_n8814_, new_n8811_ );
or   ( new_n9036_, new_n8825_, new_n8822_ );
or   ( new_n9037_, new_n8836_, new_n8833_ );
or   ( new_n9038_, new_n8847_, new_n8844_ );
or   ( new_n9039_, new_n8858_, new_n8855_ );
or   ( new_n9040_, new_n8869_, new_n8866_ );
or   ( new_n9041_, new_n8880_, new_n8877_ );
or   ( new_n9042_, new_n8891_, new_n8888_ );
or   ( new_n9043_, new_n8902_, new_n8899_ );
or   ( new_n9044_, new_n8913_, new_n8910_ );
or   ( new_n9045_, new_n8924_, new_n8921_ );
or   ( new_n9046_, new_n8935_, new_n8932_ );
or   ( new_n9047_, new_n8946_, new_n8943_ );
or   ( new_n9048_, new_n8962_, new_n8959_ );
and  ( new_n9049_, new_n8730_, new_n8728_ );
or   ( new_n9050_, new_n9049_, new_n8643_ );
or   ( new_n9051_, new_n8706_, new_n3548_ );
or   ( new_n9052_, new_n9051_, new_n9050_ );
and  ( new_n9053_, new_n8962_, new_n8959_ );
or   ( new_n9054_, new_n9053_, new_n8953_ );
or   ( new_n9055_, new_n9054_, new_n9052_ );
and  ( new_n9056_, new_n9055_, new_n9048_ );
and  ( new_n9057_, new_n8946_, new_n8943_ );
or   ( new_n9058_, new_n9057_, new_n8942_ );
or   ( new_n9059_, new_n9058_, new_n9056_ );
and  ( new_n9060_, new_n9059_, new_n9047_ );
and  ( new_n9061_, new_n8935_, new_n8932_ );
or   ( new_n9062_, new_n9061_, new_n8931_ );
or   ( new_n9063_, new_n9062_, new_n9060_ );
and  ( new_n9064_, new_n9063_, new_n9046_ );
and  ( new_n9065_, new_n8924_, new_n8921_ );
or   ( new_n9066_, new_n9065_, new_n8920_ );
or   ( new_n9067_, new_n9066_, new_n9064_ );
and  ( new_n9068_, new_n9067_, new_n9045_ );
and  ( new_n9069_, new_n8913_, new_n8910_ );
or   ( new_n9070_, new_n9069_, new_n8909_ );
or   ( new_n9071_, new_n9070_, new_n9068_ );
and  ( new_n9072_, new_n9071_, new_n9044_ );
and  ( new_n9073_, new_n8902_, new_n8899_ );
or   ( new_n9074_, new_n9073_, new_n8898_ );
or   ( new_n9075_, new_n9074_, new_n9072_ );
and  ( new_n9076_, new_n9075_, new_n9043_ );
and  ( new_n9077_, new_n8891_, new_n8888_ );
or   ( new_n9078_, new_n9077_, new_n8887_ );
or   ( new_n9079_, new_n9078_, new_n9076_ );
and  ( new_n9080_, new_n9079_, new_n9042_ );
and  ( new_n9081_, new_n8880_, new_n8877_ );
or   ( new_n9082_, new_n9081_, new_n8876_ );
or   ( new_n9083_, new_n9082_, new_n9080_ );
and  ( new_n9084_, new_n9083_, new_n9041_ );
and  ( new_n9085_, new_n8869_, new_n8866_ );
or   ( new_n9086_, new_n9085_, new_n8865_ );
or   ( new_n9087_, new_n9086_, new_n9084_ );
and  ( new_n9088_, new_n9087_, new_n9040_ );
and  ( new_n9089_, new_n8858_, new_n8855_ );
or   ( new_n9090_, new_n9089_, new_n8854_ );
or   ( new_n9091_, new_n9090_, new_n9088_ );
and  ( new_n9092_, new_n9091_, new_n9039_ );
and  ( new_n9093_, new_n8847_, new_n8844_ );
or   ( new_n9094_, new_n9093_, new_n8843_ );
or   ( new_n9095_, new_n9094_, new_n9092_ );
and  ( new_n9096_, new_n9095_, new_n9038_ );
and  ( new_n9097_, new_n8836_, new_n8833_ );
or   ( new_n9098_, new_n9097_, new_n8832_ );
or   ( new_n9099_, new_n9098_, new_n9096_ );
and  ( new_n9100_, new_n9099_, new_n9037_ );
and  ( new_n9101_, new_n8825_, new_n8822_ );
or   ( new_n9102_, new_n9101_, new_n8821_ );
or   ( new_n9103_, new_n9102_, new_n9100_ );
and  ( new_n9104_, new_n9103_, new_n9036_ );
and  ( new_n9105_, new_n8814_, new_n8811_ );
or   ( new_n9106_, new_n9105_, new_n8810_ );
or   ( new_n9107_, new_n9106_, new_n9104_ );
and  ( new_n9108_, new_n9107_, new_n9035_ );
and  ( new_n9109_, new_n8803_, new_n8800_ );
or   ( new_n9110_, new_n9109_, new_n8799_ );
or   ( new_n9111_, new_n9110_, new_n9108_ );
and  ( new_n9112_, new_n9111_, new_n9034_ );
and  ( new_n9113_, new_n8792_, new_n8707_ );
or   ( new_n9114_, new_n9113_, new_n8705_ );
or   ( new_n9115_, new_n9114_, new_n9112_ );
and  ( new_n9116_, new_n9115_, new_n9033_ );
and  ( new_n9117_, new_n9116_, new_n9028_ );
or   ( new_n9118_, new_n9117_, new_n9032_ );
and  ( new_n9119_, new_n9112_, new_n8794_ );
and  ( new_n9120_, new_n9114_, new_n8994_ );
or   ( new_n9121_, new_n9120_, new_n9119_ );
and  ( new_n9122_, new_n9027_, new_n3143_ );
and  ( new_n9123_, new_n9122_, new_n9121_ );
or   ( new_n9124_, new_n9030_, new_n2297_ );
and  ( new_n9125_, new_n9124_, new_n9121_ );
and  ( new_n9126_, new_n9114_, new_n9112_ );
or   ( new_n9127_, new_n9126_, new_n8995_ );
and  ( new_n9128_, new_n9127_, new_n9122_ );
or   ( new_n9129_, new_n9128_, new_n9125_ );
and  ( new_n9130_, new_n9108_, new_n8805_ );
and  ( new_n9131_, new_n9110_, new_n8992_ );
or   ( new_n9132_, new_n9131_, new_n9130_ );
and  ( new_n9133_, new_n9027_, new_n2420_ );
and  ( new_n9134_, new_n9133_, new_n9132_ );
or   ( new_n9135_, new_n9030_, new_n2288_ );
and  ( new_n9136_, new_n9135_, new_n9132_ );
and  ( new_n9137_, new_n9110_, new_n9108_ );
or   ( new_n9138_, new_n9137_, new_n8993_ );
and  ( new_n9139_, new_n9138_, new_n9133_ );
or   ( new_n9140_, new_n9139_, new_n9136_ );
and  ( new_n9141_, new_n9104_, new_n8816_ );
and  ( new_n9142_, new_n9106_, new_n8990_ );
or   ( new_n9143_, new_n9142_, new_n9141_ );
and  ( new_n9144_, new_n9027_, new_n3734_ );
and  ( new_n9145_, new_n9144_, new_n9143_ );
or   ( new_n9146_, new_n9030_, new_n2304_ );
and  ( new_n9147_, new_n9146_, new_n9143_ );
and  ( new_n9148_, new_n9106_, new_n9104_ );
or   ( new_n9149_, new_n9148_, new_n8991_ );
and  ( new_n9150_, new_n9149_, new_n9144_ );
or   ( new_n9151_, new_n9150_, new_n9147_ );
and  ( new_n9152_, new_n9100_, new_n8827_ );
and  ( new_n9153_, new_n9102_, new_n8988_ );
or   ( new_n9154_, new_n9153_, new_n9152_ );
and  ( new_n9155_, new_n9027_, new_n2441_ );
and  ( new_n9156_, new_n9155_, new_n9154_ );
or   ( new_n9157_, new_n9030_, new_n2440_ );
and  ( new_n9158_, new_n9157_, new_n9154_ );
and  ( new_n9159_, new_n9102_, new_n9100_ );
or   ( new_n9160_, new_n9159_, new_n8989_ );
and  ( new_n9161_, new_n9160_, new_n9155_ );
or   ( new_n9162_, new_n9161_, new_n9158_ );
and  ( new_n9163_, new_n9096_, new_n8838_ );
and  ( new_n9164_, new_n9098_, new_n8986_ );
or   ( new_n9165_, new_n9164_, new_n9163_ );
and  ( new_n9166_, new_n9027_, new_n6342_ );
and  ( new_n9167_, new_n9166_, new_n9165_ );
or   ( new_n9168_, new_n9030_, new_n2566_ );
and  ( new_n9169_, new_n9168_, new_n9165_ );
and  ( new_n9170_, new_n9098_, new_n9096_ );
or   ( new_n9171_, new_n9170_, new_n8987_ );
and  ( new_n9172_, new_n9171_, new_n9166_ );
or   ( new_n9173_, new_n9172_, new_n9169_ );
and  ( new_n9174_, new_n9092_, new_n8849_ );
and  ( new_n9175_, new_n9094_, new_n8984_ );
or   ( new_n9176_, new_n9175_, new_n9174_ );
and  ( new_n9177_, new_n9027_, new_n3693_ );
and  ( new_n9178_, new_n9177_, new_n9176_ );
or   ( new_n9179_, new_n9030_, new_n2705_ );
and  ( new_n9180_, new_n9179_, new_n9176_ );
and  ( new_n9181_, new_n9094_, new_n9092_ );
or   ( new_n9182_, new_n9181_, new_n8985_ );
and  ( new_n9183_, new_n9182_, new_n9177_ );
or   ( new_n9184_, new_n9183_, new_n9180_ );
and  ( new_n9185_, new_n9088_, new_n8860_ );
and  ( new_n9186_, new_n9090_, new_n8982_ );
or   ( new_n9187_, new_n9186_, new_n9185_ );
and  ( new_n9188_, new_n9027_, new_n4017_ );
and  ( new_n9189_, new_n9188_, new_n9187_ );
or   ( new_n9190_, new_n9030_, new_n2723_ );
and  ( new_n9191_, new_n9190_, new_n9187_ );
and  ( new_n9192_, new_n9090_, new_n9088_ );
or   ( new_n9193_, new_n9192_, new_n8983_ );
and  ( new_n9194_, new_n9193_, new_n9188_ );
or   ( new_n9195_, new_n9194_, new_n9191_ );
and  ( new_n9196_, new_n9084_, new_n8871_ );
and  ( new_n9197_, new_n9086_, new_n8980_ );
or   ( new_n9198_, new_n9197_, new_n9196_ );
and  ( new_n9199_, new_n9027_, new_n4085_ );
and  ( new_n9200_, new_n9199_, new_n9198_ );
or   ( new_n9201_, new_n9030_, new_n2760_ );
and  ( new_n9202_, new_n9201_, new_n9198_ );
and  ( new_n9203_, new_n9086_, new_n9084_ );
or   ( new_n9204_, new_n9203_, new_n8981_ );
and  ( new_n9205_, new_n9204_, new_n9199_ );
or   ( new_n9206_, new_n9205_, new_n9202_ );
and  ( new_n9207_, new_n9080_, new_n8882_ );
and  ( new_n9208_, new_n9082_, new_n8978_ );
or   ( new_n9209_, new_n9208_, new_n9207_ );
and  ( new_n9210_, new_n9027_, new_n2924_ );
and  ( new_n9211_, new_n9210_, new_n9209_ );
or   ( new_n9212_, new_n9030_, new_n2923_ );
and  ( new_n9213_, new_n9212_, new_n9209_ );
and  ( new_n9214_, new_n9082_, new_n9080_ );
or   ( new_n9215_, new_n9214_, new_n8979_ );
and  ( new_n9216_, new_n9215_, new_n9210_ );
or   ( new_n9217_, new_n9216_, new_n9213_ );
and  ( new_n9218_, new_n9076_, new_n8893_ );
and  ( new_n9219_, new_n9078_, new_n8976_ );
or   ( new_n9220_, new_n9219_, new_n9218_ );
and  ( new_n9221_, new_n9027_, new_n4177_ );
and  ( new_n9222_, new_n9221_, new_n9220_ );
or   ( new_n9223_, new_n9030_, new_n3066_ );
and  ( new_n9224_, new_n9223_, new_n9220_ );
and  ( new_n9225_, new_n9078_, new_n9076_ );
or   ( new_n9226_, new_n9225_, new_n8977_ );
and  ( new_n9227_, new_n9226_, new_n9221_ );
or   ( new_n9228_, new_n9227_, new_n9224_ );
and  ( new_n9229_, new_n9072_, new_n8904_ );
and  ( new_n9230_, new_n9074_, new_n8974_ );
or   ( new_n9231_, new_n9230_, new_n9229_ );
and  ( new_n9232_, new_n9027_, new_n3109_ );
and  ( new_n9233_, new_n9232_, new_n9231_ );
or   ( new_n9234_, new_n9030_, new_n3108_ );
and  ( new_n9235_, new_n9234_, new_n9231_ );
and  ( new_n9236_, new_n9074_, new_n9072_ );
or   ( new_n9237_, new_n9236_, new_n8975_ );
and  ( new_n9238_, new_n9237_, new_n9232_ );
or   ( new_n9239_, new_n9238_, new_n9235_ );
and  ( new_n9240_, new_n9068_, new_n8915_ );
and  ( new_n9241_, new_n9070_, new_n8972_ );
or   ( new_n9242_, new_n9241_, new_n9240_ );
and  ( new_n9243_, new_n9027_, new_n4257_ );
and  ( new_n9244_, new_n9243_, new_n9242_ );
or   ( new_n9245_, new_n9030_, new_n3244_ );
and  ( new_n9246_, new_n9245_, new_n9242_ );
and  ( new_n9247_, new_n9070_, new_n9068_ );
or   ( new_n9248_, new_n9247_, new_n8973_ );
and  ( new_n9249_, new_n9248_, new_n9243_ );
or   ( new_n9250_, new_n9249_, new_n9246_ );
and  ( new_n9251_, new_n9064_, new_n8926_ );
and  ( new_n9252_, new_n9066_, new_n8970_ );
or   ( new_n9253_, new_n9252_, new_n9251_ );
and  ( new_n9254_, new_n9027_, new_n4275_ );
and  ( new_n9255_, new_n9254_, new_n9253_ );
or   ( new_n9256_, new_n9030_, new_n3306_ );
and  ( new_n9257_, new_n9256_, new_n9253_ );
and  ( new_n9258_, new_n9066_, new_n9064_ );
or   ( new_n9259_, new_n9258_, new_n8971_ );
and  ( new_n9260_, new_n9259_, new_n9254_ );
or   ( new_n9261_, new_n9260_, new_n9257_ );
and  ( new_n9262_, new_n9060_, new_n8937_ );
and  ( new_n9263_, new_n9062_, new_n8968_ );
or   ( new_n9264_, new_n9263_, new_n9262_ );
and  ( new_n9265_, new_n9027_, new_n3407_ );
and  ( new_n9266_, new_n9265_, new_n9264_ );
or   ( new_n9267_, new_n9030_, new_n3406_ );
and  ( new_n9268_, new_n9267_, new_n9264_ );
and  ( new_n9269_, new_n9062_, new_n9060_ );
or   ( new_n9270_, new_n9269_, new_n8969_ );
and  ( new_n9271_, new_n9270_, new_n9265_ );
or   ( new_n9272_, new_n9271_, new_n9268_ );
and  ( new_n9273_, new_n9056_, new_n8948_ );
and  ( new_n9274_, new_n9058_, new_n8966_ );
or   ( new_n9275_, new_n9274_, new_n9273_ );
and  ( new_n9276_, new_n9027_, new_n4311_ );
and  ( new_n9277_, new_n9276_, new_n9275_ );
and  ( new_n9278_, new_n9052_, new_n8964_ );
and  ( new_n9279_, new_n9054_, new_n8958_ );
or   ( new_n9280_, new_n9279_, new_n9278_ );
and  ( new_n9281_, new_n9027_, new_n3547_ );
and  ( new_n9282_, new_n9281_, new_n9280_ );
or   ( new_n9283_, new_n9030_, new_n3507_ );
and  ( new_n9284_, new_n9283_, new_n9275_ );
and  ( new_n9285_, new_n9058_, new_n9056_ );
or   ( new_n9286_, new_n9285_, new_n8967_ );
and  ( new_n9287_, new_n9286_, new_n9276_ );
or   ( new_n9288_, new_n9287_, new_n9284_ );
and  ( new_n9289_, new_n9288_, new_n9282_ );
or   ( new_n9290_, new_n9289_, new_n9277_ );
and  ( new_n9291_, new_n9290_, new_n9272_ );
or   ( new_n9292_, new_n9291_, new_n9266_ );
and  ( new_n9293_, new_n9292_, new_n9261_ );
or   ( new_n9294_, new_n9293_, new_n9255_ );
and  ( new_n9295_, new_n9294_, new_n9250_ );
or   ( new_n9296_, new_n9295_, new_n9244_ );
and  ( new_n9297_, new_n9296_, new_n9239_ );
or   ( new_n9298_, new_n9297_, new_n9233_ );
and  ( new_n9299_, new_n9298_, new_n9228_ );
or   ( new_n9300_, new_n9299_, new_n9222_ );
and  ( new_n9301_, new_n9300_, new_n9217_ );
or   ( new_n9302_, new_n9301_, new_n9211_ );
and  ( new_n9303_, new_n9302_, new_n9206_ );
or   ( new_n9304_, new_n9303_, new_n9200_ );
and  ( new_n9305_, new_n9304_, new_n9195_ );
or   ( new_n9306_, new_n9305_, new_n9189_ );
and  ( new_n9307_, new_n9306_, new_n9184_ );
or   ( new_n9308_, new_n9307_, new_n9178_ );
and  ( new_n9309_, new_n9308_, new_n9173_ );
or   ( new_n9310_, new_n9309_, new_n9167_ );
and  ( new_n9311_, new_n9310_, new_n9162_ );
or   ( new_n9312_, new_n9311_, new_n9156_ );
and  ( new_n9313_, new_n9312_, new_n9151_ );
or   ( new_n9314_, new_n9313_, new_n9145_ );
and  ( new_n9315_, new_n9314_, new_n9140_ );
or   ( new_n9316_, new_n9315_, new_n9134_ );
and  ( new_n9317_, new_n9316_, new_n9129_ );
or   ( new_n9318_, new_n9317_, new_n9123_ );
and  ( new_n9319_, new_n9318_, new_n9118_ );
or   ( new_n9320_, new_n9319_, new_n9029_ );
and  ( new_n9321_, new_n5083_, new_n2343_ );
not  ( new_n9322_, new_n9321_ );
xor  ( new_n9323_, new_n5434_, new_n389_ );
and  ( new_n9324_, new_n9323_, new_n5098_ );
and  ( new_n9325_, new_n5102_, new_n2355_ );
nor  ( new_n9326_, new_n9325_, new_n9324_ );
and  ( new_n9327_, new_n9326_, new_n9322_ );
and  ( new_n9328_, new_n5110_, \a[11]  );
and  ( new_n9329_, new_n5092_, \c[11]  );
nor  ( new_n9330_, new_n9329_, new_n9328_ );
and  ( new_n9331_, new_n5076_, new_n2350_ );
and  ( new_n9332_, new_n5080_, new_n2374_ );
nor  ( new_n9333_, new_n9332_, new_n9331_ );
and  ( new_n9334_, new_n9333_, new_n9330_ );
and  ( new_n9335_, new_n9334_, new_n9327_ );
and  ( new_n9336_, new_n5064_, \c[11]  );
nor  ( new_n9337_, new_n9336_, new_n5116_ );
nor  ( new_n9338_, new_n9337_, new_n1154_ );
not  ( new_n9339_, new_n9338_ );
xor  ( new_n9340_, new_n5973_, new_n1206_ );
and  ( new_n9341_, new_n9340_, new_n5052_ );
not  ( new_n9342_, new_n9341_ );
and  ( new_n9343_, new_n5072_, \d[11]  );
and  ( new_n9344_, new_n5056_, new_n2358_ );
nor  ( new_n9345_, new_n9344_, new_n9343_ );
and  ( new_n9346_, new_n9345_, new_n9342_ );
and  ( new_n9347_, new_n9346_, new_n9339_ );
and  ( new_n9348_, new_n9347_, new_n9335_ );
not  ( new_n9349_, new_n9348_ );
and  ( new_n9350_, new_n9349_, new_n2407_ );
and  ( new_n9351_, new_n9350_, new_n9320_ );
and  ( new_n9352_, new_n9348_, new_n5120_ );
or   ( new_n9353_, new_n9352_, new_n2906_ );
and  ( new_n9354_, new_n9353_, new_n9320_ );
or   ( new_n9355_, new_n9116_, new_n9031_ );
or   ( new_n9356_, new_n9127_, new_n9124_ );
or   ( new_n9357_, new_n9138_, new_n9135_ );
or   ( new_n9358_, new_n9149_, new_n9146_ );
or   ( new_n9359_, new_n9160_, new_n9157_ );
or   ( new_n9360_, new_n9171_, new_n9168_ );
or   ( new_n9361_, new_n9182_, new_n9179_ );
or   ( new_n9362_, new_n9193_, new_n9190_ );
or   ( new_n9363_, new_n9204_, new_n9201_ );
or   ( new_n9364_, new_n9215_, new_n9212_ );
or   ( new_n9365_, new_n9226_, new_n9223_ );
or   ( new_n9366_, new_n9237_, new_n9234_ );
or   ( new_n9367_, new_n9248_, new_n9245_ );
or   ( new_n9368_, new_n9259_, new_n9256_ );
or   ( new_n9369_, new_n9270_, new_n9267_ );
or   ( new_n9370_, new_n9286_, new_n9283_ );
and  ( new_n9371_, new_n9054_, new_n9052_ );
or   ( new_n9372_, new_n9371_, new_n8965_ );
or   ( new_n9373_, new_n9030_, new_n3548_ );
or   ( new_n9374_, new_n9373_, new_n9372_ );
and  ( new_n9375_, new_n9286_, new_n9283_ );
or   ( new_n9376_, new_n9375_, new_n9277_ );
or   ( new_n9377_, new_n9376_, new_n9374_ );
and  ( new_n9378_, new_n9377_, new_n9370_ );
and  ( new_n9379_, new_n9270_, new_n9267_ );
or   ( new_n9380_, new_n9379_, new_n9266_ );
or   ( new_n9381_, new_n9380_, new_n9378_ );
and  ( new_n9382_, new_n9381_, new_n9369_ );
and  ( new_n9383_, new_n9259_, new_n9256_ );
or   ( new_n9384_, new_n9383_, new_n9255_ );
or   ( new_n9385_, new_n9384_, new_n9382_ );
and  ( new_n9386_, new_n9385_, new_n9368_ );
and  ( new_n9387_, new_n9248_, new_n9245_ );
or   ( new_n9388_, new_n9387_, new_n9244_ );
or   ( new_n9389_, new_n9388_, new_n9386_ );
and  ( new_n9390_, new_n9389_, new_n9367_ );
and  ( new_n9391_, new_n9237_, new_n9234_ );
or   ( new_n9392_, new_n9391_, new_n9233_ );
or   ( new_n9393_, new_n9392_, new_n9390_ );
and  ( new_n9394_, new_n9393_, new_n9366_ );
and  ( new_n9395_, new_n9226_, new_n9223_ );
or   ( new_n9396_, new_n9395_, new_n9222_ );
or   ( new_n9397_, new_n9396_, new_n9394_ );
and  ( new_n9398_, new_n9397_, new_n9365_ );
and  ( new_n9399_, new_n9215_, new_n9212_ );
or   ( new_n9400_, new_n9399_, new_n9211_ );
or   ( new_n9401_, new_n9400_, new_n9398_ );
and  ( new_n9402_, new_n9401_, new_n9364_ );
and  ( new_n9403_, new_n9204_, new_n9201_ );
or   ( new_n9404_, new_n9403_, new_n9200_ );
or   ( new_n9405_, new_n9404_, new_n9402_ );
and  ( new_n9406_, new_n9405_, new_n9363_ );
and  ( new_n9407_, new_n9193_, new_n9190_ );
or   ( new_n9408_, new_n9407_, new_n9189_ );
or   ( new_n9409_, new_n9408_, new_n9406_ );
and  ( new_n9410_, new_n9409_, new_n9362_ );
and  ( new_n9411_, new_n9182_, new_n9179_ );
or   ( new_n9412_, new_n9411_, new_n9178_ );
or   ( new_n9413_, new_n9412_, new_n9410_ );
and  ( new_n9414_, new_n9413_, new_n9361_ );
and  ( new_n9415_, new_n9171_, new_n9168_ );
or   ( new_n9416_, new_n9415_, new_n9167_ );
or   ( new_n9417_, new_n9416_, new_n9414_ );
and  ( new_n9418_, new_n9417_, new_n9360_ );
and  ( new_n9419_, new_n9160_, new_n9157_ );
or   ( new_n9420_, new_n9419_, new_n9156_ );
or   ( new_n9421_, new_n9420_, new_n9418_ );
and  ( new_n9422_, new_n9421_, new_n9359_ );
and  ( new_n9423_, new_n9149_, new_n9146_ );
or   ( new_n9424_, new_n9423_, new_n9145_ );
or   ( new_n9425_, new_n9424_, new_n9422_ );
and  ( new_n9426_, new_n9425_, new_n9358_ );
and  ( new_n9427_, new_n9138_, new_n9135_ );
or   ( new_n9428_, new_n9427_, new_n9134_ );
or   ( new_n9429_, new_n9428_, new_n9426_ );
and  ( new_n9430_, new_n9429_, new_n9357_ );
and  ( new_n9431_, new_n9127_, new_n9124_ );
or   ( new_n9432_, new_n9431_, new_n9123_ );
or   ( new_n9433_, new_n9432_, new_n9430_ );
and  ( new_n9434_, new_n9433_, new_n9356_ );
and  ( new_n9435_, new_n9116_, new_n9031_ );
or   ( new_n9436_, new_n9435_, new_n9029_ );
or   ( new_n9437_, new_n9436_, new_n9434_ );
and  ( new_n9438_, new_n9437_, new_n9355_ );
and  ( new_n9439_, new_n9438_, new_n9350_ );
or   ( new_n9440_, new_n9439_, new_n9354_ );
and  ( new_n9441_, new_n9434_, new_n9118_ );
and  ( new_n9442_, new_n9436_, new_n9318_ );
or   ( new_n9443_, new_n9442_, new_n9441_ );
and  ( new_n9444_, new_n9349_, new_n3143_ );
and  ( new_n9445_, new_n9444_, new_n9443_ );
or   ( new_n9446_, new_n9352_, new_n2297_ );
and  ( new_n9447_, new_n9446_, new_n9443_ );
and  ( new_n9448_, new_n9436_, new_n9434_ );
or   ( new_n9449_, new_n9448_, new_n9319_ );
and  ( new_n9450_, new_n9449_, new_n9444_ );
or   ( new_n9451_, new_n9450_, new_n9447_ );
and  ( new_n9452_, new_n9430_, new_n9129_ );
and  ( new_n9453_, new_n9432_, new_n9316_ );
or   ( new_n9454_, new_n9453_, new_n9452_ );
and  ( new_n9455_, new_n9349_, new_n2420_ );
and  ( new_n9456_, new_n9455_, new_n9454_ );
or   ( new_n9457_, new_n9352_, new_n2288_ );
and  ( new_n9458_, new_n9457_, new_n9454_ );
and  ( new_n9459_, new_n9432_, new_n9430_ );
or   ( new_n9460_, new_n9459_, new_n9317_ );
and  ( new_n9461_, new_n9460_, new_n9455_ );
or   ( new_n9462_, new_n9461_, new_n9458_ );
and  ( new_n9463_, new_n9426_, new_n9140_ );
and  ( new_n9464_, new_n9428_, new_n9314_ );
or   ( new_n9465_, new_n9464_, new_n9463_ );
and  ( new_n9466_, new_n9349_, new_n3734_ );
and  ( new_n9467_, new_n9466_, new_n9465_ );
or   ( new_n9468_, new_n9352_, new_n2304_ );
and  ( new_n9469_, new_n9468_, new_n9465_ );
and  ( new_n9470_, new_n9428_, new_n9426_ );
or   ( new_n9471_, new_n9470_, new_n9315_ );
and  ( new_n9472_, new_n9471_, new_n9466_ );
or   ( new_n9473_, new_n9472_, new_n9469_ );
and  ( new_n9474_, new_n9422_, new_n9151_ );
and  ( new_n9475_, new_n9424_, new_n9312_ );
or   ( new_n9476_, new_n9475_, new_n9474_ );
and  ( new_n9477_, new_n9349_, new_n2441_ );
and  ( new_n9478_, new_n9477_, new_n9476_ );
or   ( new_n9479_, new_n9352_, new_n2440_ );
and  ( new_n9480_, new_n9479_, new_n9476_ );
and  ( new_n9481_, new_n9424_, new_n9422_ );
or   ( new_n9482_, new_n9481_, new_n9313_ );
and  ( new_n9483_, new_n9482_, new_n9477_ );
or   ( new_n9484_, new_n9483_, new_n9480_ );
and  ( new_n9485_, new_n9418_, new_n9162_ );
and  ( new_n9486_, new_n9420_, new_n9310_ );
or   ( new_n9487_, new_n9486_, new_n9485_ );
and  ( new_n9488_, new_n9349_, new_n6342_ );
and  ( new_n9489_, new_n9488_, new_n9487_ );
or   ( new_n9490_, new_n9352_, new_n2566_ );
and  ( new_n9491_, new_n9490_, new_n9487_ );
and  ( new_n9492_, new_n9420_, new_n9418_ );
or   ( new_n9493_, new_n9492_, new_n9311_ );
and  ( new_n9494_, new_n9493_, new_n9488_ );
or   ( new_n9495_, new_n9494_, new_n9491_ );
and  ( new_n9496_, new_n9414_, new_n9173_ );
and  ( new_n9497_, new_n9416_, new_n9308_ );
or   ( new_n9498_, new_n9497_, new_n9496_ );
and  ( new_n9499_, new_n9349_, new_n3693_ );
and  ( new_n9500_, new_n9499_, new_n9498_ );
or   ( new_n9501_, new_n9352_, new_n2705_ );
and  ( new_n9502_, new_n9501_, new_n9498_ );
and  ( new_n9503_, new_n9416_, new_n9414_ );
or   ( new_n9504_, new_n9503_, new_n9309_ );
and  ( new_n9505_, new_n9504_, new_n9499_ );
or   ( new_n9506_, new_n9505_, new_n9502_ );
and  ( new_n9507_, new_n9410_, new_n9184_ );
and  ( new_n9508_, new_n9412_, new_n9306_ );
or   ( new_n9509_, new_n9508_, new_n9507_ );
and  ( new_n9510_, new_n9349_, new_n4017_ );
and  ( new_n9511_, new_n9510_, new_n9509_ );
or   ( new_n9512_, new_n9352_, new_n2723_ );
and  ( new_n9513_, new_n9512_, new_n9509_ );
and  ( new_n9514_, new_n9412_, new_n9410_ );
or   ( new_n9515_, new_n9514_, new_n9307_ );
and  ( new_n9516_, new_n9515_, new_n9510_ );
or   ( new_n9517_, new_n9516_, new_n9513_ );
and  ( new_n9518_, new_n9406_, new_n9195_ );
and  ( new_n9519_, new_n9408_, new_n9304_ );
or   ( new_n9520_, new_n9519_, new_n9518_ );
and  ( new_n9521_, new_n9349_, new_n4085_ );
and  ( new_n9522_, new_n9521_, new_n9520_ );
or   ( new_n9523_, new_n9352_, new_n2760_ );
and  ( new_n9524_, new_n9523_, new_n9520_ );
and  ( new_n9525_, new_n9408_, new_n9406_ );
or   ( new_n9526_, new_n9525_, new_n9305_ );
and  ( new_n9527_, new_n9526_, new_n9521_ );
or   ( new_n9528_, new_n9527_, new_n9524_ );
and  ( new_n9529_, new_n9402_, new_n9206_ );
and  ( new_n9530_, new_n9404_, new_n9302_ );
or   ( new_n9531_, new_n9530_, new_n9529_ );
and  ( new_n9532_, new_n9349_, new_n2924_ );
and  ( new_n9533_, new_n9532_, new_n9531_ );
or   ( new_n9534_, new_n9352_, new_n2923_ );
and  ( new_n9535_, new_n9534_, new_n9531_ );
and  ( new_n9536_, new_n9404_, new_n9402_ );
or   ( new_n9537_, new_n9536_, new_n9303_ );
and  ( new_n9538_, new_n9537_, new_n9532_ );
or   ( new_n9539_, new_n9538_, new_n9535_ );
and  ( new_n9540_, new_n9398_, new_n9217_ );
and  ( new_n9541_, new_n9400_, new_n9300_ );
or   ( new_n9542_, new_n9541_, new_n9540_ );
and  ( new_n9543_, new_n9349_, new_n4177_ );
and  ( new_n9544_, new_n9543_, new_n9542_ );
or   ( new_n9545_, new_n9352_, new_n3066_ );
and  ( new_n9546_, new_n9545_, new_n9542_ );
and  ( new_n9547_, new_n9400_, new_n9398_ );
or   ( new_n9548_, new_n9547_, new_n9301_ );
and  ( new_n9549_, new_n9548_, new_n9543_ );
or   ( new_n9550_, new_n9549_, new_n9546_ );
and  ( new_n9551_, new_n9394_, new_n9228_ );
and  ( new_n9552_, new_n9396_, new_n9298_ );
or   ( new_n9553_, new_n9552_, new_n9551_ );
and  ( new_n9554_, new_n9349_, new_n3109_ );
and  ( new_n9555_, new_n9554_, new_n9553_ );
or   ( new_n9556_, new_n9352_, new_n3108_ );
and  ( new_n9557_, new_n9556_, new_n9553_ );
and  ( new_n9558_, new_n9396_, new_n9394_ );
or   ( new_n9559_, new_n9558_, new_n9299_ );
and  ( new_n9560_, new_n9559_, new_n9554_ );
or   ( new_n9561_, new_n9560_, new_n9557_ );
and  ( new_n9562_, new_n9390_, new_n9239_ );
and  ( new_n9563_, new_n9392_, new_n9296_ );
or   ( new_n9564_, new_n9563_, new_n9562_ );
and  ( new_n9565_, new_n9349_, new_n4257_ );
and  ( new_n9566_, new_n9565_, new_n9564_ );
or   ( new_n9567_, new_n9352_, new_n3244_ );
and  ( new_n9568_, new_n9567_, new_n9564_ );
and  ( new_n9569_, new_n9392_, new_n9390_ );
or   ( new_n9570_, new_n9569_, new_n9297_ );
and  ( new_n9571_, new_n9570_, new_n9565_ );
or   ( new_n9572_, new_n9571_, new_n9568_ );
and  ( new_n9573_, new_n9386_, new_n9250_ );
and  ( new_n9574_, new_n9388_, new_n9294_ );
or   ( new_n9575_, new_n9574_, new_n9573_ );
and  ( new_n9576_, new_n9349_, new_n4275_ );
and  ( new_n9577_, new_n9576_, new_n9575_ );
or   ( new_n9578_, new_n9352_, new_n3306_ );
and  ( new_n9579_, new_n9578_, new_n9575_ );
and  ( new_n9580_, new_n9388_, new_n9386_ );
or   ( new_n9581_, new_n9580_, new_n9295_ );
and  ( new_n9582_, new_n9581_, new_n9576_ );
or   ( new_n9583_, new_n9582_, new_n9579_ );
and  ( new_n9584_, new_n9382_, new_n9261_ );
and  ( new_n9585_, new_n9384_, new_n9292_ );
or   ( new_n9586_, new_n9585_, new_n9584_ );
and  ( new_n9587_, new_n9349_, new_n3407_ );
and  ( new_n9588_, new_n9587_, new_n9586_ );
or   ( new_n9589_, new_n9352_, new_n3406_ );
and  ( new_n9590_, new_n9589_, new_n9586_ );
and  ( new_n9591_, new_n9384_, new_n9382_ );
or   ( new_n9592_, new_n9591_, new_n9293_ );
and  ( new_n9593_, new_n9592_, new_n9587_ );
or   ( new_n9594_, new_n9593_, new_n9590_ );
and  ( new_n9595_, new_n9378_, new_n9272_ );
and  ( new_n9596_, new_n9380_, new_n9290_ );
or   ( new_n9597_, new_n9596_, new_n9595_ );
and  ( new_n9598_, new_n9349_, new_n4311_ );
and  ( new_n9599_, new_n9598_, new_n9597_ );
and  ( new_n9600_, new_n9374_, new_n9288_ );
and  ( new_n9601_, new_n9376_, new_n9282_ );
or   ( new_n9602_, new_n9601_, new_n9600_ );
and  ( new_n9603_, new_n9349_, new_n3547_ );
and  ( new_n9604_, new_n9603_, new_n9602_ );
or   ( new_n9605_, new_n9352_, new_n3507_ );
and  ( new_n9606_, new_n9605_, new_n9597_ );
and  ( new_n9607_, new_n9380_, new_n9378_ );
or   ( new_n9608_, new_n9607_, new_n9291_ );
and  ( new_n9609_, new_n9608_, new_n9598_ );
or   ( new_n9610_, new_n9609_, new_n9606_ );
and  ( new_n9611_, new_n9610_, new_n9604_ );
or   ( new_n9612_, new_n9611_, new_n9599_ );
and  ( new_n9613_, new_n9612_, new_n9594_ );
or   ( new_n9614_, new_n9613_, new_n9588_ );
and  ( new_n9615_, new_n9614_, new_n9583_ );
or   ( new_n9616_, new_n9615_, new_n9577_ );
and  ( new_n9617_, new_n9616_, new_n9572_ );
or   ( new_n9618_, new_n9617_, new_n9566_ );
and  ( new_n9619_, new_n9618_, new_n9561_ );
or   ( new_n9620_, new_n9619_, new_n9555_ );
and  ( new_n9621_, new_n9620_, new_n9550_ );
or   ( new_n9622_, new_n9621_, new_n9544_ );
and  ( new_n9623_, new_n9622_, new_n9539_ );
or   ( new_n9624_, new_n9623_, new_n9533_ );
and  ( new_n9625_, new_n9624_, new_n9528_ );
or   ( new_n9626_, new_n9625_, new_n9522_ );
and  ( new_n9627_, new_n9626_, new_n9517_ );
or   ( new_n9628_, new_n9627_, new_n9511_ );
and  ( new_n9629_, new_n9628_, new_n9506_ );
or   ( new_n9630_, new_n9629_, new_n9500_ );
and  ( new_n9631_, new_n9630_, new_n9495_ );
or   ( new_n9632_, new_n9631_, new_n9489_ );
and  ( new_n9633_, new_n9632_, new_n9484_ );
or   ( new_n9634_, new_n9633_, new_n9478_ );
and  ( new_n9635_, new_n9634_, new_n9473_ );
or   ( new_n9636_, new_n9635_, new_n9467_ );
and  ( new_n9637_, new_n9636_, new_n9462_ );
or   ( new_n9638_, new_n9637_, new_n9456_ );
and  ( new_n9639_, new_n9638_, new_n9451_ );
or   ( new_n9640_, new_n9639_, new_n9445_ );
and  ( new_n9641_, new_n9640_, new_n9440_ );
or   ( new_n9642_, new_n9641_, new_n9351_ );
xor  ( new_n9643_, new_n6037_, new_n968_ );
and  ( new_n9644_, new_n9643_, new_n5052_ );
not  ( new_n9645_, new_n9644_ );
and  ( new_n9646_, new_n5116_, \b[12]  );
not  ( new_n9647_, new_n2120_ );
and  ( new_n9648_, new_n5083_, new_n9647_ );
nor  ( new_n9649_, new_n9648_, new_n9646_ );
and  ( new_n9650_, new_n9649_, new_n9645_ );
nor  ( new_n9651_, new_n6500_, new_n2322_ );
nor  ( new_n9652_, new_n6503_, new_n2314_ );
nor  ( new_n9653_, new_n9652_, new_n9651_ );
and  ( new_n9654_, \c[12] , \b[12]  );
and  ( new_n9655_, new_n9654_, new_n5064_ );
and  ( new_n9656_, new_n5110_, \a[12]  );
nor  ( new_n9657_, new_n9656_, new_n9655_ );
and  ( new_n9658_, new_n9657_, new_n9653_ );
and  ( new_n9659_, new_n5056_, new_n2439_ );
not  ( new_n9660_, new_n9659_ );
xor  ( new_n9661_, new_n5498_, new_n275_ );
and  ( new_n9662_, new_n9661_, new_n5098_ );
or   ( new_n9663_, \b[12] , \a[12]  );
and  ( new_n9664_, new_n9663_, new_n5102_ );
nor  ( new_n9665_, new_n9664_, new_n9662_ );
and  ( new_n9666_, new_n9665_, new_n9660_ );
and  ( new_n9667_, new_n5072_, \d[12]  );
and  ( new_n9668_, new_n5092_, \c[12]  );
nor  ( new_n9669_, new_n9668_, new_n9667_ );
and  ( new_n9670_, new_n9669_, new_n9666_ );
and  ( new_n9671_, new_n9670_, new_n9658_ );
and  ( new_n9672_, new_n9671_, new_n9650_ );
not  ( new_n9673_, new_n9672_ );
and  ( new_n9674_, new_n9673_, new_n2407_ );
and  ( new_n9675_, new_n9674_, new_n9642_ );
and  ( new_n9676_, new_n9672_, new_n5120_ );
or   ( new_n9677_, new_n9676_, new_n2906_ );
and  ( new_n9678_, new_n9677_, new_n9642_ );
or   ( new_n9679_, new_n9438_, new_n9353_ );
or   ( new_n9680_, new_n9449_, new_n9446_ );
or   ( new_n9681_, new_n9460_, new_n9457_ );
or   ( new_n9682_, new_n9471_, new_n9468_ );
or   ( new_n9683_, new_n9482_, new_n9479_ );
or   ( new_n9684_, new_n9493_, new_n9490_ );
or   ( new_n9685_, new_n9504_, new_n9501_ );
or   ( new_n9686_, new_n9515_, new_n9512_ );
or   ( new_n9687_, new_n9526_, new_n9523_ );
or   ( new_n9688_, new_n9537_, new_n9534_ );
or   ( new_n9689_, new_n9548_, new_n9545_ );
or   ( new_n9690_, new_n9559_, new_n9556_ );
or   ( new_n9691_, new_n9570_, new_n9567_ );
or   ( new_n9692_, new_n9581_, new_n9578_ );
or   ( new_n9693_, new_n9592_, new_n9589_ );
or   ( new_n9694_, new_n9608_, new_n9605_ );
and  ( new_n9695_, new_n9376_, new_n9374_ );
or   ( new_n9696_, new_n9695_, new_n9289_ );
or   ( new_n9697_, new_n9352_, new_n3548_ );
or   ( new_n9698_, new_n9697_, new_n9696_ );
and  ( new_n9699_, new_n9608_, new_n9605_ );
or   ( new_n9700_, new_n9699_, new_n9599_ );
or   ( new_n9701_, new_n9700_, new_n9698_ );
and  ( new_n9702_, new_n9701_, new_n9694_ );
and  ( new_n9703_, new_n9592_, new_n9589_ );
or   ( new_n9704_, new_n9703_, new_n9588_ );
or   ( new_n9705_, new_n9704_, new_n9702_ );
and  ( new_n9706_, new_n9705_, new_n9693_ );
and  ( new_n9707_, new_n9581_, new_n9578_ );
or   ( new_n9708_, new_n9707_, new_n9577_ );
or   ( new_n9709_, new_n9708_, new_n9706_ );
and  ( new_n9710_, new_n9709_, new_n9692_ );
and  ( new_n9711_, new_n9570_, new_n9567_ );
or   ( new_n9712_, new_n9711_, new_n9566_ );
or   ( new_n9713_, new_n9712_, new_n9710_ );
and  ( new_n9714_, new_n9713_, new_n9691_ );
and  ( new_n9715_, new_n9559_, new_n9556_ );
or   ( new_n9716_, new_n9715_, new_n9555_ );
or   ( new_n9717_, new_n9716_, new_n9714_ );
and  ( new_n9718_, new_n9717_, new_n9690_ );
and  ( new_n9719_, new_n9548_, new_n9545_ );
or   ( new_n9720_, new_n9719_, new_n9544_ );
or   ( new_n9721_, new_n9720_, new_n9718_ );
and  ( new_n9722_, new_n9721_, new_n9689_ );
and  ( new_n9723_, new_n9537_, new_n9534_ );
or   ( new_n9724_, new_n9723_, new_n9533_ );
or   ( new_n9725_, new_n9724_, new_n9722_ );
and  ( new_n9726_, new_n9725_, new_n9688_ );
and  ( new_n9727_, new_n9526_, new_n9523_ );
or   ( new_n9728_, new_n9727_, new_n9522_ );
or   ( new_n9729_, new_n9728_, new_n9726_ );
and  ( new_n9730_, new_n9729_, new_n9687_ );
and  ( new_n9731_, new_n9515_, new_n9512_ );
or   ( new_n9732_, new_n9731_, new_n9511_ );
or   ( new_n9733_, new_n9732_, new_n9730_ );
and  ( new_n9734_, new_n9733_, new_n9686_ );
and  ( new_n9735_, new_n9504_, new_n9501_ );
or   ( new_n9736_, new_n9735_, new_n9500_ );
or   ( new_n9737_, new_n9736_, new_n9734_ );
and  ( new_n9738_, new_n9737_, new_n9685_ );
and  ( new_n9739_, new_n9493_, new_n9490_ );
or   ( new_n9740_, new_n9739_, new_n9489_ );
or   ( new_n9741_, new_n9740_, new_n9738_ );
and  ( new_n9742_, new_n9741_, new_n9684_ );
and  ( new_n9743_, new_n9482_, new_n9479_ );
or   ( new_n9744_, new_n9743_, new_n9478_ );
or   ( new_n9745_, new_n9744_, new_n9742_ );
and  ( new_n9746_, new_n9745_, new_n9683_ );
and  ( new_n9747_, new_n9471_, new_n9468_ );
or   ( new_n9748_, new_n9747_, new_n9467_ );
or   ( new_n9749_, new_n9748_, new_n9746_ );
and  ( new_n9750_, new_n9749_, new_n9682_ );
and  ( new_n9751_, new_n9460_, new_n9457_ );
or   ( new_n9752_, new_n9751_, new_n9456_ );
or   ( new_n9753_, new_n9752_, new_n9750_ );
and  ( new_n9754_, new_n9753_, new_n9681_ );
and  ( new_n9755_, new_n9449_, new_n9446_ );
or   ( new_n9756_, new_n9755_, new_n9445_ );
or   ( new_n9757_, new_n9756_, new_n9754_ );
and  ( new_n9758_, new_n9757_, new_n9680_ );
and  ( new_n9759_, new_n9438_, new_n9353_ );
or   ( new_n9760_, new_n9759_, new_n9351_ );
or   ( new_n9761_, new_n9760_, new_n9758_ );
and  ( new_n9762_, new_n9761_, new_n9679_ );
and  ( new_n9763_, new_n9762_, new_n9674_ );
or   ( new_n9764_, new_n9763_, new_n9678_ );
and  ( new_n9765_, new_n9758_, new_n9440_ );
and  ( new_n9766_, new_n9760_, new_n9640_ );
or   ( new_n9767_, new_n9766_, new_n9765_ );
and  ( new_n9768_, new_n9673_, new_n3143_ );
and  ( new_n9769_, new_n9768_, new_n9767_ );
or   ( new_n9770_, new_n9676_, new_n2297_ );
and  ( new_n9771_, new_n9770_, new_n9767_ );
and  ( new_n9772_, new_n9760_, new_n9758_ );
or   ( new_n9773_, new_n9772_, new_n9641_ );
and  ( new_n9774_, new_n9773_, new_n9768_ );
or   ( new_n9775_, new_n9774_, new_n9771_ );
and  ( new_n9776_, new_n9754_, new_n9451_ );
and  ( new_n9777_, new_n9756_, new_n9638_ );
or   ( new_n9778_, new_n9777_, new_n9776_ );
and  ( new_n9779_, new_n9673_, new_n2420_ );
and  ( new_n9780_, new_n9779_, new_n9778_ );
or   ( new_n9781_, new_n9676_, new_n2288_ );
and  ( new_n9782_, new_n9781_, new_n9778_ );
and  ( new_n9783_, new_n9756_, new_n9754_ );
or   ( new_n9784_, new_n9783_, new_n9639_ );
and  ( new_n9785_, new_n9784_, new_n9779_ );
or   ( new_n9786_, new_n9785_, new_n9782_ );
and  ( new_n9787_, new_n9750_, new_n9462_ );
and  ( new_n9788_, new_n9752_, new_n9636_ );
or   ( new_n9789_, new_n9788_, new_n9787_ );
and  ( new_n9790_, new_n9673_, new_n3734_ );
and  ( new_n9791_, new_n9790_, new_n9789_ );
or   ( new_n9792_, new_n9676_, new_n2304_ );
and  ( new_n9793_, new_n9792_, new_n9789_ );
and  ( new_n9794_, new_n9752_, new_n9750_ );
or   ( new_n9795_, new_n9794_, new_n9637_ );
and  ( new_n9796_, new_n9795_, new_n9790_ );
or   ( new_n9797_, new_n9796_, new_n9793_ );
and  ( new_n9798_, new_n9746_, new_n9473_ );
and  ( new_n9799_, new_n9748_, new_n9634_ );
or   ( new_n9800_, new_n9799_, new_n9798_ );
and  ( new_n9801_, new_n9673_, new_n2441_ );
and  ( new_n9802_, new_n9801_, new_n9800_ );
or   ( new_n9803_, new_n9676_, new_n2440_ );
and  ( new_n9804_, new_n9803_, new_n9800_ );
and  ( new_n9805_, new_n9748_, new_n9746_ );
or   ( new_n9806_, new_n9805_, new_n9635_ );
and  ( new_n9807_, new_n9806_, new_n9801_ );
or   ( new_n9808_, new_n9807_, new_n9804_ );
and  ( new_n9809_, new_n9742_, new_n9484_ );
and  ( new_n9810_, new_n9744_, new_n9632_ );
or   ( new_n9811_, new_n9810_, new_n9809_ );
and  ( new_n9812_, new_n9673_, new_n6342_ );
and  ( new_n9813_, new_n9812_, new_n9811_ );
or   ( new_n9814_, new_n9676_, new_n2566_ );
and  ( new_n9815_, new_n9814_, new_n9811_ );
and  ( new_n9816_, new_n9744_, new_n9742_ );
or   ( new_n9817_, new_n9816_, new_n9633_ );
and  ( new_n9818_, new_n9817_, new_n9812_ );
or   ( new_n9819_, new_n9818_, new_n9815_ );
and  ( new_n9820_, new_n9738_, new_n9495_ );
and  ( new_n9821_, new_n9740_, new_n9630_ );
or   ( new_n9822_, new_n9821_, new_n9820_ );
and  ( new_n9823_, new_n9673_, new_n3693_ );
and  ( new_n9824_, new_n9823_, new_n9822_ );
or   ( new_n9825_, new_n9676_, new_n2705_ );
and  ( new_n9826_, new_n9825_, new_n9822_ );
and  ( new_n9827_, new_n9740_, new_n9738_ );
or   ( new_n9828_, new_n9827_, new_n9631_ );
and  ( new_n9829_, new_n9828_, new_n9823_ );
or   ( new_n9830_, new_n9829_, new_n9826_ );
and  ( new_n9831_, new_n9734_, new_n9506_ );
and  ( new_n9832_, new_n9736_, new_n9628_ );
or   ( new_n9833_, new_n9832_, new_n9831_ );
and  ( new_n9834_, new_n9673_, new_n4017_ );
and  ( new_n9835_, new_n9834_, new_n9833_ );
or   ( new_n9836_, new_n9676_, new_n2723_ );
and  ( new_n9837_, new_n9836_, new_n9833_ );
and  ( new_n9838_, new_n9736_, new_n9734_ );
or   ( new_n9839_, new_n9838_, new_n9629_ );
and  ( new_n9840_, new_n9839_, new_n9834_ );
or   ( new_n9841_, new_n9840_, new_n9837_ );
and  ( new_n9842_, new_n9730_, new_n9517_ );
and  ( new_n9843_, new_n9732_, new_n9626_ );
or   ( new_n9844_, new_n9843_, new_n9842_ );
and  ( new_n9845_, new_n9673_, new_n4085_ );
and  ( new_n9846_, new_n9845_, new_n9844_ );
or   ( new_n9847_, new_n9676_, new_n2760_ );
and  ( new_n9848_, new_n9847_, new_n9844_ );
and  ( new_n9849_, new_n9732_, new_n9730_ );
or   ( new_n9850_, new_n9849_, new_n9627_ );
and  ( new_n9851_, new_n9850_, new_n9845_ );
or   ( new_n9852_, new_n9851_, new_n9848_ );
and  ( new_n9853_, new_n9726_, new_n9528_ );
and  ( new_n9854_, new_n9728_, new_n9624_ );
or   ( new_n9855_, new_n9854_, new_n9853_ );
and  ( new_n9856_, new_n9673_, new_n2924_ );
and  ( new_n9857_, new_n9856_, new_n9855_ );
or   ( new_n9858_, new_n9676_, new_n2923_ );
and  ( new_n9859_, new_n9858_, new_n9855_ );
and  ( new_n9860_, new_n9728_, new_n9726_ );
or   ( new_n9861_, new_n9860_, new_n9625_ );
and  ( new_n9862_, new_n9861_, new_n9856_ );
or   ( new_n9863_, new_n9862_, new_n9859_ );
and  ( new_n9864_, new_n9722_, new_n9539_ );
and  ( new_n9865_, new_n9724_, new_n9622_ );
or   ( new_n9866_, new_n9865_, new_n9864_ );
and  ( new_n9867_, new_n9673_, new_n4177_ );
and  ( new_n9868_, new_n9867_, new_n9866_ );
or   ( new_n9869_, new_n9676_, new_n3066_ );
and  ( new_n9870_, new_n9869_, new_n9866_ );
and  ( new_n9871_, new_n9724_, new_n9722_ );
or   ( new_n9872_, new_n9871_, new_n9623_ );
and  ( new_n9873_, new_n9872_, new_n9867_ );
or   ( new_n9874_, new_n9873_, new_n9870_ );
and  ( new_n9875_, new_n9718_, new_n9550_ );
and  ( new_n9876_, new_n9720_, new_n9620_ );
or   ( new_n9877_, new_n9876_, new_n9875_ );
and  ( new_n9878_, new_n9673_, new_n3109_ );
and  ( new_n9879_, new_n9878_, new_n9877_ );
or   ( new_n9880_, new_n9676_, new_n3108_ );
and  ( new_n9881_, new_n9880_, new_n9877_ );
and  ( new_n9882_, new_n9720_, new_n9718_ );
or   ( new_n9883_, new_n9882_, new_n9621_ );
and  ( new_n9884_, new_n9883_, new_n9878_ );
or   ( new_n9885_, new_n9884_, new_n9881_ );
and  ( new_n9886_, new_n9714_, new_n9561_ );
and  ( new_n9887_, new_n9716_, new_n9618_ );
or   ( new_n9888_, new_n9887_, new_n9886_ );
and  ( new_n9889_, new_n9673_, new_n4257_ );
and  ( new_n9890_, new_n9889_, new_n9888_ );
or   ( new_n9891_, new_n9676_, new_n3244_ );
and  ( new_n9892_, new_n9891_, new_n9888_ );
and  ( new_n9893_, new_n9716_, new_n9714_ );
or   ( new_n9894_, new_n9893_, new_n9619_ );
and  ( new_n9895_, new_n9894_, new_n9889_ );
or   ( new_n9896_, new_n9895_, new_n9892_ );
and  ( new_n9897_, new_n9710_, new_n9572_ );
and  ( new_n9898_, new_n9712_, new_n9616_ );
or   ( new_n9899_, new_n9898_, new_n9897_ );
and  ( new_n9900_, new_n9673_, new_n4275_ );
and  ( new_n9901_, new_n9900_, new_n9899_ );
or   ( new_n9902_, new_n9676_, new_n3306_ );
and  ( new_n9903_, new_n9902_, new_n9899_ );
and  ( new_n9904_, new_n9712_, new_n9710_ );
or   ( new_n9905_, new_n9904_, new_n9617_ );
and  ( new_n9906_, new_n9905_, new_n9900_ );
or   ( new_n9907_, new_n9906_, new_n9903_ );
and  ( new_n9908_, new_n9706_, new_n9583_ );
and  ( new_n9909_, new_n9708_, new_n9614_ );
or   ( new_n9910_, new_n9909_, new_n9908_ );
and  ( new_n9911_, new_n9673_, new_n3407_ );
and  ( new_n9912_, new_n9911_, new_n9910_ );
or   ( new_n9913_, new_n9676_, new_n3406_ );
and  ( new_n9914_, new_n9913_, new_n9910_ );
and  ( new_n9915_, new_n9708_, new_n9706_ );
or   ( new_n9916_, new_n9915_, new_n9615_ );
and  ( new_n9917_, new_n9916_, new_n9911_ );
or   ( new_n9918_, new_n9917_, new_n9914_ );
and  ( new_n9919_, new_n9702_, new_n9594_ );
and  ( new_n9920_, new_n9704_, new_n9612_ );
or   ( new_n9921_, new_n9920_, new_n9919_ );
and  ( new_n9922_, new_n9673_, new_n4311_ );
and  ( new_n9923_, new_n9922_, new_n9921_ );
and  ( new_n9924_, new_n9698_, new_n9610_ );
and  ( new_n9925_, new_n9700_, new_n9604_ );
or   ( new_n9926_, new_n9925_, new_n9924_ );
and  ( new_n9927_, new_n9673_, new_n3547_ );
and  ( new_n9928_, new_n9927_, new_n9926_ );
or   ( new_n9929_, new_n9676_, new_n3507_ );
and  ( new_n9930_, new_n9929_, new_n9921_ );
and  ( new_n9931_, new_n9704_, new_n9702_ );
or   ( new_n9932_, new_n9931_, new_n9613_ );
and  ( new_n9933_, new_n9932_, new_n9922_ );
or   ( new_n9934_, new_n9933_, new_n9930_ );
and  ( new_n9935_, new_n9934_, new_n9928_ );
or   ( new_n9936_, new_n9935_, new_n9923_ );
and  ( new_n9937_, new_n9936_, new_n9918_ );
or   ( new_n9938_, new_n9937_, new_n9912_ );
and  ( new_n9939_, new_n9938_, new_n9907_ );
or   ( new_n9940_, new_n9939_, new_n9901_ );
and  ( new_n9941_, new_n9940_, new_n9896_ );
or   ( new_n9942_, new_n9941_, new_n9890_ );
and  ( new_n9943_, new_n9942_, new_n9885_ );
or   ( new_n9944_, new_n9943_, new_n9879_ );
and  ( new_n9945_, new_n9944_, new_n9874_ );
or   ( new_n9946_, new_n9945_, new_n9868_ );
and  ( new_n9947_, new_n9946_, new_n9863_ );
or   ( new_n9948_, new_n9947_, new_n9857_ );
and  ( new_n9949_, new_n9948_, new_n9852_ );
or   ( new_n9950_, new_n9949_, new_n9846_ );
and  ( new_n9951_, new_n9950_, new_n9841_ );
or   ( new_n9952_, new_n9951_, new_n9835_ );
and  ( new_n9953_, new_n9952_, new_n9830_ );
or   ( new_n9954_, new_n9953_, new_n9824_ );
and  ( new_n9955_, new_n9954_, new_n9819_ );
or   ( new_n9956_, new_n9955_, new_n9813_ );
and  ( new_n9957_, new_n9956_, new_n9808_ );
or   ( new_n9958_, new_n9957_, new_n9802_ );
and  ( new_n9959_, new_n9958_, new_n9797_ );
or   ( new_n9960_, new_n9959_, new_n9791_ );
and  ( new_n9961_, new_n9960_, new_n9786_ );
or   ( new_n9962_, new_n9961_, new_n9780_ );
and  ( new_n9963_, new_n9962_, new_n9775_ );
or   ( new_n9964_, new_n9963_, new_n9769_ );
and  ( new_n9965_, new_n9964_, new_n9764_ );
or   ( new_n9966_, new_n9965_, new_n9675_ );
and  ( new_n9967_, new_n5083_, new_n2147_ );
not  ( new_n9968_, new_n9967_ );
xor  ( new_n9969_, new_n5568_, new_n277_ );
and  ( new_n9970_, new_n9969_, new_n5098_ );
or   ( new_n9971_, \b[13] , \a[13]  );
and  ( new_n9972_, new_n9971_, new_n5102_ );
nor  ( new_n9973_, new_n9972_, new_n9970_ );
and  ( new_n9974_, new_n9973_, new_n9968_ );
and  ( new_n9975_, new_n5110_, \a[13]  );
and  ( new_n9976_, new_n5092_, \c[13]  );
nor  ( new_n9977_, new_n9976_, new_n9975_ );
and  ( new_n9978_, new_n5076_, new_n2173_ );
and  ( new_n9979_, new_n5080_, new_n2169_ );
nor  ( new_n9980_, new_n9979_, new_n9978_ );
and  ( new_n9981_, new_n9980_, new_n9977_ );
and  ( new_n9982_, new_n9981_, new_n9974_ );
and  ( new_n9983_, new_n5064_, \c[13]  );
nor  ( new_n9984_, new_n9983_, new_n5116_ );
nor  ( new_n9985_, new_n9984_, new_n992_ );
not  ( new_n9986_, new_n9985_ );
xor  ( new_n9987_, new_n6107_, new_n972_ );
and  ( new_n9988_, new_n9987_, new_n5052_ );
not  ( new_n9989_, new_n9988_ );
and  ( new_n9990_, new_n5072_, \d[13]  );
and  ( new_n9991_, new_n5056_, new_n2157_ );
nor  ( new_n9992_, new_n9991_, new_n9990_ );
and  ( new_n9993_, new_n9992_, new_n9989_ );
and  ( new_n9994_, new_n9993_, new_n9986_ );
and  ( new_n9995_, new_n9994_, new_n9982_ );
not  ( new_n9996_, new_n9995_ );
and  ( new_n9997_, new_n9996_, new_n2407_ );
and  ( new_n9998_, new_n9997_, new_n9966_ );
and  ( new_n9999_, new_n9995_, new_n5120_ );
or   ( new_n10000_, new_n9999_, new_n2906_ );
and  ( new_n10001_, new_n10000_, new_n9966_ );
or   ( new_n10002_, new_n9762_, new_n9677_ );
or   ( new_n10003_, new_n9773_, new_n9770_ );
or   ( new_n10004_, new_n9784_, new_n9781_ );
or   ( new_n10005_, new_n9795_, new_n9792_ );
or   ( new_n10006_, new_n9806_, new_n9803_ );
or   ( new_n10007_, new_n9817_, new_n9814_ );
or   ( new_n10008_, new_n9828_, new_n9825_ );
or   ( new_n10009_, new_n9839_, new_n9836_ );
or   ( new_n10010_, new_n9850_, new_n9847_ );
or   ( new_n10011_, new_n9861_, new_n9858_ );
or   ( new_n10012_, new_n9872_, new_n9869_ );
or   ( new_n10013_, new_n9883_, new_n9880_ );
or   ( new_n10014_, new_n9894_, new_n9891_ );
or   ( new_n10015_, new_n9905_, new_n9902_ );
or   ( new_n10016_, new_n9916_, new_n9913_ );
or   ( new_n10017_, new_n9932_, new_n9929_ );
and  ( new_n10018_, new_n9700_, new_n9698_ );
or   ( new_n10019_, new_n10018_, new_n9611_ );
or   ( new_n10020_, new_n9676_, new_n3548_ );
or   ( new_n10021_, new_n10020_, new_n10019_ );
and  ( new_n10022_, new_n9932_, new_n9929_ );
or   ( new_n10023_, new_n10022_, new_n9923_ );
or   ( new_n10024_, new_n10023_, new_n10021_ );
and  ( new_n10025_, new_n10024_, new_n10017_ );
and  ( new_n10026_, new_n9916_, new_n9913_ );
or   ( new_n10027_, new_n10026_, new_n9912_ );
or   ( new_n10028_, new_n10027_, new_n10025_ );
and  ( new_n10029_, new_n10028_, new_n10016_ );
and  ( new_n10030_, new_n9905_, new_n9902_ );
or   ( new_n10031_, new_n10030_, new_n9901_ );
or   ( new_n10032_, new_n10031_, new_n10029_ );
and  ( new_n10033_, new_n10032_, new_n10015_ );
and  ( new_n10034_, new_n9894_, new_n9891_ );
or   ( new_n10035_, new_n10034_, new_n9890_ );
or   ( new_n10036_, new_n10035_, new_n10033_ );
and  ( new_n10037_, new_n10036_, new_n10014_ );
and  ( new_n10038_, new_n9883_, new_n9880_ );
or   ( new_n10039_, new_n10038_, new_n9879_ );
or   ( new_n10040_, new_n10039_, new_n10037_ );
and  ( new_n10041_, new_n10040_, new_n10013_ );
and  ( new_n10042_, new_n9872_, new_n9869_ );
or   ( new_n10043_, new_n10042_, new_n9868_ );
or   ( new_n10044_, new_n10043_, new_n10041_ );
and  ( new_n10045_, new_n10044_, new_n10012_ );
and  ( new_n10046_, new_n9861_, new_n9858_ );
or   ( new_n10047_, new_n10046_, new_n9857_ );
or   ( new_n10048_, new_n10047_, new_n10045_ );
and  ( new_n10049_, new_n10048_, new_n10011_ );
and  ( new_n10050_, new_n9850_, new_n9847_ );
or   ( new_n10051_, new_n10050_, new_n9846_ );
or   ( new_n10052_, new_n10051_, new_n10049_ );
and  ( new_n10053_, new_n10052_, new_n10010_ );
and  ( new_n10054_, new_n9839_, new_n9836_ );
or   ( new_n10055_, new_n10054_, new_n9835_ );
or   ( new_n10056_, new_n10055_, new_n10053_ );
and  ( new_n10057_, new_n10056_, new_n10009_ );
and  ( new_n10058_, new_n9828_, new_n9825_ );
or   ( new_n10059_, new_n10058_, new_n9824_ );
or   ( new_n10060_, new_n10059_, new_n10057_ );
and  ( new_n10061_, new_n10060_, new_n10008_ );
and  ( new_n10062_, new_n9817_, new_n9814_ );
or   ( new_n10063_, new_n10062_, new_n9813_ );
or   ( new_n10064_, new_n10063_, new_n10061_ );
and  ( new_n10065_, new_n10064_, new_n10007_ );
and  ( new_n10066_, new_n9806_, new_n9803_ );
or   ( new_n10067_, new_n10066_, new_n9802_ );
or   ( new_n10068_, new_n10067_, new_n10065_ );
and  ( new_n10069_, new_n10068_, new_n10006_ );
and  ( new_n10070_, new_n9795_, new_n9792_ );
or   ( new_n10071_, new_n10070_, new_n9791_ );
or   ( new_n10072_, new_n10071_, new_n10069_ );
and  ( new_n10073_, new_n10072_, new_n10005_ );
and  ( new_n10074_, new_n9784_, new_n9781_ );
or   ( new_n10075_, new_n10074_, new_n9780_ );
or   ( new_n10076_, new_n10075_, new_n10073_ );
and  ( new_n10077_, new_n10076_, new_n10004_ );
and  ( new_n10078_, new_n9773_, new_n9770_ );
or   ( new_n10079_, new_n10078_, new_n9769_ );
or   ( new_n10080_, new_n10079_, new_n10077_ );
and  ( new_n10081_, new_n10080_, new_n10003_ );
and  ( new_n10082_, new_n9762_, new_n9677_ );
or   ( new_n10083_, new_n10082_, new_n9675_ );
or   ( new_n10084_, new_n10083_, new_n10081_ );
and  ( new_n10085_, new_n10084_, new_n10002_ );
and  ( new_n10086_, new_n10085_, new_n9997_ );
or   ( new_n10087_, new_n10086_, new_n10001_ );
and  ( new_n10088_, new_n10081_, new_n9764_ );
and  ( new_n10089_, new_n10083_, new_n9964_ );
or   ( new_n10090_, new_n10089_, new_n10088_ );
and  ( new_n10091_, new_n9996_, new_n3143_ );
and  ( new_n10092_, new_n10091_, new_n10090_ );
or   ( new_n10093_, new_n9999_, new_n2297_ );
and  ( new_n10094_, new_n10093_, new_n10090_ );
and  ( new_n10095_, new_n10083_, new_n10081_ );
or   ( new_n10096_, new_n10095_, new_n9965_ );
and  ( new_n10097_, new_n10096_, new_n10091_ );
or   ( new_n10098_, new_n10097_, new_n10094_ );
and  ( new_n10099_, new_n10077_, new_n9775_ );
and  ( new_n10100_, new_n10079_, new_n9962_ );
or   ( new_n10101_, new_n10100_, new_n10099_ );
and  ( new_n10102_, new_n9996_, new_n2420_ );
and  ( new_n10103_, new_n10102_, new_n10101_ );
or   ( new_n10104_, new_n9999_, new_n2288_ );
and  ( new_n10105_, new_n10104_, new_n10101_ );
and  ( new_n10106_, new_n10079_, new_n10077_ );
or   ( new_n10107_, new_n10106_, new_n9963_ );
and  ( new_n10108_, new_n10107_, new_n10102_ );
or   ( new_n10109_, new_n10108_, new_n10105_ );
and  ( new_n10110_, new_n10073_, new_n9786_ );
and  ( new_n10111_, new_n10075_, new_n9960_ );
or   ( new_n10112_, new_n10111_, new_n10110_ );
and  ( new_n10113_, new_n9996_, new_n3734_ );
and  ( new_n10114_, new_n10113_, new_n10112_ );
or   ( new_n10115_, new_n9999_, new_n2304_ );
and  ( new_n10116_, new_n10115_, new_n10112_ );
and  ( new_n10117_, new_n10075_, new_n10073_ );
or   ( new_n10118_, new_n10117_, new_n9961_ );
and  ( new_n10119_, new_n10118_, new_n10113_ );
or   ( new_n10120_, new_n10119_, new_n10116_ );
and  ( new_n10121_, new_n10069_, new_n9797_ );
and  ( new_n10122_, new_n10071_, new_n9958_ );
or   ( new_n10123_, new_n10122_, new_n10121_ );
and  ( new_n10124_, new_n9996_, new_n2441_ );
and  ( new_n10125_, new_n10124_, new_n10123_ );
or   ( new_n10126_, new_n9999_, new_n2440_ );
and  ( new_n10127_, new_n10126_, new_n10123_ );
and  ( new_n10128_, new_n10071_, new_n10069_ );
or   ( new_n10129_, new_n10128_, new_n9959_ );
and  ( new_n10130_, new_n10129_, new_n10124_ );
or   ( new_n10131_, new_n10130_, new_n10127_ );
and  ( new_n10132_, new_n10065_, new_n9808_ );
and  ( new_n10133_, new_n10067_, new_n9956_ );
or   ( new_n10134_, new_n10133_, new_n10132_ );
and  ( new_n10135_, new_n9996_, new_n6342_ );
and  ( new_n10136_, new_n10135_, new_n10134_ );
or   ( new_n10137_, new_n9999_, new_n2566_ );
and  ( new_n10138_, new_n10137_, new_n10134_ );
and  ( new_n10139_, new_n10067_, new_n10065_ );
or   ( new_n10140_, new_n10139_, new_n9957_ );
and  ( new_n10141_, new_n10140_, new_n10135_ );
or   ( new_n10142_, new_n10141_, new_n10138_ );
and  ( new_n10143_, new_n10061_, new_n9819_ );
and  ( new_n10144_, new_n10063_, new_n9954_ );
or   ( new_n10145_, new_n10144_, new_n10143_ );
and  ( new_n10146_, new_n9996_, new_n3693_ );
and  ( new_n10147_, new_n10146_, new_n10145_ );
or   ( new_n10148_, new_n9999_, new_n2705_ );
and  ( new_n10149_, new_n10148_, new_n10145_ );
and  ( new_n10150_, new_n10063_, new_n10061_ );
or   ( new_n10151_, new_n10150_, new_n9955_ );
and  ( new_n10152_, new_n10151_, new_n10146_ );
or   ( new_n10153_, new_n10152_, new_n10149_ );
and  ( new_n10154_, new_n10057_, new_n9830_ );
and  ( new_n10155_, new_n10059_, new_n9952_ );
or   ( new_n10156_, new_n10155_, new_n10154_ );
and  ( new_n10157_, new_n9996_, new_n4017_ );
and  ( new_n10158_, new_n10157_, new_n10156_ );
or   ( new_n10159_, new_n9999_, new_n2723_ );
and  ( new_n10160_, new_n10159_, new_n10156_ );
and  ( new_n10161_, new_n10059_, new_n10057_ );
or   ( new_n10162_, new_n10161_, new_n9953_ );
and  ( new_n10163_, new_n10162_, new_n10157_ );
or   ( new_n10164_, new_n10163_, new_n10160_ );
and  ( new_n10165_, new_n10053_, new_n9841_ );
and  ( new_n10166_, new_n10055_, new_n9950_ );
or   ( new_n10167_, new_n10166_, new_n10165_ );
and  ( new_n10168_, new_n9996_, new_n4085_ );
and  ( new_n10169_, new_n10168_, new_n10167_ );
or   ( new_n10170_, new_n9999_, new_n2760_ );
and  ( new_n10171_, new_n10170_, new_n10167_ );
and  ( new_n10172_, new_n10055_, new_n10053_ );
or   ( new_n10173_, new_n10172_, new_n9951_ );
and  ( new_n10174_, new_n10173_, new_n10168_ );
or   ( new_n10175_, new_n10174_, new_n10171_ );
and  ( new_n10176_, new_n10049_, new_n9852_ );
and  ( new_n10177_, new_n10051_, new_n9948_ );
or   ( new_n10178_, new_n10177_, new_n10176_ );
and  ( new_n10179_, new_n9996_, new_n2924_ );
and  ( new_n10180_, new_n10179_, new_n10178_ );
or   ( new_n10181_, new_n9999_, new_n2923_ );
and  ( new_n10182_, new_n10181_, new_n10178_ );
and  ( new_n10183_, new_n10051_, new_n10049_ );
or   ( new_n10184_, new_n10183_, new_n9949_ );
and  ( new_n10185_, new_n10184_, new_n10179_ );
or   ( new_n10186_, new_n10185_, new_n10182_ );
and  ( new_n10187_, new_n10045_, new_n9863_ );
and  ( new_n10188_, new_n10047_, new_n9946_ );
or   ( new_n10189_, new_n10188_, new_n10187_ );
and  ( new_n10190_, new_n9996_, new_n4177_ );
and  ( new_n10191_, new_n10190_, new_n10189_ );
or   ( new_n10192_, new_n9999_, new_n3066_ );
and  ( new_n10193_, new_n10192_, new_n10189_ );
and  ( new_n10194_, new_n10047_, new_n10045_ );
or   ( new_n10195_, new_n10194_, new_n9947_ );
and  ( new_n10196_, new_n10195_, new_n10190_ );
or   ( new_n10197_, new_n10196_, new_n10193_ );
and  ( new_n10198_, new_n10041_, new_n9874_ );
and  ( new_n10199_, new_n10043_, new_n9944_ );
or   ( new_n10200_, new_n10199_, new_n10198_ );
and  ( new_n10201_, new_n9996_, new_n3109_ );
and  ( new_n10202_, new_n10201_, new_n10200_ );
or   ( new_n10203_, new_n9999_, new_n3108_ );
and  ( new_n10204_, new_n10203_, new_n10200_ );
and  ( new_n10205_, new_n10043_, new_n10041_ );
or   ( new_n10206_, new_n10205_, new_n9945_ );
and  ( new_n10207_, new_n10206_, new_n10201_ );
or   ( new_n10208_, new_n10207_, new_n10204_ );
and  ( new_n10209_, new_n10037_, new_n9885_ );
and  ( new_n10210_, new_n10039_, new_n9942_ );
or   ( new_n10211_, new_n10210_, new_n10209_ );
and  ( new_n10212_, new_n9996_, new_n4257_ );
and  ( new_n10213_, new_n10212_, new_n10211_ );
or   ( new_n10214_, new_n9999_, new_n3244_ );
and  ( new_n10215_, new_n10214_, new_n10211_ );
and  ( new_n10216_, new_n10039_, new_n10037_ );
or   ( new_n10217_, new_n10216_, new_n9943_ );
and  ( new_n10218_, new_n10217_, new_n10212_ );
or   ( new_n10219_, new_n10218_, new_n10215_ );
and  ( new_n10220_, new_n10033_, new_n9896_ );
and  ( new_n10221_, new_n10035_, new_n9940_ );
or   ( new_n10222_, new_n10221_, new_n10220_ );
and  ( new_n10223_, new_n9996_, new_n4275_ );
and  ( new_n10224_, new_n10223_, new_n10222_ );
or   ( new_n10225_, new_n9999_, new_n3306_ );
and  ( new_n10226_, new_n10225_, new_n10222_ );
and  ( new_n10227_, new_n10035_, new_n10033_ );
or   ( new_n10228_, new_n10227_, new_n9941_ );
and  ( new_n10229_, new_n10228_, new_n10223_ );
or   ( new_n10230_, new_n10229_, new_n10226_ );
and  ( new_n10231_, new_n10029_, new_n9907_ );
and  ( new_n10232_, new_n10031_, new_n9938_ );
or   ( new_n10233_, new_n10232_, new_n10231_ );
and  ( new_n10234_, new_n9996_, new_n3407_ );
and  ( new_n10235_, new_n10234_, new_n10233_ );
or   ( new_n10236_, new_n9999_, new_n3406_ );
and  ( new_n10237_, new_n10236_, new_n10233_ );
and  ( new_n10238_, new_n10031_, new_n10029_ );
or   ( new_n10239_, new_n10238_, new_n9939_ );
and  ( new_n10240_, new_n10239_, new_n10234_ );
or   ( new_n10241_, new_n10240_, new_n10237_ );
and  ( new_n10242_, new_n10025_, new_n9918_ );
and  ( new_n10243_, new_n10027_, new_n9936_ );
or   ( new_n10244_, new_n10243_, new_n10242_ );
and  ( new_n10245_, new_n9996_, new_n4311_ );
and  ( new_n10246_, new_n10245_, new_n10244_ );
and  ( new_n10247_, new_n10021_, new_n9934_ );
and  ( new_n10248_, new_n10023_, new_n9928_ );
or   ( new_n10249_, new_n10248_, new_n10247_ );
and  ( new_n10250_, new_n9996_, new_n3547_ );
and  ( new_n10251_, new_n10250_, new_n10249_ );
or   ( new_n10252_, new_n9999_, new_n3507_ );
and  ( new_n10253_, new_n10252_, new_n10244_ );
and  ( new_n10254_, new_n10027_, new_n10025_ );
or   ( new_n10255_, new_n10254_, new_n9937_ );
and  ( new_n10256_, new_n10255_, new_n10245_ );
or   ( new_n10257_, new_n10256_, new_n10253_ );
and  ( new_n10258_, new_n10257_, new_n10251_ );
or   ( new_n10259_, new_n10258_, new_n10246_ );
and  ( new_n10260_, new_n10259_, new_n10241_ );
or   ( new_n10261_, new_n10260_, new_n10235_ );
and  ( new_n10262_, new_n10261_, new_n10230_ );
or   ( new_n10263_, new_n10262_, new_n10224_ );
and  ( new_n10264_, new_n10263_, new_n10219_ );
or   ( new_n10265_, new_n10264_, new_n10213_ );
and  ( new_n10266_, new_n10265_, new_n10208_ );
or   ( new_n10267_, new_n10266_, new_n10202_ );
and  ( new_n10268_, new_n10267_, new_n10197_ );
or   ( new_n10269_, new_n10268_, new_n10191_ );
and  ( new_n10270_, new_n10269_, new_n10186_ );
or   ( new_n10271_, new_n10270_, new_n10180_ );
and  ( new_n10272_, new_n10271_, new_n10175_ );
or   ( new_n10273_, new_n10272_, new_n10169_ );
and  ( new_n10274_, new_n10273_, new_n10164_ );
or   ( new_n10275_, new_n10274_, new_n10158_ );
and  ( new_n10276_, new_n10275_, new_n10153_ );
or   ( new_n10277_, new_n10276_, new_n10147_ );
and  ( new_n10278_, new_n10277_, new_n10142_ );
or   ( new_n10279_, new_n10278_, new_n10136_ );
and  ( new_n10280_, new_n10279_, new_n10131_ );
or   ( new_n10281_, new_n10280_, new_n10125_ );
and  ( new_n10282_, new_n10281_, new_n10120_ );
or   ( new_n10283_, new_n10282_, new_n10114_ );
and  ( new_n10284_, new_n10283_, new_n10109_ );
or   ( new_n10285_, new_n10284_, new_n10103_ );
and  ( new_n10286_, new_n10285_, new_n10098_ );
or   ( new_n10287_, new_n10286_, new_n10092_ );
and  ( new_n10288_, new_n10287_, new_n10087_ );
or   ( new_n10289_, new_n10288_, new_n9998_ );
and  ( new_n10290_, new_n10289_, new_n6196_ );
or   ( new_n10291_, new_n10085_, new_n10000_ );
or   ( new_n10292_, new_n10096_, new_n10093_ );
or   ( new_n10293_, new_n10107_, new_n10104_ );
or   ( new_n10294_, new_n10118_, new_n10115_ );
or   ( new_n10295_, new_n10129_, new_n10126_ );
or   ( new_n10296_, new_n10140_, new_n10137_ );
or   ( new_n10297_, new_n10151_, new_n10148_ );
or   ( new_n10298_, new_n10162_, new_n10159_ );
or   ( new_n10299_, new_n10173_, new_n10170_ );
or   ( new_n10300_, new_n10184_, new_n10181_ );
or   ( new_n10301_, new_n10195_, new_n10192_ );
or   ( new_n10302_, new_n10206_, new_n10203_ );
or   ( new_n10303_, new_n10217_, new_n10214_ );
or   ( new_n10304_, new_n10228_, new_n10225_ );
or   ( new_n10305_, new_n10239_, new_n10236_ );
or   ( new_n10306_, new_n10255_, new_n10252_ );
and  ( new_n10307_, new_n10023_, new_n10021_ );
or   ( new_n10308_, new_n10307_, new_n9935_ );
or   ( new_n10309_, new_n9999_, new_n3548_ );
or   ( new_n10310_, new_n10309_, new_n10308_ );
and  ( new_n10311_, new_n10255_, new_n10252_ );
or   ( new_n10312_, new_n10311_, new_n10246_ );
or   ( new_n10313_, new_n10312_, new_n10310_ );
and  ( new_n10314_, new_n10313_, new_n10306_ );
and  ( new_n10315_, new_n10239_, new_n10236_ );
or   ( new_n10316_, new_n10315_, new_n10235_ );
or   ( new_n10317_, new_n10316_, new_n10314_ );
and  ( new_n10318_, new_n10317_, new_n10305_ );
and  ( new_n10319_, new_n10228_, new_n10225_ );
or   ( new_n10320_, new_n10319_, new_n10224_ );
or   ( new_n10321_, new_n10320_, new_n10318_ );
and  ( new_n10322_, new_n10321_, new_n10304_ );
and  ( new_n10323_, new_n10217_, new_n10214_ );
or   ( new_n10324_, new_n10323_, new_n10213_ );
or   ( new_n10325_, new_n10324_, new_n10322_ );
and  ( new_n10326_, new_n10325_, new_n10303_ );
and  ( new_n10327_, new_n10206_, new_n10203_ );
or   ( new_n10328_, new_n10327_, new_n10202_ );
or   ( new_n10329_, new_n10328_, new_n10326_ );
and  ( new_n10330_, new_n10329_, new_n10302_ );
and  ( new_n10331_, new_n10195_, new_n10192_ );
or   ( new_n10332_, new_n10331_, new_n10191_ );
or   ( new_n10333_, new_n10332_, new_n10330_ );
and  ( new_n10334_, new_n10333_, new_n10301_ );
and  ( new_n10335_, new_n10184_, new_n10181_ );
or   ( new_n10336_, new_n10335_, new_n10180_ );
or   ( new_n10337_, new_n10336_, new_n10334_ );
and  ( new_n10338_, new_n10337_, new_n10300_ );
and  ( new_n10339_, new_n10173_, new_n10170_ );
or   ( new_n10340_, new_n10339_, new_n10169_ );
or   ( new_n10341_, new_n10340_, new_n10338_ );
and  ( new_n10342_, new_n10341_, new_n10299_ );
and  ( new_n10343_, new_n10162_, new_n10159_ );
or   ( new_n10344_, new_n10343_, new_n10158_ );
or   ( new_n10345_, new_n10344_, new_n10342_ );
and  ( new_n10346_, new_n10345_, new_n10298_ );
and  ( new_n10347_, new_n10151_, new_n10148_ );
or   ( new_n10348_, new_n10347_, new_n10147_ );
or   ( new_n10349_, new_n10348_, new_n10346_ );
and  ( new_n10350_, new_n10349_, new_n10297_ );
and  ( new_n10351_, new_n10140_, new_n10137_ );
or   ( new_n10352_, new_n10351_, new_n10136_ );
or   ( new_n10353_, new_n10352_, new_n10350_ );
and  ( new_n10354_, new_n10353_, new_n10296_ );
and  ( new_n10355_, new_n10129_, new_n10126_ );
or   ( new_n10356_, new_n10355_, new_n10125_ );
or   ( new_n10357_, new_n10356_, new_n10354_ );
and  ( new_n10358_, new_n10357_, new_n10295_ );
and  ( new_n10359_, new_n10118_, new_n10115_ );
or   ( new_n10360_, new_n10359_, new_n10114_ );
or   ( new_n10361_, new_n10360_, new_n10358_ );
and  ( new_n10362_, new_n10361_, new_n10294_ );
and  ( new_n10363_, new_n10107_, new_n10104_ );
or   ( new_n10364_, new_n10363_, new_n10103_ );
or   ( new_n10365_, new_n10364_, new_n10362_ );
and  ( new_n10366_, new_n10365_, new_n10293_ );
and  ( new_n10367_, new_n10096_, new_n10093_ );
or   ( new_n10368_, new_n10367_, new_n10092_ );
or   ( new_n10369_, new_n10368_, new_n10366_ );
and  ( new_n10370_, new_n10369_, new_n10292_ );
and  ( new_n10371_, new_n10085_, new_n10000_ );
or   ( new_n10372_, new_n10371_, new_n9998_ );
or   ( new_n10373_, new_n10372_, new_n10370_ );
and  ( new_n10374_, new_n10373_, new_n10291_ );
not  ( new_n10375_, new_n6194_ );
and  ( new_n10376_, new_n10375_, new_n2407_ );
and  ( new_n10377_, new_n10376_, new_n10374_ );
or   ( new_n10378_, new_n10377_, new_n10290_ );
and  ( new_n10379_, new_n10370_, new_n10087_ );
and  ( new_n10380_, new_n10372_, new_n10287_ );
or   ( new_n10381_, new_n10380_, new_n10379_ );
and  ( new_n10382_, new_n10375_, new_n3143_ );
and  ( new_n10383_, new_n10382_, new_n10381_ );
or   ( new_n10384_, new_n6195_, new_n2297_ );
and  ( new_n10385_, new_n10384_, new_n10381_ );
and  ( new_n10386_, new_n10372_, new_n10370_ );
or   ( new_n10387_, new_n10386_, new_n10288_ );
and  ( new_n10388_, new_n10387_, new_n10382_ );
or   ( new_n10389_, new_n10388_, new_n10385_ );
and  ( new_n10390_, new_n10366_, new_n10098_ );
and  ( new_n10391_, new_n10368_, new_n10285_ );
or   ( new_n10392_, new_n10391_, new_n10390_ );
and  ( new_n10393_, new_n10375_, new_n2420_ );
and  ( new_n10394_, new_n10393_, new_n10392_ );
or   ( new_n10395_, new_n6195_, new_n2288_ );
and  ( new_n10396_, new_n10395_, new_n10392_ );
and  ( new_n10397_, new_n10368_, new_n10366_ );
or   ( new_n10398_, new_n10397_, new_n10286_ );
and  ( new_n10399_, new_n10398_, new_n10393_ );
or   ( new_n10400_, new_n10399_, new_n10396_ );
and  ( new_n10401_, new_n10362_, new_n10109_ );
and  ( new_n10402_, new_n10364_, new_n10283_ );
or   ( new_n10403_, new_n10402_, new_n10401_ );
and  ( new_n10404_, new_n10375_, new_n3734_ );
and  ( new_n10405_, new_n10404_, new_n10403_ );
or   ( new_n10406_, new_n6195_, new_n2304_ );
and  ( new_n10407_, new_n10406_, new_n10403_ );
and  ( new_n10408_, new_n10364_, new_n10362_ );
or   ( new_n10409_, new_n10408_, new_n10284_ );
and  ( new_n10410_, new_n10409_, new_n10404_ );
or   ( new_n10411_, new_n10410_, new_n10407_ );
and  ( new_n10412_, new_n10358_, new_n10120_ );
and  ( new_n10413_, new_n10360_, new_n10281_ );
or   ( new_n10414_, new_n10413_, new_n10412_ );
and  ( new_n10415_, new_n10375_, new_n2441_ );
and  ( new_n10416_, new_n10415_, new_n10414_ );
or   ( new_n10417_, new_n6195_, new_n2440_ );
and  ( new_n10418_, new_n10417_, new_n10414_ );
and  ( new_n10419_, new_n10360_, new_n10358_ );
or   ( new_n10420_, new_n10419_, new_n10282_ );
and  ( new_n10421_, new_n10420_, new_n10415_ );
or   ( new_n10422_, new_n10421_, new_n10418_ );
and  ( new_n10423_, new_n10354_, new_n10131_ );
and  ( new_n10424_, new_n10356_, new_n10279_ );
or   ( new_n10425_, new_n10424_, new_n10423_ );
and  ( new_n10426_, new_n10375_, new_n6342_ );
and  ( new_n10427_, new_n10426_, new_n10425_ );
or   ( new_n10428_, new_n6195_, new_n2566_ );
and  ( new_n10429_, new_n10428_, new_n10425_ );
and  ( new_n10430_, new_n10356_, new_n10354_ );
or   ( new_n10431_, new_n10430_, new_n10280_ );
and  ( new_n10432_, new_n10431_, new_n10426_ );
or   ( new_n10433_, new_n10432_, new_n10429_ );
and  ( new_n10434_, new_n10350_, new_n10142_ );
and  ( new_n10435_, new_n10352_, new_n10277_ );
or   ( new_n10436_, new_n10435_, new_n10434_ );
and  ( new_n10437_, new_n10375_, new_n3693_ );
and  ( new_n10438_, new_n10437_, new_n10436_ );
or   ( new_n10439_, new_n6195_, new_n2705_ );
and  ( new_n10440_, new_n10439_, new_n10436_ );
and  ( new_n10441_, new_n10352_, new_n10350_ );
or   ( new_n10442_, new_n10441_, new_n10278_ );
and  ( new_n10443_, new_n10442_, new_n10437_ );
or   ( new_n10444_, new_n10443_, new_n10440_ );
and  ( new_n10445_, new_n10346_, new_n10153_ );
and  ( new_n10446_, new_n10348_, new_n10275_ );
or   ( new_n10447_, new_n10446_, new_n10445_ );
and  ( new_n10448_, new_n10375_, new_n4017_ );
and  ( new_n10449_, new_n10448_, new_n10447_ );
or   ( new_n10450_, new_n6195_, new_n2723_ );
and  ( new_n10451_, new_n10450_, new_n10447_ );
and  ( new_n10452_, new_n10348_, new_n10346_ );
or   ( new_n10453_, new_n10452_, new_n10276_ );
and  ( new_n10454_, new_n10453_, new_n10448_ );
or   ( new_n10455_, new_n10454_, new_n10451_ );
and  ( new_n10456_, new_n10342_, new_n10164_ );
and  ( new_n10457_, new_n10344_, new_n10273_ );
or   ( new_n10458_, new_n10457_, new_n10456_ );
and  ( new_n10459_, new_n10375_, new_n4085_ );
and  ( new_n10460_, new_n10459_, new_n10458_ );
or   ( new_n10461_, new_n6195_, new_n2760_ );
and  ( new_n10462_, new_n10461_, new_n10458_ );
and  ( new_n10463_, new_n10344_, new_n10342_ );
or   ( new_n10464_, new_n10463_, new_n10274_ );
and  ( new_n10465_, new_n10464_, new_n10459_ );
or   ( new_n10466_, new_n10465_, new_n10462_ );
and  ( new_n10467_, new_n10338_, new_n10175_ );
and  ( new_n10468_, new_n10340_, new_n10271_ );
or   ( new_n10469_, new_n10468_, new_n10467_ );
and  ( new_n10470_, new_n10375_, new_n2924_ );
and  ( new_n10471_, new_n10470_, new_n10469_ );
or   ( new_n10472_, new_n6195_, new_n2923_ );
and  ( new_n10473_, new_n10472_, new_n10469_ );
and  ( new_n10474_, new_n10340_, new_n10338_ );
or   ( new_n10475_, new_n10474_, new_n10272_ );
and  ( new_n10476_, new_n10475_, new_n10470_ );
or   ( new_n10477_, new_n10476_, new_n10473_ );
and  ( new_n10478_, new_n10334_, new_n10186_ );
and  ( new_n10479_, new_n10336_, new_n10269_ );
or   ( new_n10480_, new_n10479_, new_n10478_ );
and  ( new_n10481_, new_n10375_, new_n4177_ );
and  ( new_n10482_, new_n10481_, new_n10480_ );
or   ( new_n10483_, new_n6195_, new_n3066_ );
and  ( new_n10484_, new_n10483_, new_n10480_ );
and  ( new_n10485_, new_n10336_, new_n10334_ );
or   ( new_n10486_, new_n10485_, new_n10270_ );
and  ( new_n10487_, new_n10486_, new_n10481_ );
or   ( new_n10488_, new_n10487_, new_n10484_ );
and  ( new_n10489_, new_n10330_, new_n10197_ );
and  ( new_n10490_, new_n10332_, new_n10267_ );
or   ( new_n10491_, new_n10490_, new_n10489_ );
and  ( new_n10492_, new_n10375_, new_n3109_ );
and  ( new_n10493_, new_n10492_, new_n10491_ );
or   ( new_n10494_, new_n6195_, new_n3108_ );
and  ( new_n10495_, new_n10494_, new_n10491_ );
and  ( new_n10496_, new_n10332_, new_n10330_ );
or   ( new_n10497_, new_n10496_, new_n10268_ );
and  ( new_n10498_, new_n10497_, new_n10492_ );
or   ( new_n10499_, new_n10498_, new_n10495_ );
and  ( new_n10500_, new_n10326_, new_n10208_ );
and  ( new_n10501_, new_n10328_, new_n10265_ );
or   ( new_n10502_, new_n10501_, new_n10500_ );
and  ( new_n10503_, new_n10375_, new_n4257_ );
and  ( new_n10504_, new_n10503_, new_n10502_ );
or   ( new_n10505_, new_n6195_, new_n3244_ );
and  ( new_n10506_, new_n10505_, new_n10502_ );
and  ( new_n10507_, new_n10328_, new_n10326_ );
or   ( new_n10508_, new_n10507_, new_n10266_ );
and  ( new_n10509_, new_n10508_, new_n10503_ );
or   ( new_n10510_, new_n10509_, new_n10506_ );
and  ( new_n10511_, new_n10322_, new_n10219_ );
and  ( new_n10512_, new_n10324_, new_n10263_ );
or   ( new_n10513_, new_n10512_, new_n10511_ );
and  ( new_n10514_, new_n10375_, new_n4275_ );
and  ( new_n10515_, new_n10514_, new_n10513_ );
or   ( new_n10516_, new_n6195_, new_n3306_ );
and  ( new_n10517_, new_n10516_, new_n10513_ );
and  ( new_n10518_, new_n10324_, new_n10322_ );
or   ( new_n10519_, new_n10518_, new_n10264_ );
and  ( new_n10520_, new_n10519_, new_n10514_ );
or   ( new_n10521_, new_n10520_, new_n10517_ );
and  ( new_n10522_, new_n10318_, new_n10230_ );
and  ( new_n10523_, new_n10320_, new_n10261_ );
or   ( new_n10524_, new_n10523_, new_n10522_ );
and  ( new_n10525_, new_n10375_, new_n3407_ );
and  ( new_n10526_, new_n10525_, new_n10524_ );
or   ( new_n10527_, new_n6195_, new_n3406_ );
and  ( new_n10528_, new_n10527_, new_n10524_ );
and  ( new_n10529_, new_n10320_, new_n10318_ );
or   ( new_n10530_, new_n10529_, new_n10262_ );
and  ( new_n10531_, new_n10530_, new_n10525_ );
or   ( new_n10532_, new_n10531_, new_n10528_ );
and  ( new_n10533_, new_n10314_, new_n10241_ );
and  ( new_n10534_, new_n10316_, new_n10259_ );
or   ( new_n10535_, new_n10534_, new_n10533_ );
and  ( new_n10536_, new_n10375_, new_n4311_ );
and  ( new_n10537_, new_n10536_, new_n10535_ );
and  ( new_n10538_, new_n10310_, new_n10257_ );
and  ( new_n10539_, new_n10312_, new_n10251_ );
or   ( new_n10540_, new_n10539_, new_n10538_ );
and  ( new_n10541_, new_n10375_, new_n3547_ );
and  ( new_n10542_, new_n10541_, new_n10540_ );
or   ( new_n10543_, new_n6195_, new_n3507_ );
and  ( new_n10544_, new_n10543_, new_n10535_ );
and  ( new_n10545_, new_n10316_, new_n10314_ );
or   ( new_n10546_, new_n10545_, new_n10260_ );
and  ( new_n10547_, new_n10546_, new_n10536_ );
or   ( new_n10548_, new_n10547_, new_n10544_ );
and  ( new_n10549_, new_n10548_, new_n10542_ );
or   ( new_n10550_, new_n10549_, new_n10537_ );
and  ( new_n10551_, new_n10550_, new_n10532_ );
or   ( new_n10552_, new_n10551_, new_n10526_ );
and  ( new_n10553_, new_n10552_, new_n10521_ );
or   ( new_n10554_, new_n10553_, new_n10515_ );
and  ( new_n10555_, new_n10554_, new_n10510_ );
or   ( new_n10556_, new_n10555_, new_n10504_ );
and  ( new_n10557_, new_n10556_, new_n10499_ );
or   ( new_n10558_, new_n10557_, new_n10493_ );
and  ( new_n10559_, new_n10558_, new_n10488_ );
or   ( new_n10560_, new_n10559_, new_n10482_ );
and  ( new_n10561_, new_n10560_, new_n10477_ );
or   ( new_n10562_, new_n10561_, new_n10471_ );
and  ( new_n10563_, new_n10562_, new_n10466_ );
or   ( new_n10564_, new_n10563_, new_n10460_ );
and  ( new_n10565_, new_n10564_, new_n10455_ );
or   ( new_n10566_, new_n10565_, new_n10449_ );
and  ( new_n10567_, new_n10566_, new_n10444_ );
or   ( new_n10568_, new_n10567_, new_n10438_ );
and  ( new_n10569_, new_n10568_, new_n10433_ );
or   ( new_n10570_, new_n10569_, new_n10427_ );
and  ( new_n10571_, new_n10570_, new_n10422_ );
or   ( new_n10572_, new_n10571_, new_n10416_ );
and  ( new_n10573_, new_n10572_, new_n10411_ );
or   ( new_n10574_, new_n10573_, new_n10405_ );
and  ( new_n10575_, new_n10574_, new_n10400_ );
or   ( new_n10576_, new_n10575_, new_n10394_ );
and  ( new_n10577_, new_n10576_, new_n10389_ );
or   ( new_n10578_, new_n10577_, new_n10383_ );
and  ( new_n10579_, new_n10578_, new_n10378_ );
and  ( new_n10580_, new_n10374_, new_n6196_ );
and  ( new_n10581_, new_n10376_, new_n10289_ );
or   ( new_n10582_, new_n10581_, new_n10580_ );
or   ( new_n10583_, new_n10387_, new_n10384_ );
or   ( new_n10584_, new_n10398_, new_n10395_ );
or   ( new_n10585_, new_n10409_, new_n10406_ );
or   ( new_n10586_, new_n10420_, new_n10417_ );
or   ( new_n10587_, new_n10431_, new_n10428_ );
or   ( new_n10588_, new_n10442_, new_n10439_ );
or   ( new_n10589_, new_n10453_, new_n10450_ );
or   ( new_n10590_, new_n10464_, new_n10461_ );
or   ( new_n10591_, new_n10475_, new_n10472_ );
or   ( new_n10592_, new_n10486_, new_n10483_ );
or   ( new_n10593_, new_n10497_, new_n10494_ );
or   ( new_n10594_, new_n10508_, new_n10505_ );
or   ( new_n10595_, new_n10519_, new_n10516_ );
or   ( new_n10596_, new_n10530_, new_n10527_ );
or   ( new_n10597_, new_n10546_, new_n10543_ );
and  ( new_n10598_, new_n10312_, new_n10310_ );
or   ( new_n10599_, new_n10598_, new_n10258_ );
or   ( new_n10600_, new_n6195_, new_n3548_ );
or   ( new_n10601_, new_n10600_, new_n10599_ );
and  ( new_n10602_, new_n10546_, new_n10543_ );
or   ( new_n10603_, new_n10602_, new_n10537_ );
or   ( new_n10604_, new_n10603_, new_n10601_ );
and  ( new_n10605_, new_n10604_, new_n10597_ );
and  ( new_n10606_, new_n10530_, new_n10527_ );
or   ( new_n10607_, new_n10606_, new_n10526_ );
or   ( new_n10608_, new_n10607_, new_n10605_ );
and  ( new_n10609_, new_n10608_, new_n10596_ );
and  ( new_n10610_, new_n10519_, new_n10516_ );
or   ( new_n10611_, new_n10610_, new_n10515_ );
or   ( new_n10612_, new_n10611_, new_n10609_ );
and  ( new_n10613_, new_n10612_, new_n10595_ );
and  ( new_n10614_, new_n10508_, new_n10505_ );
or   ( new_n10615_, new_n10614_, new_n10504_ );
or   ( new_n10616_, new_n10615_, new_n10613_ );
and  ( new_n10617_, new_n10616_, new_n10594_ );
and  ( new_n10618_, new_n10497_, new_n10494_ );
or   ( new_n10619_, new_n10618_, new_n10493_ );
or   ( new_n10620_, new_n10619_, new_n10617_ );
and  ( new_n10621_, new_n10620_, new_n10593_ );
and  ( new_n10622_, new_n10486_, new_n10483_ );
or   ( new_n10623_, new_n10622_, new_n10482_ );
or   ( new_n10624_, new_n10623_, new_n10621_ );
and  ( new_n10625_, new_n10624_, new_n10592_ );
and  ( new_n10626_, new_n10475_, new_n10472_ );
or   ( new_n10627_, new_n10626_, new_n10471_ );
or   ( new_n10628_, new_n10627_, new_n10625_ );
and  ( new_n10629_, new_n10628_, new_n10591_ );
and  ( new_n10630_, new_n10464_, new_n10461_ );
or   ( new_n10631_, new_n10630_, new_n10460_ );
or   ( new_n10632_, new_n10631_, new_n10629_ );
and  ( new_n10633_, new_n10632_, new_n10590_ );
and  ( new_n10634_, new_n10453_, new_n10450_ );
or   ( new_n10635_, new_n10634_, new_n10449_ );
or   ( new_n10636_, new_n10635_, new_n10633_ );
and  ( new_n10637_, new_n10636_, new_n10589_ );
and  ( new_n10638_, new_n10442_, new_n10439_ );
or   ( new_n10639_, new_n10638_, new_n10438_ );
or   ( new_n10640_, new_n10639_, new_n10637_ );
and  ( new_n10641_, new_n10640_, new_n10588_ );
and  ( new_n10642_, new_n10431_, new_n10428_ );
or   ( new_n10643_, new_n10642_, new_n10427_ );
or   ( new_n10644_, new_n10643_, new_n10641_ );
and  ( new_n10645_, new_n10644_, new_n10587_ );
and  ( new_n10646_, new_n10420_, new_n10417_ );
or   ( new_n10647_, new_n10646_, new_n10416_ );
or   ( new_n10648_, new_n10647_, new_n10645_ );
and  ( new_n10649_, new_n10648_, new_n10586_ );
and  ( new_n10650_, new_n10409_, new_n10406_ );
or   ( new_n10651_, new_n10650_, new_n10405_ );
or   ( new_n10652_, new_n10651_, new_n10649_ );
and  ( new_n10653_, new_n10652_, new_n10585_ );
and  ( new_n10654_, new_n10398_, new_n10395_ );
or   ( new_n10655_, new_n10654_, new_n10394_ );
or   ( new_n10656_, new_n10655_, new_n10653_ );
and  ( new_n10657_, new_n10656_, new_n10584_ );
and  ( new_n10658_, new_n10387_, new_n10384_ );
or   ( new_n10659_, new_n10658_, new_n10383_ );
or   ( new_n10660_, new_n10659_, new_n10657_ );
and  ( new_n10661_, new_n10660_, new_n10583_ );
and  ( new_n10662_, new_n10661_, new_n10582_ );
or   ( new_n10663_, new_n10662_, new_n10579_ );
and  ( new_n10664_, \c[14] , \b[1]  );
or   ( new_n10665_, new_n969_, new_n815_ );
or   ( new_n10666_, new_n1127_, new_n847_ );
or   ( new_n10667_, new_n1010_, new_n1023_ );
or   ( new_n10668_, new_n1373_, new_n1296_ );
or   ( new_n10669_, new_n1468_, new_n1154_ );
or   ( new_n10670_, new_n1104_, new_n2206_ );
and  ( new_n10671_, \c[2] , \b[13]  );
xor  ( new_n10672_, new_n10671_, new_n10670_ );
xor  ( new_n10673_, new_n10672_, new_n10669_ );
xor  ( new_n10674_, new_n10673_, new_n10668_ );
xor  ( new_n10675_, new_n10674_, new_n10667_ );
xor  ( new_n10676_, new_n10675_, new_n10666_ );
xor  ( new_n10677_, new_n10676_, new_n10665_ );
xnor ( new_n10678_, new_n10677_, new_n10664_ );
not  ( new_n10679_, new_n10678_ );
and  ( new_n10680_, new_n6183_, new_n6109_ );
and  ( new_n10681_, new_n6184_, new_n6108_ );
nor  ( new_n10682_, new_n10681_, new_n10680_ );
and  ( new_n10683_, new_n6179_, new_n6117_ );
and  ( new_n10684_, new_n6180_, new_n6116_ );
or   ( new_n10685_, new_n10684_, new_n10683_ );
and  ( new_n10686_, new_n6175_, new_n6125_ );
and  ( new_n10687_, new_n6176_, new_n6124_ );
or   ( new_n10688_, new_n10687_, new_n10686_ );
and  ( new_n10689_, new_n6171_, new_n6133_ );
and  ( new_n10690_, new_n6172_, new_n6132_ );
or   ( new_n10691_, new_n10690_, new_n10689_ );
and  ( new_n10692_, new_n6167_, new_n6141_ );
and  ( new_n10693_, new_n6168_, new_n6140_ );
or   ( new_n10694_, new_n10693_, new_n10692_ );
and  ( new_n10695_, new_n6163_, new_n6149_ );
and  ( new_n10696_, new_n6164_, new_n6148_ );
or   ( new_n10697_, new_n10696_, new_n10695_ );
nand ( new_n10698_, new_n6159_, new_n1056_ );
nand ( new_n10699_, new_n6160_, new_n6158_ );
and  ( new_n10700_, new_n10699_, new_n10698_ );
xor  ( new_n10701_, new_n10700_, new_n10697_ );
xor  ( new_n10702_, new_n10701_, new_n10694_ );
xor  ( new_n10703_, new_n10702_, new_n10691_ );
xor  ( new_n10704_, new_n10703_, new_n10688_ );
xor  ( new_n10705_, new_n10704_, new_n10685_ );
xnor ( new_n10706_, new_n10705_, new_n10682_ );
nand ( new_n10707_, new_n6185_, new_n1627_ );
and  ( new_n10708_, new_n6181_, new_n6113_ );
and  ( new_n10709_, new_n6182_, new_n6112_ );
or   ( new_n10710_, new_n10709_, new_n10708_ );
and  ( new_n10711_, new_n6177_, new_n6121_ );
and  ( new_n10712_, new_n6178_, new_n6120_ );
or   ( new_n10713_, new_n10712_, new_n10711_ );
and  ( new_n10714_, new_n6173_, new_n6129_ );
and  ( new_n10715_, new_n6174_, new_n6128_ );
or   ( new_n10716_, new_n10715_, new_n10714_ );
and  ( new_n10717_, new_n6169_, new_n6137_ );
and  ( new_n10718_, new_n6170_, new_n6136_ );
or   ( new_n10719_, new_n10718_, new_n10717_ );
and  ( new_n10720_, new_n6165_, new_n6145_ );
and  ( new_n10721_, new_n6166_, new_n6144_ );
or   ( new_n10722_, new_n10721_, new_n10720_ );
nand ( new_n10723_, new_n6161_, new_n6154_ );
nand ( new_n10724_, new_n6162_, new_n6153_ );
and  ( new_n10725_, new_n10724_, new_n10723_ );
xor  ( new_n10726_, new_n10725_, new_n10722_ );
xor  ( new_n10727_, new_n10726_, new_n10719_ );
xor  ( new_n10728_, new_n10727_, new_n10716_ );
xor  ( new_n10729_, new_n10728_, new_n10713_ );
xor  ( new_n10730_, new_n10729_, new_n10710_ );
xor  ( new_n10731_, new_n10730_, new_n10707_ );
xor  ( new_n10732_, new_n10731_, new_n10706_ );
or   ( new_n10733_, new_n1653_, new_n804_ );
or   ( new_n10734_, new_n1066_, new_n865_ );
or   ( new_n10735_, new_n952_, new_n832_ );
or   ( new_n10736_, new_n1003_, new_n1019_ );
or   ( new_n10737_, new_n1000_, new_n1328_ );
or   ( new_n10738_, new_n943_, new_n1038_ );
or   ( new_n10739_, new_n978_, new_n1053_ );
xor  ( new_n10740_, new_n1620_, new_n10739_ );
xor  ( new_n10741_, new_n10740_, new_n10738_ );
xor  ( new_n10742_, new_n10741_, new_n10737_ );
xor  ( new_n10743_, new_n10742_, new_n10736_ );
xor  ( new_n10744_, new_n10743_, new_n10735_ );
xor  ( new_n10745_, new_n10744_, new_n10734_ );
xor  ( new_n10746_, new_n10745_, new_n10733_ );
xnor ( new_n10747_, new_n10746_, new_n10732_ );
not  ( new_n10748_, new_n10747_ );
and  ( new_n10749_, new_n10748_, new_n10679_ );
not  ( new_n10750_, new_n10749_ );
or   ( new_n10751_, new_n10748_, new_n10679_ );
and  ( new_n10752_, new_n10751_, new_n5052_ );
and  ( new_n10753_, new_n10752_, new_n10750_ );
not  ( new_n10754_, new_n10753_ );
and  ( new_n10755_, \d[14] , \a[1]  );
or   ( new_n10756_, new_n99_, new_n163_ );
or   ( new_n10757_, new_n326_, new_n176_ );
or   ( new_n10758_, new_n179_, new_n185_ );
or   ( new_n10759_, new_n563_, new_n137_ );
or   ( new_n10760_, new_n660_, new_n354_ );
or   ( new_n10761_, new_n90_, new_n2116_ );
and  ( new_n10762_, \d[2] , \a[13]  );
xor  ( new_n10763_, new_n10762_, new_n10761_ );
xor  ( new_n10764_, new_n10763_, new_n10760_ );
xor  ( new_n10765_, new_n10764_, new_n10759_ );
xor  ( new_n10766_, new_n10765_, new_n10758_ );
xor  ( new_n10767_, new_n10766_, new_n10757_ );
xor  ( new_n10768_, new_n10767_, new_n10756_ );
xnor ( new_n10769_, new_n10768_, new_n10755_ );
not  ( new_n10770_, new_n10769_ );
and  ( new_n10771_, new_n5644_, new_n5570_ );
and  ( new_n10772_, new_n5645_, new_n5569_ );
nor  ( new_n10773_, new_n10772_, new_n10771_ );
and  ( new_n10774_, new_n5640_, new_n5578_ );
and  ( new_n10775_, new_n5641_, new_n5577_ );
or   ( new_n10776_, new_n10775_, new_n10774_ );
and  ( new_n10777_, new_n5636_, new_n5586_ );
and  ( new_n10778_, new_n5637_, new_n5585_ );
or   ( new_n10779_, new_n10778_, new_n10777_ );
and  ( new_n10780_, new_n5632_, new_n5594_ );
and  ( new_n10781_, new_n5633_, new_n5593_ );
or   ( new_n10782_, new_n10781_, new_n10780_ );
and  ( new_n10783_, new_n5628_, new_n5602_ );
and  ( new_n10784_, new_n5629_, new_n5601_ );
or   ( new_n10785_, new_n10784_, new_n10783_ );
and  ( new_n10786_, new_n5624_, new_n5610_ );
and  ( new_n10787_, new_n5625_, new_n5609_ );
or   ( new_n10788_, new_n10787_, new_n10786_ );
nand ( new_n10789_, new_n5620_, new_n93_ );
nand ( new_n10790_, new_n5621_, new_n5619_ );
and  ( new_n10791_, new_n10790_, new_n10789_ );
xor  ( new_n10792_, new_n10791_, new_n10788_ );
xor  ( new_n10793_, new_n10792_, new_n10785_ );
xor  ( new_n10794_, new_n10793_, new_n10782_ );
xor  ( new_n10795_, new_n10794_, new_n10779_ );
xor  ( new_n10796_, new_n10795_, new_n10776_ );
xnor ( new_n10797_, new_n10796_, new_n10773_ );
nand ( new_n10798_, new_n5646_, new_n259_ );
and  ( new_n10799_, new_n5642_, new_n5574_ );
and  ( new_n10800_, new_n5643_, new_n5573_ );
or   ( new_n10801_, new_n10800_, new_n10799_ );
and  ( new_n10802_, new_n5638_, new_n5582_ );
and  ( new_n10803_, new_n5639_, new_n5581_ );
or   ( new_n10804_, new_n10803_, new_n10802_ );
and  ( new_n10805_, new_n5634_, new_n5590_ );
and  ( new_n10806_, new_n5635_, new_n5589_ );
or   ( new_n10807_, new_n10806_, new_n10805_ );
and  ( new_n10808_, new_n5630_, new_n5598_ );
and  ( new_n10809_, new_n5631_, new_n5597_ );
or   ( new_n10810_, new_n10809_, new_n10808_ );
and  ( new_n10811_, new_n5626_, new_n5606_ );
and  ( new_n10812_, new_n5627_, new_n5605_ );
or   ( new_n10813_, new_n10812_, new_n10811_ );
nand ( new_n10814_, new_n5622_, new_n5615_ );
nand ( new_n10815_, new_n5623_, new_n5614_ );
and  ( new_n10816_, new_n10815_, new_n10814_ );
xor  ( new_n10817_, new_n10816_, new_n10813_ );
xor  ( new_n10818_, new_n10817_, new_n10810_ );
xor  ( new_n10819_, new_n10818_, new_n10807_ );
xor  ( new_n10820_, new_n10819_, new_n10804_ );
xor  ( new_n10821_, new_n10820_, new_n10801_ );
xor  ( new_n10822_, new_n10821_, new_n10798_ );
xor  ( new_n10823_, new_n10822_, new_n10797_ );
or   ( new_n10824_, new_n255_, new_n98_ );
or   ( new_n10825_, new_n103_, new_n115_ );
or   ( new_n10826_, new_n75_, new_n231_ );
or   ( new_n10827_, new_n171_, new_n212_ );
or   ( new_n10828_, new_n128_, new_n133_ );
or   ( new_n10829_, new_n66_, new_n352_ );
or   ( new_n10830_, new_n150_, new_n85_ );
xor  ( new_n10831_, new_n200_, new_n10830_ );
xor  ( new_n10832_, new_n10831_, new_n10829_ );
xor  ( new_n10833_, new_n10832_, new_n10828_ );
xor  ( new_n10834_, new_n10833_, new_n10827_ );
xor  ( new_n10835_, new_n10834_, new_n10826_ );
xor  ( new_n10836_, new_n10835_, new_n10825_ );
xor  ( new_n10837_, new_n10836_, new_n10824_ );
xnor ( new_n10838_, new_n10837_, new_n10823_ );
not  ( new_n10839_, new_n10838_ );
and  ( new_n10840_, new_n10839_, new_n10770_ );
not  ( new_n10841_, new_n10840_ );
or   ( new_n10842_, new_n10839_, new_n10770_ );
and  ( new_n10843_, new_n10842_, new_n5098_ );
and  ( new_n10844_, new_n10843_, new_n10841_ );
not  ( new_n10845_, new_n10844_ );
not  ( new_n10846_, new_n2101_ );
and  ( new_n10847_, new_n5083_, new_n10846_ );
or   ( new_n10848_, \b[15] , \a[15]  );
and  ( new_n10849_, new_n10848_, new_n5102_ );
nor  ( new_n10850_, new_n10849_, new_n10847_ );
and  ( new_n10851_, new_n10850_, new_n10845_ );
and  ( new_n10852_, new_n10851_, new_n10754_ );
and  ( new_n10853_, \c[15] , \b[15]  );
and  ( new_n10854_, new_n10853_, new_n5064_ );
and  ( new_n10855_, new_n5110_, \a[15]  );
nor  ( new_n10856_, new_n10855_, new_n10854_ );
and  ( new_n10857_, new_n5056_, new_n2296_ );
and  ( new_n10858_, new_n5116_, \b[15]  );
nor  ( new_n10859_, new_n10858_, new_n10857_ );
and  ( new_n10860_, new_n10859_, new_n10856_ );
and  ( new_n10861_, new_n5072_, \d[15]  );
and  ( new_n10862_, new_n5092_, \c[15]  );
nor  ( new_n10863_, new_n10862_, new_n10861_ );
and  ( new_n10864_, new_n5076_, new_n1842_ );
and  ( new_n10865_, new_n5080_, new_n1778_ );
nor  ( new_n10866_, new_n10865_, new_n10864_ );
and  ( new_n10867_, new_n10866_, new_n10863_ );
and  ( new_n10868_, new_n10867_, new_n10860_ );
and  ( new_n10869_, new_n10868_, new_n10852_ );
and  ( new_n10870_, new_n10869_, new_n5120_ );
or   ( new_n10871_, new_n10870_, new_n2297_ );
or   ( new_n10872_, new_n10871_, new_n10663_ );
and  ( new_n10873_, new_n10871_, new_n10663_ );
and  ( new_n10874_, new_n10661_, new_n10378_ );
and  ( new_n10875_, new_n10582_, new_n10578_ );
or   ( new_n10876_, new_n10875_, new_n10874_ );
not  ( new_n10877_, new_n10869_ );
and  ( new_n10878_, new_n10877_, new_n3143_ );
and  ( new_n10879_, new_n10878_, new_n10876_ );
or   ( new_n10880_, new_n10879_, new_n10873_ );
or   ( new_n10881_, new_n10870_, new_n2288_ );
and  ( new_n10882_, new_n10659_, new_n10657_ );
or   ( new_n10883_, new_n10882_, new_n10577_ );
or   ( new_n10884_, new_n10883_, new_n10881_ );
and  ( new_n10885_, new_n10883_, new_n10881_ );
and  ( new_n10886_, new_n10657_, new_n10389_ );
and  ( new_n10887_, new_n10659_, new_n10576_ );
or   ( new_n10888_, new_n10887_, new_n10886_ );
and  ( new_n10889_, new_n10877_, new_n2420_ );
and  ( new_n10890_, new_n10889_, new_n10888_ );
or   ( new_n10891_, new_n10890_, new_n10885_ );
or   ( new_n10892_, new_n10870_, new_n2304_ );
and  ( new_n10893_, new_n10655_, new_n10653_ );
or   ( new_n10894_, new_n10893_, new_n10575_ );
or   ( new_n10895_, new_n10894_, new_n10892_ );
and  ( new_n10896_, new_n10894_, new_n10892_ );
and  ( new_n10897_, new_n10653_, new_n10400_ );
and  ( new_n10898_, new_n10655_, new_n10574_ );
or   ( new_n10899_, new_n10898_, new_n10897_ );
and  ( new_n10900_, new_n10877_, new_n3734_ );
and  ( new_n10901_, new_n10900_, new_n10899_ );
or   ( new_n10902_, new_n10901_, new_n10896_ );
or   ( new_n10903_, new_n10870_, new_n2440_ );
and  ( new_n10904_, new_n10651_, new_n10649_ );
or   ( new_n10905_, new_n10904_, new_n10573_ );
or   ( new_n10906_, new_n10905_, new_n10903_ );
and  ( new_n10907_, new_n10905_, new_n10903_ );
and  ( new_n10908_, new_n10649_, new_n10411_ );
and  ( new_n10909_, new_n10651_, new_n10572_ );
or   ( new_n10910_, new_n10909_, new_n10908_ );
and  ( new_n10911_, new_n10877_, new_n2441_ );
and  ( new_n10912_, new_n10911_, new_n10910_ );
or   ( new_n10913_, new_n10912_, new_n10907_ );
or   ( new_n10914_, new_n10870_, new_n2566_ );
and  ( new_n10915_, new_n10647_, new_n10645_ );
or   ( new_n10916_, new_n10915_, new_n10571_ );
or   ( new_n10917_, new_n10916_, new_n10914_ );
and  ( new_n10918_, new_n10916_, new_n10914_ );
and  ( new_n10919_, new_n10645_, new_n10422_ );
and  ( new_n10920_, new_n10647_, new_n10570_ );
or   ( new_n10921_, new_n10920_, new_n10919_ );
and  ( new_n10922_, new_n10877_, new_n6342_ );
and  ( new_n10923_, new_n10922_, new_n10921_ );
or   ( new_n10924_, new_n10923_, new_n10918_ );
or   ( new_n10925_, new_n10870_, new_n2705_ );
and  ( new_n10926_, new_n10643_, new_n10641_ );
or   ( new_n10927_, new_n10926_, new_n10569_ );
or   ( new_n10928_, new_n10927_, new_n10925_ );
and  ( new_n10929_, new_n10927_, new_n10925_ );
and  ( new_n10930_, new_n10641_, new_n10433_ );
and  ( new_n10931_, new_n10643_, new_n10568_ );
or   ( new_n10932_, new_n10931_, new_n10930_ );
and  ( new_n10933_, new_n10877_, new_n3693_ );
and  ( new_n10934_, new_n10933_, new_n10932_ );
or   ( new_n10935_, new_n10934_, new_n10929_ );
or   ( new_n10936_, new_n10870_, new_n2723_ );
and  ( new_n10937_, new_n10639_, new_n10637_ );
or   ( new_n10938_, new_n10937_, new_n10567_ );
or   ( new_n10939_, new_n10938_, new_n10936_ );
and  ( new_n10940_, new_n10938_, new_n10936_ );
and  ( new_n10941_, new_n10637_, new_n10444_ );
and  ( new_n10942_, new_n10639_, new_n10566_ );
or   ( new_n10943_, new_n10942_, new_n10941_ );
and  ( new_n10944_, new_n10877_, new_n4017_ );
and  ( new_n10945_, new_n10944_, new_n10943_ );
or   ( new_n10946_, new_n10945_, new_n10940_ );
or   ( new_n10947_, new_n10870_, new_n2760_ );
and  ( new_n10948_, new_n10635_, new_n10633_ );
or   ( new_n10949_, new_n10948_, new_n10565_ );
or   ( new_n10950_, new_n10949_, new_n10947_ );
and  ( new_n10951_, new_n10949_, new_n10947_ );
and  ( new_n10952_, new_n10633_, new_n10455_ );
and  ( new_n10953_, new_n10635_, new_n10564_ );
or   ( new_n10954_, new_n10953_, new_n10952_ );
and  ( new_n10955_, new_n10877_, new_n4085_ );
and  ( new_n10956_, new_n10955_, new_n10954_ );
or   ( new_n10957_, new_n10956_, new_n10951_ );
or   ( new_n10958_, new_n10870_, new_n2923_ );
and  ( new_n10959_, new_n10631_, new_n10629_ );
or   ( new_n10960_, new_n10959_, new_n10563_ );
or   ( new_n10961_, new_n10960_, new_n10958_ );
and  ( new_n10962_, new_n10960_, new_n10958_ );
and  ( new_n10963_, new_n10629_, new_n10466_ );
and  ( new_n10964_, new_n10631_, new_n10562_ );
or   ( new_n10965_, new_n10964_, new_n10963_ );
and  ( new_n10966_, new_n10877_, new_n2924_ );
and  ( new_n10967_, new_n10966_, new_n10965_ );
or   ( new_n10968_, new_n10967_, new_n10962_ );
or   ( new_n10969_, new_n10870_, new_n3066_ );
and  ( new_n10970_, new_n10627_, new_n10625_ );
or   ( new_n10971_, new_n10970_, new_n10561_ );
or   ( new_n10972_, new_n10971_, new_n10969_ );
and  ( new_n10973_, new_n10971_, new_n10969_ );
and  ( new_n10974_, new_n10625_, new_n10477_ );
and  ( new_n10975_, new_n10627_, new_n10560_ );
or   ( new_n10976_, new_n10975_, new_n10974_ );
and  ( new_n10977_, new_n10877_, new_n4177_ );
and  ( new_n10978_, new_n10977_, new_n10976_ );
or   ( new_n10979_, new_n10978_, new_n10973_ );
or   ( new_n10980_, new_n10870_, new_n3108_ );
and  ( new_n10981_, new_n10623_, new_n10621_ );
or   ( new_n10982_, new_n10981_, new_n10559_ );
or   ( new_n10983_, new_n10982_, new_n10980_ );
and  ( new_n10984_, new_n10982_, new_n10980_ );
and  ( new_n10985_, new_n10621_, new_n10488_ );
and  ( new_n10986_, new_n10623_, new_n10558_ );
or   ( new_n10987_, new_n10986_, new_n10985_ );
and  ( new_n10988_, new_n10877_, new_n3109_ );
and  ( new_n10989_, new_n10988_, new_n10987_ );
or   ( new_n10990_, new_n10989_, new_n10984_ );
or   ( new_n10991_, new_n10870_, new_n3244_ );
and  ( new_n10992_, new_n10619_, new_n10617_ );
or   ( new_n10993_, new_n10992_, new_n10557_ );
or   ( new_n10994_, new_n10993_, new_n10991_ );
and  ( new_n10995_, new_n10993_, new_n10991_ );
and  ( new_n10996_, new_n10617_, new_n10499_ );
and  ( new_n10997_, new_n10619_, new_n10556_ );
or   ( new_n10998_, new_n10997_, new_n10996_ );
and  ( new_n10999_, new_n10877_, new_n4257_ );
and  ( new_n11000_, new_n10999_, new_n10998_ );
or   ( new_n11001_, new_n11000_, new_n10995_ );
or   ( new_n11002_, new_n10870_, new_n3306_ );
and  ( new_n11003_, new_n10615_, new_n10613_ );
or   ( new_n11004_, new_n11003_, new_n10555_ );
or   ( new_n11005_, new_n11004_, new_n11002_ );
and  ( new_n11006_, new_n11004_, new_n11002_ );
and  ( new_n11007_, new_n10613_, new_n10510_ );
and  ( new_n11008_, new_n10615_, new_n10554_ );
or   ( new_n11009_, new_n11008_, new_n11007_ );
and  ( new_n11010_, new_n10877_, new_n4275_ );
and  ( new_n11011_, new_n11010_, new_n11009_ );
or   ( new_n11012_, new_n11011_, new_n11006_ );
or   ( new_n11013_, new_n10870_, new_n3406_ );
and  ( new_n11014_, new_n10611_, new_n10609_ );
or   ( new_n11015_, new_n11014_, new_n10553_ );
or   ( new_n11016_, new_n11015_, new_n11013_ );
and  ( new_n11017_, new_n11015_, new_n11013_ );
and  ( new_n11018_, new_n10609_, new_n10521_ );
and  ( new_n11019_, new_n10611_, new_n10552_ );
or   ( new_n11020_, new_n11019_, new_n11018_ );
and  ( new_n11021_, new_n10877_, new_n3407_ );
and  ( new_n11022_, new_n11021_, new_n11020_ );
or   ( new_n11023_, new_n11022_, new_n11017_ );
or   ( new_n11024_, new_n10870_, new_n3507_ );
and  ( new_n11025_, new_n10607_, new_n10605_ );
or   ( new_n11026_, new_n11025_, new_n10551_ );
or   ( new_n11027_, new_n11026_, new_n11024_ );
and  ( new_n11028_, new_n11026_, new_n11024_ );
and  ( new_n11029_, new_n10605_, new_n10532_ );
and  ( new_n11030_, new_n10607_, new_n10550_ );
or   ( new_n11031_, new_n11030_, new_n11029_ );
and  ( new_n11032_, new_n10877_, new_n4311_ );
and  ( new_n11033_, new_n11032_, new_n11031_ );
or   ( new_n11034_, new_n11033_, new_n11028_ );
and  ( new_n11035_, new_n10603_, new_n10601_ );
or   ( new_n11036_, new_n11035_, new_n10549_ );
or   ( new_n11037_, new_n10870_, new_n3548_ );
or   ( new_n11038_, new_n11037_, new_n11036_ );
or   ( new_n11039_, new_n11038_, new_n11034_ );
and  ( new_n11040_, new_n11039_, new_n11027_ );
or   ( new_n11041_, new_n11040_, new_n11023_ );
and  ( new_n11042_, new_n11041_, new_n11016_ );
or   ( new_n11043_, new_n11042_, new_n11012_ );
and  ( new_n11044_, new_n11043_, new_n11005_ );
or   ( new_n11045_, new_n11044_, new_n11001_ );
and  ( new_n11046_, new_n11045_, new_n10994_ );
or   ( new_n11047_, new_n11046_, new_n10990_ );
and  ( new_n11048_, new_n11047_, new_n10983_ );
or   ( new_n11049_, new_n11048_, new_n10979_ );
and  ( new_n11050_, new_n11049_, new_n10972_ );
or   ( new_n11051_, new_n11050_, new_n10968_ );
and  ( new_n11052_, new_n11051_, new_n10961_ );
or   ( new_n11053_, new_n11052_, new_n10957_ );
and  ( new_n11054_, new_n11053_, new_n10950_ );
or   ( new_n11055_, new_n11054_, new_n10946_ );
and  ( new_n11056_, new_n11055_, new_n10939_ );
or   ( new_n11057_, new_n11056_, new_n10935_ );
and  ( new_n11058_, new_n11057_, new_n10928_ );
or   ( new_n11059_, new_n11058_, new_n10924_ );
and  ( new_n11060_, new_n11059_, new_n10917_ );
or   ( new_n11061_, new_n11060_, new_n10913_ );
and  ( new_n11062_, new_n11061_, new_n10906_ );
or   ( new_n11063_, new_n11062_, new_n10902_ );
and  ( new_n11064_, new_n11063_, new_n10895_ );
or   ( new_n11065_, new_n11064_, new_n10891_ );
and  ( new_n11066_, new_n11065_, new_n10884_ );
or   ( new_n11067_, new_n11066_, new_n10880_ );
and  ( new_n11068_, new_n11067_, new_n10872_ );
or   ( new_n11069_, new_n10870_, new_n2906_ );
or   ( new_n11070_, new_n10374_, new_n6196_ );
or   ( new_n11071_, new_n10661_, new_n10582_ );
and  ( new_n11072_, new_n11071_, new_n11070_ );
and  ( new_n11073_, new_n11072_, new_n11069_ );
or   ( new_n11074_, new_n10581_, new_n10579_ );
and  ( new_n11075_, new_n10877_, new_n2407_ );
and  ( new_n11076_, new_n11075_, new_n11074_ );
or   ( new_n11077_, new_n11076_, new_n11073_ );
and  ( new_n11078_, new_n11077_, new_n11068_ );
and  ( new_n11079_, new_n11074_, new_n11069_ );
and  ( new_n11080_, new_n11075_, new_n11072_ );
or   ( new_n11081_, new_n11080_, new_n11079_ );
and  ( new_n11082_, new_n10876_, new_n10871_ );
and  ( new_n11083_, new_n10878_, new_n10663_ );
or   ( new_n11084_, new_n11083_, new_n11082_ );
and  ( new_n11085_, new_n10888_, new_n10881_ );
and  ( new_n11086_, new_n10889_, new_n10883_ );
or   ( new_n11087_, new_n11086_, new_n11085_ );
and  ( new_n11088_, new_n10899_, new_n10892_ );
and  ( new_n11089_, new_n10900_, new_n10894_ );
or   ( new_n11090_, new_n11089_, new_n11088_ );
and  ( new_n11091_, new_n10910_, new_n10903_ );
and  ( new_n11092_, new_n10911_, new_n10905_ );
or   ( new_n11093_, new_n11092_, new_n11091_ );
and  ( new_n11094_, new_n10921_, new_n10914_ );
and  ( new_n11095_, new_n10922_, new_n10916_ );
or   ( new_n11096_, new_n11095_, new_n11094_ );
and  ( new_n11097_, new_n10932_, new_n10925_ );
and  ( new_n11098_, new_n10933_, new_n10927_ );
or   ( new_n11099_, new_n11098_, new_n11097_ );
and  ( new_n11100_, new_n10943_, new_n10936_ );
and  ( new_n11101_, new_n10944_, new_n10938_ );
or   ( new_n11102_, new_n11101_, new_n11100_ );
and  ( new_n11103_, new_n10954_, new_n10947_ );
and  ( new_n11104_, new_n10955_, new_n10949_ );
or   ( new_n11105_, new_n11104_, new_n11103_ );
and  ( new_n11106_, new_n10965_, new_n10958_ );
and  ( new_n11107_, new_n10966_, new_n10960_ );
or   ( new_n11108_, new_n11107_, new_n11106_ );
and  ( new_n11109_, new_n10976_, new_n10969_ );
and  ( new_n11110_, new_n10977_, new_n10971_ );
or   ( new_n11111_, new_n11110_, new_n11109_ );
and  ( new_n11112_, new_n10987_, new_n10980_ );
and  ( new_n11113_, new_n10988_, new_n10982_ );
or   ( new_n11114_, new_n11113_, new_n11112_ );
and  ( new_n11115_, new_n10998_, new_n10991_ );
and  ( new_n11116_, new_n10999_, new_n10993_ );
or   ( new_n11117_, new_n11116_, new_n11115_ );
and  ( new_n11118_, new_n11009_, new_n11002_ );
and  ( new_n11119_, new_n11010_, new_n11004_ );
or   ( new_n11120_, new_n11119_, new_n11118_ );
and  ( new_n11121_, new_n11020_, new_n11013_ );
and  ( new_n11122_, new_n11021_, new_n11015_ );
or   ( new_n11123_, new_n11122_, new_n11121_ );
and  ( new_n11124_, new_n10601_, new_n10548_ );
and  ( new_n11125_, new_n10603_, new_n10542_ );
or   ( new_n11126_, new_n11125_, new_n11124_ );
and  ( new_n11127_, new_n10877_, new_n3547_ );
and  ( new_n11128_, new_n11127_, new_n11126_ );
and  ( new_n11129_, new_n11031_, new_n11024_ );
and  ( new_n11130_, new_n11032_, new_n11026_ );
or   ( new_n11131_, new_n11130_, new_n11129_ );
and  ( new_n11132_, new_n11131_, new_n11128_ );
or   ( new_n11133_, new_n11132_, new_n11033_ );
and  ( new_n11134_, new_n11133_, new_n11123_ );
or   ( new_n11135_, new_n11134_, new_n11022_ );
and  ( new_n11136_, new_n11135_, new_n11120_ );
or   ( new_n11137_, new_n11136_, new_n11011_ );
and  ( new_n11138_, new_n11137_, new_n11117_ );
or   ( new_n11139_, new_n11138_, new_n11000_ );
and  ( new_n11140_, new_n11139_, new_n11114_ );
or   ( new_n11141_, new_n11140_, new_n10989_ );
and  ( new_n11142_, new_n11141_, new_n11111_ );
or   ( new_n11143_, new_n11142_, new_n10978_ );
and  ( new_n11144_, new_n11143_, new_n11108_ );
or   ( new_n11145_, new_n11144_, new_n10967_ );
and  ( new_n11146_, new_n11145_, new_n11105_ );
or   ( new_n11147_, new_n11146_, new_n10956_ );
and  ( new_n11148_, new_n11147_, new_n11102_ );
or   ( new_n11149_, new_n11148_, new_n10945_ );
and  ( new_n11150_, new_n11149_, new_n11099_ );
or   ( new_n11151_, new_n11150_, new_n10934_ );
and  ( new_n11152_, new_n11151_, new_n11096_ );
or   ( new_n11153_, new_n11152_, new_n10923_ );
and  ( new_n11154_, new_n11153_, new_n11093_ );
or   ( new_n11155_, new_n11154_, new_n10912_ );
and  ( new_n11156_, new_n11155_, new_n11090_ );
or   ( new_n11157_, new_n11156_, new_n10901_ );
and  ( new_n11158_, new_n11157_, new_n11087_ );
or   ( new_n11159_, new_n11158_, new_n10890_ );
and  ( new_n11160_, new_n11159_, new_n11084_ );
or   ( new_n11161_, new_n11160_, new_n10879_ );
and  ( new_n11162_, new_n11161_, new_n11081_ );
or   ( new_n11163_, new_n11162_, new_n11078_ );
and  ( new_n11164_, new_n11163_, new_n4388_ );
and  ( new_n11165_, new_n11081_, new_n11068_ );
and  ( new_n11166_, new_n11161_, new_n11077_ );
nor  ( new_n11167_, new_n11166_, new_n11165_ );
nor  ( new_n11168_, new_n11167_, new_n4388_ );
and  ( new_n11169_, new_n11066_, new_n10880_ );
not  ( new_n11170_, new_n11160_ );
xor  ( new_n11171_, new_n2586_, new_n2585_ );
xnor ( new_n11172_, new_n11171_, new_n4385_ );
nand ( new_n11173_, new_n11172_, new_n11170_ );
or   ( new_n11174_, new_n11173_, new_n11169_ );
and  ( new_n11175_, new_n11159_, new_n10880_ );
and  ( new_n11176_, new_n11084_, new_n11066_ );
or   ( new_n11177_, new_n11176_, new_n11172_ );
or   ( new_n11178_, new_n11177_, new_n11175_ );
and  ( new_n11179_, new_n11178_, new_n11174_ );
and  ( new_n11180_, new_n11064_, new_n10891_ );
not  ( new_n11181_, new_n11158_ );
xor  ( new_n11182_, new_n2700_, new_n2589_ );
xnor ( new_n11183_, new_n11182_, new_n4383_ );
nand ( new_n11184_, new_n11183_, new_n11181_ );
or   ( new_n11185_, new_n11184_, new_n11180_ );
and  ( new_n11186_, new_n11157_, new_n10891_ );
and  ( new_n11187_, new_n11087_, new_n11064_ );
or   ( new_n11188_, new_n11187_, new_n11183_ );
or   ( new_n11189_, new_n11188_, new_n11186_ );
and  ( new_n11190_, new_n11189_, new_n11185_ );
and  ( new_n11191_, new_n11155_, new_n10902_ );
nand ( new_n11192_, new_n11090_, new_n11062_ );
xor  ( new_n11193_, new_n2752_, new_n2704_ );
xor  ( new_n11194_, new_n11193_, new_n4381_ );
nand ( new_n11195_, new_n11194_, new_n11192_ );
or   ( new_n11196_, new_n11195_, new_n11191_ );
and  ( new_n11197_, new_n11062_, new_n10902_ );
or   ( new_n11198_, new_n11194_, new_n11156_ );
or   ( new_n11199_, new_n11198_, new_n11197_ );
and  ( new_n11200_, new_n11199_, new_n11196_ );
and  ( new_n11201_, new_n11153_, new_n10913_ );
nand ( new_n11202_, new_n11093_, new_n11060_ );
xor  ( new_n11203_, new_n2880_, new_n2878_ );
xnor ( new_n11204_, new_n11203_, new_n4378_ );
nand ( new_n11205_, new_n11204_, new_n11202_ );
or   ( new_n11206_, new_n11205_, new_n11201_ );
and  ( new_n11207_, new_n11060_, new_n10913_ );
or   ( new_n11208_, new_n11204_, new_n11154_ );
or   ( new_n11209_, new_n11208_, new_n11207_ );
and  ( new_n11210_, new_n11209_, new_n11206_ );
and  ( new_n11211_, new_n11058_, new_n10924_ );
not  ( new_n11212_, new_n11152_ );
xor  ( new_n11213_, new_n2938_, new_n2937_ );
xor  ( new_n11214_, new_n11213_, new_n4376_ );
nand ( new_n11215_, new_n11214_, new_n11212_ );
or   ( new_n11216_, new_n11215_, new_n11211_ );
and  ( new_n11217_, new_n11151_, new_n10924_ );
and  ( new_n11218_, new_n11096_, new_n11058_ );
or   ( new_n11219_, new_n11218_, new_n11214_ );
or   ( new_n11220_, new_n11219_, new_n11217_ );
and  ( new_n11221_, new_n11220_, new_n11216_ );
and  ( new_n11222_, new_n11056_, new_n10935_ );
not  ( new_n11223_, new_n11150_ );
xor  ( new_n11224_, new_n3130_, new_n3129_ );
xnor ( new_n11225_, new_n11224_, new_n4373_ );
nand ( new_n11226_, new_n11225_, new_n11223_ );
or   ( new_n11227_, new_n11226_, new_n11222_ );
and  ( new_n11228_, new_n11149_, new_n10935_ );
and  ( new_n11229_, new_n11099_, new_n11056_ );
or   ( new_n11230_, new_n11229_, new_n11225_ );
or   ( new_n11231_, new_n11230_, new_n11228_ );
and  ( new_n11232_, new_n11231_, new_n11227_ );
and  ( new_n11233_, new_n11147_, new_n10946_ );
nand ( new_n11234_, new_n11102_, new_n11054_ );
xor  ( new_n11235_, new_n3296_, new_n3133_ );
xor  ( new_n11236_, new_n11235_, new_n4371_ );
nand ( new_n11237_, new_n11236_, new_n11234_ );
or   ( new_n11238_, new_n11237_, new_n11233_ );
and  ( new_n11239_, new_n11054_, new_n10946_ );
or   ( new_n11240_, new_n11236_, new_n11148_ );
or   ( new_n11241_, new_n11240_, new_n11239_ );
and  ( new_n11242_, new_n11241_, new_n11238_ );
and  ( new_n11243_, new_n11145_, new_n10957_ );
nand ( new_n11244_, new_n11105_, new_n11052_ );
xor  ( new_n11245_, new_n3354_, new_n3352_ );
xnor ( new_n11246_, new_n11245_, new_n4368_ );
nand ( new_n11247_, new_n11246_, new_n11244_ );
or   ( new_n11248_, new_n11247_, new_n11243_ );
and  ( new_n11249_, new_n11052_, new_n10957_ );
or   ( new_n11250_, new_n11246_, new_n11146_ );
or   ( new_n11251_, new_n11250_, new_n11249_ );
and  ( new_n11252_, new_n11251_, new_n11248_ );
and  ( new_n11253_, new_n11143_, new_n10968_ );
nand ( new_n11254_, new_n11108_, new_n11050_ );
xor  ( new_n11255_, new_n3445_, new_n3444_ );
xnor ( new_n11256_, new_n11255_, new_n4366_ );
nand ( new_n11257_, new_n11256_, new_n11254_ );
or   ( new_n11258_, new_n11257_, new_n11253_ );
and  ( new_n11259_, new_n11050_, new_n10968_ );
or   ( new_n11260_, new_n11256_, new_n11144_ );
or   ( new_n11261_, new_n11260_, new_n11259_ );
and  ( new_n11262_, new_n11261_, new_n11258_ );
and  ( new_n11263_, new_n11141_, new_n10979_ );
nand ( new_n11264_, new_n11111_, new_n11048_ );
xor  ( new_n11265_, new_n3610_, new_n3609_ );
xnor ( new_n11266_, new_n11265_, new_n4364_ );
nand ( new_n11267_, new_n11266_, new_n11264_ );
or   ( new_n11268_, new_n11267_, new_n11263_ );
and  ( new_n11269_, new_n11048_, new_n10979_ );
or   ( new_n11270_, new_n11266_, new_n11142_ );
or   ( new_n11271_, new_n11270_, new_n11269_ );
and  ( new_n11272_, new_n11271_, new_n11268_ );
and  ( new_n11273_, new_n11139_, new_n10990_ );
nand ( new_n11274_, new_n11114_, new_n11046_ );
xor  ( new_n11275_, new_n3642_, new_n3640_ );
xnor ( new_n11276_, new_n11275_, new_n4362_ );
nand ( new_n11277_, new_n11276_, new_n11274_ );
or   ( new_n11278_, new_n11277_, new_n11273_ );
and  ( new_n11279_, new_n11046_, new_n10990_ );
or   ( new_n11280_, new_n11276_, new_n11140_ );
or   ( new_n11281_, new_n11280_, new_n11279_ );
and  ( new_n11282_, new_n11281_, new_n11278_ );
and  ( new_n11283_, new_n11044_, new_n11001_ );
not  ( new_n11284_, new_n11138_ );
xor  ( new_n11285_, new_n3719_, new_n3645_ );
xor  ( new_n11286_, new_n11285_, new_n4360_ );
nand ( new_n11287_, new_n11286_, new_n11284_ );
or   ( new_n11288_, new_n11287_, new_n11283_ );
and  ( new_n11289_, new_n11137_, new_n11001_ );
and  ( new_n11290_, new_n11117_, new_n11044_ );
or   ( new_n11291_, new_n11290_, new_n11286_ );
or   ( new_n11292_, new_n11291_, new_n11289_ );
and  ( new_n11293_, new_n11292_, new_n11288_ );
and  ( new_n11294_, new_n11135_, new_n11012_ );
nand ( new_n11295_, new_n11120_, new_n11042_ );
xor  ( new_n11296_, new_n3801_, new_n3723_ );
xor  ( new_n11297_, new_n11296_, new_n4357_ );
nand ( new_n11298_, new_n11297_, new_n11295_ );
or   ( new_n11299_, new_n11298_, new_n11294_ );
and  ( new_n11300_, new_n11042_, new_n11012_ );
or   ( new_n11301_, new_n11297_, new_n11136_ );
or   ( new_n11302_, new_n11301_, new_n11300_ );
and  ( new_n11303_, new_n11302_, new_n11299_ );
and  ( new_n11304_, new_n11133_, new_n11023_ );
nand ( new_n11305_, new_n11123_, new_n11040_ );
xor  ( new_n11306_, new_n3860_, new_n3858_ );
xnor ( new_n11307_, new_n11306_, new_n4354_ );
nand ( new_n11308_, new_n11307_, new_n11305_ );
or   ( new_n11309_, new_n11308_, new_n11304_ );
and  ( new_n11310_, new_n11040_, new_n11023_ );
or   ( new_n11311_, new_n11307_, new_n11134_ );
or   ( new_n11312_, new_n11311_, new_n11310_ );
and  ( new_n11313_, new_n11312_, new_n11309_ );
and  ( new_n11314_, new_n11128_, new_n11034_ );
nand ( new_n11315_, new_n11131_, new_n11038_ );
xor  ( new_n11316_, new_n3914_, new_n3913_ );
xnor ( new_n11317_, new_n11316_, new_n4352_ );
nand ( new_n11318_, new_n11317_, new_n11315_ );
or   ( new_n11319_, new_n11318_, new_n11314_ );
and  ( new_n11320_, new_n11038_, new_n11034_ );
or   ( new_n11321_, new_n11317_, new_n11132_ );
or   ( new_n11322_, new_n11321_, new_n11320_ );
and  ( new_n11323_, new_n11322_, new_n11319_ );
xor  ( new_n11324_, new_n3972_, new_n3971_ );
xnor ( new_n11325_, new_n11324_, new_n4350_ );
and  ( new_n11326_, new_n11037_, new_n11036_ );
nor  ( new_n11327_, new_n11326_, new_n11128_ );
nor  ( new_n11328_, new_n11327_, new_n11325_ );
and  ( new_n11329_, new_n11126_, new_n11037_ );
and  ( new_n11330_, new_n11127_, new_n11036_ );
or   ( new_n11331_, new_n11330_, new_n11329_ );
and  ( new_n11332_, new_n11331_, new_n11325_ );
and  ( new_n11333_, new_n10600_, new_n10540_ );
nand ( new_n11334_, new_n10599_, new_n10541_ );
xor  ( new_n11335_, new_n4006_, new_n3975_ );
xor  ( new_n11336_, new_n11335_, new_n4347_ );
nand ( new_n11337_, new_n11336_, new_n11334_ );
or   ( new_n11338_, new_n11337_, new_n11333_ );
and  ( new_n11339_, new_n10600_, new_n10599_ );
or   ( new_n11340_, new_n11336_, new_n10542_ );
or   ( new_n11341_, new_n11340_, new_n11339_ );
and  ( new_n11342_, new_n11341_, new_n11338_ );
and  ( new_n11343_, new_n10309_, new_n10249_ );
and  ( new_n11344_, new_n10308_, new_n10250_ );
xor  ( new_n11345_, new_n4055_, new_n4053_ );
xnor ( new_n11346_, new_n11345_, new_n4345_ );
or   ( new_n11347_, new_n11346_, new_n11344_ );
or   ( new_n11348_, new_n11347_, new_n11343_ );
and  ( new_n11349_, new_n10309_, new_n10308_ );
not  ( new_n11350_, new_n10251_ );
nand ( new_n11351_, new_n11346_, new_n11350_ );
or   ( new_n11352_, new_n11351_, new_n11349_ );
and  ( new_n11353_, new_n11352_, new_n11348_ );
and  ( new_n11354_, new_n10020_, new_n9926_ );
and  ( new_n11355_, new_n10019_, new_n9927_ );
xor  ( new_n11356_, new_n4101_, new_n4099_ );
xnor ( new_n11357_, new_n11356_, new_n4343_ );
or   ( new_n11358_, new_n11357_, new_n11355_ );
or   ( new_n11359_, new_n11358_, new_n11354_ );
and  ( new_n11360_, new_n10020_, new_n10019_ );
not  ( new_n11361_, new_n9928_ );
nand ( new_n11362_, new_n11357_, new_n11361_ );
or   ( new_n11363_, new_n11362_, new_n11360_ );
and  ( new_n11364_, new_n11363_, new_n11359_ );
and  ( new_n11365_, new_n9697_, new_n9602_ );
and  ( new_n11366_, new_n9696_, new_n9603_ );
xor  ( new_n11367_, new_n4138_, new_n4105_ );
xnor ( new_n11368_, new_n11367_, new_n4341_ );
or   ( new_n11369_, new_n11368_, new_n11366_ );
or   ( new_n11370_, new_n11369_, new_n11365_ );
and  ( new_n11371_, new_n9697_, new_n9696_ );
not  ( new_n11372_, new_n9604_ );
nand ( new_n11373_, new_n11368_, new_n11372_ );
or   ( new_n11374_, new_n11373_, new_n11371_ );
and  ( new_n11375_, new_n11374_, new_n11370_ );
and  ( new_n11376_, new_n9373_, new_n9280_ );
and  ( new_n11377_, new_n9372_, new_n9281_ );
xor  ( new_n11378_, new_n4170_, new_n4168_ );
xnor ( new_n11379_, new_n11378_, new_n4339_ );
or   ( new_n11380_, new_n11379_, new_n11377_ );
or   ( new_n11381_, new_n11380_, new_n11376_ );
and  ( new_n11382_, new_n9373_, new_n9372_ );
not  ( new_n11383_, new_n9282_ );
nand ( new_n11384_, new_n11379_, new_n11383_ );
or   ( new_n11385_, new_n11384_, new_n11382_ );
and  ( new_n11386_, new_n11385_, new_n11381_ );
and  ( new_n11387_, new_n9051_, new_n8956_ );
and  ( new_n11388_, new_n9050_, new_n8957_ );
xor  ( new_n11389_, new_n4199_, new_n4198_ );
xnor ( new_n11390_, new_n11389_, new_n4337_ );
or   ( new_n11391_, new_n11390_, new_n11388_ );
or   ( new_n11392_, new_n11391_, new_n11387_ );
and  ( new_n11393_, new_n9051_, new_n9050_ );
not  ( new_n11394_, new_n8958_ );
nand ( new_n11395_, new_n11390_, new_n11394_ );
or   ( new_n11396_, new_n11395_, new_n11393_ );
and  ( new_n11397_, new_n11396_, new_n11392_ );
and  ( new_n11398_, new_n8727_, new_n8634_ );
and  ( new_n11399_, new_n8726_, new_n8635_ );
xor  ( new_n11400_, new_n4222_, new_n4221_ );
xnor ( new_n11401_, new_n11400_, new_n4335_ );
or   ( new_n11402_, new_n11401_, new_n11399_ );
or   ( new_n11403_, new_n11402_, new_n11398_ );
and  ( new_n11404_, new_n8727_, new_n8726_ );
not  ( new_n11405_, new_n8636_ );
nand ( new_n11406_, new_n11401_, new_n11405_ );
or   ( new_n11407_, new_n11406_, new_n11404_ );
and  ( new_n11408_, new_n11407_, new_n11403_ );
and  ( new_n11409_, new_n8405_, new_n8310_ );
and  ( new_n11410_, new_n8404_, new_n8311_ );
xor  ( new_n11411_, new_n4333_, new_n4246_ );
or   ( new_n11412_, new_n11411_, new_n11410_ );
or   ( new_n11413_, new_n11412_, new_n11409_ );
and  ( new_n11414_, new_n8405_, new_n8404_ );
not  ( new_n11415_, new_n8312_ );
nand ( new_n11416_, new_n11411_, new_n11415_ );
or   ( new_n11417_, new_n11416_, new_n11414_ );
and  ( new_n11418_, new_n11417_, new_n11413_ );
and  ( new_n11419_, new_n8081_, new_n7986_ );
and  ( new_n11420_, new_n8080_, new_n7987_ );
xor  ( new_n11421_, new_n4268_, new_n4266_ );
xnor ( new_n11422_, new_n11421_, new_n4331_ );
or   ( new_n11423_, new_n11422_, new_n11420_ );
or   ( new_n11424_, new_n11423_, new_n11419_ );
and  ( new_n11425_, new_n8081_, new_n8080_ );
not  ( new_n11426_, new_n7988_ );
nand ( new_n11427_, new_n11422_, new_n11426_ );
or   ( new_n11428_, new_n11427_, new_n11425_ );
and  ( new_n11429_, new_n11428_, new_n11424_ );
xor  ( new_n11430_, new_n4289_, new_n4287_ );
xnor ( new_n11431_, new_n11430_, new_n4329_ );
and  ( new_n11432_, new_n7757_, new_n7756_ );
or   ( new_n11433_, new_n11432_, new_n7664_ );
and  ( new_n11434_, new_n11433_, new_n11431_ );
and  ( new_n11435_, new_n7757_, new_n7662_ );
and  ( new_n11436_, new_n7756_, new_n7663_ );
nor  ( new_n11437_, new_n11436_, new_n11435_ );
nor  ( new_n11438_, new_n11437_, new_n11431_ );
and  ( new_n11439_, new_n7433_, new_n7337_ );
nand ( new_n11440_, new_n7432_, new_n7338_ );
xor  ( new_n11441_, new_n4301_, new_n4299_ );
xor  ( new_n11442_, new_n11441_, new_n4327_ );
nand ( new_n11443_, new_n11442_, new_n11440_ );
or   ( new_n11444_, new_n11443_, new_n11439_ );
and  ( new_n11445_, new_n7433_, new_n7432_ );
or   ( new_n11446_, new_n11442_, new_n7339_ );
or   ( new_n11447_, new_n11446_, new_n11445_ );
and  ( new_n11448_, new_n11447_, new_n11444_ );
and  ( new_n11449_, new_n7108_, new_n7013_ );
and  ( new_n11450_, new_n7107_, new_n7014_ );
xor  ( new_n11451_, new_n4325_, new_n4324_ );
or   ( new_n11452_, new_n11451_, new_n11450_ );
or   ( new_n11453_, new_n11452_, new_n11449_ );
and  ( new_n11454_, new_n7108_, new_n7107_ );
not  ( new_n11455_, new_n7015_ );
nand ( new_n11456_, new_n11451_, new_n11455_ );
or   ( new_n11457_, new_n11456_, new_n11454_ );
and  ( new_n11458_, new_n11457_, new_n11453_ );
and  ( new_n11459_, new_n6782_, new_n6684_ );
nand ( new_n11460_, new_n6781_, new_n6685_ );
xor  ( new_n11461_, new_n4308_, new_n4307_ );
xnor ( new_n11462_, new_n11461_, new_n4315_ );
nand ( new_n11463_, new_n11462_, new_n11460_ );
or   ( new_n11464_, new_n11463_, new_n11459_ );
and  ( new_n11465_, new_n6782_, new_n6781_ );
or   ( new_n11466_, new_n11462_, new_n6686_ );
or   ( new_n11467_, new_n11466_, new_n11465_ );
and  ( new_n11468_, new_n11467_, new_n11464_ );
or   ( new_n11469_, new_n6255_, new_n3488_ );
or   ( new_n11470_, new_n6258_, new_n3552_ );
or   ( new_n11471_, new_n3547_, new_n4311_ );
and  ( new_n11472_, new_n11471_, new_n11470_ );
and  ( new_n11473_, new_n11472_, new_n11469_ );
or   ( new_n11474_, new_n6258_, new_n3507_ );
and  ( new_n11475_, new_n11474_, new_n3230_ );
or   ( new_n11476_, new_n11475_, new_n5120_ );
nand ( new_n11477_, new_n6221_, new_n3230_ );
or   ( new_n11478_, new_n6221_, new_n3230_ );
and  ( new_n11479_, new_n11478_, new_n3547_ );
and  ( new_n11480_, new_n11479_, new_n11477_ );
and  ( new_n11481_, new_n11480_, new_n11476_ );
or   ( new_n11482_, new_n11481_, new_n11473_ );
or   ( new_n11483_, new_n11482_, new_n11468_ );
or   ( new_n11484_, new_n11483_, new_n11458_ );
or   ( new_n11485_, new_n11484_, new_n11448_ );
or   ( new_n11486_, new_n11485_, new_n11438_ );
or   ( new_n11487_, new_n11486_, new_n11434_ );
or   ( new_n11488_, new_n11487_, new_n11429_ );
or   ( new_n11489_, new_n11488_, new_n11418_ );
or   ( new_n11490_, new_n11489_, new_n11408_ );
or   ( new_n11491_, new_n11490_, new_n11397_ );
or   ( new_n11492_, new_n11491_, new_n11386_ );
or   ( new_n11493_, new_n11492_, new_n11375_ );
or   ( new_n11494_, new_n11493_, new_n11364_ );
or   ( new_n11495_, new_n11494_, new_n11353_ );
or   ( new_n11496_, new_n11495_, new_n11342_ );
or   ( new_n11497_, new_n11496_, new_n11332_ );
or   ( new_n11498_, new_n11497_, new_n11328_ );
or   ( new_n11499_, new_n11498_, new_n11323_ );
or   ( new_n11500_, new_n11499_, new_n11313_ );
or   ( new_n11501_, new_n11500_, new_n11303_ );
or   ( new_n11502_, new_n11501_, new_n11293_ );
or   ( new_n11503_, new_n11502_, new_n11282_ );
or   ( new_n11504_, new_n11503_, new_n11272_ );
or   ( new_n11505_, new_n11504_, new_n11262_ );
or   ( new_n11506_, new_n11505_, new_n11252_ );
or   ( new_n11507_, new_n11506_, new_n11242_ );
or   ( new_n11508_, new_n11507_, new_n11232_ );
or   ( new_n11509_, new_n11508_, new_n11221_ );
or   ( new_n11510_, new_n11509_, new_n11210_ );
or   ( new_n11511_, new_n11510_, new_n11200_ );
or   ( new_n11512_, new_n11511_, new_n11190_ );
or   ( new_n11513_, new_n11512_, new_n11179_ );
or   ( new_n11514_, new_n11513_, new_n11168_ );
or   ( eq, new_n11514_, new_n11164_ );
endmodule


