module miter ( 
    \A[2][9] , \A[2][8] , \A[2][7] , \A[2][6] , \A[2][5] , \A[2][4] ,
    \A[2][3] , \A[2][2] , \A[2][1] , \A[2][0] , \A[1][9] , \A[1][8] ,
    \A[1][7] , \A[1][6] , \A[1][5] , \A[1][4] , \A[1][3] , \A[1][2] ,
    \A[1][1] , \A[1][0] , \A[0][9] , \A[0][8] , \A[0][7] , \A[0][6] ,
    \A[0][5] , \A[0][4] , \A[0][3] , \A[0][2] , \A[0][1] , \A[0][0] ,
    \B[9] , \B[8] , \B[7] , \B[6] , \B[5] , \B[4] , \B[3] , \B[2] , \B[1] ,
    \B[0] , \I[7] , \I[6] , \I[5] , \I[4] , \I[3] , \I[2] , \I[1] , \I[0] ,
    eq  );
  input  \A[2][9] , \A[2][8] , \A[2][7] , \A[2][6] , \A[2][5] ,
    \A[2][4] , \A[2][3] , \A[2][2] , \A[2][1] , \A[2][0] , \A[1][9] ,
    \A[1][8] , \A[1][7] , \A[1][6] , \A[1][5] , \A[1][4] , \A[1][3] ,
    \A[1][2] , \A[1][1] , \A[1][0] , \A[0][9] , \A[0][8] , \A[0][7] ,
    \A[0][6] , \A[0][5] , \A[0][4] , \A[0][3] , \A[0][2] , \A[0][1] ,
    \A[0][0] , \B[9] , \B[8] , \B[7] , \B[6] , \B[5] , \B[4] , \B[3] ,
    \B[2] , \B[1] , \B[0] , \I[7] , \I[6] , \I[5] , \I[4] , \I[3] , \I[2] ,
    \I[1] , \I[0] ;
  output eq;
  wire new_n50_, new_n51_, new_n52_, new_n53_, new_n54_, new_n55_, new_n56_,
    new_n57_, new_n58_, new_n59_, new_n60_, new_n61_, new_n62_, new_n63_,
    new_n64_, new_n65_, new_n66_, new_n67_, new_n68_, new_n69_, new_n70_,
    new_n71_, new_n72_, new_n73_, new_n74_, new_n75_, new_n76_, new_n77_,
    new_n78_, new_n79_, new_n80_, new_n81_, new_n82_, new_n83_, new_n84_,
    new_n85_, new_n86_, new_n87_, new_n88_, new_n89_, new_n90_, new_n91_,
    new_n92_, new_n93_, new_n94_, new_n95_, new_n96_, new_n97_, new_n98_,
    new_n99_, new_n100_, new_n101_, new_n102_, new_n103_, new_n104_,
    new_n105_, new_n106_, new_n107_, new_n108_, new_n109_, new_n110_,
    new_n111_, new_n112_, new_n113_, new_n114_, new_n115_, new_n116_,
    new_n117_, new_n118_, new_n119_, new_n120_, new_n121_, new_n122_,
    new_n123_, new_n124_, new_n125_, new_n126_, new_n127_, new_n128_,
    new_n129_, new_n130_, new_n131_, new_n132_, new_n133_, new_n134_,
    new_n135_, new_n136_, new_n137_, new_n138_, new_n139_, new_n140_,
    new_n141_, new_n142_, new_n143_, new_n144_, new_n145_, new_n146_,
    new_n147_, new_n148_, new_n149_, new_n150_, new_n151_, new_n152_,
    new_n153_, new_n154_, new_n155_, new_n156_, new_n157_, new_n158_,
    new_n159_, new_n160_, new_n161_, new_n162_, new_n163_, new_n164_,
    new_n165_, new_n166_, new_n167_, new_n168_, new_n169_, new_n170_,
    new_n171_, new_n172_, new_n173_, new_n174_, new_n175_, new_n176_,
    new_n177_, new_n178_, new_n179_, new_n180_, new_n181_, new_n182_,
    new_n183_, new_n184_, new_n185_, new_n186_, new_n187_, new_n188_,
    new_n189_, new_n190_, new_n191_, new_n192_, new_n193_, new_n194_,
    new_n195_, new_n196_, new_n197_, new_n198_, new_n199_, new_n200_,
    new_n201_, new_n202_, new_n203_, new_n204_, new_n205_, new_n206_,
    new_n207_, new_n208_, new_n209_, new_n210_, new_n211_, new_n212_,
    new_n213_, new_n214_, new_n215_, new_n216_, new_n217_, new_n218_,
    new_n219_, new_n220_, new_n221_, new_n222_, new_n223_, new_n224_,
    new_n225_, new_n226_, new_n227_, new_n228_, new_n229_, new_n230_,
    new_n231_, new_n232_, new_n233_, new_n234_, new_n235_, new_n236_,
    new_n237_, new_n238_, new_n239_, new_n240_, new_n241_, new_n242_,
    new_n243_, new_n244_, new_n245_, new_n246_, new_n247_, new_n248_,
    new_n249_, new_n250_, new_n251_, new_n252_, new_n253_, new_n254_,
    new_n255_, new_n256_, new_n257_, new_n258_, new_n259_, new_n260_,
    new_n261_, new_n262_, new_n263_, new_n264_, new_n265_, new_n266_,
    new_n267_, new_n268_, new_n269_, new_n270_, new_n271_, new_n272_,
    new_n273_, new_n274_, new_n275_, new_n276_, new_n277_, new_n278_,
    new_n279_, new_n280_, new_n281_, new_n282_, new_n283_, new_n284_,
    new_n285_, new_n286_, new_n287_, new_n288_, new_n289_, new_n290_,
    new_n291_, new_n292_, new_n293_, new_n294_, new_n295_, new_n296_,
    new_n297_, new_n298_, new_n299_, new_n300_, new_n301_, new_n302_,
    new_n303_, new_n304_, new_n305_, new_n306_, new_n307_, new_n308_,
    new_n309_, new_n310_, new_n311_, new_n312_, new_n313_, new_n314_,
    new_n315_, new_n316_, new_n317_, new_n318_, new_n319_, new_n320_,
    new_n321_, new_n322_, new_n323_, new_n324_, new_n325_, new_n326_,
    new_n327_, new_n328_, new_n329_, new_n330_, new_n331_, new_n332_,
    new_n333_, new_n334_, new_n335_, new_n336_, new_n337_, new_n338_,
    new_n339_, new_n340_, new_n341_, new_n342_, new_n343_, new_n344_,
    new_n345_, new_n346_, new_n347_, new_n348_, new_n349_, new_n350_,
    new_n351_, new_n352_, new_n353_, new_n354_, new_n355_, new_n356_,
    new_n357_, new_n358_, new_n359_, new_n360_, new_n361_, new_n362_,
    new_n363_, new_n364_, new_n365_, new_n366_, new_n367_, new_n368_,
    new_n369_, new_n370_, new_n371_, new_n372_, new_n373_, new_n374_,
    new_n375_, new_n376_, new_n377_, new_n378_, new_n379_, new_n380_,
    new_n381_, new_n382_, new_n383_, new_n384_, new_n385_, new_n386_,
    new_n387_, new_n388_, new_n389_, new_n390_, new_n391_, new_n392_,
    new_n393_, new_n394_, new_n395_, new_n396_, new_n397_, new_n398_,
    new_n399_, new_n400_, new_n401_, new_n402_, new_n403_, new_n404_,
    new_n405_, new_n406_, new_n407_, new_n408_, new_n409_, new_n410_,
    new_n411_, new_n412_, new_n413_, new_n414_, new_n415_, new_n416_,
    new_n417_, new_n418_, new_n419_, new_n420_, new_n421_, new_n422_,
    new_n423_, new_n424_, new_n425_, new_n426_, new_n427_, new_n428_,
    new_n429_, new_n430_, new_n431_, new_n432_, new_n433_, new_n434_,
    new_n435_, new_n436_, new_n437_, new_n438_, new_n439_, new_n440_,
    new_n441_, new_n442_, new_n443_, new_n444_, new_n445_, new_n446_,
    new_n447_, new_n448_, new_n449_, new_n450_, new_n451_, new_n452_,
    new_n453_, new_n454_, new_n455_, new_n456_, new_n457_, new_n458_,
    new_n459_, new_n460_, new_n461_, new_n462_, new_n463_, new_n464_,
    new_n465_, new_n466_, new_n467_, new_n468_, new_n469_, new_n470_,
    new_n471_, new_n472_, new_n473_, new_n474_, new_n475_, new_n476_,
    new_n477_, new_n478_, new_n479_, new_n480_, new_n481_, new_n482_,
    new_n483_, new_n484_, new_n485_, new_n486_, new_n487_, new_n488_,
    new_n489_, new_n490_, new_n491_, new_n492_, new_n493_, new_n494_,
    new_n495_, new_n496_, new_n497_, new_n498_, new_n499_, new_n500_,
    new_n501_, new_n502_, new_n503_, new_n504_, new_n505_, new_n506_,
    new_n507_, new_n508_, new_n509_, new_n510_, new_n511_, new_n512_,
    new_n513_, new_n514_, new_n515_, new_n516_, new_n517_, new_n518_,
    new_n519_, new_n520_, new_n521_, new_n522_, new_n523_, new_n524_,
    new_n525_, new_n526_, new_n527_, new_n528_, new_n529_, new_n530_,
    new_n531_, new_n532_, new_n533_, new_n534_, new_n535_, new_n536_,
    new_n537_, new_n538_, new_n539_, new_n540_, new_n541_, new_n542_,
    new_n543_, new_n544_, new_n545_, new_n546_, new_n547_, new_n548_,
    new_n549_, new_n550_, new_n551_, new_n552_, new_n553_, new_n554_,
    new_n555_, new_n556_, new_n557_, new_n558_, new_n559_, new_n560_,
    new_n561_, new_n562_, new_n563_, new_n564_, new_n565_, new_n566_,
    new_n567_, new_n568_, new_n569_, new_n570_, new_n571_, new_n572_,
    new_n573_, new_n574_, new_n575_, new_n576_, new_n577_, new_n578_,
    new_n579_, new_n580_, new_n581_, new_n582_, new_n583_, new_n584_,
    new_n585_, new_n586_, new_n587_, new_n588_, new_n589_, new_n590_,
    new_n591_, new_n592_, new_n593_, new_n594_, new_n595_, new_n596_,
    new_n597_, new_n598_, new_n599_, new_n600_, new_n601_, new_n602_,
    new_n603_, new_n604_, new_n605_, new_n606_, new_n607_, new_n608_,
    new_n609_, new_n610_, new_n611_, new_n612_, new_n613_, new_n614_,
    new_n615_, new_n616_, new_n617_, new_n618_, new_n619_, new_n620_,
    new_n621_, new_n622_, new_n623_, new_n624_, new_n625_, new_n626_,
    new_n627_, new_n628_, new_n629_, new_n630_, new_n631_, new_n632_,
    new_n633_, new_n634_, new_n635_, new_n636_, new_n637_, new_n638_,
    new_n639_, new_n640_, new_n641_, new_n642_, new_n643_, new_n644_,
    new_n645_, new_n646_, new_n647_, new_n648_, new_n649_, new_n650_,
    new_n651_, new_n652_, new_n653_, new_n654_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n749_, new_n750_, new_n751_, new_n752_,
    new_n753_, new_n754_, new_n755_, new_n756_, new_n757_, new_n758_,
    new_n759_, new_n760_, new_n761_, new_n762_, new_n763_, new_n764_,
    new_n765_, new_n766_, new_n767_, new_n768_, new_n769_, new_n770_,
    new_n771_, new_n772_, new_n773_, new_n774_, new_n775_, new_n776_,
    new_n777_, new_n778_, new_n779_, new_n780_, new_n781_, new_n782_,
    new_n783_, new_n784_, new_n785_, new_n786_, new_n787_, new_n788_,
    new_n789_, new_n790_, new_n791_, new_n792_, new_n793_, new_n794_,
    new_n795_, new_n796_, new_n797_, new_n798_, new_n799_, new_n800_,
    new_n801_, new_n802_, new_n803_, new_n804_, new_n805_, new_n806_,
    new_n807_, new_n808_, new_n809_, new_n810_, new_n811_, new_n812_,
    new_n813_, new_n814_, new_n815_, new_n816_, new_n817_, new_n818_,
    new_n819_, new_n820_, new_n821_, new_n822_, new_n823_, new_n824_,
    new_n825_, new_n826_, new_n827_, new_n828_, new_n829_, new_n830_,
    new_n831_, new_n832_, new_n833_, new_n834_, new_n835_, new_n836_,
    new_n837_, new_n838_, new_n839_, new_n840_, new_n841_, new_n842_,
    new_n843_, new_n844_, new_n845_, new_n846_, new_n847_, new_n848_,
    new_n849_, new_n850_, new_n851_, new_n852_, new_n853_, new_n854_,
    new_n855_, new_n856_, new_n857_, new_n858_, new_n859_, new_n860_,
    new_n861_, new_n862_, new_n863_, new_n864_, new_n865_, new_n866_,
    new_n867_, new_n868_, new_n869_, new_n870_, new_n871_, new_n872_,
    new_n873_, new_n874_, new_n875_, new_n876_, new_n877_, new_n878_,
    new_n879_, new_n880_, new_n881_, new_n882_, new_n883_, new_n884_,
    new_n885_, new_n886_, new_n887_, new_n888_, new_n889_, new_n890_,
    new_n891_, new_n892_, new_n893_, new_n894_, new_n895_, new_n896_,
    new_n897_, new_n898_, new_n899_, new_n900_, new_n901_, new_n902_,
    new_n903_, new_n904_, new_n905_, new_n906_, new_n907_, new_n908_,
    new_n909_, new_n910_, new_n911_, new_n912_, new_n913_, new_n914_,
    new_n915_, new_n916_, new_n917_, new_n918_, new_n919_, new_n920_,
    new_n921_, new_n922_, new_n923_, new_n924_, new_n925_, new_n926_,
    new_n927_, new_n928_, new_n929_, new_n930_, new_n931_, new_n932_,
    new_n933_, new_n934_, new_n935_, new_n936_, new_n937_, new_n938_,
    new_n939_, new_n940_, new_n941_, new_n942_, new_n943_, new_n944_,
    new_n945_, new_n946_, new_n947_, new_n948_, new_n949_, new_n950_,
    new_n951_, new_n952_, new_n953_, new_n954_, new_n955_, new_n956_,
    new_n957_, new_n958_, new_n959_, new_n960_, new_n961_, new_n962_,
    new_n963_, new_n964_, new_n965_, new_n966_, new_n967_, new_n968_,
    new_n969_, new_n970_, new_n971_, new_n972_, new_n973_, new_n974_,
    new_n975_, new_n976_, new_n977_, new_n978_, new_n979_, new_n980_,
    new_n981_, new_n982_, new_n983_, new_n984_, new_n985_, new_n986_,
    new_n987_, new_n988_, new_n989_, new_n990_, new_n991_, new_n992_,
    new_n993_, new_n994_, new_n995_, new_n996_, new_n997_, new_n998_,
    new_n999_, new_n1000_, new_n1001_, new_n1002_, new_n1003_, new_n1004_,
    new_n1005_, new_n1006_, new_n1007_, new_n1008_, new_n1009_, new_n1010_,
    new_n1011_, new_n1012_, new_n1013_, new_n1014_, new_n1015_, new_n1016_,
    new_n1017_, new_n1018_, new_n1019_, new_n1020_, new_n1021_, new_n1022_,
    new_n1023_, new_n1024_, new_n1025_, new_n1026_, new_n1027_, new_n1028_,
    new_n1029_, new_n1030_, new_n1031_, new_n1032_, new_n1033_, new_n1034_,
    new_n1035_, new_n1036_, new_n1037_, new_n1038_, new_n1039_, new_n1040_,
    new_n1041_, new_n1042_, new_n1043_, new_n1044_, new_n1045_, new_n1046_,
    new_n1047_, new_n1048_, new_n1049_, new_n1050_, new_n1051_, new_n1052_,
    new_n1053_, new_n1054_, new_n1055_, new_n1056_, new_n1057_, new_n1058_,
    new_n1059_, new_n1060_, new_n1061_, new_n1062_, new_n1063_, new_n1064_,
    new_n1065_, new_n1066_, new_n1067_, new_n1068_, new_n1069_, new_n1070_,
    new_n1071_, new_n1072_, new_n1073_, new_n1074_, new_n1075_, new_n1076_,
    new_n1077_, new_n1078_, new_n1079_, new_n1080_, new_n1081_, new_n1082_,
    new_n1083_, new_n1084_, new_n1085_, new_n1086_, new_n1087_, new_n1088_,
    new_n1089_, new_n1090_, new_n1091_, new_n1092_, new_n1093_, new_n1094_,
    new_n1095_, new_n1096_, new_n1097_, new_n1098_, new_n1099_, new_n1100_,
    new_n1101_, new_n1102_, new_n1103_, new_n1104_, new_n1105_, new_n1106_,
    new_n1107_, new_n1108_, new_n1109_, new_n1110_, new_n1111_, new_n1112_,
    new_n1113_, new_n1114_, new_n1115_, new_n1116_, new_n1117_, new_n1118_,
    new_n1119_, new_n1120_, new_n1121_, new_n1122_, new_n1123_, new_n1124_,
    new_n1125_, new_n1126_, new_n1127_, new_n1128_, new_n1129_, new_n1130_,
    new_n1131_, new_n1132_, new_n1133_, new_n1134_, new_n1135_, new_n1136_,
    new_n1137_, new_n1138_, new_n1139_, new_n1140_, new_n1141_, new_n1142_,
    new_n1143_, new_n1144_, new_n1145_, new_n1146_, new_n1147_, new_n1148_,
    new_n1149_, new_n1150_, new_n1151_, new_n1152_, new_n1153_, new_n1154_,
    new_n1155_, new_n1156_, new_n1157_, new_n1158_, new_n1159_, new_n1160_,
    new_n1161_, new_n1162_, new_n1163_, new_n1164_, new_n1165_, new_n1166_,
    new_n1167_, new_n1168_, new_n1169_, new_n1170_, new_n1171_, new_n1172_,
    new_n1173_, new_n1174_, new_n1175_, new_n1176_, new_n1177_, new_n1178_,
    new_n1179_, new_n1180_, new_n1181_, new_n1182_, new_n1183_, new_n1184_,
    new_n1185_, new_n1186_, new_n1187_, new_n1188_, new_n1189_, new_n1190_,
    new_n1191_, new_n1192_, new_n1193_, new_n1194_, new_n1195_, new_n1196_,
    new_n1197_, new_n1198_, new_n1199_, new_n1200_, new_n1201_, new_n1202_,
    new_n1203_, new_n1204_, new_n1205_, new_n1206_, new_n1207_, new_n1208_,
    new_n1209_, new_n1210_, new_n1211_, new_n1212_, new_n1213_, new_n1214_,
    new_n1215_, new_n1216_, new_n1217_, new_n1218_, new_n1219_, new_n1220_,
    new_n1221_, new_n1222_, new_n1223_, new_n1224_, new_n1225_, new_n1226_,
    new_n1227_, new_n1228_, new_n1229_, new_n1230_, new_n1231_, new_n1232_,
    new_n1233_, new_n1234_, new_n1235_, new_n1236_, new_n1237_, new_n1238_,
    new_n1239_, new_n1240_, new_n1241_, new_n1242_, new_n1243_, new_n1244_,
    new_n1245_, new_n1246_, new_n1247_, new_n1248_, new_n1249_, new_n1250_,
    new_n1251_, new_n1252_, new_n1253_, new_n1254_, new_n1255_, new_n1256_,
    new_n1257_, new_n1258_, new_n1259_, new_n1260_, new_n1261_, new_n1262_,
    new_n1263_, new_n1264_, new_n1265_, new_n1266_, new_n1267_, new_n1268_,
    new_n1269_, new_n1270_, new_n1271_, new_n1272_, new_n1273_, new_n1274_,
    new_n1275_, new_n1276_, new_n1277_, new_n1278_, new_n1279_, new_n1280_,
    new_n1281_, new_n1282_, new_n1283_, new_n1284_, new_n1285_, new_n1286_,
    new_n1287_, new_n1288_, new_n1289_, new_n1290_, new_n1291_, new_n1292_,
    new_n1293_, new_n1294_, new_n1295_, new_n1296_, new_n1297_, new_n1298_,
    new_n1299_, new_n1300_, new_n1301_, new_n1302_, new_n1303_, new_n1304_,
    new_n1305_, new_n1306_, new_n1307_, new_n1308_, new_n1309_, new_n1310_,
    new_n1311_, new_n1312_, new_n1313_, new_n1314_, new_n1315_, new_n1316_,
    new_n1317_, new_n1318_, new_n1319_, new_n1320_, new_n1321_, new_n1322_,
    new_n1323_, new_n1324_, new_n1325_, new_n1326_, new_n1327_, new_n1328_,
    new_n1329_, new_n1330_, new_n1331_, new_n1332_, new_n1333_, new_n1334_,
    new_n1335_, new_n1336_, new_n1337_, new_n1338_, new_n1339_, new_n1340_,
    new_n1341_, new_n1342_, new_n1343_, new_n1344_, new_n1345_, new_n1346_,
    new_n1347_, new_n1348_, new_n1349_, new_n1350_, new_n1351_, new_n1352_,
    new_n1353_, new_n1354_, new_n1355_, new_n1356_, new_n1357_, new_n1358_,
    new_n1359_, new_n1360_, new_n1361_, new_n1362_, new_n1363_, new_n1364_,
    new_n1365_, new_n1366_, new_n1367_, new_n1368_, new_n1369_, new_n1370_,
    new_n1371_, new_n1372_, new_n1373_, new_n1374_, new_n1375_, new_n1376_,
    new_n1377_, new_n1378_, new_n1379_, new_n1380_, new_n1381_, new_n1382_,
    new_n1383_, new_n1384_, new_n1385_, new_n1386_, new_n1387_, new_n1388_,
    new_n1389_, new_n1390_, new_n1391_, new_n1392_, new_n1393_, new_n1394_,
    new_n1395_, new_n1396_, new_n1397_, new_n1398_, new_n1399_, new_n1400_,
    new_n1401_, new_n1402_, new_n1403_, new_n1404_, new_n1405_, new_n1406_,
    new_n1407_, new_n1408_, new_n1409_, new_n1410_, new_n1411_, new_n1412_,
    new_n1413_, new_n1414_, new_n1415_, new_n1416_, new_n1417_, new_n1418_,
    new_n1419_, new_n1420_, new_n1421_, new_n1422_, new_n1423_, new_n1424_,
    new_n1425_, new_n1426_, new_n1427_, new_n1428_, new_n1429_, new_n1430_,
    new_n1431_, new_n1432_, new_n1433_, new_n1434_, new_n1435_, new_n1436_,
    new_n1437_, new_n1438_, new_n1439_, new_n1440_, new_n1441_, new_n1442_,
    new_n1443_, new_n1444_, new_n1445_, new_n1446_, new_n1447_, new_n1448_,
    new_n1449_, new_n1450_, new_n1451_, new_n1452_, new_n1453_, new_n1454_,
    new_n1455_, new_n1456_, new_n1457_, new_n1458_, new_n1459_, new_n1460_,
    new_n1461_, new_n1462_, new_n1463_, new_n1464_, new_n1465_, new_n1466_,
    new_n1467_, new_n1468_, new_n1469_, new_n1470_, new_n1471_, new_n1472_,
    new_n1473_, new_n1474_, new_n1475_, new_n1476_, new_n1477_, new_n1478_,
    new_n1479_, new_n1480_, new_n1481_, new_n1482_, new_n1483_, new_n1484_,
    new_n1485_, new_n1486_, new_n1487_, new_n1488_, new_n1489_, new_n1490_,
    new_n1491_, new_n1492_, new_n1493_, new_n1494_, new_n1495_, new_n1496_,
    new_n1497_, new_n1498_, new_n1499_, new_n1500_, new_n1501_, new_n1502_,
    new_n1503_, new_n1504_, new_n1505_, new_n1506_, new_n1507_, new_n1508_,
    new_n1509_, new_n1510_, new_n1511_, new_n1512_, new_n1513_, new_n1514_,
    new_n1515_, new_n1516_, new_n1517_, new_n1518_, new_n1519_, new_n1520_,
    new_n1521_, new_n1522_, new_n1523_, new_n1524_, new_n1525_, new_n1526_,
    new_n1527_, new_n1528_, new_n1529_, new_n1530_, new_n1531_, new_n1532_,
    new_n1533_, new_n1534_, new_n1535_, new_n1536_, new_n1537_, new_n1538_,
    new_n1539_, new_n1540_, new_n1541_, new_n1542_, new_n1543_, new_n1544_,
    new_n1545_, new_n1546_, new_n1547_, new_n1548_, new_n1549_, new_n1550_,
    new_n1551_, new_n1552_, new_n1553_, new_n1554_, new_n1555_, new_n1556_,
    new_n1557_, new_n1558_, new_n1559_, new_n1560_, new_n1561_, new_n1562_,
    new_n1563_, new_n1564_, new_n1565_, new_n1566_, new_n1567_, new_n1568_,
    new_n1569_, new_n1570_, new_n1571_, new_n1572_, new_n1573_, new_n1574_,
    new_n1575_, new_n1576_, new_n1577_, new_n1578_, new_n1579_, new_n1580_,
    new_n1581_, new_n1582_, new_n1583_, new_n1584_, new_n1585_, new_n1586_,
    new_n1587_, new_n1588_, new_n1589_, new_n1590_, new_n1591_, new_n1592_,
    new_n1593_, new_n1594_, new_n1595_, new_n1596_, new_n1597_, new_n1598_,
    new_n1599_, new_n1600_, new_n1601_, new_n1602_, new_n1603_, new_n1604_,
    new_n1605_, new_n1606_, new_n1607_, new_n1608_, new_n1609_, new_n1610_,
    new_n1611_, new_n1612_, new_n1613_, new_n1614_, new_n1615_, new_n1616_,
    new_n1617_, new_n1618_, new_n1619_, new_n1620_, new_n1621_, new_n1622_,
    new_n1623_, new_n1624_, new_n1625_, new_n1626_, new_n1627_, new_n1628_,
    new_n1629_, new_n1630_, new_n1631_, new_n1632_, new_n1633_, new_n1634_,
    new_n1635_, new_n1636_, new_n1637_, new_n1638_, new_n1639_, new_n1640_,
    new_n1641_, new_n1642_, new_n1643_, new_n1644_, new_n1645_, new_n1646_,
    new_n1647_, new_n1648_, new_n1649_, new_n1650_, new_n1651_, new_n1652_,
    new_n1653_, new_n1654_, new_n1655_, new_n1656_, new_n1657_, new_n1658_,
    new_n1659_, new_n1660_, new_n1661_, new_n1662_, new_n1663_, new_n1664_,
    new_n1665_, new_n1666_, new_n1667_, new_n1668_, new_n1669_, new_n1670_,
    new_n1671_, new_n1672_, new_n1673_, new_n1674_, new_n1675_, new_n1676_,
    new_n1677_, new_n1678_, new_n1679_, new_n1680_, new_n1681_, new_n1682_,
    new_n1683_, new_n1684_, new_n1685_, new_n1686_, new_n1687_, new_n1688_,
    new_n1689_, new_n1690_, new_n1691_, new_n1692_, new_n1693_, new_n1694_,
    new_n1695_, new_n1696_, new_n1697_, new_n1698_, new_n1699_, new_n1700_,
    new_n1701_, new_n1702_, new_n1703_, new_n1704_, new_n1705_, new_n1706_,
    new_n1707_, new_n1708_, new_n1709_, new_n1710_, new_n1711_, new_n1712_,
    new_n1713_, new_n1714_, new_n1715_, new_n1716_, new_n1717_, new_n1718_,
    new_n1719_, new_n1720_, new_n1721_, new_n1722_, new_n1723_, new_n1724_,
    new_n1725_, new_n1726_, new_n1727_, new_n1728_, new_n1729_, new_n1730_,
    new_n1731_, new_n1732_, new_n1733_, new_n1734_, new_n1735_, new_n1736_,
    new_n1737_, new_n1738_, new_n1739_, new_n1740_, new_n1741_, new_n1742_,
    new_n1743_, new_n1744_, new_n1745_, new_n1746_, new_n1747_, new_n1748_,
    new_n1749_, new_n1750_, new_n1751_, new_n1752_, new_n1753_, new_n1754_,
    new_n1755_, new_n1756_, new_n1757_, new_n1758_, new_n1759_, new_n1760_,
    new_n1761_, new_n1762_, new_n1763_, new_n1764_, new_n1765_, new_n1766_,
    new_n1767_, new_n1768_, new_n1769_, new_n1770_, new_n1771_, new_n1772_,
    new_n1773_, new_n1774_, new_n1775_, new_n1776_, new_n1777_, new_n1778_,
    new_n1779_, new_n1780_, new_n1781_, new_n1782_, new_n1783_, new_n1784_,
    new_n1785_, new_n1786_, new_n1787_, new_n1788_, new_n1789_, new_n1790_,
    new_n1791_, new_n1792_, new_n1793_, new_n1794_, new_n1795_, new_n1796_,
    new_n1797_, new_n1798_, new_n1799_, new_n1800_, new_n1801_, new_n1802_,
    new_n1803_, new_n1804_, new_n1805_, new_n1806_, new_n1807_, new_n1808_,
    new_n1809_, new_n1810_, new_n1811_, new_n1812_, new_n1813_, new_n1814_,
    new_n1815_, new_n1816_, new_n1817_, new_n1818_, new_n1819_, new_n1820_,
    new_n1821_, new_n1822_, new_n1823_, new_n1824_, new_n1825_, new_n1826_,
    new_n1827_, new_n1828_, new_n1829_, new_n1830_, new_n1831_, new_n1832_,
    new_n1833_, new_n1834_, new_n1835_, new_n1836_, new_n1837_, new_n1838_,
    new_n1839_, new_n1840_, new_n1841_, new_n1842_, new_n1843_, new_n1844_,
    new_n1845_, new_n1846_, new_n1847_, new_n1848_, new_n1849_, new_n1850_,
    new_n1851_, new_n1852_, new_n1853_, new_n1854_, new_n1855_, new_n1856_,
    new_n1857_, new_n1858_, new_n1859_, new_n1860_, new_n1861_, new_n1862_,
    new_n1863_, new_n1864_, new_n1865_, new_n1866_, new_n1867_, new_n1868_,
    new_n1869_, new_n1870_, new_n1871_, new_n1872_, new_n1873_, new_n1874_,
    new_n1875_, new_n1876_, new_n1877_, new_n1878_, new_n1879_, new_n1880_,
    new_n1881_, new_n1882_, new_n1883_, new_n1884_, new_n1885_, new_n1886_,
    new_n1887_, new_n1888_, new_n1889_, new_n1890_, new_n1891_, new_n1892_,
    new_n1893_, new_n1894_, new_n1895_, new_n1896_, new_n1897_, new_n1898_,
    new_n1899_, new_n1900_, new_n1901_, new_n1902_, new_n1903_, new_n1904_,
    new_n1905_, new_n1906_, new_n1907_, new_n1908_, new_n1909_, new_n1910_,
    new_n1911_, new_n1912_, new_n1913_, new_n1914_, new_n1915_, new_n1916_,
    new_n1917_, new_n1918_, new_n1919_, new_n1920_, new_n1921_, new_n1922_,
    new_n1923_, new_n1924_, new_n1925_, new_n1926_, new_n1927_, new_n1928_,
    new_n1929_, new_n1930_, new_n1931_, new_n1932_, new_n1933_, new_n1934_,
    new_n1935_, new_n1936_, new_n1937_, new_n1938_, new_n1939_, new_n1940_,
    new_n1941_, new_n1942_, new_n1943_, new_n1944_, new_n1945_, new_n1946_,
    new_n1947_, new_n1948_, new_n1949_, new_n1950_, new_n1951_, new_n1952_,
    new_n1953_, new_n1954_, new_n1955_, new_n1956_, new_n1957_, new_n1958_,
    new_n1959_, new_n1960_, new_n1961_, new_n1962_, new_n1963_, new_n1964_,
    new_n1965_, new_n1966_, new_n1967_, new_n1968_, new_n1969_, new_n1970_,
    new_n1971_, new_n1972_, new_n1973_, new_n1974_, new_n1975_, new_n1976_,
    new_n1977_, new_n1978_, new_n1979_, new_n1980_, new_n1981_, new_n1982_,
    new_n1983_, new_n1984_, new_n1985_, new_n1986_, new_n1987_, new_n1988_,
    new_n1989_, new_n1990_, new_n1991_, new_n1992_, new_n1993_, new_n1994_,
    new_n1995_, new_n1996_, new_n1997_, new_n1998_, new_n1999_, new_n2000_,
    new_n2001_, new_n2002_, new_n2003_, new_n2004_, new_n2005_, new_n2006_,
    new_n2007_, new_n2008_, new_n2009_, new_n2010_, new_n2011_, new_n2012_,
    new_n2013_, new_n2014_, new_n2015_, new_n2016_, new_n2017_, new_n2018_,
    new_n2019_, new_n2020_, new_n2021_, new_n2022_, new_n2023_, new_n2024_,
    new_n2025_, new_n2026_, new_n2027_, new_n2028_, new_n2029_, new_n2030_,
    new_n2031_, new_n2032_, new_n2033_, new_n2034_, new_n2035_, new_n2036_,
    new_n2037_, new_n2038_, new_n2039_, new_n2040_, new_n2041_, new_n2042_,
    new_n2043_, new_n2044_, new_n2045_, new_n2046_, new_n2047_, new_n2048_,
    new_n2049_, new_n2050_, new_n2051_, new_n2052_, new_n2053_, new_n2054_,
    new_n2055_, new_n2056_, new_n2057_, new_n2058_, new_n2059_, new_n2060_,
    new_n2061_, new_n2062_, new_n2063_, new_n2064_, new_n2065_, new_n2066_,
    new_n2067_, new_n2068_, new_n2069_, new_n2070_, new_n2071_, new_n2072_,
    new_n2073_, new_n2074_, new_n2075_, new_n2076_, new_n2077_, new_n2078_,
    new_n2079_, new_n2080_, new_n2081_, new_n2082_, new_n2083_, new_n2084_,
    new_n2085_, new_n2086_, new_n2087_, new_n2088_, new_n2089_, new_n2090_,
    new_n2091_, new_n2092_, new_n2093_, new_n2094_, new_n2095_, new_n2096_,
    new_n2097_, new_n2098_, new_n2099_, new_n2100_, new_n2101_, new_n2102_,
    new_n2103_, new_n2104_, new_n2105_, new_n2106_, new_n2107_, new_n2108_,
    new_n2109_, new_n2110_, new_n2111_, new_n2112_, new_n2113_, new_n2114_,
    new_n2115_, new_n2116_, new_n2117_, new_n2118_, new_n2119_, new_n2120_,
    new_n2121_, new_n2122_, new_n2123_, new_n2124_, new_n2125_, new_n2126_,
    new_n2127_, new_n2128_, new_n2129_, new_n2130_, new_n2131_, new_n2132_,
    new_n2133_, new_n2134_, new_n2135_, new_n2136_, new_n2137_, new_n2138_,
    new_n2139_, new_n2140_, new_n2141_, new_n2142_, new_n2143_, new_n2144_,
    new_n2145_, new_n2146_, new_n2147_, new_n2148_, new_n2149_, new_n2150_,
    new_n2151_, new_n2152_, new_n2153_, new_n2154_, new_n2155_, new_n2156_,
    new_n2157_, new_n2158_, new_n2159_, new_n2160_, new_n2161_, new_n2162_,
    new_n2163_, new_n2164_, new_n2165_, new_n2166_, new_n2167_, new_n2168_,
    new_n2169_, new_n2170_, new_n2171_, new_n2172_, new_n2173_, new_n2174_,
    new_n2175_, new_n2176_, new_n2177_, new_n2178_, new_n2179_, new_n2180_,
    new_n2181_, new_n2182_, new_n2183_, new_n2184_, new_n2185_, new_n2186_,
    new_n2187_, new_n2188_, new_n2189_, new_n2190_, new_n2191_, new_n2192_,
    new_n2193_, new_n2194_, new_n2195_, new_n2196_, new_n2197_, new_n2198_,
    new_n2199_, new_n2200_, new_n2201_, new_n2202_, new_n2203_, new_n2204_,
    new_n2205_, new_n2206_, new_n2207_, new_n2208_, new_n2209_, new_n2210_,
    new_n2211_, new_n2212_, new_n2213_, new_n2214_, new_n2215_, new_n2216_,
    new_n2217_, new_n2218_, new_n2219_, new_n2220_, new_n2221_, new_n2222_,
    new_n2223_, new_n2224_, new_n2225_, new_n2226_, new_n2227_, new_n2228_,
    new_n2229_, new_n2230_, new_n2231_, new_n2232_, new_n2233_, new_n2234_,
    new_n2235_, new_n2236_, new_n2237_, new_n2238_, new_n2239_, new_n2240_,
    new_n2241_, new_n2242_, new_n2243_, new_n2244_, new_n2245_, new_n2246_,
    new_n2247_, new_n2248_, new_n2249_, new_n2250_, new_n2251_, new_n2252_,
    new_n2253_, new_n2254_, new_n2255_, new_n2256_, new_n2257_, new_n2258_,
    new_n2259_, new_n2260_, new_n2261_, new_n2262_, new_n2263_, new_n2264_,
    new_n2265_, new_n2266_, new_n2267_, new_n2268_, new_n2269_, new_n2270_,
    new_n2271_, new_n2272_, new_n2273_, new_n2274_, new_n2275_, new_n2276_,
    new_n2277_, new_n2278_, new_n2279_, new_n2280_, new_n2281_, new_n2282_,
    new_n2283_, new_n2284_, new_n2285_, new_n2286_, new_n2287_, new_n2288_,
    new_n2289_, new_n2290_, new_n2291_, new_n2292_, new_n2293_, new_n2294_,
    new_n2295_, new_n2296_, new_n2297_, new_n2298_, new_n2299_, new_n2300_,
    new_n2301_, new_n2302_, new_n2303_, new_n2304_, new_n2305_, new_n2306_,
    new_n2307_, new_n2308_, new_n2309_, new_n2310_, new_n2311_, new_n2312_,
    new_n2313_, new_n2314_, new_n2315_, new_n2316_, new_n2317_, new_n2318_,
    new_n2319_, new_n2320_, new_n2321_, new_n2322_, new_n2323_, new_n2324_,
    new_n2325_, new_n2326_, new_n2327_, new_n2328_, new_n2329_, new_n2330_,
    new_n2331_, new_n2332_, new_n2333_, new_n2334_, new_n2335_, new_n2336_,
    new_n2337_, new_n2338_, new_n2339_, new_n2340_, new_n2341_, new_n2342_,
    new_n2343_, new_n2344_, new_n2345_, new_n2346_, new_n2347_, new_n2348_,
    new_n2349_, new_n2350_, new_n2351_, new_n2352_, new_n2353_, new_n2354_,
    new_n2355_, new_n2356_, new_n2357_, new_n2358_, new_n2359_, new_n2360_,
    new_n2361_, new_n2362_, new_n2363_, new_n2364_, new_n2365_, new_n2366_,
    new_n2367_, new_n2368_, new_n2369_, new_n2370_, new_n2371_, new_n2372_,
    new_n2373_, new_n2374_, new_n2375_, new_n2376_, new_n2377_, new_n2378_,
    new_n2379_, new_n2380_, new_n2381_, new_n2382_, new_n2383_, new_n2384_,
    new_n2385_, new_n2386_, new_n2387_, new_n2388_, new_n2389_, new_n2390_,
    new_n2391_, new_n2392_, new_n2393_, new_n2394_, new_n2395_, new_n2396_,
    new_n2397_, new_n2398_, new_n2399_, new_n2400_, new_n2401_, new_n2402_,
    new_n2403_, new_n2404_, new_n2405_, new_n2406_, new_n2407_, new_n2408_,
    new_n2409_, new_n2410_, new_n2411_, new_n2412_, new_n2413_, new_n2414_,
    new_n2415_, new_n2416_, new_n2417_, new_n2418_, new_n2419_, new_n2420_,
    new_n2421_, new_n2422_, new_n2423_, new_n2424_, new_n2425_, new_n2426_,
    new_n2427_, new_n2428_, new_n2429_, new_n2430_, new_n2431_, new_n2432_,
    new_n2433_, new_n2434_, new_n2435_, new_n2436_, new_n2437_, new_n2438_,
    new_n2439_, new_n2440_, new_n2441_, new_n2442_, new_n2443_, new_n2444_,
    new_n2445_, new_n2446_, new_n2447_, new_n2448_, new_n2449_, new_n2450_,
    new_n2451_, new_n2452_, new_n2453_, new_n2454_, new_n2455_, new_n2456_,
    new_n2457_, new_n2458_, new_n2459_, new_n2460_, new_n2461_, new_n2462_,
    new_n2463_, new_n2464_, new_n2465_, new_n2466_, new_n2467_, new_n2468_,
    new_n2469_, new_n2470_, new_n2471_;
not  ( new_n50_, \B[9]  );
not  ( new_n51_, \I[1]  );
not  ( new_n52_, \I[0]  );
or   ( new_n53_, new_n52_, new_n51_ );
nor  ( new_n54_, \I[4] , \I[5]  );
nor  ( new_n55_, \I[2] , \I[3]  );
and  ( new_n56_, new_n55_, new_n54_ );
nor  ( new_n57_, \I[6] , \I[7]  );
and  ( new_n58_, new_n57_, new_n56_ );
and  ( new_n59_, new_n58_, new_n53_ );
and  ( new_n60_, new_n52_, \I[1]  );
and  ( new_n61_, new_n60_, new_n58_ );
and  ( new_n62_, new_n61_, \A[2][8]  );
not  ( new_n63_, new_n62_ );
and  ( new_n64_, new_n52_, new_n51_ );
and  ( new_n65_, new_n64_, \A[0][8]  );
and  ( new_n66_, new_n65_, new_n58_ );
and  ( new_n67_, \I[0] , new_n51_ );
and  ( new_n68_, new_n67_, new_n57_ );
and  ( new_n69_, new_n68_, new_n56_ );
and  ( new_n70_, new_n69_, \A[1][8]  );
nor  ( new_n71_, new_n70_, new_n66_ );
and  ( new_n72_, new_n71_, new_n63_ );
and  ( new_n73_, new_n72_, new_n59_ );
or   ( new_n74_, new_n73_, new_n50_ );
not  ( new_n75_, \B[7]  );
and  ( new_n76_, new_n61_, \A[2][9]  );
not  ( new_n77_, new_n76_ );
and  ( new_n78_, new_n64_, \A[0][9]  );
and  ( new_n79_, new_n78_, new_n58_ );
and  ( new_n80_, new_n69_, \A[1][9]  );
nor  ( new_n81_, new_n80_, new_n79_ );
and  ( new_n82_, new_n81_, new_n77_ );
and  ( new_n83_, new_n82_, new_n59_ );
or   ( new_n84_, new_n83_, new_n75_ );
not  ( new_n85_, new_n82_ );
and  ( new_n86_, new_n59_, \B[1]  );
and  ( new_n87_, new_n86_, new_n85_ );
not  ( new_n88_, \B[1]  );
and  ( new_n89_, new_n61_, \A[2][2]  );
not  ( new_n90_, new_n89_ );
and  ( new_n91_, new_n69_, \A[1][2]  );
and  ( new_n92_, new_n64_, \A[0][2]  );
and  ( new_n93_, new_n92_, new_n58_ );
nor  ( new_n94_, new_n93_, new_n91_ );
and  ( new_n95_, new_n94_, new_n90_ );
and  ( new_n96_, new_n95_, new_n59_ );
or   ( new_n97_, new_n96_, new_n88_ );
not  ( new_n98_, \B[0]  );
and  ( new_n99_, new_n61_, \A[2][3]  );
not  ( new_n100_, new_n99_ );
and  ( new_n101_, new_n64_, \A[0][3]  );
and  ( new_n102_, new_n101_, new_n58_ );
and  ( new_n103_, new_n69_, \A[1][3]  );
nor  ( new_n104_, new_n103_, new_n102_ );
and  ( new_n105_, new_n104_, new_n100_ );
and  ( new_n106_, new_n105_, new_n59_ );
or   ( new_n107_, new_n106_, new_n98_ );
and  ( new_n108_, new_n107_, new_n97_ );
not  ( new_n109_, new_n59_ );
nor  ( new_n110_, new_n95_, new_n109_ );
and  ( new_n111_, new_n110_, \B[0]  );
not  ( new_n112_, new_n105_ );
and  ( new_n113_, new_n112_, new_n86_ );
and  ( new_n114_, new_n113_, new_n111_ );
or   ( new_n115_, new_n114_, new_n108_ );
and  ( new_n116_, new_n61_, \A[2][1]  );
not  ( new_n117_, new_n116_ );
and  ( new_n118_, new_n69_, \A[1][1]  );
and  ( new_n119_, new_n64_, \A[0][1]  );
and  ( new_n120_, new_n119_, new_n58_ );
nor  ( new_n121_, new_n120_, new_n118_ );
and  ( new_n122_, new_n121_, new_n117_ );
and  ( new_n123_, new_n122_, new_n59_ );
or   ( new_n124_, new_n123_, new_n88_ );
or   ( new_n125_, new_n96_, new_n98_ );
and  ( new_n126_, new_n125_, new_n124_ );
not  ( new_n127_, new_n122_ );
and  ( new_n128_, new_n127_, new_n86_ );
and  ( new_n129_, new_n128_, new_n111_ );
or   ( new_n130_, new_n129_, new_n126_ );
or   ( new_n131_, new_n123_, new_n98_ );
and  ( new_n132_, new_n61_, \A[2][0]  );
not  ( new_n133_, new_n132_ );
and  ( new_n134_, new_n64_, \A[0][0]  );
and  ( new_n135_, new_n134_, new_n58_ );
and  ( new_n136_, new_n69_, \A[1][0]  );
nor  ( new_n137_, new_n136_, new_n135_ );
and  ( new_n138_, new_n137_, new_n133_ );
and  ( new_n139_, new_n138_, new_n59_ );
or   ( new_n140_, new_n139_, new_n88_ );
or   ( new_n141_, new_n140_, new_n131_ );
or   ( new_n142_, new_n141_, new_n130_ );
or   ( new_n143_, new_n131_, new_n97_ );
and  ( new_n144_, new_n143_, new_n142_ );
or   ( new_n145_, new_n144_, new_n115_ );
or   ( new_n146_, new_n107_, new_n97_ );
and  ( new_n147_, new_n146_, new_n145_ );
or   ( new_n148_, new_n106_, new_n88_ );
and  ( new_n149_, new_n61_, \A[2][4]  );
not  ( new_n150_, new_n149_ );
and  ( new_n151_, new_n64_, \A[0][4]  );
and  ( new_n152_, new_n151_, new_n58_ );
and  ( new_n153_, new_n69_, \A[1][4]  );
nor  ( new_n154_, new_n153_, new_n152_ );
and  ( new_n155_, new_n154_, new_n150_ );
and  ( new_n156_, new_n155_, new_n59_ );
or   ( new_n157_, new_n156_, new_n98_ );
and  ( new_n158_, new_n157_, new_n148_ );
and  ( new_n159_, new_n112_, new_n59_ );
and  ( new_n160_, new_n159_, \B[0]  );
not  ( new_n161_, new_n155_ );
and  ( new_n162_, new_n161_, new_n86_ );
and  ( new_n163_, new_n162_, new_n160_ );
or   ( new_n164_, new_n163_, new_n158_ );
or   ( new_n165_, new_n164_, new_n147_ );
or   ( new_n166_, new_n157_, new_n148_ );
and  ( new_n167_, new_n166_, new_n165_ );
or   ( new_n168_, new_n156_, new_n88_ );
and  ( new_n169_, new_n61_, \A[2][5]  );
not  ( new_n170_, new_n169_ );
and  ( new_n171_, new_n64_, \A[0][5]  );
and  ( new_n172_, new_n171_, new_n58_ );
and  ( new_n173_, new_n69_, \A[1][5]  );
nor  ( new_n174_, new_n173_, new_n172_ );
and  ( new_n175_, new_n174_, new_n170_ );
and  ( new_n176_, new_n175_, new_n59_ );
or   ( new_n177_, new_n176_, new_n98_ );
and  ( new_n178_, new_n177_, new_n168_ );
and  ( new_n179_, new_n161_, new_n59_ );
and  ( new_n180_, new_n179_, \B[0]  );
not  ( new_n181_, new_n175_ );
and  ( new_n182_, new_n181_, new_n86_ );
and  ( new_n183_, new_n182_, new_n180_ );
or   ( new_n184_, new_n183_, new_n178_ );
or   ( new_n185_, new_n184_, new_n167_ );
or   ( new_n186_, new_n177_, new_n168_ );
and  ( new_n187_, new_n186_, new_n185_ );
or   ( new_n188_, new_n176_, new_n88_ );
and  ( new_n189_, new_n61_, \A[2][6]  );
not  ( new_n190_, new_n189_ );
and  ( new_n191_, new_n64_, \A[0][6]  );
and  ( new_n192_, new_n191_, new_n58_ );
and  ( new_n193_, new_n69_, \A[1][6]  );
nor  ( new_n194_, new_n193_, new_n192_ );
and  ( new_n195_, new_n194_, new_n190_ );
and  ( new_n196_, new_n195_, new_n59_ );
or   ( new_n197_, new_n196_, new_n98_ );
and  ( new_n198_, new_n197_, new_n188_ );
and  ( new_n199_, new_n181_, new_n59_ );
and  ( new_n200_, new_n199_, \B[0]  );
not  ( new_n201_, new_n195_ );
and  ( new_n202_, new_n201_, new_n86_ );
and  ( new_n203_, new_n202_, new_n200_ );
or   ( new_n204_, new_n203_, new_n198_ );
or   ( new_n205_, new_n204_, new_n187_ );
or   ( new_n206_, new_n197_, new_n188_ );
and  ( new_n207_, new_n206_, new_n205_ );
or   ( new_n208_, new_n196_, new_n88_ );
and  ( new_n209_, new_n61_, \A[2][7]  );
not  ( new_n210_, new_n209_ );
and  ( new_n211_, new_n64_, \A[0][7]  );
and  ( new_n212_, new_n211_, new_n58_ );
and  ( new_n213_, new_n69_, \A[1][7]  );
nor  ( new_n214_, new_n213_, new_n212_ );
and  ( new_n215_, new_n214_, new_n210_ );
and  ( new_n216_, new_n215_, new_n59_ );
or   ( new_n217_, new_n216_, new_n98_ );
and  ( new_n218_, new_n217_, new_n208_ );
and  ( new_n219_, new_n201_, new_n59_ );
and  ( new_n220_, new_n219_, \B[0]  );
not  ( new_n221_, new_n215_ );
and  ( new_n222_, new_n221_, new_n86_ );
and  ( new_n223_, new_n222_, new_n220_ );
or   ( new_n224_, new_n223_, new_n218_ );
or   ( new_n225_, new_n224_, new_n207_ );
or   ( new_n226_, new_n217_, new_n208_ );
and  ( new_n227_, new_n226_, new_n225_ );
or   ( new_n228_, new_n216_, new_n88_ );
or   ( new_n229_, new_n73_, new_n98_ );
and  ( new_n230_, new_n229_, new_n228_ );
and  ( new_n231_, new_n221_, new_n59_ );
and  ( new_n232_, new_n231_, \B[0]  );
not  ( new_n233_, new_n72_ );
and  ( new_n234_, new_n86_, new_n233_ );
and  ( new_n235_, new_n234_, new_n232_ );
or   ( new_n236_, new_n235_, new_n230_ );
or   ( new_n237_, new_n236_, new_n227_ );
or   ( new_n238_, new_n229_, new_n228_ );
and  ( new_n239_, new_n238_, new_n237_ );
or   ( new_n240_, new_n73_, new_n88_ );
or   ( new_n241_, new_n83_, new_n98_ );
and  ( new_n242_, new_n241_, new_n240_ );
and  ( new_n243_, new_n233_, new_n59_ );
and  ( new_n244_, new_n243_, \B[0]  );
and  ( new_n245_, new_n244_, new_n87_ );
or   ( new_n246_, new_n245_, new_n242_ );
or   ( new_n247_, new_n246_, new_n239_ );
or   ( new_n248_, new_n241_, new_n240_ );
and  ( new_n249_, new_n248_, new_n247_ );
and  ( new_n250_, new_n249_, new_n87_ );
or   ( new_n251_, new_n83_, new_n88_ );
and  ( new_n252_, new_n244_, new_n228_ );
and  ( new_n253_, new_n229_, new_n222_ );
or   ( new_n254_, new_n253_, new_n252_ );
and  ( new_n255_, new_n232_, new_n208_ );
and  ( new_n256_, new_n217_, new_n202_ );
or   ( new_n257_, new_n256_, new_n255_ );
and  ( new_n258_, new_n220_, new_n188_ );
and  ( new_n259_, new_n197_, new_n182_ );
or   ( new_n260_, new_n259_, new_n258_ );
and  ( new_n261_, new_n200_, new_n168_ );
and  ( new_n262_, new_n177_, new_n162_ );
or   ( new_n263_, new_n262_, new_n261_ );
and  ( new_n264_, new_n180_, new_n148_ );
and  ( new_n265_, new_n157_, new_n113_ );
or   ( new_n266_, new_n265_, new_n264_ );
and  ( new_n267_, new_n124_, new_n111_ );
and  ( new_n268_, new_n128_, new_n125_ );
or   ( new_n269_, new_n268_, new_n267_ );
and  ( new_n270_, new_n127_, new_n59_ );
not  ( new_n271_, new_n138_ );
and  ( new_n272_, \B[0] , \B[1]  );
and  ( new_n273_, new_n272_, new_n271_ );
and  ( new_n274_, new_n273_, new_n270_ );
and  ( new_n275_, new_n274_, new_n269_ );
or   ( new_n276_, new_n275_, new_n129_ );
and  ( new_n277_, new_n160_, new_n97_ );
and  ( new_n278_, new_n110_, \B[1]  );
and  ( new_n279_, new_n278_, new_n107_ );
or   ( new_n280_, new_n279_, new_n277_ );
and  ( new_n281_, new_n280_, new_n276_ );
or   ( new_n282_, new_n281_, new_n114_ );
and  ( new_n283_, new_n282_, new_n266_ );
or   ( new_n284_, new_n283_, new_n163_ );
and  ( new_n285_, new_n284_, new_n263_ );
or   ( new_n286_, new_n285_, new_n183_ );
and  ( new_n287_, new_n286_, new_n260_ );
or   ( new_n288_, new_n287_, new_n203_ );
and  ( new_n289_, new_n288_, new_n257_ );
or   ( new_n290_, new_n289_, new_n223_ );
and  ( new_n291_, new_n290_, new_n254_ );
or   ( new_n292_, new_n291_, new_n235_ );
and  ( new_n293_, new_n241_, new_n234_ );
and  ( new_n294_, new_n85_, new_n59_ );
and  ( new_n295_, new_n294_, \B[0]  );
and  ( new_n296_, new_n295_, new_n240_ );
or   ( new_n297_, new_n296_, new_n293_ );
and  ( new_n298_, new_n297_, new_n292_ );
or   ( new_n299_, new_n298_, new_n245_ );
and  ( new_n300_, new_n299_, new_n251_ );
or   ( new_n301_, new_n300_, new_n250_ );
and  ( new_n302_, new_n243_, \B[2]  );
and  ( new_n303_, new_n302_, new_n301_ );
not  ( new_n304_, \B[2]  );
or   ( new_n305_, new_n73_, new_n304_ );
and  ( new_n306_, new_n305_, new_n301_ );
and  ( new_n307_, new_n299_, new_n87_ );
and  ( new_n308_, new_n251_, new_n247_ );
or   ( new_n309_, new_n308_, new_n307_ );
and  ( new_n310_, new_n309_, new_n302_ );
or   ( new_n311_, new_n310_, new_n306_ );
and  ( new_n312_, new_n297_, new_n239_ );
and  ( new_n313_, new_n292_, new_n246_ );
or   ( new_n314_, new_n313_, new_n312_ );
and  ( new_n315_, new_n231_, \B[2]  );
and  ( new_n316_, new_n315_, new_n314_ );
or   ( new_n317_, new_n216_, new_n304_ );
and  ( new_n318_, new_n317_, new_n314_ );
and  ( new_n319_, new_n246_, new_n239_ );
or   ( new_n320_, new_n319_, new_n298_ );
and  ( new_n321_, new_n320_, new_n315_ );
or   ( new_n322_, new_n321_, new_n318_ );
and  ( new_n323_, new_n254_, new_n227_ );
and  ( new_n324_, new_n290_, new_n236_ );
or   ( new_n325_, new_n324_, new_n323_ );
and  ( new_n326_, new_n219_, \B[2]  );
and  ( new_n327_, new_n326_, new_n325_ );
or   ( new_n328_, new_n196_, new_n304_ );
and  ( new_n329_, new_n328_, new_n325_ );
and  ( new_n330_, new_n236_, new_n227_ );
or   ( new_n331_, new_n330_, new_n291_ );
and  ( new_n332_, new_n331_, new_n326_ );
or   ( new_n333_, new_n332_, new_n329_ );
and  ( new_n334_, new_n257_, new_n207_ );
and  ( new_n335_, new_n288_, new_n224_ );
or   ( new_n336_, new_n335_, new_n334_ );
and  ( new_n337_, new_n199_, \B[2]  );
and  ( new_n338_, new_n337_, new_n336_ );
or   ( new_n339_, new_n176_, new_n304_ );
and  ( new_n340_, new_n339_, new_n336_ );
and  ( new_n341_, new_n224_, new_n207_ );
or   ( new_n342_, new_n341_, new_n289_ );
and  ( new_n343_, new_n342_, new_n337_ );
or   ( new_n344_, new_n343_, new_n340_ );
and  ( new_n345_, new_n260_, new_n187_ );
and  ( new_n346_, new_n286_, new_n204_ );
or   ( new_n347_, new_n346_, new_n345_ );
and  ( new_n348_, new_n179_, \B[2]  );
and  ( new_n349_, new_n348_, new_n347_ );
or   ( new_n350_, new_n156_, new_n304_ );
and  ( new_n351_, new_n350_, new_n347_ );
and  ( new_n352_, new_n204_, new_n187_ );
or   ( new_n353_, new_n352_, new_n287_ );
and  ( new_n354_, new_n353_, new_n348_ );
or   ( new_n355_, new_n354_, new_n351_ );
and  ( new_n356_, new_n263_, new_n167_ );
and  ( new_n357_, new_n284_, new_n184_ );
or   ( new_n358_, new_n357_, new_n356_ );
and  ( new_n359_, new_n159_, \B[2]  );
and  ( new_n360_, new_n359_, new_n358_ );
or   ( new_n361_, new_n106_, new_n304_ );
and  ( new_n362_, new_n361_, new_n358_ );
and  ( new_n363_, new_n184_, new_n167_ );
or   ( new_n364_, new_n363_, new_n285_ );
and  ( new_n365_, new_n364_, new_n359_ );
or   ( new_n366_, new_n365_, new_n362_ );
and  ( new_n367_, new_n266_, new_n147_ );
and  ( new_n368_, new_n282_, new_n164_ );
or   ( new_n369_, new_n368_, new_n367_ );
and  ( new_n370_, new_n110_, \B[2]  );
and  ( new_n371_, new_n370_, new_n369_ );
or   ( new_n372_, new_n96_, new_n304_ );
and  ( new_n373_, new_n372_, new_n369_ );
and  ( new_n374_, new_n164_, new_n147_ );
or   ( new_n375_, new_n374_, new_n283_ );
and  ( new_n376_, new_n375_, new_n370_ );
or   ( new_n377_, new_n376_, new_n373_ );
and  ( new_n378_, new_n280_, new_n144_ );
and  ( new_n379_, new_n276_, new_n115_ );
or   ( new_n380_, new_n379_, new_n378_ );
and  ( new_n381_, new_n270_, \B[2]  );
and  ( new_n382_, new_n381_, new_n380_ );
and  ( new_n383_, new_n269_, new_n141_ );
and  ( new_n384_, new_n274_, new_n130_ );
or   ( new_n385_, new_n384_, new_n383_ );
and  ( new_n386_, new_n271_, new_n59_ );
and  ( new_n387_, new_n386_, \B[2]  );
and  ( new_n388_, new_n387_, new_n385_ );
or   ( new_n389_, new_n123_, new_n304_ );
and  ( new_n390_, new_n389_, new_n380_ );
and  ( new_n391_, new_n144_, new_n115_ );
or   ( new_n392_, new_n391_, new_n281_ );
and  ( new_n393_, new_n392_, new_n381_ );
or   ( new_n394_, new_n393_, new_n390_ );
and  ( new_n395_, new_n394_, new_n388_ );
or   ( new_n396_, new_n395_, new_n382_ );
and  ( new_n397_, new_n396_, new_n377_ );
or   ( new_n398_, new_n397_, new_n371_ );
and  ( new_n399_, new_n398_, new_n366_ );
or   ( new_n400_, new_n399_, new_n360_ );
and  ( new_n401_, new_n400_, new_n355_ );
or   ( new_n402_, new_n401_, new_n349_ );
and  ( new_n403_, new_n402_, new_n344_ );
or   ( new_n404_, new_n403_, new_n338_ );
and  ( new_n405_, new_n404_, new_n333_ );
or   ( new_n406_, new_n405_, new_n327_ );
and  ( new_n407_, new_n406_, new_n322_ );
or   ( new_n408_, new_n407_, new_n316_ );
and  ( new_n409_, new_n408_, new_n311_ );
or   ( new_n410_, new_n409_, new_n303_ );
or   ( new_n411_, new_n83_, new_n304_ );
and  ( new_n412_, new_n411_, new_n307_ );
or   ( new_n413_, new_n251_, new_n249_ );
and  ( new_n414_, new_n294_, \B[2]  );
and  ( new_n415_, new_n414_, new_n413_ );
or   ( new_n416_, new_n415_, new_n412_ );
and  ( new_n417_, new_n416_, new_n410_ );
and  ( new_n418_, new_n307_, \B[2]  );
or   ( new_n419_, new_n418_, new_n417_ );
and  ( new_n420_, new_n294_, \B[3]  );
and  ( new_n421_, new_n420_, new_n419_ );
not  ( new_n422_, \B[3]  );
or   ( new_n423_, new_n83_, new_n422_ );
and  ( new_n424_, new_n423_, new_n419_ );
or   ( new_n425_, new_n309_, new_n305_ );
or   ( new_n426_, new_n320_, new_n317_ );
or   ( new_n427_, new_n331_, new_n328_ );
or   ( new_n428_, new_n342_, new_n339_ );
or   ( new_n429_, new_n353_, new_n350_ );
or   ( new_n430_, new_n364_, new_n361_ );
or   ( new_n431_, new_n375_, new_n372_ );
or   ( new_n432_, new_n392_, new_n389_ );
and  ( new_n433_, new_n141_, new_n130_ );
or   ( new_n434_, new_n433_, new_n275_ );
or   ( new_n435_, new_n139_, new_n304_ );
or   ( new_n436_, new_n435_, new_n434_ );
and  ( new_n437_, new_n392_, new_n389_ );
or   ( new_n438_, new_n437_, new_n382_ );
or   ( new_n439_, new_n438_, new_n436_ );
and  ( new_n440_, new_n439_, new_n432_ );
and  ( new_n441_, new_n375_, new_n372_ );
or   ( new_n442_, new_n441_, new_n371_ );
or   ( new_n443_, new_n442_, new_n440_ );
and  ( new_n444_, new_n443_, new_n431_ );
and  ( new_n445_, new_n364_, new_n361_ );
or   ( new_n446_, new_n445_, new_n360_ );
or   ( new_n447_, new_n446_, new_n444_ );
and  ( new_n448_, new_n447_, new_n430_ );
and  ( new_n449_, new_n353_, new_n350_ );
or   ( new_n450_, new_n449_, new_n349_ );
or   ( new_n451_, new_n450_, new_n448_ );
and  ( new_n452_, new_n451_, new_n429_ );
and  ( new_n453_, new_n342_, new_n339_ );
or   ( new_n454_, new_n453_, new_n338_ );
or   ( new_n455_, new_n454_, new_n452_ );
and  ( new_n456_, new_n455_, new_n428_ );
and  ( new_n457_, new_n331_, new_n328_ );
or   ( new_n458_, new_n457_, new_n327_ );
or   ( new_n459_, new_n458_, new_n456_ );
and  ( new_n460_, new_n459_, new_n427_ );
and  ( new_n461_, new_n320_, new_n317_ );
or   ( new_n462_, new_n461_, new_n316_ );
or   ( new_n463_, new_n462_, new_n460_ );
and  ( new_n464_, new_n463_, new_n426_ );
and  ( new_n465_, new_n309_, new_n305_ );
or   ( new_n466_, new_n465_, new_n303_ );
or   ( new_n467_, new_n466_, new_n464_ );
and  ( new_n468_, new_n467_, new_n425_ );
and  ( new_n469_, new_n413_, new_n411_ );
or   ( new_n470_, new_n469_, new_n418_ );
or   ( new_n471_, new_n470_, new_n468_ );
or   ( new_n472_, new_n413_, new_n304_ );
and  ( new_n473_, new_n472_, new_n471_ );
and  ( new_n474_, new_n473_, new_n420_ );
or   ( new_n475_, new_n474_, new_n424_ );
and  ( new_n476_, new_n468_, new_n416_ );
and  ( new_n477_, new_n470_, new_n410_ );
or   ( new_n478_, new_n477_, new_n476_ );
and  ( new_n479_, new_n243_, \B[3]  );
and  ( new_n480_, new_n479_, new_n478_ );
or   ( new_n481_, new_n73_, new_n422_ );
and  ( new_n482_, new_n481_, new_n478_ );
and  ( new_n483_, new_n470_, new_n468_ );
or   ( new_n484_, new_n483_, new_n417_ );
and  ( new_n485_, new_n484_, new_n479_ );
or   ( new_n486_, new_n485_, new_n482_ );
and  ( new_n487_, new_n464_, new_n311_ );
and  ( new_n488_, new_n466_, new_n408_ );
or   ( new_n489_, new_n488_, new_n487_ );
and  ( new_n490_, new_n231_, \B[3]  );
and  ( new_n491_, new_n490_, new_n489_ );
or   ( new_n492_, new_n216_, new_n422_ );
and  ( new_n493_, new_n492_, new_n489_ );
and  ( new_n494_, new_n466_, new_n464_ );
or   ( new_n495_, new_n494_, new_n409_ );
and  ( new_n496_, new_n495_, new_n490_ );
or   ( new_n497_, new_n496_, new_n493_ );
and  ( new_n498_, new_n460_, new_n322_ );
and  ( new_n499_, new_n462_, new_n406_ );
or   ( new_n500_, new_n499_, new_n498_ );
and  ( new_n501_, new_n219_, \B[3]  );
and  ( new_n502_, new_n501_, new_n500_ );
or   ( new_n503_, new_n196_, new_n422_ );
and  ( new_n504_, new_n503_, new_n500_ );
and  ( new_n505_, new_n462_, new_n460_ );
or   ( new_n506_, new_n505_, new_n407_ );
and  ( new_n507_, new_n506_, new_n501_ );
or   ( new_n508_, new_n507_, new_n504_ );
and  ( new_n509_, new_n456_, new_n333_ );
and  ( new_n510_, new_n458_, new_n404_ );
or   ( new_n511_, new_n510_, new_n509_ );
and  ( new_n512_, new_n199_, \B[3]  );
and  ( new_n513_, new_n512_, new_n511_ );
or   ( new_n514_, new_n176_, new_n422_ );
and  ( new_n515_, new_n514_, new_n511_ );
and  ( new_n516_, new_n458_, new_n456_ );
or   ( new_n517_, new_n516_, new_n405_ );
and  ( new_n518_, new_n517_, new_n512_ );
or   ( new_n519_, new_n518_, new_n515_ );
and  ( new_n520_, new_n452_, new_n344_ );
and  ( new_n521_, new_n454_, new_n402_ );
or   ( new_n522_, new_n521_, new_n520_ );
and  ( new_n523_, new_n179_, \B[3]  );
and  ( new_n524_, new_n523_, new_n522_ );
or   ( new_n525_, new_n156_, new_n422_ );
and  ( new_n526_, new_n525_, new_n522_ );
and  ( new_n527_, new_n454_, new_n452_ );
or   ( new_n528_, new_n527_, new_n403_ );
and  ( new_n529_, new_n528_, new_n523_ );
or   ( new_n530_, new_n529_, new_n526_ );
and  ( new_n531_, new_n448_, new_n355_ );
and  ( new_n532_, new_n450_, new_n400_ );
or   ( new_n533_, new_n532_, new_n531_ );
and  ( new_n534_, new_n159_, \B[3]  );
and  ( new_n535_, new_n534_, new_n533_ );
or   ( new_n536_, new_n106_, new_n422_ );
and  ( new_n537_, new_n536_, new_n533_ );
and  ( new_n538_, new_n450_, new_n448_ );
or   ( new_n539_, new_n538_, new_n401_ );
and  ( new_n540_, new_n539_, new_n534_ );
or   ( new_n541_, new_n540_, new_n537_ );
and  ( new_n542_, new_n444_, new_n366_ );
and  ( new_n543_, new_n446_, new_n398_ );
or   ( new_n544_, new_n543_, new_n542_ );
and  ( new_n545_, new_n110_, \B[3]  );
and  ( new_n546_, new_n545_, new_n544_ );
or   ( new_n547_, new_n96_, new_n422_ );
and  ( new_n548_, new_n547_, new_n544_ );
and  ( new_n549_, new_n446_, new_n444_ );
or   ( new_n550_, new_n549_, new_n399_ );
and  ( new_n551_, new_n550_, new_n545_ );
or   ( new_n552_, new_n551_, new_n548_ );
and  ( new_n553_, new_n440_, new_n377_ );
and  ( new_n554_, new_n442_, new_n396_ );
or   ( new_n555_, new_n554_, new_n553_ );
and  ( new_n556_, new_n270_, \B[3]  );
and  ( new_n557_, new_n556_, new_n555_ );
and  ( new_n558_, new_n436_, new_n394_ );
and  ( new_n559_, new_n438_, new_n388_ );
or   ( new_n560_, new_n559_, new_n558_ );
and  ( new_n561_, new_n386_, \B[3]  );
and  ( new_n562_, new_n561_, new_n560_ );
or   ( new_n563_, new_n123_, new_n422_ );
and  ( new_n564_, new_n563_, new_n555_ );
and  ( new_n565_, new_n442_, new_n440_ );
or   ( new_n566_, new_n565_, new_n397_ );
and  ( new_n567_, new_n566_, new_n556_ );
or   ( new_n568_, new_n567_, new_n564_ );
and  ( new_n569_, new_n568_, new_n562_ );
or   ( new_n570_, new_n569_, new_n557_ );
and  ( new_n571_, new_n570_, new_n552_ );
or   ( new_n572_, new_n571_, new_n546_ );
and  ( new_n573_, new_n572_, new_n541_ );
or   ( new_n574_, new_n573_, new_n535_ );
and  ( new_n575_, new_n574_, new_n530_ );
or   ( new_n576_, new_n575_, new_n524_ );
and  ( new_n577_, new_n576_, new_n519_ );
or   ( new_n578_, new_n577_, new_n513_ );
and  ( new_n579_, new_n578_, new_n508_ );
or   ( new_n580_, new_n579_, new_n502_ );
and  ( new_n581_, new_n580_, new_n497_ );
or   ( new_n582_, new_n581_, new_n491_ );
and  ( new_n583_, new_n582_, new_n486_ );
or   ( new_n584_, new_n583_, new_n480_ );
and  ( new_n585_, new_n584_, new_n475_ );
or   ( new_n586_, new_n585_, new_n421_ );
and  ( new_n587_, new_n294_, \B[4]  );
and  ( new_n588_, new_n587_, new_n586_ );
not  ( new_n589_, \B[4]  );
or   ( new_n590_, new_n83_, new_n589_ );
and  ( new_n591_, new_n590_, new_n586_ );
or   ( new_n592_, new_n473_, new_n423_ );
or   ( new_n593_, new_n484_, new_n481_ );
or   ( new_n594_, new_n495_, new_n492_ );
or   ( new_n595_, new_n506_, new_n503_ );
or   ( new_n596_, new_n517_, new_n514_ );
or   ( new_n597_, new_n528_, new_n525_ );
or   ( new_n598_, new_n539_, new_n536_ );
or   ( new_n599_, new_n550_, new_n547_ );
or   ( new_n600_, new_n566_, new_n563_ );
and  ( new_n601_, new_n438_, new_n436_ );
or   ( new_n602_, new_n601_, new_n395_ );
or   ( new_n603_, new_n139_, new_n422_ );
or   ( new_n604_, new_n603_, new_n602_ );
and  ( new_n605_, new_n566_, new_n563_ );
or   ( new_n606_, new_n605_, new_n557_ );
or   ( new_n607_, new_n606_, new_n604_ );
and  ( new_n608_, new_n607_, new_n600_ );
and  ( new_n609_, new_n550_, new_n547_ );
or   ( new_n610_, new_n609_, new_n546_ );
or   ( new_n611_, new_n610_, new_n608_ );
and  ( new_n612_, new_n611_, new_n599_ );
and  ( new_n613_, new_n539_, new_n536_ );
or   ( new_n614_, new_n613_, new_n535_ );
or   ( new_n615_, new_n614_, new_n612_ );
and  ( new_n616_, new_n615_, new_n598_ );
and  ( new_n617_, new_n528_, new_n525_ );
or   ( new_n618_, new_n617_, new_n524_ );
or   ( new_n619_, new_n618_, new_n616_ );
and  ( new_n620_, new_n619_, new_n597_ );
and  ( new_n621_, new_n517_, new_n514_ );
or   ( new_n622_, new_n621_, new_n513_ );
or   ( new_n623_, new_n622_, new_n620_ );
and  ( new_n624_, new_n623_, new_n596_ );
and  ( new_n625_, new_n506_, new_n503_ );
or   ( new_n626_, new_n625_, new_n502_ );
or   ( new_n627_, new_n626_, new_n624_ );
and  ( new_n628_, new_n627_, new_n595_ );
and  ( new_n629_, new_n495_, new_n492_ );
or   ( new_n630_, new_n629_, new_n491_ );
or   ( new_n631_, new_n630_, new_n628_ );
and  ( new_n632_, new_n631_, new_n594_ );
and  ( new_n633_, new_n484_, new_n481_ );
or   ( new_n634_, new_n633_, new_n480_ );
or   ( new_n635_, new_n634_, new_n632_ );
and  ( new_n636_, new_n635_, new_n593_ );
and  ( new_n637_, new_n473_, new_n423_ );
or   ( new_n638_, new_n637_, new_n421_ );
or   ( new_n639_, new_n638_, new_n636_ );
and  ( new_n640_, new_n639_, new_n592_ );
and  ( new_n641_, new_n640_, new_n587_ );
or   ( new_n642_, new_n641_, new_n591_ );
and  ( new_n643_, new_n636_, new_n475_ );
and  ( new_n644_, new_n638_, new_n584_ );
or   ( new_n645_, new_n644_, new_n643_ );
and  ( new_n646_, new_n243_, \B[4]  );
and  ( new_n647_, new_n646_, new_n645_ );
or   ( new_n648_, new_n73_, new_n589_ );
and  ( new_n649_, new_n648_, new_n645_ );
and  ( new_n650_, new_n638_, new_n636_ );
or   ( new_n651_, new_n650_, new_n585_ );
and  ( new_n652_, new_n651_, new_n646_ );
or   ( new_n653_, new_n652_, new_n649_ );
and  ( new_n654_, new_n632_, new_n486_ );
and  ( new_n655_, new_n634_, new_n582_ );
or   ( new_n656_, new_n655_, new_n654_ );
and  ( new_n657_, new_n231_, \B[4]  );
and  ( new_n658_, new_n657_, new_n656_ );
or   ( new_n659_, new_n216_, new_n589_ );
and  ( new_n660_, new_n659_, new_n656_ );
and  ( new_n661_, new_n634_, new_n632_ );
or   ( new_n662_, new_n661_, new_n583_ );
and  ( new_n663_, new_n662_, new_n657_ );
or   ( new_n664_, new_n663_, new_n660_ );
and  ( new_n665_, new_n628_, new_n497_ );
and  ( new_n666_, new_n630_, new_n580_ );
or   ( new_n667_, new_n666_, new_n665_ );
and  ( new_n668_, new_n219_, \B[4]  );
and  ( new_n669_, new_n668_, new_n667_ );
or   ( new_n670_, new_n196_, new_n589_ );
and  ( new_n671_, new_n670_, new_n667_ );
and  ( new_n672_, new_n630_, new_n628_ );
or   ( new_n673_, new_n672_, new_n581_ );
and  ( new_n674_, new_n673_, new_n668_ );
or   ( new_n675_, new_n674_, new_n671_ );
and  ( new_n676_, new_n624_, new_n508_ );
and  ( new_n677_, new_n626_, new_n578_ );
or   ( new_n678_, new_n677_, new_n676_ );
and  ( new_n679_, new_n199_, \B[4]  );
and  ( new_n680_, new_n679_, new_n678_ );
or   ( new_n681_, new_n176_, new_n589_ );
and  ( new_n682_, new_n681_, new_n678_ );
and  ( new_n683_, new_n626_, new_n624_ );
or   ( new_n684_, new_n683_, new_n579_ );
and  ( new_n685_, new_n684_, new_n679_ );
or   ( new_n686_, new_n685_, new_n682_ );
and  ( new_n687_, new_n620_, new_n519_ );
and  ( new_n688_, new_n622_, new_n576_ );
or   ( new_n689_, new_n688_, new_n687_ );
and  ( new_n690_, new_n179_, \B[4]  );
and  ( new_n691_, new_n690_, new_n689_ );
or   ( new_n692_, new_n156_, new_n589_ );
and  ( new_n693_, new_n692_, new_n689_ );
and  ( new_n694_, new_n622_, new_n620_ );
or   ( new_n695_, new_n694_, new_n577_ );
and  ( new_n696_, new_n695_, new_n690_ );
or   ( new_n697_, new_n696_, new_n693_ );
and  ( new_n698_, new_n616_, new_n530_ );
and  ( new_n699_, new_n618_, new_n574_ );
or   ( new_n700_, new_n699_, new_n698_ );
and  ( new_n701_, new_n159_, \B[4]  );
and  ( new_n702_, new_n701_, new_n700_ );
or   ( new_n703_, new_n106_, new_n589_ );
and  ( new_n704_, new_n703_, new_n700_ );
and  ( new_n705_, new_n618_, new_n616_ );
or   ( new_n706_, new_n705_, new_n575_ );
and  ( new_n707_, new_n706_, new_n701_ );
or   ( new_n708_, new_n707_, new_n704_ );
and  ( new_n709_, new_n612_, new_n541_ );
and  ( new_n710_, new_n614_, new_n572_ );
or   ( new_n711_, new_n710_, new_n709_ );
and  ( new_n712_, new_n110_, \B[4]  );
and  ( new_n713_, new_n712_, new_n711_ );
or   ( new_n714_, new_n96_, new_n589_ );
and  ( new_n715_, new_n714_, new_n711_ );
and  ( new_n716_, new_n614_, new_n612_ );
or   ( new_n717_, new_n716_, new_n573_ );
and  ( new_n718_, new_n717_, new_n712_ );
or   ( new_n719_, new_n718_, new_n715_ );
and  ( new_n720_, new_n608_, new_n552_ );
and  ( new_n721_, new_n610_, new_n570_ );
or   ( new_n722_, new_n721_, new_n720_ );
and  ( new_n723_, new_n270_, \B[4]  );
and  ( new_n724_, new_n723_, new_n722_ );
and  ( new_n725_, new_n604_, new_n568_ );
and  ( new_n726_, new_n606_, new_n562_ );
or   ( new_n727_, new_n726_, new_n725_ );
and  ( new_n728_, new_n386_, \B[4]  );
and  ( new_n729_, new_n728_, new_n727_ );
or   ( new_n730_, new_n123_, new_n589_ );
and  ( new_n731_, new_n730_, new_n722_ );
and  ( new_n732_, new_n610_, new_n608_ );
or   ( new_n733_, new_n732_, new_n571_ );
and  ( new_n734_, new_n733_, new_n723_ );
or   ( new_n735_, new_n734_, new_n731_ );
and  ( new_n736_, new_n735_, new_n729_ );
or   ( new_n737_, new_n736_, new_n724_ );
and  ( new_n738_, new_n737_, new_n719_ );
or   ( new_n739_, new_n738_, new_n713_ );
and  ( new_n740_, new_n739_, new_n708_ );
or   ( new_n741_, new_n740_, new_n702_ );
and  ( new_n742_, new_n741_, new_n697_ );
or   ( new_n743_, new_n742_, new_n691_ );
and  ( new_n744_, new_n743_, new_n686_ );
or   ( new_n745_, new_n744_, new_n680_ );
and  ( new_n746_, new_n745_, new_n675_ );
or   ( new_n747_, new_n746_, new_n669_ );
and  ( new_n748_, new_n747_, new_n664_ );
or   ( new_n749_, new_n748_, new_n658_ );
and  ( new_n750_, new_n749_, new_n653_ );
or   ( new_n751_, new_n750_, new_n647_ );
and  ( new_n752_, new_n751_, new_n642_ );
or   ( new_n753_, new_n752_, new_n588_ );
and  ( new_n754_, new_n294_, \B[5]  );
and  ( new_n755_, new_n754_, new_n753_ );
not  ( new_n756_, \B[5]  );
or   ( new_n757_, new_n83_, new_n756_ );
and  ( new_n758_, new_n757_, new_n753_ );
or   ( new_n759_, new_n640_, new_n590_ );
or   ( new_n760_, new_n651_, new_n648_ );
or   ( new_n761_, new_n662_, new_n659_ );
or   ( new_n762_, new_n673_, new_n670_ );
or   ( new_n763_, new_n684_, new_n681_ );
or   ( new_n764_, new_n695_, new_n692_ );
or   ( new_n765_, new_n706_, new_n703_ );
or   ( new_n766_, new_n717_, new_n714_ );
or   ( new_n767_, new_n733_, new_n730_ );
and  ( new_n768_, new_n606_, new_n604_ );
or   ( new_n769_, new_n768_, new_n569_ );
or   ( new_n770_, new_n139_, new_n589_ );
or   ( new_n771_, new_n770_, new_n769_ );
and  ( new_n772_, new_n733_, new_n730_ );
or   ( new_n773_, new_n772_, new_n724_ );
or   ( new_n774_, new_n773_, new_n771_ );
and  ( new_n775_, new_n774_, new_n767_ );
and  ( new_n776_, new_n717_, new_n714_ );
or   ( new_n777_, new_n776_, new_n713_ );
or   ( new_n778_, new_n777_, new_n775_ );
and  ( new_n779_, new_n778_, new_n766_ );
and  ( new_n780_, new_n706_, new_n703_ );
or   ( new_n781_, new_n780_, new_n702_ );
or   ( new_n782_, new_n781_, new_n779_ );
and  ( new_n783_, new_n782_, new_n765_ );
and  ( new_n784_, new_n695_, new_n692_ );
or   ( new_n785_, new_n784_, new_n691_ );
or   ( new_n786_, new_n785_, new_n783_ );
and  ( new_n787_, new_n786_, new_n764_ );
and  ( new_n788_, new_n684_, new_n681_ );
or   ( new_n789_, new_n788_, new_n680_ );
or   ( new_n790_, new_n789_, new_n787_ );
and  ( new_n791_, new_n790_, new_n763_ );
and  ( new_n792_, new_n673_, new_n670_ );
or   ( new_n793_, new_n792_, new_n669_ );
or   ( new_n794_, new_n793_, new_n791_ );
and  ( new_n795_, new_n794_, new_n762_ );
and  ( new_n796_, new_n662_, new_n659_ );
or   ( new_n797_, new_n796_, new_n658_ );
or   ( new_n798_, new_n797_, new_n795_ );
and  ( new_n799_, new_n798_, new_n761_ );
and  ( new_n800_, new_n651_, new_n648_ );
or   ( new_n801_, new_n800_, new_n647_ );
or   ( new_n802_, new_n801_, new_n799_ );
and  ( new_n803_, new_n802_, new_n760_ );
and  ( new_n804_, new_n640_, new_n590_ );
or   ( new_n805_, new_n804_, new_n588_ );
or   ( new_n806_, new_n805_, new_n803_ );
and  ( new_n807_, new_n806_, new_n759_ );
and  ( new_n808_, new_n807_, new_n754_ );
or   ( new_n809_, new_n808_, new_n758_ );
and  ( new_n810_, new_n803_, new_n642_ );
and  ( new_n811_, new_n805_, new_n751_ );
or   ( new_n812_, new_n811_, new_n810_ );
and  ( new_n813_, new_n243_, \B[5]  );
and  ( new_n814_, new_n813_, new_n812_ );
or   ( new_n815_, new_n73_, new_n756_ );
and  ( new_n816_, new_n815_, new_n812_ );
and  ( new_n817_, new_n805_, new_n803_ );
or   ( new_n818_, new_n817_, new_n752_ );
and  ( new_n819_, new_n818_, new_n813_ );
or   ( new_n820_, new_n819_, new_n816_ );
and  ( new_n821_, new_n799_, new_n653_ );
and  ( new_n822_, new_n801_, new_n749_ );
or   ( new_n823_, new_n822_, new_n821_ );
and  ( new_n824_, new_n231_, \B[5]  );
and  ( new_n825_, new_n824_, new_n823_ );
or   ( new_n826_, new_n216_, new_n756_ );
and  ( new_n827_, new_n826_, new_n823_ );
and  ( new_n828_, new_n801_, new_n799_ );
or   ( new_n829_, new_n828_, new_n750_ );
and  ( new_n830_, new_n829_, new_n824_ );
or   ( new_n831_, new_n830_, new_n827_ );
and  ( new_n832_, new_n795_, new_n664_ );
and  ( new_n833_, new_n797_, new_n747_ );
or   ( new_n834_, new_n833_, new_n832_ );
and  ( new_n835_, new_n219_, \B[5]  );
and  ( new_n836_, new_n835_, new_n834_ );
or   ( new_n837_, new_n196_, new_n756_ );
and  ( new_n838_, new_n837_, new_n834_ );
and  ( new_n839_, new_n797_, new_n795_ );
or   ( new_n840_, new_n839_, new_n748_ );
and  ( new_n841_, new_n840_, new_n835_ );
or   ( new_n842_, new_n841_, new_n838_ );
and  ( new_n843_, new_n791_, new_n675_ );
and  ( new_n844_, new_n793_, new_n745_ );
or   ( new_n845_, new_n844_, new_n843_ );
and  ( new_n846_, new_n199_, \B[5]  );
and  ( new_n847_, new_n846_, new_n845_ );
or   ( new_n848_, new_n176_, new_n756_ );
and  ( new_n849_, new_n848_, new_n845_ );
and  ( new_n850_, new_n793_, new_n791_ );
or   ( new_n851_, new_n850_, new_n746_ );
and  ( new_n852_, new_n851_, new_n846_ );
or   ( new_n853_, new_n852_, new_n849_ );
and  ( new_n854_, new_n787_, new_n686_ );
and  ( new_n855_, new_n789_, new_n743_ );
or   ( new_n856_, new_n855_, new_n854_ );
and  ( new_n857_, new_n179_, \B[5]  );
and  ( new_n858_, new_n857_, new_n856_ );
or   ( new_n859_, new_n156_, new_n756_ );
and  ( new_n860_, new_n859_, new_n856_ );
and  ( new_n861_, new_n789_, new_n787_ );
or   ( new_n862_, new_n861_, new_n744_ );
and  ( new_n863_, new_n862_, new_n857_ );
or   ( new_n864_, new_n863_, new_n860_ );
and  ( new_n865_, new_n783_, new_n697_ );
and  ( new_n866_, new_n785_, new_n741_ );
or   ( new_n867_, new_n866_, new_n865_ );
and  ( new_n868_, new_n159_, \B[5]  );
and  ( new_n869_, new_n868_, new_n867_ );
or   ( new_n870_, new_n106_, new_n756_ );
and  ( new_n871_, new_n870_, new_n867_ );
and  ( new_n872_, new_n785_, new_n783_ );
or   ( new_n873_, new_n872_, new_n742_ );
and  ( new_n874_, new_n873_, new_n868_ );
or   ( new_n875_, new_n874_, new_n871_ );
and  ( new_n876_, new_n779_, new_n708_ );
and  ( new_n877_, new_n781_, new_n739_ );
or   ( new_n878_, new_n877_, new_n876_ );
and  ( new_n879_, new_n110_, \B[5]  );
and  ( new_n880_, new_n879_, new_n878_ );
or   ( new_n881_, new_n96_, new_n756_ );
and  ( new_n882_, new_n881_, new_n878_ );
and  ( new_n883_, new_n781_, new_n779_ );
or   ( new_n884_, new_n883_, new_n740_ );
and  ( new_n885_, new_n884_, new_n879_ );
or   ( new_n886_, new_n885_, new_n882_ );
and  ( new_n887_, new_n775_, new_n719_ );
and  ( new_n888_, new_n777_, new_n737_ );
or   ( new_n889_, new_n888_, new_n887_ );
and  ( new_n890_, new_n270_, \B[5]  );
and  ( new_n891_, new_n890_, new_n889_ );
and  ( new_n892_, new_n771_, new_n735_ );
and  ( new_n893_, new_n773_, new_n729_ );
or   ( new_n894_, new_n893_, new_n892_ );
and  ( new_n895_, new_n386_, \B[5]  );
and  ( new_n896_, new_n895_, new_n894_ );
or   ( new_n897_, new_n123_, new_n756_ );
and  ( new_n898_, new_n897_, new_n889_ );
and  ( new_n899_, new_n777_, new_n775_ );
or   ( new_n900_, new_n899_, new_n738_ );
and  ( new_n901_, new_n900_, new_n890_ );
or   ( new_n902_, new_n901_, new_n898_ );
and  ( new_n903_, new_n902_, new_n896_ );
or   ( new_n904_, new_n903_, new_n891_ );
and  ( new_n905_, new_n904_, new_n886_ );
or   ( new_n906_, new_n905_, new_n880_ );
and  ( new_n907_, new_n906_, new_n875_ );
or   ( new_n908_, new_n907_, new_n869_ );
and  ( new_n909_, new_n908_, new_n864_ );
or   ( new_n910_, new_n909_, new_n858_ );
and  ( new_n911_, new_n910_, new_n853_ );
or   ( new_n912_, new_n911_, new_n847_ );
and  ( new_n913_, new_n912_, new_n842_ );
or   ( new_n914_, new_n913_, new_n836_ );
and  ( new_n915_, new_n914_, new_n831_ );
or   ( new_n916_, new_n915_, new_n825_ );
and  ( new_n917_, new_n916_, new_n820_ );
or   ( new_n918_, new_n917_, new_n814_ );
and  ( new_n919_, new_n918_, new_n809_ );
or   ( new_n920_, new_n919_, new_n755_ );
and  ( new_n921_, new_n294_, \B[6]  );
and  ( new_n922_, new_n921_, new_n920_ );
not  ( new_n923_, \B[6]  );
or   ( new_n924_, new_n83_, new_n923_ );
and  ( new_n925_, new_n924_, new_n920_ );
or   ( new_n926_, new_n807_, new_n757_ );
or   ( new_n927_, new_n818_, new_n815_ );
or   ( new_n928_, new_n829_, new_n826_ );
or   ( new_n929_, new_n840_, new_n837_ );
or   ( new_n930_, new_n851_, new_n848_ );
or   ( new_n931_, new_n862_, new_n859_ );
or   ( new_n932_, new_n873_, new_n870_ );
or   ( new_n933_, new_n884_, new_n881_ );
or   ( new_n934_, new_n900_, new_n897_ );
and  ( new_n935_, new_n773_, new_n771_ );
or   ( new_n936_, new_n935_, new_n736_ );
or   ( new_n937_, new_n139_, new_n756_ );
or   ( new_n938_, new_n937_, new_n936_ );
and  ( new_n939_, new_n900_, new_n897_ );
or   ( new_n940_, new_n939_, new_n891_ );
or   ( new_n941_, new_n940_, new_n938_ );
and  ( new_n942_, new_n941_, new_n934_ );
and  ( new_n943_, new_n884_, new_n881_ );
or   ( new_n944_, new_n943_, new_n880_ );
or   ( new_n945_, new_n944_, new_n942_ );
and  ( new_n946_, new_n945_, new_n933_ );
and  ( new_n947_, new_n873_, new_n870_ );
or   ( new_n948_, new_n947_, new_n869_ );
or   ( new_n949_, new_n948_, new_n946_ );
and  ( new_n950_, new_n949_, new_n932_ );
and  ( new_n951_, new_n862_, new_n859_ );
or   ( new_n952_, new_n951_, new_n858_ );
or   ( new_n953_, new_n952_, new_n950_ );
and  ( new_n954_, new_n953_, new_n931_ );
and  ( new_n955_, new_n851_, new_n848_ );
or   ( new_n956_, new_n955_, new_n847_ );
or   ( new_n957_, new_n956_, new_n954_ );
and  ( new_n958_, new_n957_, new_n930_ );
and  ( new_n959_, new_n840_, new_n837_ );
or   ( new_n960_, new_n959_, new_n836_ );
or   ( new_n961_, new_n960_, new_n958_ );
and  ( new_n962_, new_n961_, new_n929_ );
and  ( new_n963_, new_n829_, new_n826_ );
or   ( new_n964_, new_n963_, new_n825_ );
or   ( new_n965_, new_n964_, new_n962_ );
and  ( new_n966_, new_n965_, new_n928_ );
and  ( new_n967_, new_n818_, new_n815_ );
or   ( new_n968_, new_n967_, new_n814_ );
or   ( new_n969_, new_n968_, new_n966_ );
and  ( new_n970_, new_n969_, new_n927_ );
and  ( new_n971_, new_n807_, new_n757_ );
or   ( new_n972_, new_n971_, new_n755_ );
or   ( new_n973_, new_n972_, new_n970_ );
and  ( new_n974_, new_n973_, new_n926_ );
and  ( new_n975_, new_n974_, new_n921_ );
or   ( new_n976_, new_n975_, new_n925_ );
and  ( new_n977_, new_n970_, new_n809_ );
and  ( new_n978_, new_n972_, new_n918_ );
or   ( new_n979_, new_n978_, new_n977_ );
and  ( new_n980_, new_n243_, \B[6]  );
and  ( new_n981_, new_n980_, new_n979_ );
or   ( new_n982_, new_n73_, new_n923_ );
and  ( new_n983_, new_n982_, new_n979_ );
and  ( new_n984_, new_n972_, new_n970_ );
or   ( new_n985_, new_n984_, new_n919_ );
and  ( new_n986_, new_n985_, new_n980_ );
or   ( new_n987_, new_n986_, new_n983_ );
and  ( new_n988_, new_n966_, new_n820_ );
and  ( new_n989_, new_n968_, new_n916_ );
or   ( new_n990_, new_n989_, new_n988_ );
and  ( new_n991_, new_n231_, \B[6]  );
and  ( new_n992_, new_n991_, new_n990_ );
or   ( new_n993_, new_n216_, new_n923_ );
and  ( new_n994_, new_n993_, new_n990_ );
and  ( new_n995_, new_n968_, new_n966_ );
or   ( new_n996_, new_n995_, new_n917_ );
and  ( new_n997_, new_n996_, new_n991_ );
or   ( new_n998_, new_n997_, new_n994_ );
and  ( new_n999_, new_n962_, new_n831_ );
and  ( new_n1000_, new_n964_, new_n914_ );
or   ( new_n1001_, new_n1000_, new_n999_ );
and  ( new_n1002_, new_n219_, \B[6]  );
and  ( new_n1003_, new_n1002_, new_n1001_ );
or   ( new_n1004_, new_n196_, new_n923_ );
and  ( new_n1005_, new_n1004_, new_n1001_ );
and  ( new_n1006_, new_n964_, new_n962_ );
or   ( new_n1007_, new_n1006_, new_n915_ );
and  ( new_n1008_, new_n1007_, new_n1002_ );
or   ( new_n1009_, new_n1008_, new_n1005_ );
and  ( new_n1010_, new_n958_, new_n842_ );
and  ( new_n1011_, new_n960_, new_n912_ );
or   ( new_n1012_, new_n1011_, new_n1010_ );
and  ( new_n1013_, new_n199_, \B[6]  );
and  ( new_n1014_, new_n1013_, new_n1012_ );
or   ( new_n1015_, new_n176_, new_n923_ );
and  ( new_n1016_, new_n1015_, new_n1012_ );
and  ( new_n1017_, new_n960_, new_n958_ );
or   ( new_n1018_, new_n1017_, new_n913_ );
and  ( new_n1019_, new_n1018_, new_n1013_ );
or   ( new_n1020_, new_n1019_, new_n1016_ );
and  ( new_n1021_, new_n954_, new_n853_ );
and  ( new_n1022_, new_n956_, new_n910_ );
or   ( new_n1023_, new_n1022_, new_n1021_ );
and  ( new_n1024_, new_n179_, \B[6]  );
and  ( new_n1025_, new_n1024_, new_n1023_ );
or   ( new_n1026_, new_n156_, new_n923_ );
and  ( new_n1027_, new_n1026_, new_n1023_ );
and  ( new_n1028_, new_n956_, new_n954_ );
or   ( new_n1029_, new_n1028_, new_n911_ );
and  ( new_n1030_, new_n1029_, new_n1024_ );
or   ( new_n1031_, new_n1030_, new_n1027_ );
and  ( new_n1032_, new_n950_, new_n864_ );
and  ( new_n1033_, new_n952_, new_n908_ );
or   ( new_n1034_, new_n1033_, new_n1032_ );
and  ( new_n1035_, new_n159_, \B[6]  );
and  ( new_n1036_, new_n1035_, new_n1034_ );
or   ( new_n1037_, new_n106_, new_n923_ );
and  ( new_n1038_, new_n1037_, new_n1034_ );
and  ( new_n1039_, new_n952_, new_n950_ );
or   ( new_n1040_, new_n1039_, new_n909_ );
and  ( new_n1041_, new_n1040_, new_n1035_ );
or   ( new_n1042_, new_n1041_, new_n1038_ );
and  ( new_n1043_, new_n946_, new_n875_ );
and  ( new_n1044_, new_n948_, new_n906_ );
or   ( new_n1045_, new_n1044_, new_n1043_ );
and  ( new_n1046_, new_n110_, \B[6]  );
and  ( new_n1047_, new_n1046_, new_n1045_ );
or   ( new_n1048_, new_n96_, new_n923_ );
and  ( new_n1049_, new_n1048_, new_n1045_ );
and  ( new_n1050_, new_n948_, new_n946_ );
or   ( new_n1051_, new_n1050_, new_n907_ );
and  ( new_n1052_, new_n1051_, new_n1046_ );
or   ( new_n1053_, new_n1052_, new_n1049_ );
and  ( new_n1054_, new_n942_, new_n886_ );
and  ( new_n1055_, new_n944_, new_n904_ );
or   ( new_n1056_, new_n1055_, new_n1054_ );
and  ( new_n1057_, new_n270_, \B[6]  );
and  ( new_n1058_, new_n1057_, new_n1056_ );
and  ( new_n1059_, new_n938_, new_n902_ );
and  ( new_n1060_, new_n940_, new_n896_ );
or   ( new_n1061_, new_n1060_, new_n1059_ );
and  ( new_n1062_, new_n386_, \B[6]  );
and  ( new_n1063_, new_n1062_, new_n1061_ );
or   ( new_n1064_, new_n123_, new_n923_ );
and  ( new_n1065_, new_n1064_, new_n1056_ );
and  ( new_n1066_, new_n944_, new_n942_ );
or   ( new_n1067_, new_n1066_, new_n905_ );
and  ( new_n1068_, new_n1067_, new_n1057_ );
or   ( new_n1069_, new_n1068_, new_n1065_ );
and  ( new_n1070_, new_n1069_, new_n1063_ );
or   ( new_n1071_, new_n1070_, new_n1058_ );
and  ( new_n1072_, new_n1071_, new_n1053_ );
or   ( new_n1073_, new_n1072_, new_n1047_ );
and  ( new_n1074_, new_n1073_, new_n1042_ );
or   ( new_n1075_, new_n1074_, new_n1036_ );
and  ( new_n1076_, new_n1075_, new_n1031_ );
or   ( new_n1077_, new_n1076_, new_n1025_ );
and  ( new_n1078_, new_n1077_, new_n1020_ );
or   ( new_n1079_, new_n1078_, new_n1014_ );
and  ( new_n1080_, new_n1079_, new_n1009_ );
or   ( new_n1081_, new_n1080_, new_n1003_ );
and  ( new_n1082_, new_n1081_, new_n998_ );
or   ( new_n1083_, new_n1082_, new_n992_ );
and  ( new_n1084_, new_n1083_, new_n987_ );
or   ( new_n1085_, new_n1084_, new_n981_ );
and  ( new_n1086_, new_n1085_, new_n976_ );
or   ( new_n1087_, new_n1086_, new_n922_ );
and  ( new_n1088_, new_n1087_, new_n84_ );
or   ( new_n1089_, new_n974_, new_n924_ );
or   ( new_n1090_, new_n985_, new_n982_ );
or   ( new_n1091_, new_n996_, new_n993_ );
or   ( new_n1092_, new_n1007_, new_n1004_ );
or   ( new_n1093_, new_n1018_, new_n1015_ );
or   ( new_n1094_, new_n1029_, new_n1026_ );
or   ( new_n1095_, new_n1040_, new_n1037_ );
or   ( new_n1096_, new_n1051_, new_n1048_ );
or   ( new_n1097_, new_n1067_, new_n1064_ );
and  ( new_n1098_, new_n940_, new_n938_ );
or   ( new_n1099_, new_n1098_, new_n903_ );
or   ( new_n1100_, new_n139_, new_n923_ );
or   ( new_n1101_, new_n1100_, new_n1099_ );
and  ( new_n1102_, new_n1067_, new_n1064_ );
or   ( new_n1103_, new_n1102_, new_n1058_ );
or   ( new_n1104_, new_n1103_, new_n1101_ );
and  ( new_n1105_, new_n1104_, new_n1097_ );
and  ( new_n1106_, new_n1051_, new_n1048_ );
or   ( new_n1107_, new_n1106_, new_n1047_ );
or   ( new_n1108_, new_n1107_, new_n1105_ );
and  ( new_n1109_, new_n1108_, new_n1096_ );
and  ( new_n1110_, new_n1040_, new_n1037_ );
or   ( new_n1111_, new_n1110_, new_n1036_ );
or   ( new_n1112_, new_n1111_, new_n1109_ );
and  ( new_n1113_, new_n1112_, new_n1095_ );
and  ( new_n1114_, new_n1029_, new_n1026_ );
or   ( new_n1115_, new_n1114_, new_n1025_ );
or   ( new_n1116_, new_n1115_, new_n1113_ );
and  ( new_n1117_, new_n1116_, new_n1094_ );
and  ( new_n1118_, new_n1018_, new_n1015_ );
or   ( new_n1119_, new_n1118_, new_n1014_ );
or   ( new_n1120_, new_n1119_, new_n1117_ );
and  ( new_n1121_, new_n1120_, new_n1093_ );
and  ( new_n1122_, new_n1007_, new_n1004_ );
or   ( new_n1123_, new_n1122_, new_n1003_ );
or   ( new_n1124_, new_n1123_, new_n1121_ );
and  ( new_n1125_, new_n1124_, new_n1092_ );
and  ( new_n1126_, new_n996_, new_n993_ );
or   ( new_n1127_, new_n1126_, new_n992_ );
or   ( new_n1128_, new_n1127_, new_n1125_ );
and  ( new_n1129_, new_n1128_, new_n1091_ );
and  ( new_n1130_, new_n985_, new_n982_ );
or   ( new_n1131_, new_n1130_, new_n981_ );
or   ( new_n1132_, new_n1131_, new_n1129_ );
and  ( new_n1133_, new_n1132_, new_n1090_ );
and  ( new_n1134_, new_n974_, new_n924_ );
or   ( new_n1135_, new_n1134_, new_n922_ );
or   ( new_n1136_, new_n1135_, new_n1133_ );
and  ( new_n1137_, new_n1136_, new_n1089_ );
and  ( new_n1138_, new_n294_, \B[7]  );
and  ( new_n1139_, new_n1138_, new_n1137_ );
or   ( new_n1140_, new_n1139_, new_n1088_ );
and  ( new_n1141_, new_n1133_, new_n976_ );
and  ( new_n1142_, new_n1135_, new_n1085_ );
or   ( new_n1143_, new_n1142_, new_n1141_ );
and  ( new_n1144_, new_n243_, \B[7]  );
and  ( new_n1145_, new_n1144_, new_n1143_ );
or   ( new_n1146_, new_n73_, new_n75_ );
and  ( new_n1147_, new_n1146_, new_n1143_ );
and  ( new_n1148_, new_n1135_, new_n1133_ );
or   ( new_n1149_, new_n1148_, new_n1086_ );
and  ( new_n1150_, new_n1149_, new_n1144_ );
or   ( new_n1151_, new_n1150_, new_n1147_ );
and  ( new_n1152_, new_n1129_, new_n987_ );
and  ( new_n1153_, new_n1131_, new_n1083_ );
or   ( new_n1154_, new_n1153_, new_n1152_ );
and  ( new_n1155_, new_n231_, \B[7]  );
and  ( new_n1156_, new_n1155_, new_n1154_ );
or   ( new_n1157_, new_n216_, new_n75_ );
and  ( new_n1158_, new_n1157_, new_n1154_ );
and  ( new_n1159_, new_n1131_, new_n1129_ );
or   ( new_n1160_, new_n1159_, new_n1084_ );
and  ( new_n1161_, new_n1160_, new_n1155_ );
or   ( new_n1162_, new_n1161_, new_n1158_ );
and  ( new_n1163_, new_n1125_, new_n998_ );
and  ( new_n1164_, new_n1127_, new_n1081_ );
or   ( new_n1165_, new_n1164_, new_n1163_ );
and  ( new_n1166_, new_n219_, \B[7]  );
and  ( new_n1167_, new_n1166_, new_n1165_ );
or   ( new_n1168_, new_n196_, new_n75_ );
and  ( new_n1169_, new_n1168_, new_n1165_ );
and  ( new_n1170_, new_n1127_, new_n1125_ );
or   ( new_n1171_, new_n1170_, new_n1082_ );
and  ( new_n1172_, new_n1171_, new_n1166_ );
or   ( new_n1173_, new_n1172_, new_n1169_ );
and  ( new_n1174_, new_n1121_, new_n1009_ );
and  ( new_n1175_, new_n1123_, new_n1079_ );
or   ( new_n1176_, new_n1175_, new_n1174_ );
and  ( new_n1177_, new_n199_, \B[7]  );
and  ( new_n1178_, new_n1177_, new_n1176_ );
or   ( new_n1179_, new_n176_, new_n75_ );
and  ( new_n1180_, new_n1179_, new_n1176_ );
and  ( new_n1181_, new_n1123_, new_n1121_ );
or   ( new_n1182_, new_n1181_, new_n1080_ );
and  ( new_n1183_, new_n1182_, new_n1177_ );
or   ( new_n1184_, new_n1183_, new_n1180_ );
and  ( new_n1185_, new_n1117_, new_n1020_ );
and  ( new_n1186_, new_n1119_, new_n1077_ );
or   ( new_n1187_, new_n1186_, new_n1185_ );
and  ( new_n1188_, new_n179_, \B[7]  );
and  ( new_n1189_, new_n1188_, new_n1187_ );
or   ( new_n1190_, new_n156_, new_n75_ );
and  ( new_n1191_, new_n1190_, new_n1187_ );
and  ( new_n1192_, new_n1119_, new_n1117_ );
or   ( new_n1193_, new_n1192_, new_n1078_ );
and  ( new_n1194_, new_n1193_, new_n1188_ );
or   ( new_n1195_, new_n1194_, new_n1191_ );
and  ( new_n1196_, new_n1113_, new_n1031_ );
and  ( new_n1197_, new_n1115_, new_n1075_ );
or   ( new_n1198_, new_n1197_, new_n1196_ );
and  ( new_n1199_, new_n159_, \B[7]  );
and  ( new_n1200_, new_n1199_, new_n1198_ );
or   ( new_n1201_, new_n106_, new_n75_ );
and  ( new_n1202_, new_n1201_, new_n1198_ );
and  ( new_n1203_, new_n1115_, new_n1113_ );
or   ( new_n1204_, new_n1203_, new_n1076_ );
and  ( new_n1205_, new_n1204_, new_n1199_ );
or   ( new_n1206_, new_n1205_, new_n1202_ );
and  ( new_n1207_, new_n1109_, new_n1042_ );
and  ( new_n1208_, new_n1111_, new_n1073_ );
or   ( new_n1209_, new_n1208_, new_n1207_ );
and  ( new_n1210_, new_n110_, \B[7]  );
and  ( new_n1211_, new_n1210_, new_n1209_ );
or   ( new_n1212_, new_n96_, new_n75_ );
and  ( new_n1213_, new_n1212_, new_n1209_ );
and  ( new_n1214_, new_n1111_, new_n1109_ );
or   ( new_n1215_, new_n1214_, new_n1074_ );
and  ( new_n1216_, new_n1215_, new_n1210_ );
or   ( new_n1217_, new_n1216_, new_n1213_ );
and  ( new_n1218_, new_n1105_, new_n1053_ );
and  ( new_n1219_, new_n1107_, new_n1071_ );
or   ( new_n1220_, new_n1219_, new_n1218_ );
and  ( new_n1221_, new_n270_, \B[7]  );
and  ( new_n1222_, new_n1221_, new_n1220_ );
and  ( new_n1223_, new_n1101_, new_n1069_ );
and  ( new_n1224_, new_n1103_, new_n1063_ );
or   ( new_n1225_, new_n1224_, new_n1223_ );
and  ( new_n1226_, new_n386_, \B[7]  );
and  ( new_n1227_, new_n1226_, new_n1225_ );
or   ( new_n1228_, new_n123_, new_n75_ );
and  ( new_n1229_, new_n1228_, new_n1220_ );
and  ( new_n1230_, new_n1107_, new_n1105_ );
or   ( new_n1231_, new_n1230_, new_n1072_ );
and  ( new_n1232_, new_n1231_, new_n1221_ );
or   ( new_n1233_, new_n1232_, new_n1229_ );
and  ( new_n1234_, new_n1233_, new_n1227_ );
or   ( new_n1235_, new_n1234_, new_n1222_ );
and  ( new_n1236_, new_n1235_, new_n1217_ );
or   ( new_n1237_, new_n1236_, new_n1211_ );
and  ( new_n1238_, new_n1237_, new_n1206_ );
or   ( new_n1239_, new_n1238_, new_n1200_ );
and  ( new_n1240_, new_n1239_, new_n1195_ );
or   ( new_n1241_, new_n1240_, new_n1189_ );
and  ( new_n1242_, new_n1241_, new_n1184_ );
or   ( new_n1243_, new_n1242_, new_n1178_ );
and  ( new_n1244_, new_n1243_, new_n1173_ );
or   ( new_n1245_, new_n1244_, new_n1167_ );
and  ( new_n1246_, new_n1245_, new_n1162_ );
or   ( new_n1247_, new_n1246_, new_n1156_ );
and  ( new_n1248_, new_n1247_, new_n1151_ );
or   ( new_n1249_, new_n1248_, new_n1145_ );
and  ( new_n1250_, new_n1249_, new_n1140_ );
and  ( new_n1251_, new_n1138_, new_n1087_ );
or   ( new_n1252_, new_n1251_, new_n1250_ );
not  ( new_n1253_, \B[8]  );
or   ( new_n1254_, new_n83_, new_n1253_ );
and  ( new_n1255_, new_n1254_, new_n1252_ );
and  ( new_n1256_, new_n294_, \B[8]  );
or   ( new_n1257_, new_n1137_, new_n84_ );
or   ( new_n1258_, new_n1149_, new_n1146_ );
or   ( new_n1259_, new_n1160_, new_n1157_ );
or   ( new_n1260_, new_n1171_, new_n1168_ );
or   ( new_n1261_, new_n1182_, new_n1179_ );
or   ( new_n1262_, new_n1193_, new_n1190_ );
or   ( new_n1263_, new_n1204_, new_n1201_ );
or   ( new_n1264_, new_n1215_, new_n1212_ );
or   ( new_n1265_, new_n1231_, new_n1228_ );
and  ( new_n1266_, new_n1103_, new_n1101_ );
or   ( new_n1267_, new_n1266_, new_n1070_ );
or   ( new_n1268_, new_n139_, new_n75_ );
or   ( new_n1269_, new_n1268_, new_n1267_ );
and  ( new_n1270_, new_n1231_, new_n1228_ );
or   ( new_n1271_, new_n1270_, new_n1222_ );
or   ( new_n1272_, new_n1271_, new_n1269_ );
and  ( new_n1273_, new_n1272_, new_n1265_ );
and  ( new_n1274_, new_n1215_, new_n1212_ );
or   ( new_n1275_, new_n1274_, new_n1211_ );
or   ( new_n1276_, new_n1275_, new_n1273_ );
and  ( new_n1277_, new_n1276_, new_n1264_ );
and  ( new_n1278_, new_n1204_, new_n1201_ );
or   ( new_n1279_, new_n1278_, new_n1200_ );
or   ( new_n1280_, new_n1279_, new_n1277_ );
and  ( new_n1281_, new_n1280_, new_n1263_ );
and  ( new_n1282_, new_n1193_, new_n1190_ );
or   ( new_n1283_, new_n1282_, new_n1189_ );
or   ( new_n1284_, new_n1283_, new_n1281_ );
and  ( new_n1285_, new_n1284_, new_n1262_ );
and  ( new_n1286_, new_n1182_, new_n1179_ );
or   ( new_n1287_, new_n1286_, new_n1178_ );
or   ( new_n1288_, new_n1287_, new_n1285_ );
and  ( new_n1289_, new_n1288_, new_n1261_ );
and  ( new_n1290_, new_n1171_, new_n1168_ );
or   ( new_n1291_, new_n1290_, new_n1167_ );
or   ( new_n1292_, new_n1291_, new_n1289_ );
and  ( new_n1293_, new_n1292_, new_n1260_ );
and  ( new_n1294_, new_n1160_, new_n1157_ );
or   ( new_n1295_, new_n1294_, new_n1156_ );
or   ( new_n1296_, new_n1295_, new_n1293_ );
and  ( new_n1297_, new_n1296_, new_n1259_ );
and  ( new_n1298_, new_n1149_, new_n1146_ );
or   ( new_n1299_, new_n1298_, new_n1145_ );
or   ( new_n1300_, new_n1299_, new_n1297_ );
and  ( new_n1301_, new_n1300_, new_n1258_ );
and  ( new_n1302_, new_n1137_, new_n84_ );
or   ( new_n1303_, new_n1302_, new_n1251_ );
or   ( new_n1304_, new_n1303_, new_n1301_ );
and  ( new_n1305_, new_n1304_, new_n1257_ );
and  ( new_n1306_, new_n1305_, new_n1256_ );
or   ( new_n1307_, new_n1306_, new_n1255_ );
or   ( new_n1308_, new_n73_, new_n1253_ );
and  ( new_n1309_, new_n1303_, new_n1301_ );
or   ( new_n1310_, new_n1309_, new_n1250_ );
or   ( new_n1311_, new_n1310_, new_n1308_ );
or   ( new_n1312_, new_n216_, new_n1253_ );
and  ( new_n1313_, new_n1299_, new_n1297_ );
or   ( new_n1314_, new_n1313_, new_n1248_ );
or   ( new_n1315_, new_n1314_, new_n1312_ );
or   ( new_n1316_, new_n196_, new_n1253_ );
and  ( new_n1317_, new_n1295_, new_n1293_ );
or   ( new_n1318_, new_n1317_, new_n1246_ );
or   ( new_n1319_, new_n1318_, new_n1316_ );
or   ( new_n1320_, new_n176_, new_n1253_ );
and  ( new_n1321_, new_n1291_, new_n1289_ );
or   ( new_n1322_, new_n1321_, new_n1244_ );
or   ( new_n1323_, new_n1322_, new_n1320_ );
or   ( new_n1324_, new_n156_, new_n1253_ );
and  ( new_n1325_, new_n1287_, new_n1285_ );
or   ( new_n1326_, new_n1325_, new_n1242_ );
or   ( new_n1327_, new_n1326_, new_n1324_ );
or   ( new_n1328_, new_n106_, new_n1253_ );
and  ( new_n1329_, new_n1283_, new_n1281_ );
or   ( new_n1330_, new_n1329_, new_n1240_ );
or   ( new_n1331_, new_n1330_, new_n1328_ );
or   ( new_n1332_, new_n96_, new_n1253_ );
and  ( new_n1333_, new_n1279_, new_n1277_ );
or   ( new_n1334_, new_n1333_, new_n1238_ );
or   ( new_n1335_, new_n1334_, new_n1332_ );
or   ( new_n1336_, new_n123_, new_n1253_ );
and  ( new_n1337_, new_n1275_, new_n1273_ );
or   ( new_n1338_, new_n1337_, new_n1236_ );
or   ( new_n1339_, new_n1338_, new_n1336_ );
and  ( new_n1340_, new_n1271_, new_n1269_ );
or   ( new_n1341_, new_n1340_, new_n1234_ );
or   ( new_n1342_, new_n139_, new_n1253_ );
or   ( new_n1343_, new_n1342_, new_n1341_ );
and  ( new_n1344_, new_n1273_, new_n1217_ );
and  ( new_n1345_, new_n1275_, new_n1235_ );
or   ( new_n1346_, new_n1345_, new_n1344_ );
and  ( new_n1347_, new_n270_, \B[8]  );
and  ( new_n1348_, new_n1347_, new_n1346_ );
and  ( new_n1349_, new_n1338_, new_n1336_ );
or   ( new_n1350_, new_n1349_, new_n1348_ );
or   ( new_n1351_, new_n1350_, new_n1343_ );
and  ( new_n1352_, new_n1351_, new_n1339_ );
and  ( new_n1353_, new_n1277_, new_n1206_ );
and  ( new_n1354_, new_n1279_, new_n1237_ );
or   ( new_n1355_, new_n1354_, new_n1353_ );
and  ( new_n1356_, new_n110_, \B[8]  );
and  ( new_n1357_, new_n1356_, new_n1355_ );
and  ( new_n1358_, new_n1334_, new_n1332_ );
or   ( new_n1359_, new_n1358_, new_n1357_ );
or   ( new_n1360_, new_n1359_, new_n1352_ );
and  ( new_n1361_, new_n1360_, new_n1335_ );
and  ( new_n1362_, new_n1281_, new_n1195_ );
and  ( new_n1363_, new_n1283_, new_n1239_ );
or   ( new_n1364_, new_n1363_, new_n1362_ );
and  ( new_n1365_, new_n159_, \B[8]  );
and  ( new_n1366_, new_n1365_, new_n1364_ );
and  ( new_n1367_, new_n1330_, new_n1328_ );
or   ( new_n1368_, new_n1367_, new_n1366_ );
or   ( new_n1369_, new_n1368_, new_n1361_ );
and  ( new_n1370_, new_n1369_, new_n1331_ );
and  ( new_n1371_, new_n1285_, new_n1184_ );
and  ( new_n1372_, new_n1287_, new_n1241_ );
or   ( new_n1373_, new_n1372_, new_n1371_ );
and  ( new_n1374_, new_n179_, \B[8]  );
and  ( new_n1375_, new_n1374_, new_n1373_ );
and  ( new_n1376_, new_n1326_, new_n1324_ );
or   ( new_n1377_, new_n1376_, new_n1375_ );
or   ( new_n1378_, new_n1377_, new_n1370_ );
and  ( new_n1379_, new_n1378_, new_n1327_ );
and  ( new_n1380_, new_n1289_, new_n1173_ );
and  ( new_n1381_, new_n1291_, new_n1243_ );
or   ( new_n1382_, new_n1381_, new_n1380_ );
and  ( new_n1383_, new_n199_, \B[8]  );
and  ( new_n1384_, new_n1383_, new_n1382_ );
and  ( new_n1385_, new_n1322_, new_n1320_ );
or   ( new_n1386_, new_n1385_, new_n1384_ );
or   ( new_n1387_, new_n1386_, new_n1379_ );
and  ( new_n1388_, new_n1387_, new_n1323_ );
and  ( new_n1389_, new_n1293_, new_n1162_ );
and  ( new_n1390_, new_n1295_, new_n1245_ );
or   ( new_n1391_, new_n1390_, new_n1389_ );
and  ( new_n1392_, new_n219_, \B[8]  );
and  ( new_n1393_, new_n1392_, new_n1391_ );
and  ( new_n1394_, new_n1318_, new_n1316_ );
or   ( new_n1395_, new_n1394_, new_n1393_ );
or   ( new_n1396_, new_n1395_, new_n1388_ );
and  ( new_n1397_, new_n1396_, new_n1319_ );
and  ( new_n1398_, new_n1297_, new_n1151_ );
and  ( new_n1399_, new_n1299_, new_n1247_ );
or   ( new_n1400_, new_n1399_, new_n1398_ );
and  ( new_n1401_, new_n231_, \B[8]  );
and  ( new_n1402_, new_n1401_, new_n1400_ );
and  ( new_n1403_, new_n1314_, new_n1312_ );
or   ( new_n1404_, new_n1403_, new_n1402_ );
or   ( new_n1405_, new_n1404_, new_n1397_ );
and  ( new_n1406_, new_n1405_, new_n1315_ );
and  ( new_n1407_, new_n1301_, new_n1140_ );
and  ( new_n1408_, new_n1303_, new_n1249_ );
or   ( new_n1409_, new_n1408_, new_n1407_ );
and  ( new_n1410_, new_n243_, \B[8]  );
and  ( new_n1411_, new_n1410_, new_n1409_ );
and  ( new_n1412_, new_n1310_, new_n1308_ );
or   ( new_n1413_, new_n1412_, new_n1411_ );
or   ( new_n1414_, new_n1413_, new_n1406_ );
and  ( new_n1415_, new_n1414_, new_n1311_ );
and  ( new_n1416_, new_n1415_, new_n1307_ );
and  ( new_n1417_, new_n1409_, new_n1308_ );
and  ( new_n1418_, new_n1410_, new_n1310_ );
or   ( new_n1419_, new_n1418_, new_n1417_ );
and  ( new_n1420_, new_n1400_, new_n1312_ );
and  ( new_n1421_, new_n1401_, new_n1314_ );
or   ( new_n1422_, new_n1421_, new_n1420_ );
and  ( new_n1423_, new_n1391_, new_n1316_ );
and  ( new_n1424_, new_n1392_, new_n1318_ );
or   ( new_n1425_, new_n1424_, new_n1423_ );
and  ( new_n1426_, new_n1382_, new_n1320_ );
and  ( new_n1427_, new_n1383_, new_n1322_ );
or   ( new_n1428_, new_n1427_, new_n1426_ );
and  ( new_n1429_, new_n1373_, new_n1324_ );
and  ( new_n1430_, new_n1374_, new_n1326_ );
or   ( new_n1431_, new_n1430_, new_n1429_ );
and  ( new_n1432_, new_n1364_, new_n1328_ );
and  ( new_n1433_, new_n1365_, new_n1330_ );
or   ( new_n1434_, new_n1433_, new_n1432_ );
and  ( new_n1435_, new_n1355_, new_n1332_ );
and  ( new_n1436_, new_n1356_, new_n1334_ );
or   ( new_n1437_, new_n1436_, new_n1435_ );
and  ( new_n1438_, new_n1269_, new_n1233_ );
and  ( new_n1439_, new_n1271_, new_n1227_ );
or   ( new_n1440_, new_n1439_, new_n1438_ );
and  ( new_n1441_, new_n386_, \B[8]  );
and  ( new_n1442_, new_n1441_, new_n1440_ );
and  ( new_n1443_, new_n1346_, new_n1336_ );
and  ( new_n1444_, new_n1347_, new_n1338_ );
or   ( new_n1445_, new_n1444_, new_n1443_ );
and  ( new_n1446_, new_n1445_, new_n1442_ );
or   ( new_n1447_, new_n1446_, new_n1348_ );
and  ( new_n1448_, new_n1447_, new_n1437_ );
or   ( new_n1449_, new_n1448_, new_n1357_ );
and  ( new_n1450_, new_n1449_, new_n1434_ );
or   ( new_n1451_, new_n1450_, new_n1366_ );
and  ( new_n1452_, new_n1451_, new_n1431_ );
or   ( new_n1453_, new_n1452_, new_n1375_ );
and  ( new_n1454_, new_n1453_, new_n1428_ );
or   ( new_n1455_, new_n1454_, new_n1384_ );
and  ( new_n1456_, new_n1455_, new_n1425_ );
or   ( new_n1457_, new_n1456_, new_n1393_ );
and  ( new_n1458_, new_n1457_, new_n1422_ );
or   ( new_n1459_, new_n1458_, new_n1402_ );
and  ( new_n1460_, new_n1459_, new_n1419_ );
or   ( new_n1461_, new_n1460_, new_n1411_ );
and  ( new_n1462_, new_n1256_, new_n1252_ );
and  ( new_n1463_, new_n1305_, new_n1254_ );
or   ( new_n1464_, new_n1463_, new_n1462_ );
and  ( new_n1465_, new_n1464_, new_n1461_ );
or   ( new_n1466_, new_n1465_, new_n1416_ );
and  ( new_n1467_, new_n1466_, new_n74_ );
and  ( new_n1468_, new_n1461_, new_n1307_ );
and  ( new_n1469_, new_n1464_, new_n1415_ );
or   ( new_n1470_, new_n1469_, new_n1468_ );
and  ( new_n1471_, new_n243_, \B[9]  );
and  ( new_n1472_, new_n1471_, new_n1470_ );
or   ( new_n1473_, new_n1472_, new_n1467_ );
or   ( new_n1474_, new_n216_, new_n50_ );
and  ( new_n1475_, new_n1413_, new_n1406_ );
or   ( new_n1476_, new_n1475_, new_n1460_ );
or   ( new_n1477_, new_n1476_, new_n1474_ );
and  ( new_n1478_, new_n1419_, new_n1406_ );
and  ( new_n1479_, new_n1459_, new_n1413_ );
or   ( new_n1480_, new_n1479_, new_n1478_ );
and  ( new_n1481_, new_n231_, \B[9]  );
and  ( new_n1482_, new_n1481_, new_n1480_ );
and  ( new_n1483_, new_n1476_, new_n1474_ );
or   ( new_n1484_, new_n1483_, new_n1482_ );
or   ( new_n1485_, new_n196_, new_n50_ );
and  ( new_n1486_, new_n1404_, new_n1397_ );
or   ( new_n1487_, new_n1486_, new_n1458_ );
or   ( new_n1488_, new_n1487_, new_n1485_ );
and  ( new_n1489_, new_n1422_, new_n1397_ );
and  ( new_n1490_, new_n1457_, new_n1404_ );
or   ( new_n1491_, new_n1490_, new_n1489_ );
and  ( new_n1492_, new_n219_, \B[9]  );
and  ( new_n1493_, new_n1492_, new_n1491_ );
and  ( new_n1494_, new_n1487_, new_n1485_ );
or   ( new_n1495_, new_n1494_, new_n1493_ );
or   ( new_n1496_, new_n176_, new_n50_ );
and  ( new_n1497_, new_n1395_, new_n1388_ );
or   ( new_n1498_, new_n1497_, new_n1456_ );
or   ( new_n1499_, new_n1498_, new_n1496_ );
and  ( new_n1500_, new_n1425_, new_n1388_ );
and  ( new_n1501_, new_n1455_, new_n1395_ );
or   ( new_n1502_, new_n1501_, new_n1500_ );
and  ( new_n1503_, new_n199_, \B[9]  );
and  ( new_n1504_, new_n1503_, new_n1502_ );
and  ( new_n1505_, new_n1498_, new_n1496_ );
or   ( new_n1506_, new_n1505_, new_n1504_ );
or   ( new_n1507_, new_n156_, new_n50_ );
and  ( new_n1508_, new_n1386_, new_n1379_ );
or   ( new_n1509_, new_n1508_, new_n1454_ );
or   ( new_n1510_, new_n1509_, new_n1507_ );
and  ( new_n1511_, new_n1428_, new_n1379_ );
and  ( new_n1512_, new_n1453_, new_n1386_ );
or   ( new_n1513_, new_n1512_, new_n1511_ );
and  ( new_n1514_, new_n179_, \B[9]  );
and  ( new_n1515_, new_n1514_, new_n1513_ );
and  ( new_n1516_, new_n1509_, new_n1507_ );
or   ( new_n1517_, new_n1516_, new_n1515_ );
or   ( new_n1518_, new_n106_, new_n50_ );
and  ( new_n1519_, new_n1377_, new_n1370_ );
or   ( new_n1520_, new_n1519_, new_n1452_ );
or   ( new_n1521_, new_n1520_, new_n1518_ );
and  ( new_n1522_, new_n1431_, new_n1370_ );
and  ( new_n1523_, new_n1451_, new_n1377_ );
or   ( new_n1524_, new_n1523_, new_n1522_ );
and  ( new_n1525_, new_n159_, \B[9]  );
and  ( new_n1526_, new_n1525_, new_n1524_ );
and  ( new_n1527_, new_n1520_, new_n1518_ );
or   ( new_n1528_, new_n1527_, new_n1526_ );
or   ( new_n1529_, new_n96_, new_n50_ );
and  ( new_n1530_, new_n1368_, new_n1361_ );
or   ( new_n1531_, new_n1530_, new_n1450_ );
or   ( new_n1532_, new_n1531_, new_n1529_ );
and  ( new_n1533_, new_n1434_, new_n1361_ );
and  ( new_n1534_, new_n1449_, new_n1368_ );
or   ( new_n1535_, new_n1534_, new_n1533_ );
and  ( new_n1536_, new_n110_, \B[9]  );
and  ( new_n1537_, new_n1536_, new_n1535_ );
and  ( new_n1538_, new_n1531_, new_n1529_ );
or   ( new_n1539_, new_n1538_, new_n1537_ );
or   ( new_n1540_, new_n123_, new_n50_ );
and  ( new_n1541_, new_n1359_, new_n1352_ );
or   ( new_n1542_, new_n1541_, new_n1448_ );
or   ( new_n1543_, new_n1542_, new_n1540_ );
and  ( new_n1544_, new_n1437_, new_n1352_ );
and  ( new_n1545_, new_n1447_, new_n1359_ );
or   ( new_n1546_, new_n1545_, new_n1544_ );
and  ( new_n1547_, new_n270_, \B[9]  );
and  ( new_n1548_, new_n1547_, new_n1546_ );
and  ( new_n1549_, new_n1542_, new_n1540_ );
or   ( new_n1550_, new_n1549_, new_n1548_ );
and  ( new_n1551_, new_n1350_, new_n1343_ );
or   ( new_n1552_, new_n1551_, new_n1446_ );
or   ( new_n1553_, new_n139_, new_n50_ );
or   ( new_n1554_, new_n1553_, new_n1552_ );
or   ( new_n1555_, new_n1554_, new_n1550_ );
and  ( new_n1556_, new_n1555_, new_n1543_ );
or   ( new_n1557_, new_n1556_, new_n1539_ );
and  ( new_n1558_, new_n1557_, new_n1532_ );
or   ( new_n1559_, new_n1558_, new_n1528_ );
and  ( new_n1560_, new_n1559_, new_n1521_ );
or   ( new_n1561_, new_n1560_, new_n1517_ );
and  ( new_n1562_, new_n1561_, new_n1510_ );
or   ( new_n1563_, new_n1562_, new_n1506_ );
and  ( new_n1564_, new_n1563_, new_n1499_ );
or   ( new_n1565_, new_n1564_, new_n1495_ );
and  ( new_n1566_, new_n1565_, new_n1488_ );
or   ( new_n1567_, new_n1566_, new_n1484_ );
and  ( new_n1568_, new_n1567_, new_n1477_ );
and  ( new_n1569_, new_n1568_, new_n1473_ );
and  ( new_n1570_, new_n1480_, new_n1474_ );
and  ( new_n1571_, new_n1481_, new_n1476_ );
or   ( new_n1572_, new_n1571_, new_n1570_ );
and  ( new_n1573_, new_n1491_, new_n1485_ );
and  ( new_n1574_, new_n1492_, new_n1487_ );
or   ( new_n1575_, new_n1574_, new_n1573_ );
and  ( new_n1576_, new_n1502_, new_n1496_ );
and  ( new_n1577_, new_n1503_, new_n1498_ );
or   ( new_n1578_, new_n1577_, new_n1576_ );
and  ( new_n1579_, new_n1513_, new_n1507_ );
and  ( new_n1580_, new_n1514_, new_n1509_ );
or   ( new_n1581_, new_n1580_, new_n1579_ );
and  ( new_n1582_, new_n1524_, new_n1518_ );
and  ( new_n1583_, new_n1525_, new_n1520_ );
or   ( new_n1584_, new_n1583_, new_n1582_ );
and  ( new_n1585_, new_n1535_, new_n1529_ );
and  ( new_n1586_, new_n1536_, new_n1531_ );
or   ( new_n1587_, new_n1586_, new_n1585_ );
and  ( new_n1588_, new_n1445_, new_n1343_ );
and  ( new_n1589_, new_n1442_, new_n1350_ );
or   ( new_n1590_, new_n1589_, new_n1588_ );
and  ( new_n1591_, new_n386_, \B[9]  );
and  ( new_n1592_, new_n1591_, new_n1590_ );
and  ( new_n1593_, new_n1546_, new_n1540_ );
and  ( new_n1594_, new_n1547_, new_n1542_ );
or   ( new_n1595_, new_n1594_, new_n1593_ );
and  ( new_n1596_, new_n1595_, new_n1592_ );
or   ( new_n1597_, new_n1596_, new_n1548_ );
and  ( new_n1598_, new_n1597_, new_n1587_ );
or   ( new_n1599_, new_n1598_, new_n1537_ );
and  ( new_n1600_, new_n1599_, new_n1584_ );
or   ( new_n1601_, new_n1600_, new_n1526_ );
and  ( new_n1602_, new_n1601_, new_n1581_ );
or   ( new_n1603_, new_n1602_, new_n1515_ );
and  ( new_n1604_, new_n1603_, new_n1578_ );
or   ( new_n1605_, new_n1604_, new_n1504_ );
and  ( new_n1606_, new_n1605_, new_n1575_ );
or   ( new_n1607_, new_n1606_, new_n1493_ );
and  ( new_n1608_, new_n1607_, new_n1572_ );
or   ( new_n1609_, new_n1608_, new_n1482_ );
and  ( new_n1610_, new_n1471_, new_n1466_ );
and  ( new_n1611_, new_n1470_, new_n74_ );
or   ( new_n1612_, new_n1611_, new_n1610_ );
and  ( new_n1613_, new_n1612_, new_n1609_ );
not  ( new_n1614_, new_n211_ );
and  ( new_n1615_, \I[0] , \A[1][7]  );
and  ( new_n1616_, \I[1] , \A[2][7]  );
nor  ( new_n1617_, new_n1616_, new_n1615_ );
and  ( new_n1618_, new_n1617_, new_n1614_ );
not  ( new_n1619_, new_n1618_ );
and  ( new_n1620_, new_n1619_, \B[7]  );
not  ( new_n1621_, new_n171_ );
and  ( new_n1622_, \I[1] , \A[2][5]  );
and  ( new_n1623_, \I[0] , \A[1][5]  );
nor  ( new_n1624_, new_n1623_, new_n1622_ );
and  ( new_n1625_, new_n1624_, new_n1621_ );
not  ( new_n1626_, new_n1625_ );
and  ( new_n1627_, new_n1626_, \B[9]  );
nor  ( new_n1628_, new_n1627_, new_n1620_ );
and  ( new_n1629_, new_n1626_, \B[8]  );
not  ( new_n1630_, new_n151_ );
and  ( new_n1631_, \I[1] , \A[2][4]  );
and  ( new_n1632_, \I[0] , \A[1][4]  );
nor  ( new_n1633_, new_n1632_, new_n1631_ );
and  ( new_n1634_, new_n1633_, new_n1630_ );
not  ( new_n1635_, new_n1634_ );
and  ( new_n1636_, new_n1635_, \B[9]  );
nor  ( new_n1637_, new_n1636_, new_n1629_ );
and  ( new_n1638_, new_n1619_, \B[6]  );
not  ( new_n1639_, new_n1638_ );
xor  ( new_n1640_, new_n1636_, new_n1629_ );
and  ( new_n1641_, new_n1640_, new_n1639_ );
nor  ( new_n1642_, new_n1641_, new_n1637_ );
not  ( new_n1643_, new_n1642_ );
xor  ( new_n1644_, new_n1627_, new_n1620_ );
and  ( new_n1645_, new_n1644_, new_n1643_ );
or   ( new_n1646_, new_n1645_, new_n1628_ );
not  ( new_n1647_, new_n191_ );
and  ( new_n1648_, \I[1] , \A[2][6]  );
and  ( new_n1649_, \I[0] , \A[1][6]  );
nor  ( new_n1650_, new_n1649_, new_n1648_ );
and  ( new_n1651_, new_n1650_, new_n1647_ );
or   ( new_n1652_, new_n1651_, new_n50_ );
not  ( new_n1653_, new_n65_ );
and  ( new_n1654_, \I[1] , \A[2][8]  );
and  ( new_n1655_, \I[0] , \A[1][8]  );
nor  ( new_n1656_, new_n1655_, new_n1654_ );
and  ( new_n1657_, new_n1656_, new_n1653_ );
not  ( new_n1658_, new_n1657_ );
and  ( new_n1659_, new_n1658_, \B[7]  );
not  ( new_n1660_, new_n78_ );
and  ( new_n1661_, \I[1] , \A[2][9]  );
and  ( new_n1662_, \I[0] , \A[1][9]  );
nor  ( new_n1663_, new_n1662_, new_n1661_ );
and  ( new_n1664_, new_n1663_, new_n1660_ );
not  ( new_n1665_, new_n1664_ );
and  ( new_n1666_, new_n1665_, \B[6]  );
xor  ( new_n1667_, new_n1666_, new_n1659_ );
xor  ( new_n1668_, new_n1667_, new_n1652_ );
and  ( new_n1669_, new_n1619_, \B[8]  );
not  ( new_n1670_, new_n1651_ );
and  ( new_n1671_, new_n1670_, \B[8]  );
and  ( new_n1672_, new_n1665_, \B[5]  );
or   ( new_n1673_, new_n1672_, new_n1671_ );
or   ( new_n1674_, new_n1657_, new_n923_ );
xor  ( new_n1675_, new_n1672_, new_n1671_ );
nand ( new_n1676_, new_n1675_, new_n1674_ );
and  ( new_n1677_, new_n1676_, new_n1673_ );
xor  ( new_n1678_, new_n1677_, new_n1669_ );
xor  ( new_n1679_, new_n1678_, new_n1668_ );
and  ( new_n1680_, new_n1679_, new_n1646_ );
xor  ( new_n1681_, new_n1679_, new_n1646_ );
and  ( new_n1682_, new_n1658_, \B[5]  );
and  ( new_n1683_, new_n1665_, \B[4]  );
nor  ( new_n1684_, new_n1683_, new_n1682_ );
and  ( new_n1685_, new_n1670_, \B[7]  );
xnor ( new_n1686_, new_n1683_, new_n1682_ );
nor  ( new_n1687_, new_n1686_, new_n1685_ );
or   ( new_n1688_, new_n1687_, new_n1684_ );
xor  ( new_n1689_, new_n1675_, new_n1674_ );
or   ( new_n1690_, new_n1689_, new_n1688_ );
and  ( new_n1691_, new_n1689_, new_n1688_ );
xor  ( new_n1692_, new_n1644_, new_n1643_ );
or   ( new_n1693_, new_n1692_, new_n1691_ );
and  ( new_n1694_, new_n1693_, new_n1690_ );
and  ( new_n1695_, new_n1694_, new_n1681_ );
or   ( new_n1696_, new_n1695_, new_n1680_ );
nor  ( new_n1697_, new_n1677_, new_n1669_ );
and  ( new_n1698_, new_n1678_, new_n1668_ );
or   ( new_n1699_, new_n1698_, new_n1697_ );
nor  ( new_n1700_, new_n1666_, new_n1659_ );
and  ( new_n1701_, new_n1667_, new_n1652_ );
or   ( new_n1702_, new_n1701_, new_n1700_ );
or   ( new_n1703_, new_n1657_, new_n1253_ );
and  ( new_n1704_, new_n1619_, \B[9]  );
and  ( new_n1705_, new_n1665_, \B[7]  );
xor  ( new_n1706_, new_n1705_, new_n1704_ );
xor  ( new_n1707_, new_n1706_, new_n1703_ );
xor  ( new_n1708_, new_n1707_, new_n1702_ );
xor  ( new_n1709_, new_n1708_, new_n1699_ );
nor  ( new_n1710_, new_n1709_, new_n1696_ );
and  ( new_n1711_, new_n1709_, new_n1696_ );
xor  ( new_n1712_, new_n1689_, new_n1688_ );
xnor ( new_n1713_, new_n1712_, new_n1692_ );
xnor ( new_n1714_, new_n1686_, new_n1685_ );
and  ( new_n1715_, new_n1635_, \B[8]  );
and  ( new_n1716_, new_n1619_, \B[5]  );
nor  ( new_n1717_, new_n1716_, new_n1715_ );
and  ( new_n1718_, new_n1626_, \B[7]  );
and  ( new_n1719_, new_n1635_, \B[5]  );
and  ( new_n1720_, new_n1719_, new_n1669_ );
nor  ( new_n1721_, new_n1720_, new_n1718_ );
nor  ( new_n1722_, new_n1721_, new_n1717_ );
or   ( new_n1723_, new_n1722_, new_n1714_ );
and  ( new_n1724_, new_n1722_, new_n1714_ );
and  ( new_n1725_, new_n1658_, \B[4]  );
and  ( new_n1726_, new_n1665_, \B[3]  );
nor  ( new_n1727_, new_n1726_, new_n1725_ );
and  ( new_n1728_, new_n1670_, \B[6]  );
and  ( new_n1729_, new_n1726_, new_n1725_ );
nor  ( new_n1730_, new_n1729_, new_n1728_ );
nor  ( new_n1731_, new_n1730_, new_n1727_ );
or   ( new_n1732_, new_n1731_, new_n1724_ );
and  ( new_n1733_, new_n1732_, new_n1723_ );
and  ( new_n1734_, new_n1733_, new_n1713_ );
xnor ( new_n1735_, new_n1733_, new_n1713_ );
xor  ( new_n1736_, new_n1640_, new_n1639_ );
xnor ( new_n1737_, new_n1722_, new_n1714_ );
xor  ( new_n1738_, new_n1737_, new_n1731_ );
or   ( new_n1739_, new_n1738_, new_n1736_ );
nand ( new_n1740_, new_n1738_, new_n1736_ );
not  ( new_n1741_, new_n101_ );
and  ( new_n1742_, \I[0] , \A[1][3]  );
and  ( new_n1743_, \I[1] , \A[2][3]  );
nor  ( new_n1744_, new_n1743_, new_n1742_ );
and  ( new_n1745_, new_n1744_, new_n1741_ );
not  ( new_n1746_, new_n1745_ );
and  ( new_n1747_, new_n1746_, \B[9]  );
and  ( new_n1748_, new_n1670_, \B[5]  );
and  ( new_n1749_, new_n1658_, \B[3]  );
or   ( new_n1750_, new_n1749_, new_n1748_ );
and  ( new_n1751_, new_n1665_, \B[2]  );
xnor ( new_n1752_, new_n1749_, new_n1748_ );
or   ( new_n1753_, new_n1752_, new_n1751_ );
and  ( new_n1754_, new_n1753_, new_n1750_ );
nor  ( new_n1755_, new_n1754_, new_n1747_ );
and  ( new_n1756_, new_n1626_, \B[6]  );
not  ( new_n1757_, new_n92_ );
and  ( new_n1758_, \I[1] , \A[2][2]  );
and  ( new_n1759_, \I[0] , \A[1][2]  );
nor  ( new_n1760_, new_n1759_, new_n1758_ );
and  ( new_n1761_, new_n1760_, new_n1757_ );
not  ( new_n1762_, new_n1761_ );
and  ( new_n1763_, new_n1762_, \B[9]  );
nor  ( new_n1764_, new_n1763_, new_n1756_ );
or   ( new_n1765_, new_n1618_, new_n589_ );
xor  ( new_n1766_, new_n1763_, new_n1756_ );
and  ( new_n1767_, new_n1766_, new_n1765_ );
nor  ( new_n1768_, new_n1767_, new_n1764_ );
xnor ( new_n1769_, new_n1754_, new_n1747_ );
nor  ( new_n1770_, new_n1769_, new_n1768_ );
nor  ( new_n1771_, new_n1770_, new_n1755_ );
nand ( new_n1772_, new_n1771_, new_n1740_ );
and  ( new_n1773_, new_n1772_, new_n1739_ );
nor  ( new_n1774_, new_n1773_, new_n1735_ );
nor  ( new_n1775_, new_n1774_, new_n1734_ );
xor  ( new_n1776_, new_n1694_, new_n1681_ );
nor  ( new_n1777_, new_n1776_, new_n1775_ );
and  ( new_n1778_, new_n1776_, new_n1775_ );
xor  ( new_n1779_, new_n1773_, new_n1735_ );
and  ( new_n1780_, new_n1746_, \B[8]  );
and  ( new_n1781_, new_n1635_, \B[7]  );
or   ( new_n1782_, new_n1781_, new_n1780_ );
xnor ( new_n1783_, new_n1781_, new_n1780_ );
and  ( new_n1784_, new_n1665_, \B[1]  );
and  ( new_n1785_, new_n1658_, \B[2]  );
and  ( new_n1786_, new_n1785_, new_n1784_ );
or   ( new_n1787_, new_n1786_, new_n1783_ );
and  ( new_n1788_, new_n1787_, new_n1782_ );
xnor ( new_n1789_, new_n1726_, new_n1725_ );
xor  ( new_n1790_, new_n1789_, new_n1728_ );
nor  ( new_n1791_, new_n1720_, new_n1717_ );
xnor ( new_n1792_, new_n1791_, new_n1718_ );
nand ( new_n1793_, new_n1792_, new_n1790_ );
and  ( new_n1794_, new_n1793_, new_n1788_ );
nor  ( new_n1795_, new_n1792_, new_n1790_ );
or   ( new_n1796_, new_n1795_, new_n1794_ );
xor  ( new_n1797_, new_n1738_, new_n1736_ );
xor  ( new_n1798_, new_n1797_, new_n1771_ );
or   ( new_n1799_, new_n1798_, new_n1796_ );
xnor ( new_n1800_, new_n1769_, new_n1768_ );
xnor ( new_n1801_, new_n1752_, new_n1751_ );
and  ( new_n1802_, new_n1670_, \B[4]  );
and  ( new_n1803_, new_n1762_, \B[8]  );
or   ( new_n1804_, new_n1803_, new_n1802_ );
not  ( new_n1805_, new_n119_ );
and  ( new_n1806_, \I[0] , \A[1][1]  );
and  ( new_n1807_, \I[1] , \A[2][1]  );
nor  ( new_n1808_, new_n1807_, new_n1806_ );
and  ( new_n1809_, new_n1808_, new_n1805_ );
not  ( new_n1810_, new_n1809_ );
and  ( new_n1811_, new_n1810_, \B[9]  );
and  ( new_n1812_, new_n1803_, new_n1802_ );
or   ( new_n1813_, new_n1812_, new_n1811_ );
and  ( new_n1814_, new_n1813_, new_n1804_ );
or   ( new_n1815_, new_n1814_, new_n1801_ );
and  ( new_n1816_, new_n1814_, new_n1801_ );
and  ( new_n1817_, new_n1635_, \B[6]  );
and  ( new_n1818_, new_n1619_, \B[3]  );
nor  ( new_n1819_, new_n1818_, new_n1817_ );
and  ( new_n1820_, new_n1626_, \B[5]  );
and  ( new_n1821_, new_n1635_, \B[3]  );
and  ( new_n1822_, new_n1821_, new_n1638_ );
nor  ( new_n1823_, new_n1822_, new_n1820_ );
nor  ( new_n1824_, new_n1823_, new_n1819_ );
or   ( new_n1825_, new_n1824_, new_n1816_ );
and  ( new_n1826_, new_n1825_, new_n1815_ );
or   ( new_n1827_, new_n1826_, new_n1800_ );
xor  ( new_n1828_, new_n1766_, new_n1765_ );
xor  ( new_n1829_, new_n1786_, new_n1783_ );
and  ( new_n1830_, new_n1829_, new_n1828_ );
and  ( new_n1831_, new_n1746_, \B[7]  );
and  ( new_n1832_, new_n1658_, \B[1]  );
and  ( new_n1833_, new_n1665_, \B[0]  );
and  ( new_n1834_, new_n1833_, new_n1832_ );
nor  ( new_n1835_, new_n1834_, new_n1831_ );
xnor ( new_n1836_, new_n1834_, new_n1831_ );
xor  ( new_n1837_, new_n1785_, new_n1784_ );
nor  ( new_n1838_, new_n1837_, new_n1836_ );
or   ( new_n1839_, new_n1838_, new_n1835_ );
xor  ( new_n1840_, new_n1829_, new_n1828_ );
and  ( new_n1841_, new_n1840_, new_n1839_ );
nor  ( new_n1842_, new_n1841_, new_n1830_ );
xnor ( new_n1843_, new_n1826_, new_n1800_ );
or   ( new_n1844_, new_n1843_, new_n1842_ );
and  ( new_n1845_, new_n1844_, new_n1827_ );
and  ( new_n1846_, new_n1798_, new_n1796_ );
or   ( new_n1847_, new_n1846_, new_n1845_ );
and  ( new_n1848_, new_n1847_, new_n1799_ );
and  ( new_n1849_, new_n1848_, new_n1779_ );
nor  ( new_n1850_, new_n1848_, new_n1779_ );
xnor ( new_n1851_, new_n1843_, new_n1842_ );
xor  ( new_n1852_, new_n1792_, new_n1790_ );
xor  ( new_n1853_, new_n1852_, new_n1788_ );
or   ( new_n1854_, new_n1853_, new_n1851_ );
and  ( new_n1855_, new_n1853_, new_n1851_ );
and  ( new_n1856_, new_n1626_, \B[4]  );
and  ( new_n1857_, new_n1619_, \B[2]  );
nor  ( new_n1858_, new_n1857_, new_n1856_ );
not  ( new_n1859_, new_n134_ );
and  ( new_n1860_, \I[1] , \A[2][0]  );
and  ( new_n1861_, \I[0] , \A[1][0]  );
nor  ( new_n1862_, new_n1861_, new_n1860_ );
and  ( new_n1863_, new_n1862_, new_n1859_ );
or   ( new_n1864_, new_n1863_, new_n50_ );
xor  ( new_n1865_, new_n1857_, new_n1856_ );
and  ( new_n1866_, new_n1865_, new_n1864_ );
nor  ( new_n1867_, new_n1866_, new_n1858_ );
nor  ( new_n1868_, new_n1822_, new_n1819_ );
xor  ( new_n1869_, new_n1868_, new_n1820_ );
nor  ( new_n1870_, new_n1869_, new_n1867_ );
xnor ( new_n1871_, new_n1869_, new_n1867_ );
and  ( new_n1872_, new_n1670_, \B[3]  );
and  ( new_n1873_, new_n1762_, \B[7]  );
or   ( new_n1874_, new_n1873_, new_n1872_ );
and  ( new_n1875_, new_n1810_, \B[8]  );
and  ( new_n1876_, new_n1873_, new_n1872_ );
or   ( new_n1877_, new_n1876_, new_n1875_ );
and  ( new_n1878_, new_n1877_, new_n1874_ );
nor  ( new_n1879_, new_n1878_, new_n1871_ );
or   ( new_n1880_, new_n1879_, new_n1870_ );
xnor ( new_n1881_, new_n1814_, new_n1801_ );
xor  ( new_n1882_, new_n1881_, new_n1824_ );
and  ( new_n1883_, new_n1882_, new_n1880_ );
and  ( new_n1884_, new_n1746_, \B[6]  );
nor  ( new_n1885_, new_n1884_, new_n1719_ );
xor  ( new_n1886_, new_n1884_, new_n1719_ );
not  ( new_n1887_, new_n1886_ );
xor  ( new_n1888_, new_n1833_, new_n1832_ );
nor  ( new_n1889_, new_n1888_, new_n1887_ );
or   ( new_n1890_, new_n1889_, new_n1885_ );
xnor ( new_n1891_, new_n1803_, new_n1802_ );
xor  ( new_n1892_, new_n1891_, new_n1811_ );
and  ( new_n1893_, new_n1892_, new_n1890_ );
and  ( new_n1894_, new_n1635_, \B[4]  );
and  ( new_n1895_, new_n1670_, \B[2]  );
nor  ( new_n1896_, new_n1895_, new_n1894_ );
and  ( new_n1897_, new_n1746_, \B[5]  );
and  ( new_n1898_, new_n1895_, new_n1894_ );
nor  ( new_n1899_, new_n1898_, new_n1897_ );
nor  ( new_n1900_, new_n1899_, new_n1896_ );
and  ( new_n1901_, new_n1619_, \B[0]  );
and  ( new_n1902_, new_n1901_, new_n1832_ );
nor  ( new_n1903_, new_n1902_, new_n1900_ );
xnor ( new_n1904_, new_n1902_, new_n1900_ );
and  ( new_n1905_, new_n1626_, \B[3]  );
and  ( new_n1906_, new_n1810_, \B[7]  );
or   ( new_n1907_, new_n1906_, new_n1905_ );
not  ( new_n1908_, new_n1863_ );
and  ( new_n1909_, new_n1908_, \B[8]  );
and  ( new_n1910_, new_n1906_, new_n1905_ );
or   ( new_n1911_, new_n1910_, new_n1909_ );
and  ( new_n1912_, new_n1911_, new_n1907_ );
nor  ( new_n1913_, new_n1912_, new_n1904_ );
or   ( new_n1914_, new_n1913_, new_n1903_ );
xor  ( new_n1915_, new_n1892_, new_n1890_ );
and  ( new_n1916_, new_n1915_, new_n1914_ );
or   ( new_n1917_, new_n1916_, new_n1893_ );
xor  ( new_n1918_, new_n1882_, new_n1880_ );
and  ( new_n1919_, new_n1918_, new_n1917_ );
nor  ( new_n1920_, new_n1919_, new_n1883_ );
or   ( new_n1921_, new_n1920_, new_n1855_ );
and  ( new_n1922_, new_n1921_, new_n1854_ );
xor  ( new_n1923_, new_n1798_, new_n1796_ );
xor  ( new_n1924_, new_n1923_, new_n1845_ );
and  ( new_n1925_, new_n1924_, new_n1922_ );
nor  ( new_n1926_, new_n1924_, new_n1922_ );
xor  ( new_n1927_, new_n1837_, new_n1836_ );
xor  ( new_n1928_, new_n1878_, new_n1871_ );
and  ( new_n1929_, new_n1928_, new_n1927_ );
and  ( new_n1930_, new_n1762_, \B[6]  );
or   ( new_n1931_, new_n1657_, new_n98_ );
or   ( new_n1932_, new_n1618_, new_n88_ );
and  ( new_n1933_, new_n1932_, new_n1931_ );
nor  ( new_n1934_, new_n1933_, new_n1902_ );
and  ( new_n1935_, new_n1934_, new_n1930_ );
xor  ( new_n1936_, new_n1934_, new_n1930_ );
and  ( new_n1937_, new_n1670_, \B[1]  );
and  ( new_n1938_, new_n1937_, new_n1901_ );
and  ( new_n1939_, new_n1938_, new_n1936_ );
nor  ( new_n1940_, new_n1939_, new_n1935_ );
xor  ( new_n1941_, new_n1865_, new_n1864_ );
xnor ( new_n1942_, new_n1873_, new_n1872_ );
xor  ( new_n1943_, new_n1942_, new_n1875_ );
and  ( new_n1944_, new_n1943_, new_n1941_ );
nor  ( new_n1945_, new_n1944_, new_n1940_ );
nor  ( new_n1946_, new_n1943_, new_n1941_ );
nor  ( new_n1947_, new_n1946_, new_n1945_ );
xor  ( new_n1948_, new_n1928_, new_n1927_ );
and  ( new_n1949_, new_n1948_, new_n1947_ );
nor  ( new_n1950_, new_n1949_, new_n1929_ );
not  ( new_n1951_, new_n1950_ );
xor  ( new_n1952_, new_n1840_, new_n1839_ );
and  ( new_n1953_, new_n1952_, new_n1951_ );
xor  ( new_n1954_, new_n1952_, new_n1951_ );
xor  ( new_n1955_, new_n1918_, new_n1917_ );
and  ( new_n1956_, new_n1955_, new_n1954_ );
or   ( new_n1957_, new_n1956_, new_n1953_ );
xnor ( new_n1958_, new_n1853_, new_n1851_ );
xor  ( new_n1959_, new_n1958_, new_n1920_ );
nor  ( new_n1960_, new_n1959_, new_n1957_ );
and  ( new_n1961_, new_n1959_, new_n1957_ );
xnor ( new_n1962_, new_n1955_, new_n1954_ );
xor  ( new_n1963_, new_n1888_, new_n1887_ );
xor  ( new_n1964_, new_n1912_, new_n1904_ );
and  ( new_n1965_, new_n1964_, new_n1963_ );
xor  ( new_n1966_, new_n1964_, new_n1963_ );
and  ( new_n1967_, new_n1908_, \B[7]  );
or   ( new_n1968_, new_n1967_, new_n1821_ );
and  ( new_n1969_, new_n1746_, \B[4]  );
and  ( new_n1970_, new_n1967_, new_n1821_ );
or   ( new_n1971_, new_n1970_, new_n1969_ );
and  ( new_n1972_, new_n1971_, new_n1968_ );
and  ( new_n1973_, new_n1626_, \B[2]  );
and  ( new_n1974_, new_n1810_, \B[6]  );
nor  ( new_n1975_, new_n1974_, new_n1973_ );
and  ( new_n1976_, new_n1762_, \B[5]  );
and  ( new_n1977_, new_n1810_, \B[2]  );
and  ( new_n1978_, new_n1977_, new_n1756_ );
nor  ( new_n1979_, new_n1978_, new_n1976_ );
nor  ( new_n1980_, new_n1979_, new_n1975_ );
nand ( new_n1981_, new_n1980_, new_n1972_ );
nor  ( new_n1982_, new_n1980_, new_n1972_ );
xor  ( new_n1983_, new_n1895_, new_n1894_ );
xnor ( new_n1984_, new_n1983_, new_n1897_ );
or   ( new_n1985_, new_n1984_, new_n1982_ );
and  ( new_n1986_, new_n1985_, new_n1981_ );
and  ( new_n1987_, new_n1986_, new_n1966_ );
or   ( new_n1988_, new_n1987_, new_n1965_ );
xor  ( new_n1989_, new_n1915_, new_n1914_ );
nand ( new_n1990_, new_n1989_, new_n1988_ );
xor  ( new_n1991_, new_n1948_, new_n1947_ );
or   ( new_n1992_, new_n1989_, new_n1988_ );
nand ( new_n1993_, new_n1992_, new_n1991_ );
and  ( new_n1994_, new_n1993_, new_n1990_ );
and  ( new_n1995_, new_n1994_, new_n1962_ );
nor  ( new_n1996_, new_n1994_, new_n1962_ );
xor  ( new_n1997_, new_n1989_, new_n1988_ );
xor  ( new_n1998_, new_n1997_, new_n1991_ );
not  ( new_n1999_, new_n1938_ );
xor  ( new_n2000_, new_n1999_, new_n1936_ );
xnor ( new_n2001_, new_n1906_, new_n1905_ );
xor  ( new_n2002_, new_n2001_, new_n1909_ );
or   ( new_n2003_, new_n2002_, new_n2000_ );
and  ( new_n2004_, new_n1670_, \B[0]  );
and  ( new_n2005_, new_n1626_, \B[1]  );
and  ( new_n2006_, new_n2005_, new_n2004_ );
and  ( new_n2007_, new_n2006_, new_n1999_ );
and  ( new_n2008_, new_n1762_, \B[4]  );
and  ( new_n2009_, new_n1746_, \B[3]  );
nor  ( new_n2010_, new_n2009_, new_n2008_ );
and  ( new_n2011_, new_n1635_, \B[2]  );
and  ( new_n2012_, new_n2009_, new_n2008_ );
nor  ( new_n2013_, new_n2012_, new_n2011_ );
nor  ( new_n2014_, new_n2013_, new_n2010_ );
or   ( new_n2015_, new_n2006_, new_n1999_ );
nor  ( new_n2016_, new_n1937_, new_n1901_ );
nor  ( new_n2017_, new_n2016_, new_n2007_ );
and  ( new_n2018_, new_n2017_, new_n2015_ );
and  ( new_n2019_, new_n2018_, new_n2014_ );
or   ( new_n2020_, new_n2019_, new_n2007_ );
xor  ( new_n2021_, new_n2002_, new_n2000_ );
nand ( new_n2022_, new_n2021_, new_n2020_ );
and  ( new_n2023_, new_n2022_, new_n2003_ );
xor  ( new_n2024_, new_n1943_, new_n1941_ );
xor  ( new_n2025_, new_n2024_, new_n1940_ );
or   ( new_n2026_, new_n2025_, new_n2023_ );
and  ( new_n2027_, new_n2025_, new_n2023_ );
xor  ( new_n2028_, new_n1986_, new_n1966_ );
or   ( new_n2029_, new_n2028_, new_n2027_ );
and  ( new_n2030_, new_n2029_, new_n2026_ );
nor  ( new_n2031_, new_n2030_, new_n1998_ );
and  ( new_n2032_, new_n2030_, new_n1998_ );
nor  ( new_n2033_, new_n1978_, new_n1975_ );
xnor ( new_n2034_, new_n2033_, new_n1976_ );
xnor ( new_n2035_, new_n1967_, new_n1821_ );
xor  ( new_n2036_, new_n2035_, new_n1969_ );
and  ( new_n2037_, new_n2036_, new_n2034_ );
and  ( new_n2038_, new_n1810_, \B[5]  );
and  ( new_n2039_, new_n1908_, \B[6]  );
nor  ( new_n2040_, new_n2039_, new_n2038_ );
and  ( new_n2041_, new_n1626_, \B[0]  );
and  ( new_n2042_, new_n1635_, \B[1]  );
and  ( new_n2043_, new_n2042_, new_n2041_ );
and  ( new_n2044_, new_n2039_, new_n2038_ );
nor  ( new_n2045_, new_n2044_, new_n2043_ );
nor  ( new_n2046_, new_n2045_, new_n2040_ );
not  ( new_n2047_, new_n2046_ );
nor  ( new_n2048_, new_n2047_, new_n2037_ );
nor  ( new_n2049_, new_n2036_, new_n2034_ );
nor  ( new_n2050_, new_n2049_, new_n2048_ );
not  ( new_n2051_, new_n2050_ );
xnor ( new_n2052_, new_n1980_, new_n1972_ );
xor  ( new_n2053_, new_n2052_, new_n1984_ );
and  ( new_n2054_, new_n2053_, new_n2051_ );
xor  ( new_n2055_, new_n2053_, new_n2051_ );
xor  ( new_n2056_, new_n2021_, new_n2020_ );
and  ( new_n2057_, new_n2056_, new_n2055_ );
or   ( new_n2058_, new_n2057_, new_n2054_ );
xnor ( new_n2059_, new_n2025_, new_n2023_ );
xor  ( new_n2060_, new_n2059_, new_n2028_ );
nor  ( new_n2061_, new_n2060_, new_n2058_ );
and  ( new_n2062_, new_n2060_, new_n2058_ );
xnor ( new_n2063_, new_n2056_, new_n2055_ );
xnor ( new_n2064_, new_n2018_, new_n2014_ );
xor  ( new_n2065_, new_n2036_, new_n2034_ );
xor  ( new_n2066_, new_n2065_, new_n2047_ );
or   ( new_n2067_, new_n2066_, new_n2064_ );
nand ( new_n2068_, new_n2066_, new_n2064_ );
and  ( new_n2069_, new_n1810_, \B[4]  );
and  ( new_n2070_, new_n1746_, \B[2]  );
or   ( new_n2071_, new_n2070_, new_n2069_ );
or   ( new_n2072_, new_n1761_, new_n422_ );
xor  ( new_n2073_, new_n2070_, new_n2069_ );
nand ( new_n2074_, new_n2073_, new_n2072_ );
and  ( new_n2075_, new_n2074_, new_n2071_ );
xor  ( new_n2076_, new_n2005_, new_n2004_ );
nor  ( new_n2077_, new_n2076_, new_n2075_ );
xor  ( new_n2078_, new_n2076_, new_n2075_ );
xnor ( new_n2079_, new_n2009_, new_n2008_ );
xor  ( new_n2080_, new_n2079_, new_n2011_ );
and  ( new_n2081_, new_n2080_, new_n2078_ );
nor  ( new_n2082_, new_n2081_, new_n2077_ );
nand ( new_n2083_, new_n2082_, new_n2068_ );
and  ( new_n2084_, new_n2083_, new_n2067_ );
nor  ( new_n2085_, new_n2084_, new_n2063_ );
and  ( new_n2086_, new_n2084_, new_n2063_ );
and  ( new_n2087_, new_n1908_, \B[5]  );
and  ( new_n2088_, new_n1635_, \B[0]  );
and  ( new_n2089_, new_n1746_, \B[1]  );
and  ( new_n2090_, new_n2089_, new_n2088_ );
nor  ( new_n2091_, new_n2090_, new_n2087_ );
not  ( new_n2092_, new_n2090_ );
xor  ( new_n2093_, new_n2092_, new_n2087_ );
xor  ( new_n2094_, new_n2042_, new_n2041_ );
nor  ( new_n2095_, new_n2094_, new_n2093_ );
or   ( new_n2096_, new_n2095_, new_n2091_ );
xnor ( new_n2097_, new_n2039_, new_n2038_ );
xor  ( new_n2098_, new_n2097_, new_n2043_ );
nand ( new_n2099_, new_n2098_, new_n2096_ );
xor  ( new_n2100_, new_n2098_, new_n2096_ );
xor  ( new_n2101_, new_n2080_, new_n2078_ );
nand ( new_n2102_, new_n2101_, new_n2100_ );
and  ( new_n2103_, new_n2102_, new_n2099_ );
xor  ( new_n2104_, new_n2066_, new_n2064_ );
xor  ( new_n2105_, new_n2104_, new_n2082_ );
and  ( new_n2106_, new_n2105_, new_n2103_ );
nor  ( new_n2107_, new_n2105_, new_n2103_ );
and  ( new_n2108_, new_n1908_, \B[4]  );
and  ( new_n2109_, new_n1762_, \B[2]  );
nor  ( new_n2110_, new_n2109_, new_n2108_ );
or   ( new_n2111_, new_n1809_, new_n422_ );
xor  ( new_n2112_, new_n2109_, new_n2108_ );
and  ( new_n2113_, new_n2112_, new_n2111_ );
or   ( new_n2114_, new_n2113_, new_n2110_ );
xor  ( new_n2115_, new_n2073_, new_n2072_ );
and  ( new_n2116_, new_n2115_, new_n2114_ );
xor  ( new_n2117_, new_n2115_, new_n2114_ );
xor  ( new_n2118_, new_n2094_, new_n2093_ );
and  ( new_n2119_, new_n2118_, new_n2117_ );
or   ( new_n2120_, new_n2119_, new_n2116_ );
xor  ( new_n2121_, new_n2101_, new_n2100_ );
nor  ( new_n2122_, new_n2121_, new_n2120_ );
and  ( new_n2123_, new_n2121_, new_n2120_ );
xor  ( new_n2124_, new_n2089_, new_n2088_ );
and  ( new_n2125_, new_n1746_, \B[0]  );
and  ( new_n2126_, new_n1762_, \B[1]  );
and  ( new_n2127_, new_n2126_, new_n2125_ );
nor  ( new_n2128_, new_n2127_, new_n2124_ );
and  ( new_n2129_, new_n2127_, new_n2092_ );
nor  ( new_n2130_, new_n2129_, new_n2128_ );
xor  ( new_n2131_, new_n2112_, new_n2111_ );
and  ( new_n2132_, new_n2131_, new_n2130_ );
or   ( new_n2133_, new_n2132_, new_n2128_ );
xor  ( new_n2134_, new_n2118_, new_n2117_ );
nor  ( new_n2135_, new_n2134_, new_n2133_ );
and  ( new_n2136_, new_n2134_, new_n2133_ );
xnor ( new_n2137_, new_n2131_, new_n2130_ );
and  ( new_n2138_, new_n1908_, \B[3]  );
nor  ( new_n2139_, new_n2138_, new_n1977_ );
xor  ( new_n2140_, new_n2126_, new_n2125_ );
and  ( new_n2141_, new_n2138_, new_n1977_ );
nor  ( new_n2142_, new_n2141_, new_n2140_ );
nor  ( new_n2143_, new_n2142_, new_n2139_ );
and  ( new_n2144_, new_n2143_, new_n2137_ );
nor  ( new_n2145_, new_n2143_, new_n2137_ );
xnor ( new_n2146_, new_n2138_, new_n1977_ );
and  ( new_n2147_, new_n2146_, new_n2140_ );
not  ( new_n2148_, new_n2139_ );
and  ( new_n2149_, new_n2142_, new_n2148_ );
or   ( new_n2150_, new_n2149_, new_n2147_ );
and  ( new_n2151_, new_n1908_, \B[2]  );
and  ( new_n2152_, new_n1762_, \B[0]  );
and  ( new_n2153_, new_n2152_, new_n2151_ );
and  ( new_n2154_, new_n2153_, new_n2150_ );
nor  ( new_n2155_, new_n2153_, new_n2150_ );
and  ( new_n2156_, new_n1810_, \B[1]  );
not  ( new_n2157_, new_n2156_ );
and  ( new_n2158_, new_n1908_, \B[0]  );
not  ( new_n2159_, new_n2158_ );
nor  ( new_n2160_, new_n2152_, new_n2151_ );
and  ( new_n2161_, new_n2160_, new_n2159_ );
nor  ( new_n2162_, new_n2161_, new_n2157_ );
not  ( new_n2163_, new_n2162_ );
nor  ( new_n2164_, new_n2163_, new_n2155_ );
nor  ( new_n2165_, new_n2164_, new_n2154_ );
nor  ( new_n2166_, new_n2165_, new_n2145_ );
nor  ( new_n2167_, new_n2166_, new_n2144_ );
nor  ( new_n2168_, new_n2167_, new_n2136_ );
nor  ( new_n2169_, new_n2168_, new_n2135_ );
nor  ( new_n2170_, new_n2169_, new_n2123_ );
nor  ( new_n2171_, new_n2170_, new_n2122_ );
nor  ( new_n2172_, new_n2171_, new_n2107_ );
nor  ( new_n2173_, new_n2172_, new_n2106_ );
nor  ( new_n2174_, new_n2173_, new_n2086_ );
nor  ( new_n2175_, new_n2174_, new_n2085_ );
not  ( new_n2176_, new_n2175_ );
nor  ( new_n2177_, new_n2176_, new_n2062_ );
nor  ( new_n2178_, new_n2177_, new_n2061_ );
not  ( new_n2179_, new_n2178_ );
nor  ( new_n2180_, new_n2179_, new_n2032_ );
nor  ( new_n2181_, new_n2180_, new_n2031_ );
nor  ( new_n2182_, new_n2181_, new_n1996_ );
nor  ( new_n2183_, new_n2182_, new_n1995_ );
nor  ( new_n2184_, new_n2183_, new_n1961_ );
nor  ( new_n2185_, new_n2184_, new_n1960_ );
nor  ( new_n2186_, new_n2185_, new_n1926_ );
nor  ( new_n2187_, new_n2186_, new_n1925_ );
nor  ( new_n2188_, new_n2187_, new_n1850_ );
nor  ( new_n2189_, new_n2188_, new_n1849_ );
nor  ( new_n2190_, new_n2189_, new_n1778_ );
nor  ( new_n2191_, new_n2190_, new_n1777_ );
nor  ( new_n2192_, new_n2191_, new_n1711_ );
nor  ( new_n2193_, new_n2192_, new_n1710_ );
and  ( new_n2194_, new_n1707_, new_n1702_ );
and  ( new_n2195_, new_n1708_, new_n1699_ );
or   ( new_n2196_, new_n2195_, new_n2194_ );
nor  ( new_n2197_, new_n1705_, new_n1704_ );
and  ( new_n2198_, new_n1706_, new_n1703_ );
or   ( new_n2199_, new_n2198_, new_n2197_ );
and  ( new_n2200_, new_n1665_, \B[8]  );
and  ( new_n2201_, new_n1658_, \B[9]  );
xor  ( new_n2202_, new_n2201_, new_n2200_ );
xor  ( new_n2203_, new_n2202_, new_n2199_ );
xnor ( new_n2204_, new_n2203_, new_n2196_ );
xor  ( new_n2205_, new_n2204_, new_n2193_ );
or   ( new_n2206_, new_n2205_, new_n1613_ );
or   ( new_n2207_, new_n2206_, new_n1569_ );
and  ( new_n2208_, new_n1612_, new_n1568_ );
and  ( new_n2209_, new_n1609_, new_n1473_ );
not  ( new_n2210_, new_n2209_ );
nand ( new_n2211_, new_n2210_, new_n2205_ );
or   ( new_n2212_, new_n2211_, new_n2208_ );
and  ( new_n2213_, new_n2212_, new_n2207_ );
or   ( new_n2214_, new_n1468_, new_n1462_ );
and  ( new_n2215_, new_n294_, \B[9]  );
and  ( new_n2216_, new_n2215_, new_n2214_ );
or   ( new_n2217_, new_n83_, new_n50_ );
or   ( new_n2218_, new_n1305_, new_n1254_ );
or   ( new_n2219_, new_n1464_, new_n1415_ );
and  ( new_n2220_, new_n2219_, new_n2218_ );
and  ( new_n2221_, new_n2220_, new_n2217_ );
or   ( new_n2222_, new_n2221_, new_n2216_ );
or   ( new_n2223_, new_n1470_, new_n74_ );
or   ( new_n2224_, new_n1612_, new_n1568_ );
and  ( new_n2225_, new_n2224_, new_n2223_ );
or   ( new_n2226_, new_n2225_, new_n2222_ );
and  ( new_n2227_, new_n1665_, \B[9]  );
or   ( new_n2228_, new_n2201_, new_n2200_ );
nand ( new_n2229_, new_n2202_, new_n2199_ );
and  ( new_n2230_, new_n2229_, new_n2228_ );
and  ( new_n2231_, new_n2230_, new_n2227_ );
nor  ( new_n2232_, new_n2230_, new_n2227_ );
nor  ( new_n2233_, new_n2203_, new_n2196_ );
and  ( new_n2234_, new_n2203_, new_n2196_ );
nor  ( new_n2235_, new_n2234_, new_n2193_ );
nor  ( new_n2236_, new_n2235_, new_n2233_ );
nor  ( new_n2237_, new_n2236_, new_n2232_ );
nor  ( new_n2238_, new_n2237_, new_n2231_ );
nor  ( new_n2239_, new_n2220_, new_n2217_ );
nor  ( new_n2240_, new_n2239_, new_n2238_ );
and  ( new_n2241_, new_n2240_, new_n2226_ );
and  ( new_n2242_, new_n1566_, new_n1484_ );
not  ( new_n2243_, new_n1608_ );
xor  ( new_n2244_, new_n1709_, new_n1696_ );
xnor ( new_n2245_, new_n2244_, new_n2191_ );
nand ( new_n2246_, new_n2245_, new_n2243_ );
or   ( new_n2247_, new_n2246_, new_n2242_ );
and  ( new_n2248_, new_n1607_, new_n1484_ );
and  ( new_n2249_, new_n1572_, new_n1566_ );
or   ( new_n2250_, new_n2249_, new_n2245_ );
or   ( new_n2251_, new_n2250_, new_n2248_ );
and  ( new_n2252_, new_n2251_, new_n2247_ );
not  ( new_n2253_, new_n2189_ );
xor  ( new_n2254_, new_n1776_, new_n1775_ );
not  ( new_n2255_, new_n2254_ );
and  ( new_n2256_, \B[4] , \B[5]  );
and  ( new_n2257_, \B[2] , \B[3]  );
and  ( new_n2258_, new_n2257_, new_n2256_ );
and  ( new_n2259_, \B[8] , \B[9]  );
and  ( new_n2260_, \B[6] , \B[7]  );
and  ( new_n2261_, new_n2260_, new_n2259_ );
and  ( new_n2262_, new_n272_, new_n64_ );
and  ( new_n2263_, new_n2262_, new_n2261_ );
and  ( new_n2264_, new_n2263_, new_n2258_ );
and  ( new_n2265_, new_n2264_, new_n58_ );
nor  ( new_n2266_, new_n2265_, new_n2255_ );
nor  ( new_n2267_, new_n2266_, new_n2253_ );
and  ( new_n2268_, new_n2254_, new_n2253_ );
nor  ( new_n2269_, new_n2268_, new_n2267_ );
and  ( new_n2270_, new_n1575_, new_n1564_ );
and  ( new_n2271_, new_n1605_, new_n1495_ );
nor  ( new_n2272_, new_n2271_, new_n2270_ );
nor  ( new_n2273_, new_n2272_, new_n2269_ );
and  ( new_n2274_, new_n1564_, new_n1495_ );
or   ( new_n2275_, new_n2274_, new_n1606_ );
and  ( new_n2276_, new_n2275_, new_n2269_ );
and  ( new_n2277_, new_n1562_, new_n1506_ );
not  ( new_n2278_, new_n1604_ );
xor  ( new_n2279_, new_n1848_, new_n1779_ );
xnor ( new_n2280_, new_n2279_, new_n2187_ );
nand ( new_n2281_, new_n2280_, new_n2278_ );
or   ( new_n2282_, new_n2281_, new_n2277_ );
and  ( new_n2283_, new_n1603_, new_n1506_ );
and  ( new_n2284_, new_n1578_, new_n1562_ );
or   ( new_n2285_, new_n2284_, new_n2280_ );
or   ( new_n2286_, new_n2285_, new_n2283_ );
and  ( new_n2287_, new_n2286_, new_n2282_ );
and  ( new_n2288_, new_n1560_, new_n1517_ );
not  ( new_n2289_, new_n1602_ );
xor  ( new_n2290_, new_n1924_, new_n1922_ );
xnor ( new_n2291_, new_n2290_, new_n2185_ );
nand ( new_n2292_, new_n2291_, new_n2289_ );
or   ( new_n2293_, new_n2292_, new_n2288_ );
and  ( new_n2294_, new_n1601_, new_n1517_ );
and  ( new_n2295_, new_n1581_, new_n1560_ );
or   ( new_n2296_, new_n2295_, new_n2291_ );
or   ( new_n2297_, new_n2296_, new_n2294_ );
and  ( new_n2298_, new_n2297_, new_n2293_ );
and  ( new_n2299_, new_n1558_, new_n1528_ );
not  ( new_n2300_, new_n1600_ );
xor  ( new_n2301_, new_n1959_, new_n1957_ );
xnor ( new_n2302_, new_n2301_, new_n2183_ );
nand ( new_n2303_, new_n2302_, new_n2300_ );
or   ( new_n2304_, new_n2303_, new_n2299_ );
and  ( new_n2305_, new_n1599_, new_n1528_ );
and  ( new_n2306_, new_n1584_, new_n1558_ );
or   ( new_n2307_, new_n2306_, new_n2302_ );
or   ( new_n2308_, new_n2307_, new_n2305_ );
and  ( new_n2309_, new_n2308_, new_n2304_ );
and  ( new_n2310_, new_n1556_, new_n1539_ );
not  ( new_n2311_, new_n1598_ );
xor  ( new_n2312_, new_n1994_, new_n1962_ );
xnor ( new_n2313_, new_n2312_, new_n2181_ );
nand ( new_n2314_, new_n2313_, new_n2311_ );
or   ( new_n2315_, new_n2314_, new_n2310_ );
and  ( new_n2316_, new_n1597_, new_n1539_ );
and  ( new_n2317_, new_n1587_, new_n1556_ );
or   ( new_n2318_, new_n2317_, new_n2313_ );
or   ( new_n2319_, new_n2318_, new_n2316_ );
and  ( new_n2320_, new_n2319_, new_n2315_ );
and  ( new_n2321_, new_n1592_, new_n1550_ );
xor  ( new_n2322_, new_n2030_, new_n1998_ );
xor  ( new_n2323_, new_n2322_, new_n2179_ );
nand ( new_n2324_, new_n1595_, new_n1554_ );
nand ( new_n2325_, new_n2324_, new_n2323_ );
or   ( new_n2326_, new_n2325_, new_n2321_ );
and  ( new_n2327_, new_n1554_, new_n1550_ );
or   ( new_n2328_, new_n2323_, new_n1596_ );
or   ( new_n2329_, new_n2328_, new_n2327_ );
and  ( new_n2330_, new_n2329_, new_n2326_ );
xor  ( new_n2331_, new_n2060_, new_n2058_ );
xor  ( new_n2332_, new_n2331_, new_n2176_ );
and  ( new_n2333_, new_n1553_, new_n1552_ );
or   ( new_n2334_, new_n2333_, new_n1592_ );
and  ( new_n2335_, new_n2334_, new_n2332_ );
and  ( new_n2336_, new_n1590_, new_n1553_ );
and  ( new_n2337_, new_n1591_, new_n1552_ );
nor  ( new_n2338_, new_n2337_, new_n2336_ );
nor  ( new_n2339_, new_n2338_, new_n2332_ );
and  ( new_n2340_, new_n1440_, new_n1342_ );
and  ( new_n2341_, new_n1441_, new_n1341_ );
xor  ( new_n2342_, new_n2084_, new_n2063_ );
xnor ( new_n2343_, new_n2342_, new_n2173_ );
or   ( new_n2344_, new_n2343_, new_n2341_ );
or   ( new_n2345_, new_n2344_, new_n2340_ );
and  ( new_n2346_, new_n1342_, new_n1341_ );
not  ( new_n2347_, new_n1442_ );
nand ( new_n2348_, new_n2343_, new_n2347_ );
or   ( new_n2349_, new_n2348_, new_n2346_ );
and  ( new_n2350_, new_n2349_, new_n2345_ );
and  ( new_n2351_, new_n1268_, new_n1225_ );
and  ( new_n2352_, new_n1267_, new_n1226_ );
xor  ( new_n2353_, new_n2105_, new_n2103_ );
xnor ( new_n2354_, new_n2353_, new_n2171_ );
or   ( new_n2355_, new_n2354_, new_n2352_ );
or   ( new_n2356_, new_n2355_, new_n2351_ );
and  ( new_n2357_, new_n1268_, new_n1267_ );
not  ( new_n2358_, new_n1227_ );
nand ( new_n2359_, new_n2354_, new_n2358_ );
or   ( new_n2360_, new_n2359_, new_n2357_ );
and  ( new_n2361_, new_n2360_, new_n2356_ );
and  ( new_n2362_, new_n1100_, new_n1061_ );
and  ( new_n2363_, new_n1099_, new_n1062_ );
xor  ( new_n2364_, new_n2121_, new_n2120_ );
xnor ( new_n2365_, new_n2364_, new_n2169_ );
or   ( new_n2366_, new_n2365_, new_n2363_ );
or   ( new_n2367_, new_n2366_, new_n2362_ );
and  ( new_n2368_, new_n1100_, new_n1099_ );
not  ( new_n2369_, new_n1063_ );
nand ( new_n2370_, new_n2365_, new_n2369_ );
or   ( new_n2371_, new_n2370_, new_n2368_ );
and  ( new_n2372_, new_n2371_, new_n2367_ );
xor  ( new_n2373_, new_n2134_, new_n2133_ );
xnor ( new_n2374_, new_n2373_, new_n2167_ );
and  ( new_n2375_, new_n937_, new_n936_ );
or   ( new_n2376_, new_n2375_, new_n896_ );
and  ( new_n2377_, new_n2376_, new_n2374_ );
and  ( new_n2378_, new_n937_, new_n894_ );
and  ( new_n2379_, new_n936_, new_n895_ );
nor  ( new_n2380_, new_n2379_, new_n2378_ );
nor  ( new_n2381_, new_n2380_, new_n2374_ );
and  ( new_n2382_, new_n770_, new_n727_ );
and  ( new_n2383_, new_n769_, new_n728_ );
xor  ( new_n2384_, new_n2143_, new_n2137_ );
xnor ( new_n2385_, new_n2384_, new_n2165_ );
or   ( new_n2386_, new_n2385_, new_n2383_ );
or   ( new_n2387_, new_n2386_, new_n2382_ );
and  ( new_n2388_, new_n770_, new_n769_ );
not  ( new_n2389_, new_n729_ );
nand ( new_n2390_, new_n2385_, new_n2389_ );
or   ( new_n2391_, new_n2390_, new_n2388_ );
and  ( new_n2392_, new_n2391_, new_n2387_ );
and  ( new_n2393_, new_n603_, new_n560_ );
and  ( new_n2394_, new_n602_, new_n561_ );
xor  ( new_n2395_, new_n2153_, new_n2150_ );
xor  ( new_n2396_, new_n2395_, new_n2162_ );
or   ( new_n2397_, new_n2396_, new_n2394_ );
or   ( new_n2398_, new_n2397_, new_n2393_ );
and  ( new_n2399_, new_n603_, new_n602_ );
not  ( new_n2400_, new_n562_ );
nand ( new_n2401_, new_n2396_, new_n2400_ );
or   ( new_n2402_, new_n2401_, new_n2399_ );
and  ( new_n2403_, new_n2402_, new_n2398_ );
and  ( new_n2404_, \B[0] , new_n88_ );
or   ( new_n2405_, new_n2404_, new_n86_ );
or   ( new_n2406_, new_n1810_, new_n270_ );
or   ( new_n2407_, new_n1809_, new_n123_ );
and  ( new_n2408_, new_n2407_, \B[0]  );
and  ( new_n2409_, new_n2408_, new_n2406_ );
and  ( new_n2410_, new_n1908_, new_n139_ );
and  ( new_n2411_, new_n1863_, new_n386_ );
or   ( new_n2412_, new_n2411_, new_n2410_ );
or   ( new_n2413_, new_n2412_, new_n2409_ );
and  ( new_n2414_, new_n2413_, new_n2405_ );
and  ( new_n2415_, new_n435_, new_n385_ );
and  ( new_n2416_, new_n434_, new_n387_ );
and  ( new_n2417_, new_n2159_, new_n2156_ );
xor  ( new_n2418_, new_n2152_, new_n2151_ );
nor  ( new_n2419_, new_n2418_, new_n2417_ );
not  ( new_n2420_, new_n2160_ );
and  ( new_n2421_, new_n2417_, new_n2420_ );
nor  ( new_n2422_, new_n2421_, new_n2419_ );
or   ( new_n2423_, new_n2422_, new_n2416_ );
or   ( new_n2424_, new_n2423_, new_n2415_ );
and  ( new_n2425_, new_n435_, new_n434_ );
not  ( new_n2426_, new_n388_ );
nand ( new_n2427_, new_n2422_, new_n2426_ );
or   ( new_n2428_, new_n2427_, new_n2425_ );
and  ( new_n2429_, new_n2428_, new_n2424_ );
or   ( new_n2430_, new_n2429_, new_n2414_ );
or   ( new_n2431_, new_n2430_, new_n2403_ );
or   ( new_n2432_, new_n2431_, new_n2392_ );
or   ( new_n2433_, new_n2432_, new_n2381_ );
or   ( new_n2434_, new_n2433_, new_n2377_ );
or   ( new_n2435_, new_n2434_, new_n2372_ );
or   ( new_n2436_, new_n2435_, new_n2361_ );
or   ( new_n2437_, new_n2436_, new_n2350_ );
or   ( new_n2438_, new_n2437_, new_n2339_ );
or   ( new_n2439_, new_n2438_, new_n2335_ );
or   ( new_n2440_, new_n2439_, new_n2330_ );
or   ( new_n2441_, new_n2440_, new_n2320_ );
or   ( new_n2442_, new_n2441_, new_n2309_ );
or   ( new_n2443_, new_n2442_, new_n2298_ );
or   ( new_n2444_, new_n2443_, new_n2287_ );
or   ( new_n2445_, new_n2444_, new_n2276_ );
or   ( new_n2446_, new_n2445_, new_n2273_ );
or   ( new_n2447_, new_n2446_, new_n2252_ );
or   ( new_n2448_, new_n2447_, new_n2241_ );
or   ( new_n2449_, new_n2448_, new_n2213_ );
xor  ( new_n2450_, new_n2230_, new_n2227_ );
not  ( new_n2451_, new_n2450_ );
and  ( new_n2452_, new_n2451_, new_n2236_ );
not  ( new_n2453_, new_n2231_ );
and  ( new_n2454_, new_n2237_, new_n2453_ );
nor  ( new_n2455_, new_n2454_, new_n2452_ );
and  ( new_n2456_, new_n2217_, new_n2214_ );
and  ( new_n2457_, new_n2220_, new_n2215_ );
or   ( new_n2458_, new_n2457_, new_n2456_ );
and  ( new_n2459_, new_n2458_, new_n2225_ );
or   ( new_n2460_, new_n2209_, new_n1610_ );
and  ( new_n2461_, new_n2460_, new_n2222_ );
nor  ( new_n2462_, new_n2461_, new_n2459_ );
nor  ( new_n2463_, new_n2462_, new_n2455_ );
and  ( new_n2464_, new_n2460_, new_n2458_ );
or   ( new_n2465_, new_n2464_, new_n2216_ );
and  ( new_n2466_, new_n2465_, new_n2238_ );
and  ( new_n2467_, new_n2225_, new_n2222_ );
or   ( new_n2468_, new_n2467_, new_n2464_ );
and  ( new_n2469_, new_n2468_, new_n2455_ );
or   ( new_n2470_, new_n2469_, new_n2466_ );
or   ( new_n2471_, new_n2470_, new_n2463_ );
or   ( eq, new_n2471_, new_n2449_ );
endmodule


